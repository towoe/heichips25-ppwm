* NGSPICE file created from tiny_wrapper.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

.subckt tiny_wrapper VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7]
X_3155_ net531 VGND VPWR _0049_ sdr_i.mac1.products_ff\[86\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_28_918 VPWR VGND sg13g2_decap_8
X_3086_ net94 VGND VPWR _0277_ ppwm_i.u_ppwm.u_mem.memory\[62\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
X_2106_ _0534_ _1232_ net512 VPWR VGND sg13g2_nand2_1
XFILLER_36_940 VPWR VGND sg13g2_decap_8
X_2037_ net771 _0484_ _0171_ VPWR VGND sg13g2_nor2b_1
XFILLER_11_807 VPWR VGND sg13g2_fill_2
XFILLER_23_667 VPWR VGND sg13g2_decap_4
XFILLER_23_689 VPWR VGND sg13g2_decap_8
X_2939_ net545 VGND VPWR _0130_ sdr_i.DP_4.matrix\[0\] clknet_leaf_16_clk sg13g2_dfrbpq_1
Xhold351 sdr_i.mac2.sum_lvl1_ff\[8\] VPWR VGND net731 sg13g2_dlygate4sd3_1
Xhold362 _0020_ VPWR VGND net742 sg13g2_dlygate4sd3_1
XFILLER_2_538 VPWR VGND sg13g2_decap_8
Xhold340 _0468_ VPWR VGND net720 sg13g2_dlygate4sd3_1
Xhold373 _0514_ VPWR VGND net753 sg13g2_dlygate4sd3_1
Xhold395 _0031_ VPWR VGND net775 sg13g2_dlygate4sd3_1
Xhold384 sdr_i.mac2.sum_lvl2_ff\[4\] VPWR VGND net764 sg13g2_dlygate4sd3_1
XFILLER_46_759 VPWR VGND sg13g2_decap_8
XFILLER_27_940 VPWR VGND sg13g2_decap_8
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_26_74 VPWR VGND sg13g2_fill_1
XFILLER_42_965 VPWR VGND sg13g2_decap_8
XFILLER_41_464 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_fill_1
XFILLER_14_667 VPWR VGND sg13g2_fill_1
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_10_895 VPWR VGND sg13g2_decap_8
XFILLER_6_877 VPWR VGND sg13g2_decap_8
XFILLER_5_343 VPWR VGND sg13g2_fill_2
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_37_726 VPWR VGND sg13g2_fill_1
XFILLER_36_247 VPWR VGND sg13g2_decap_8
XFILLER_17_472 VPWR VGND sg13g2_decap_4
XFILLER_18_995 VPWR VGND sg13g2_decap_8
XFILLER_17_494 VPWR VGND sg13g2_decap_8
XFILLER_33_965 VPWR VGND sg13g2_decap_8
XFILLER_32_453 VPWR VGND sg13g2_fill_2
X_3052__46 VPWR VGND net46 sg13g2_tiehi
X_2998__152 VPWR VGND net152 sg13g2_tiehi
X_2724_ net419 VPWR _1041_ VGND net474 ppwm_i.u_ppwm.u_mem.memory\[87\] sg13g2_o21ai_1
XFILLER_8_192 VPWR VGND sg13g2_decap_8
X_2655_ VGND VPWR net482 _1156_ _0267_ _1006_ sg13g2_a21oi_1
X_1606_ VPWR _1177_ net345 VGND sg13g2_inv_1
X_2586_ net433 VPWR _0972_ VGND net498 net697 sg13g2_o21ai_1
X_1537_ VPWR _1108_ net649 VGND sg13g2_inv_1
X_3207_ net544 VGND VPWR net758 sdr_i.mac2.sum_lvl1_ff\[1\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_28_704 VPWR VGND sg13g2_fill_2
X_3138_ net68 VGND VPWR net718 ppwm_i.u_ppwm.u_mem.bit_count\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_27_214 VPWR VGND sg13g2_decap_8
X_3069_ net162 VGND VPWR net593 ppwm_i.u_ppwm.u_mem.memory\[45\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_24_910 VPWR VGND sg13g2_decap_8
XFILLER_23_464 VPWR VGND sg13g2_fill_1
XFILLER_24_987 VPWR VGND sg13g2_decap_8
XFILLER_6_118 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_3_847 VPWR VGND sg13g2_decap_8
Xhold170 ppwm_i.u_ppwm.u_mem.memory\[27\] VPWR VGND net550 sg13g2_dlygate4sd3_1
Xhold192 ppwm_i.u_ppwm.global_counter\[15\] VPWR VGND net572 sg13g2_dlygate4sd3_1
Xhold181 ppwm_i.u_ppwm.u_mem.memory\[9\] VPWR VGND net561 sg13g2_dlygate4sd3_1
XFILLER_19_704 VPWR VGND sg13g2_fill_1
XFILLER_18_236 VPWR VGND sg13g2_decap_8
XFILLER_34_707 VPWR VGND sg13g2_fill_2
XFILLER_27_781 VPWR VGND sg13g2_decap_8
XFILLER_27_792 VPWR VGND sg13g2_fill_1
XFILLER_14_464 VPWR VGND sg13g2_decap_4
XFILLER_15_976 VPWR VGND sg13g2_decap_8
XFILLER_30_902 VPWR VGND sg13g2_decap_8
XFILLER_14_486 VPWR VGND sg13g2_decap_4
XFILLER_30_979 VPWR VGND sg13g2_decap_8
X_2440_ VGND VPWR _0691_ _0850_ _0855_ _0854_ sg13g2_a21oi_1
XFILLER_6_696 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
X_2371_ _0790_ ppwm_i.u_ppwm.global_counter\[15\] net402 VPWR VGND sg13g2_nand2_1
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_49_361 VPWR VGND sg13g2_fill_1
XFILLER_25_707 VPWR VGND sg13g2_decap_8
XFILLER_18_770 VPWR VGND sg13g2_decap_4
XFILLER_21_968 VPWR VGND sg13g2_decap_8
XFILLER_20_478 VPWR VGND sg13g2_decap_4
X_2707_ VGND VPWR net477 _1130_ _0293_ _1032_ sg13g2_a21oi_1
X_2638_ net426 VPWR _0998_ VGND net481 net356 sg13g2_o21ai_1
X_2569_ VGND VPWR net497 _1199_ _0224_ _0963_ sg13g2_a21oi_1
XFILLER_28_556 VPWR VGND sg13g2_decap_8
XFILLER_43_526 VPWR VGND sg13g2_decap_8
XFILLER_43_515 VPWR VGND sg13g2_fill_1
Xtiny_wrapper_24 VPWR VGND uo_out[4] sg13g2_tielo
XFILLER_43_548 VPWR VGND sg13g2_decap_8
XFILLER_23_261 VPWR VGND sg13g2_decap_8
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_decap_8
XFILLER_7_416 VPWR VGND sg13g2_fill_2
XFILLER_3_622 VPWR VGND sg13g2_decap_8
XFILLER_3_677 VPWR VGND sg13g2_decap_4
Xfanout491 net492 net491 VPWR VGND sg13g2_buf_8
Xfanout480 net501 net480 VPWR VGND sg13g2_buf_2
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_13 VPWR VGND sg13g2_decap_8
XFILLER_46_353 VPWR VGND sg13g2_fill_1
XFILLER_0_68 VPWR VGND sg13g2_decap_8
XFILLER_34_515 VPWR VGND sg13g2_decap_8
XFILLER_34_526 VPWR VGND sg13g2_fill_1
XFILLER_34_537 VPWR VGND sg13g2_fill_1
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_9_22 VPWR VGND sg13g2_fill_2
X_1940_ net736 sdr_i.mac1.sum_lvl1_ff\[9\] _0431_ VPWR VGND sg13g2_xor2_1
XFILLER_30_710 VPWR VGND sg13g2_fill_2
XFILLER_14_294 VPWR VGND sg13g2_decap_8
X_1871_ _0403_ _0402_ _0073_ VPWR VGND sg13g2_xor2_1
XFILLER_9_99 VPWR VGND sg13g2_fill_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
X_2423_ _0839_ ppwm_i.u_ppwm.global_counter\[18\] net402 VPWR VGND sg13g2_nand2_1
XFILLER_9_1024 VPWR VGND sg13g2_decap_4
X_2354_ _0774_ net373 _0773_ VPWR VGND sg13g2_nand2_1
X_2285_ _0708_ ppwm_i.u_ppwm.global_counter\[1\] net398 VPWR VGND sg13g2_nand2_1
XFILLER_49_191 VPWR VGND sg13g2_decap_8
XFILLER_38_854 VPWR VGND sg13g2_decap_8
XFILLER_37_353 VPWR VGND sg13g2_decap_4
XFILLER_21_710 VPWR VGND sg13g2_fill_1
XFILLER_21_721 VPWR VGND sg13g2_decap_4
XFILLER_33_570 VPWR VGND sg13g2_decap_8
XFILLER_5_909 VPWR VGND sg13g2_decap_8
XFILLER_4_419 VPWR VGND sg13g2_decap_8
XFILLER_0_625 VPWR VGND sg13g2_fill_1
XFILLER_0_658 VPWR VGND sg13g2_decap_4
XFILLER_47_128 VPWR VGND sg13g2_fill_1
XFILLER_29_843 VPWR VGND sg13g2_decap_8
XFILLER_44_802 VPWR VGND sg13g2_decap_8
XFILLER_18_97 VPWR VGND sg13g2_decap_4
XFILLER_28_386 VPWR VGND sg13g2_decap_8
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_31_507 VPWR VGND sg13g2_fill_2
XFILLER_15_1018 VPWR VGND sg13g2_decap_8
XFILLER_8_747 VPWR VGND sg13g2_decap_8
XFILLER_8_769 VPWR VGND sg13g2_decap_8
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_47_640 VPWR VGND sg13g2_decap_8
X_2070_ ppwm_i.u_ppwm.u_pwm.counter\[4\] ppwm_i.u_ppwm.u_pwm.counter\[3\] net565 _0506_
+ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[2\] sg13g2_nand4_1
XFILLER_34_323 VPWR VGND sg13g2_decap_8
XFILLER_35_857 VPWR VGND sg13g2_decap_8
XFILLER_22_507 VPWR VGND sg13g2_decap_8
X_2972_ net436 VGND VPWR net573 ppwm_i.u_ppwm.global_counter\[15\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_1923_ net291 sdr_i.mac2.sum_lvl1_ff\[8\] _0013_ VPWR VGND sg13g2_xor2_1
XFILLER_30_540 VPWR VGND sg13g2_fill_1
X_1854_ _0392_ net294 net245 VPWR VGND sg13g2_nand2_1
X_1785_ VPWR VGND _1351_ _1231_ _1349_ _1347_ _1352_ _1348_ sg13g2_a221oi_1
X_2406_ _0823_ _0822_ net376 _0676_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] VPWR VGND
+ sg13g2_a22oi_1
X_2337_ _0757_ _0716_ _0733_ VPWR VGND sg13g2_nand2_1
X_2268_ net396 _0652_ _0691_ VPWR VGND sg13g2_and2_1
XFILLER_38_640 VPWR VGND sg13g2_decap_8
XFILLER_38_662 VPWR VGND sg13g2_decap_4
XFILLER_38_673 VPWR VGND sg13g2_fill_1
XFILLER_26_857 VPWR VGND sg13g2_decap_8
X_2199_ _1229_ _0624_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0625_ VPWR VGND sg13g2_nand3_1
XFILLER_13_507 VPWR VGND sg13g2_decap_8
XFILLER_25_345 VPWR VGND sg13g2_decap_8
XFILLER_40_337 VPWR VGND sg13g2_fill_1
XFILLER_21_540 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_fill_2
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_49_916 VPWR VGND sg13g2_decap_8
Xhold30 sdr_i.mac1.products_ff\[102\] VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_0_466 VPWR VGND sg13g2_decap_8
XFILLER_1_989 VPWR VGND sg13g2_decap_8
Xhold41 sdr_i.DP_2.matrix\[19\] VPWR VGND net241 sg13g2_dlygate4sd3_1
Xhold52 sdr_i.DP_2.matrix\[1\] VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold63 sdr_i.DP_1.matrix\[37\] VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold74 sdr_i.DP_2.matrix\[9\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold96 sdr_i.DP_4.matrix\[9\] VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold85 sdr_i.DP_1.matrix\[9\] VPWR VGND net285 sg13g2_dlygate4sd3_1
XFILLER_29_651 VPWR VGND sg13g2_fill_2
XFILLER_44_610 VPWR VGND sg13g2_fill_2
XFILLER_45_95 VPWR VGND sg13g2_decap_4
XFILLER_31_304 VPWR VGND sg13g2_decap_8
XFILLER_32_849 VPWR VGND sg13g2_decap_8
XFILLER_40_871 VPWR VGND sg13g2_decap_8
XFILLER_8_544 VPWR VGND sg13g2_decap_8
X_1570_ VPWR _1141_ net574 VGND sg13g2_inv_1
XFILLER_6_67 VPWR VGND sg13g2_fill_2
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_3171_ net196 VGND VPWR _0004_ ppwm_i.u_ppwm.mem_write_done clknet_leaf_8_clk sg13g2_dfrbpq_2
X_2122_ _0548_ ppwm_i.u_ppwm.u_ex.state_q\[2\] _0547_ VPWR VGND sg13g2_nand2_1
XFILLER_48_982 VPWR VGND sg13g2_decap_8
XFILLER_47_470 VPWR VGND sg13g2_decap_8
X_2053_ _0495_ _1241_ net410 VPWR VGND sg13g2_nand2_1
XFILLER_19_183 VPWR VGND sg13g2_decap_8
XFILLER_22_315 VPWR VGND sg13g2_decap_8
X_2955_ net533 VGND VPWR _0146_ sdr_i.DP_4.matrix\[72\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2886_ net523 VGND VPWR _0077_ sdr_i.DP_1.matrix\[1\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1906_ net261 sdr_i.mac1.sum_lvl3_ff\[2\] _0030_ VPWR VGND sg13g2_xor2_1
X_1837_ _0381_ sdr_i.total_sum1\[2\] sdr_i.mac2.total_sum\[2\] VPWR VGND sg13g2_xnor2_1
X_1768_ _1335_ net448 _1180_ net453 _1159_ VPWR VGND sg13g2_a22oi_1
X_1699_ VGND VPWR _1235_ _1267_ _0003_ _1268_ sg13g2_a21oi_1
XFILLER_39_960 VPWR VGND sg13g2_decap_8
XFILLER_14_805 VPWR VGND sg13g2_decap_8
XFILLER_25_120 VPWR VGND sg13g2_decap_8
XFILLER_40_101 VPWR VGND sg13g2_decap_8
XFILLER_5_514 VPWR VGND sg13g2_fill_2
XFILLER_31_42 VPWR VGND sg13g2_decap_8
Xoutput7 net7 uio_oe[3] VPWR VGND sg13g2_buf_1
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_1_786 VPWR VGND sg13g2_decap_8
XFILLER_0_285 VPWR VGND sg13g2_decap_4
XFILLER_45_996 VPWR VGND sg13g2_decap_8
X_3049__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_13_871 VPWR VGND sg13g2_decap_8
XFILLER_31_145 VPWR VGND sg13g2_fill_1
X_2740_ net414 VPWR _1049_ VGND net468 net597 sg13g2_o21ai_1
X_2671_ VGND VPWR net465 _1148_ _0275_ _1014_ sg13g2_a21oi_1
XFILLER_8_385 VPWR VGND sg13g2_fill_1
X_1622_ VPWR _1193_ net646 VGND sg13g2_inv_1
X_1553_ VPWR _1124_ net358 VGND sg13g2_inv_1
X_3223_ net532 VGND VPWR net211 sdr_i.mac2.sum_lvl2_ff\[8\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3154_ net531 VGND VPWR _0048_ sdr_i.mac1.products_ff\[85\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_3085_ net98 VGND VPWR _0276_ ppwm_i.u_ppwm.u_mem.memory\[61\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_2105_ _0533_ net511 net451 VPWR VGND sg13g2_xnor2_1
X_2036_ VGND VPWR _1245_ net409 _0484_ net456 sg13g2_a21oi_1
XFILLER_36_996 VPWR VGND sg13g2_decap_8
XFILLER_23_646 VPWR VGND sg13g2_decap_8
X_2938_ net527 VGND VPWR _0129_ sdr_i.DP_3.matrix\[73\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2869_ net296 _0132_ VPWR VGND sg13g2_buf_1
XFILLER_11_1021 VPWR VGND sg13g2_decap_8
Xhold352 _0014_ VPWR VGND net732 sg13g2_dlygate4sd3_1
XFILLER_7_8 VPWR VGND sg13g2_fill_1
Xhold341 _0160_ VPWR VGND net721 sg13g2_dlygate4sd3_1
Xhold330 ppwm_i.u_ppwm.global_counter\[2\] VPWR VGND net710 sg13g2_dlygate4sd3_1
Xhold363 sdr_i.mac1.sum_lvl2_ff\[1\] VPWR VGND net743 sg13g2_dlygate4sd3_1
Xhold374 sdr_i.mac2.products_ff\[69\] VPWR VGND net754 sg13g2_dlygate4sd3_1
Xhold385 _0010_ VPWR VGND net765 sg13g2_dlygate4sd3_1
Xhold396 ppwm_i.u_ppwm.global_counter\[13\] VPWR VGND net776 sg13g2_dlygate4sd3_1
XFILLER_18_429 VPWR VGND sg13g2_decap_8
XFILLER_26_462 VPWR VGND sg13g2_fill_1
XFILLER_26_473 VPWR VGND sg13g2_decap_8
XFILLER_27_996 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_944 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_fill_2
XFILLER_14_679 VPWR VGND sg13g2_decap_8
XFILLER_42_30 VPWR VGND sg13g2_fill_1
XFILLER_10_830 VPWR VGND sg13g2_fill_1
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_10_874 VPWR VGND sg13g2_decap_8
XFILLER_6_856 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_1_594 VPWR VGND sg13g2_decap_8
XFILLER_49_576 VPWR VGND sg13g2_fill_1
XFILLER_3_1008 VPWR VGND sg13g2_decap_8
XFILLER_37_705 VPWR VGND sg13g2_decap_8
XFILLER_18_974 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
XFILLER_44_270 VPWR VGND sg13g2_fill_2
XFILLER_33_944 VPWR VGND sg13g2_decap_8
X_2723_ VGND VPWR net475 _1122_ _0301_ _1040_ sg13g2_a21oi_1
XFILLER_8_171 VPWR VGND sg13g2_decap_8
XFILLER_9_672 VPWR VGND sg13g2_fill_1
X_2654_ net425 VPWR _1006_ VGND net482 net657 sg13g2_o21ai_1
X_1605_ VPWR _1176_ net688 VGND sg13g2_inv_1
X_2585_ VGND VPWR net486 _1191_ _0232_ _0971_ sg13g2_a21oi_1
X_1536_ VPWR _1107_ net625 VGND sg13g2_inv_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
X_3206_ net544 VGND VPWR net255 sdr_i.mac2.sum_lvl1_ff\[0\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3137_ net100 VGND VPWR net341 ppwm_i.u_ppwm.u_mem.bit_count\[1\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_28_727 VPWR VGND sg13g2_fill_1
X_3068_ net166 VGND VPWR _0259_ ppwm_i.u_ppwm.u_mem.memory\[44\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
X_2019_ _0165_ _1253_ _0472_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_421 VPWR VGND sg13g2_fill_2
XFILLER_36_793 VPWR VGND sg13g2_decap_8
XFILLER_24_966 VPWR VGND sg13g2_decap_8
XFILLER_11_649 VPWR VGND sg13g2_fill_2
XFILLER_10_137 VPWR VGND sg13g2_fill_1
XFILLER_7_609 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
X_3003__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_12_77 VPWR VGND sg13g2_decap_8
XFILLER_3_826 VPWR VGND sg13g2_decap_8
Xhold160 ppwm_i.u_ppwm.u_mem.memory\[31\] VPWR VGND net360 sg13g2_dlygate4sd3_1
X_3114__104 VPWR VGND net104 sg13g2_tiehi
Xhold171 _0241_ VPWR VGND net551 sg13g2_dlygate4sd3_1
Xhold193 _0163_ VPWR VGND net573 sg13g2_dlygate4sd3_1
XFILLER_2_369 VPWR VGND sg13g2_fill_1
Xhold182 _0223_ VPWR VGND net562 sg13g2_dlygate4sd3_1
XFILLER_18_215 VPWR VGND sg13g2_decap_8
XFILLER_19_727 VPWR VGND sg13g2_decap_4
XFILLER_19_738 VPWR VGND sg13g2_fill_2
XFILLER_37_41 VPWR VGND sg13g2_decap_8
XFILLER_37_30 VPWR VGND sg13g2_fill_2
XFILLER_46_568 VPWR VGND sg13g2_fill_1
XFILLER_46_557 VPWR VGND sg13g2_decap_8
XFILLER_14_421 VPWR VGND sg13g2_fill_2
XFILLER_15_955 VPWR VGND sg13g2_decap_8
XFILLER_18_1016 VPWR VGND sg13g2_decap_8
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_30_958 VPWR VGND sg13g2_decap_8
XFILLER_6_620 VPWR VGND sg13g2_decap_8
XFILLER_6_675 VPWR VGND sg13g2_decap_8
X_2370_ VPWR VGND _0783_ _0788_ _0782_ net379 _0789_ _0746_ sg13g2_a221oi_1
XFILLER_21_947 VPWR VGND sg13g2_decap_8
X_2706_ net417 VPWR _1032_ VGND net477 ppwm_i.u_ppwm.u_mem.memory\[78\] sg13g2_o21ai_1
X_2637_ VGND VPWR net488 _1165_ _0258_ _0997_ sg13g2_a21oi_1
XFILLER_0_829 VPWR VGND sg13g2_decap_8
X_2568_ net431 VPWR _0963_ VGND net489 net561 sg13g2_o21ai_1
X_2499_ _0908_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] net393 VPWR VGND sg13g2_xnor2_1
Xtiny_wrapper_25 VPWR VGND uo_out[5] sg13g2_tielo
XFILLER_15_207 VPWR VGND sg13g2_decap_8
XFILLER_11_402 VPWR VGND sg13g2_fill_1
XFILLER_12_947 VPWR VGND sg13g2_decap_8
XFILLER_24_796 VPWR VGND sg13g2_fill_2
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_7_439 VPWR VGND sg13g2_fill_1
XFILLER_11_468 VPWR VGND sg13g2_decap_8
XFILLER_3_2 VPWR VGND sg13g2_fill_1
XFILLER_47_833 VPWR VGND sg13g2_decap_8
Xfanout481 net482 net481 VPWR VGND sg13g2_buf_8
Xfanout470 net501 net470 VPWR VGND sg13g2_buf_2
Xfanout492 net496 net492 VPWR VGND sg13g2_buf_8
XFILLER_0_36 VPWR VGND sg13g2_fill_2
XFILLER_14_273 VPWR VGND sg13g2_decap_4
XFILLER_42_593 VPWR VGND sg13g2_decap_8
X_1870_ _0403_ net272 net224 VPWR VGND sg13g2_nand2_1
XFILLER_31_1024 VPWR VGND sg13g2_decap_4
XFILLER_7_962 VPWR VGND sg13g2_decap_8
XFILLER_6_472 VPWR VGND sg13g2_decap_4
XFILLER_6_450 VPWR VGND sg13g2_fill_1
X_2422_ _0838_ _0836_ _0837_ _0806_ _0653_ VPWR VGND sg13g2_a22oi_1
XFILLER_9_1003 VPWR VGND sg13g2_decap_8
X_2353_ _0773_ _0772_ net376 net375 net818 VPWR VGND sg13g2_a22oi_1
X_2284_ net385 _0674_ _0707_ VPWR VGND sg13g2_nor2_1
XFILLER_49_170 VPWR VGND sg13g2_decap_8
XFILLER_38_833 VPWR VGND sg13g2_decap_8
XFILLER_25_505 VPWR VGND sg13g2_decap_8
XFILLER_37_387 VPWR VGND sg13g2_fill_2
XFILLER_40_519 VPWR VGND sg13g2_decap_4
XFILLER_33_582 VPWR VGND sg13g2_decap_8
XFILLER_21_744 VPWR VGND sg13g2_decap_4
XFILLER_21_788 VPWR VGND sg13g2_fill_2
X_1999_ _0462_ net654 _0155_ VPWR VGND sg13g2_xor2_1
XFILLER_20_276 VPWR VGND sg13g2_decap_8
XFILLER_0_604 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_47_107 VPWR VGND sg13g2_decap_8
XFILLER_29_822 VPWR VGND sg13g2_decap_8
XFILLER_28_365 VPWR VGND sg13g2_decap_8
XFILLER_29_899 VPWR VGND sg13g2_decap_8
XFILLER_44_858 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_4
XFILLER_12_711 VPWR VGND sg13g2_decap_4
XFILLER_11_210 VPWR VGND sg13g2_fill_2
XFILLER_34_75 VPWR VGND sg13g2_decap_4
XFILLER_11_298 VPWR VGND sg13g2_decap_8
XFILLER_3_420 VPWR VGND sg13g2_fill_2
XFILLER_4_965 VPWR VGND sg13g2_decap_8
XFILLER_38_107 VPWR VGND sg13g2_fill_2
XFILLER_46_140 VPWR VGND sg13g2_fill_2
XFILLER_35_836 VPWR VGND sg13g2_decap_8
XFILLER_43_880 VPWR VGND sg13g2_decap_8
X_2971_ net437 VGND VPWR _0162_ ppwm_i.u_ppwm.global_counter\[14\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_42_390 VPWR VGND sg13g2_fill_1
X_1922_ _0422_ net731 net291 VPWR VGND sg13g2_nand2_1
XFILLER_15_593 VPWR VGND sg13g2_decap_8
X_1853_ _0391_ _0390_ _0059_ VPWR VGND sg13g2_xor2_1
X_3103__191 VPWR VGND net191 sg13g2_tiehi
X_1784_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[104\] _1350_ net438 ppwm_i.u_ppwm.u_mem.memory\[97\]
+ _1351_ net442 sg13g2_a221oi_1
X_2405_ ppwm_i.u_ppwm.global_counter\[17\] ppwm_i.u_ppwm.global_counter\[7\] net399
+ _0822_ VPWR VGND sg13g2_mux2_1
XFILLER_41_0 VPWR VGND sg13g2_fill_2
X_2336_ _0714_ _0716_ _0733_ _0734_ _0756_ VPWR VGND sg13g2_and4_1
X_2267_ net457 _0688_ _0690_ _0195_ VPWR VGND sg13g2_nor3_1
XFILLER_26_825 VPWR VGND sg13g2_fill_2
XFILLER_26_836 VPWR VGND sg13g2_decap_8
X_2198_ _0624_ net507 ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] VPWR VGND sg13g2_nand2b_1
XFILLER_38_685 VPWR VGND sg13g2_fill_2
XFILLER_38_1008 VPWR VGND sg13g2_decap_8
XFILLER_25_379 VPWR VGND sg13g2_decap_8
XFILLER_40_349 VPWR VGND sg13g2_decap_8
XFILLER_5_707 VPWR VGND sg13g2_decap_4
XFILLER_4_206 VPWR VGND sg13g2_fill_2
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_20_22 VPWR VGND sg13g2_fill_2
XFILLER_0_423 VPWR VGND sg13g2_decap_4
XFILLER_1_968 VPWR VGND sg13g2_decap_8
XFILLER_29_20 VPWR VGND sg13g2_fill_2
Xhold31 _0021_ VPWR VGND net231 sg13g2_dlygate4sd3_1
Xhold20 sdr_i.DP_1.matrix\[10\] VPWR VGND net220 sg13g2_dlygate4sd3_1
Xhold64 sdr_i.DP_1.matrix\[55\] VPWR VGND net264 sg13g2_dlygate4sd3_1
XFILLER_29_75 VPWR VGND sg13g2_decap_8
Xhold42 sdr_i.DP_3.matrix\[55\] VPWR VGND net242 sg13g2_dlygate4sd3_1
Xhold53 sdr_i.DP_4.matrix\[64\] VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold86 sdr_i.DP_2.matrix\[63\] VPWR VGND net286 sg13g2_dlygate4sd3_1
XFILLER_17_803 VPWR VGND sg13g2_decap_8
Xhold75 sdr_i.DP_2.matrix\[27\] VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold97 sdr_i.mac2.sum_lvl2_ff\[0\] VPWR VGND net297 sg13g2_dlygate4sd3_1
XFILLER_29_685 VPWR VGND sg13g2_decap_8
X_2985__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_45_74 VPWR VGND sg13g2_decap_8
XFILLER_16_335 VPWR VGND sg13g2_decap_8
XFILLER_17_858 VPWR VGND sg13g2_decap_4
XFILLER_44_699 VPWR VGND sg13g2_fill_1
XFILLER_25_880 VPWR VGND sg13g2_decap_8
XFILLER_32_828 VPWR VGND sg13g2_decap_8
XFILLER_24_390 VPWR VGND sg13g2_decap_4
XFILLER_40_850 VPWR VGND sg13g2_decap_8
XFILLER_3_272 VPWR VGND sg13g2_decap_4
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1017 VPWR VGND sg13g2_decap_8
X_3170_ net195 VGND VPWR _0003_ ppwm_i.u_ppwm.u_mem.state_q\[0\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_0_990 VPWR VGND sg13g2_decap_8
X_2121_ net395 _0365_ _0547_ VPWR VGND sg13g2_and2_1
XFILLER_48_961 VPWR VGND sg13g2_decap_8
X_2052_ net456 net803 _0176_ VPWR VGND sg13g2_nor2_1
XFILLER_47_460 VPWR VGND sg13g2_fill_1
XFILLER_35_644 VPWR VGND sg13g2_decap_4
XFILLER_22_305 VPWR VGND sg13g2_fill_1
X_2954_ net538 VGND VPWR _0145_ sdr_i.DP_4.matrix\[64\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2885_ net523 VGND VPWR _0076_ sdr_i.DP_1.matrix\[0\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1905_ _0412_ net774 net261 VPWR VGND sg13g2_nand2_1
X_1836_ _0380_ sdr_i.total_sum1\[2\] sdr_i.mac2.total_sum\[2\] VPWR VGND sg13g2_nand2_1
X_1767_ VPWR VGND _1194_ _1332_ net440 _1201_ _1334_ net444 sg13g2_a221oi_1
X_1698_ net3 net324 net457 _1268_ VPWR VGND sg13g2_nor3_1
XFILLER_44_1012 VPWR VGND sg13g2_decap_8
X_2319_ _0740_ net390 net386 VPWR VGND sg13g2_nand2_1
XFILLER_26_600 VPWR VGND sg13g2_decap_4
XFILLER_26_611 VPWR VGND sg13g2_fill_2
XFILLER_38_460 VPWR VGND sg13g2_fill_1
XFILLER_26_677 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_8
XFILLER_41_636 VPWR VGND sg13g2_decap_8
XFILLER_15_55 VPWR VGND sg13g2_decap_8
XFILLER_40_157 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_21_393 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_oe[4] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_oe[6] VPWR VGND sg13g2_buf_1
X_3013__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_1_765 VPWR VGND sg13g2_decap_8
XFILLER_49_769 VPWR VGND sg13g2_decap_8
XFILLER_48_279 VPWR VGND sg13g2_decap_4
XFILLER_29_482 VPWR VGND sg13g2_decap_4
XFILLER_29_493 VPWR VGND sg13g2_fill_2
XFILLER_45_975 VPWR VGND sg13g2_decap_8
XFILLER_44_463 VPWR VGND sg13g2_decap_8
XFILLER_44_452 VPWR VGND sg13g2_fill_1
XFILLER_17_677 VPWR VGND sg13g2_decap_8
XFILLER_31_102 VPWR VGND sg13g2_decap_8
XFILLER_13_850 VPWR VGND sg13g2_fill_1
XFILLER_9_843 VPWR VGND sg13g2_fill_2
X_2670_ net412 VPWR _1014_ VGND net465 ppwm_i.u_ppwm.u_mem.memory\[60\] sg13g2_o21ai_1
XFILLER_9_898 VPWR VGND sg13g2_decap_8
X_1621_ VPWR _1192_ net352 VGND sg13g2_inv_1
X_1552_ VPWR _1123_ net634 VGND sg13g2_inv_1
X_3222_ net200 VGND VPWR _0002_ ppwm_i.u_ppwm.u_ex.state_q\[2\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
X_3153_ net529 VGND VPWR _0059_ sdr_i.mac1.products_ff\[69\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_2104_ _0532_ net511 net389 VPWR VGND sg13g2_xnor2_1
X_3084_ net102 VGND VPWR net591 ppwm_i.u_ppwm.u_mem.memory\[60\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_2035_ net770 net411 _0483_ VPWR VGND sg13g2_nor2_1
XFILLER_35_474 VPWR VGND sg13g2_decap_8
XFILLER_36_975 VPWR VGND sg13g2_decap_8
XFILLER_23_636 VPWR VGND sg13g2_decap_4
XFILLER_35_485 VPWR VGND sg13g2_fill_1
XFILLER_11_809 VPWR VGND sg13g2_fill_1
XFILLER_22_146 VPWR VGND sg13g2_decap_8
XFILLER_22_157 VPWR VGND sg13g2_fill_2
X_2937_ net533 VGND VPWR _0128_ sdr_i.DP_3.matrix\[72\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_31_691 VPWR VGND sg13g2_fill_1
X_2868_ net247 _0131_ VPWR VGND sg13g2_buf_1
XFILLER_11_1000 VPWR VGND sg13g2_decap_8
Xhold320 ppwm_i.u_ppwm.u_mem.memory\[81\] VPWR VGND net700 sg13g2_dlygate4sd3_1
X_1819_ _0368_ _0367_ _1279_ VPWR VGND sg13g2_nand2b_1
X_2799_ _1084_ _1246_ ppwm_i.u_ppwm.u_pwm.counter\[2\] _1245_ ppwm_i.u_ppwm.u_pwm.counter\[3\]
+ VPWR VGND sg13g2_a22oi_1
Xhold353 ppwm_i.u_ppwm.u_mem.memory\[21\] VPWR VGND net733 sg13g2_dlygate4sd3_1
Xhold331 _0150_ VPWR VGND net711 sg13g2_dlygate4sd3_1
Xhold342 sdr_i.mac2.sum_lvl1_ff\[17\] VPWR VGND net722 sg13g2_dlygate4sd3_1
Xhold386 ppwm_i.u_ppwm.u_pwm.counter\[8\] VPWR VGND net766 sg13g2_dlygate4sd3_1
Xhold364 _0435_ VPWR VGND net744 sg13g2_dlygate4sd3_1
Xhold375 _0409_ VPWR VGND net755 sg13g2_dlygate4sd3_1
Xhold397 _0161_ VPWR VGND net777 sg13g2_dlygate4sd3_1
XFILLER_19_909 VPWR VGND sg13g2_decap_8
XFILLER_46_728 VPWR VGND sg13g2_fill_2
XFILLER_45_249 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_42_923 VPWR VGND sg13g2_decap_8
XFILLER_14_603 VPWR VGND sg13g2_decap_4
XFILLER_27_975 VPWR VGND sg13g2_decap_8
XFILLER_41_422 VPWR VGND sg13g2_decap_8
XFILLER_14_636 VPWR VGND sg13g2_decap_8
XFILLER_41_499 VPWR VGND sg13g2_fill_1
XFILLER_6_835 VPWR VGND sg13g2_decap_8
XFILLER_5_345 VPWR VGND sg13g2_fill_1
XFILLER_3_69 VPWR VGND sg13g2_decap_8
XFILLER_1_573 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_18_953 VPWR VGND sg13g2_decap_8
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_33_923 VPWR VGND sg13g2_decap_8
XFILLER_32_411 VPWR VGND sg13g2_decap_4
XFILLER_32_488 VPWR VGND sg13g2_fill_1
XFILLER_34_1022 VPWR VGND sg13g2_decap_8
X_2722_ net419 VPWR _1040_ VGND net475 ppwm_i.u_ppwm.u_mem.memory\[86\] sg13g2_o21ai_1
X_2653_ VGND VPWR net481 _1157_ _0266_ _1005_ sg13g2_a21oi_1
X_1604_ VPWR _1175_ net675 VGND sg13g2_inv_1
X_2584_ net427 VPWR _0971_ VGND net486 net352 sg13g2_o21ai_1
X_1535_ VPWR _1106_ net594 VGND sg13g2_inv_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
X_3205_ net542 VGND VPWR _0071_ sdr_i.mac2.products_ff\[137\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_706 VPWR VGND sg13g2_fill_1
X_3136_ net131 VGND VPWR _0327_ ppwm_i.u_ppwm.u_mem.bit_count\[0\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
XFILLER_28_739 VPWR VGND sg13g2_decap_8
X_3067_ net170 VGND VPWR net357 ppwm_i.u_ppwm.u_mem.memory\[43\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2018_ _0164_ _1254_ _0471_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_945 VPWR VGND sg13g2_decap_8
XFILLER_23_433 VPWR VGND sg13g2_fill_2
XFILLER_35_293 VPWR VGND sg13g2_decap_8
XFILLER_11_617 VPWR VGND sg13g2_fill_2
XFILLER_10_127 VPWR VGND sg13g2_fill_2
XFILLER_3_805 VPWR VGND sg13g2_decap_8
Xhold161 _0245_ VPWR VGND net361 sg13g2_dlygate4sd3_1
Xhold150 _0550_ VPWR VGND net350 sg13g2_dlygate4sd3_1
Xhold194 ppwm_i.u_ppwm.u_mem.memory\[68\] VPWR VGND net574 sg13g2_dlygate4sd3_1
Xhold183 ppwm_i.u_ppwm.u_mem.memory\[58\] VPWR VGND net563 sg13g2_dlygate4sd3_1
Xhold172 sdr_i.mac1.sum_lvl3_ff\[3\] VPWR VGND net552 sg13g2_dlygate4sd3_1
XFILLER_37_20 VPWR VGND sg13g2_fill_1
XFILLER_46_536 VPWR VGND sg13g2_fill_1
XFILLER_34_709 VPWR VGND sg13g2_fill_1
XFILLER_15_934 VPWR VGND sg13g2_decap_8
XFILLER_42_797 VPWR VGND sg13g2_decap_8
XFILLER_30_937 VPWR VGND sg13g2_decap_8
XFILLER_6_654 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_fill_1
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_37_503 VPWR VGND sg13g2_fill_2
XFILLER_37_547 VPWR VGND sg13g2_decap_8
XFILLER_17_271 VPWR VGND sg13g2_decap_8
XFILLER_32_230 VPWR VGND sg13g2_fill_2
XFILLER_32_241 VPWR VGND sg13g2_fill_2
XFILLER_33_753 VPWR VGND sg13g2_decap_4
XFILLER_21_926 VPWR VGND sg13g2_decap_8
XFILLER_33_797 VPWR VGND sg13g2_decap_8
XFILLER_32_285 VPWR VGND sg13g2_decap_8
XFILLER_32_296 VPWR VGND sg13g2_fill_2
X_2705_ VGND VPWR net478 _1131_ _0292_ _1031_ sg13g2_a21oi_1
X_2636_ net430 VPWR _0997_ VGND net488 ppwm_i.u_ppwm.u_mem.memory\[43\] sg13g2_o21ai_1
XFILLER_0_808 VPWR VGND sg13g2_decap_8
X_2567_ VGND VPWR net495 _1200_ _0223_ _0962_ sg13g2_a21oi_1
X_2498_ _0906_ _0907_ _0209_ VPWR VGND sg13g2_nor2_1
XFILLER_28_514 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_26 VPWR VGND uo_out[6] sg13g2_tielo
X_3119_ net64 VGND VPWR _0310_ ppwm_i.u_ppwm.u_mem.memory\[95\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_12_926 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_11_447 VPWR VGND sg13g2_fill_2
XFILLER_2_178 VPWR VGND sg13g2_decap_4
XFILLER_47_812 VPWR VGND sg13g2_decap_8
Xfanout482 net486 net482 VPWR VGND sg13g2_buf_8
Xfanout460 _1233_ net460 VPWR VGND sg13g2_buf_8
Xfanout493 net496 net493 VPWR VGND sg13g2_buf_8
Xfanout471 net472 net471 VPWR VGND sg13g2_buf_8
XFILLER_19_525 VPWR VGND sg13g2_decap_4
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_27_580 VPWR VGND sg13g2_fill_2
XFILLER_15_764 VPWR VGND sg13g2_fill_1
XFILLER_14_252 VPWR VGND sg13g2_decap_8
XFILLER_30_712 VPWR VGND sg13g2_fill_1
XFILLER_31_1003 VPWR VGND sg13g2_decap_8
XFILLER_7_941 VPWR VGND sg13g2_decap_8
X_2995__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_6_462 VPWR VGND sg13g2_decap_4
X_2421_ VPWR VGND _0350_ _0692_ _0744_ _0661_ _0837_ _0739_ sg13g2_a221oi_1
X_2352_ _0771_ VPWR _0772_ VGND _1263_ net403 sg13g2_o21ai_1
X_2283_ _0705_ VPWR _0706_ VGND _0687_ _0704_ sg13g2_o21ai_1
XFILLER_38_812 VPWR VGND sg13g2_decap_8
X_3097__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_38_889 VPWR VGND sg13g2_decap_8
XFILLER_37_377 VPWR VGND sg13g2_decap_8
XFILLER_37_399 VPWR VGND sg13g2_decap_8
X_1998_ _0154_ net320 _0461_ VPWR VGND sg13g2_xnor2_1
X_2619_ VGND VPWR net487 _1174_ _0249_ _0988_ sg13g2_a21oi_1
XFILLER_29_801 VPWR VGND sg13g2_decap_8
XFILLER_29_878 VPWR VGND sg13g2_decap_8
XFILLER_44_837 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_11_244 VPWR VGND sg13g2_decap_8
XFILLER_7_248 VPWR VGND sg13g2_fill_2
XFILLER_4_944 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_15_8 VPWR VGND sg13g2_fill_1
XFILLER_35_815 VPWR VGND sg13g2_decap_8
XFILLER_46_185 VPWR VGND sg13g2_decap_4
XFILLER_34_358 VPWR VGND sg13g2_decap_8
XFILLER_15_572 VPWR VGND sg13g2_decap_8
X_2970_ net437 VGND VPWR net777 ppwm_i.u_ppwm.global_counter\[13\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_1921_ _0010_ _0420_ _0421_ VPWR VGND sg13g2_xnor2_1
X_1852_ _0391_ net295 net249 VPWR VGND sg13g2_nand2_1
XFILLER_30_575 VPWR VGND sg13g2_decap_8
X_1783_ _1350_ ppwm_i.u_ppwm.u_mem.memory\[111\] net515 net518 VPWR VGND sg13g2_and3_1
XFILLER_6_292 VPWR VGND sg13g2_decap_8
X_2404_ _0821_ _0819_ _0820_ _0787_ net379 VPWR VGND sg13g2_a22oi_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_2335_ _0755_ net505 net391 VPWR VGND sg13g2_xnor2_1
X_2266_ _0669_ _0677_ net371 _0689_ _0690_ VPWR VGND sg13g2_and4_1
X_2197_ net385 VPWR _0623_ VGND _0605_ _0622_ sg13g2_o21ai_1
XFILLER_26_804 VPWR VGND sg13g2_decap_8
XFILLER_37_141 VPWR VGND sg13g2_decap_4
XFILLER_41_829 VPWR VGND sg13g2_decap_8
X_3085__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_33_380 VPWR VGND sg13g2_decap_4
XFILLER_21_597 VPWR VGND sg13g2_decap_8
XFILLER_20_34 VPWR VGND sg13g2_fill_1
XFILLER_0_402 VPWR VGND sg13g2_decap_8
XFILLER_0_446 VPWR VGND sg13g2_decap_8
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold21 sdr_i.DP_1.matrix\[64\] VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold32 sdr_i.DP_1.matrix\[73\] VPWR VGND net232 sg13g2_dlygate4sd3_1
Xhold10 sdr_i.mac1.sum_lvl2_ff\[8\] VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold54 sdr_i.mac2.products_ff\[0\] VPWR VGND net254 sg13g2_dlygate4sd3_1
XFILLER_29_631 VPWR VGND sg13g2_fill_1
Xhold43 sdr_i.DP_3.matrix\[46\] VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold65 sdr_i.mac2.products_ff\[68\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold76 sdr_i.DP_1.matrix\[0\] VPWR VGND net276 sg13g2_dlygate4sd3_1
Xhold87 sdr_i.DP_2.matrix\[0\] VPWR VGND net287 sg13g2_dlygate4sd3_1
XFILLER_21_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_653 VPWR VGND sg13g2_fill_1
XFILLER_29_664 VPWR VGND sg13g2_decap_8
Xhold98 _0009_ VPWR VGND net298 sg13g2_dlygate4sd3_1
XFILLER_44_612 VPWR VGND sg13g2_fill_1
XFILLER_45_42 VPWR VGND sg13g2_decap_4
XFILLER_44_645 VPWR VGND sg13g2_fill_1
XFILLER_44_634 VPWR VGND sg13g2_decap_8
XFILLER_32_807 VPWR VGND sg13g2_decap_8
XFILLER_44_678 VPWR VGND sg13g2_decap_8
XFILLER_43_166 VPWR VGND sg13g2_decap_4
XFILLER_31_339 VPWR VGND sg13g2_decap_8
XFILLER_8_524 VPWR VGND sg13g2_fill_2
XFILLER_6_69 VPWR VGND sg13g2_fill_1
XFILLER_3_251 VPWR VGND sg13g2_decap_8
XFILLER_48_940 VPWR VGND sg13g2_decap_8
X_2120_ net458 _0546_ _0192_ VPWR VGND sg13g2_nor2_1
X_2051_ _0493_ VPWR _0494_ VGND ppwm_i.u_ppwm.pwm_value\[8\] net410 sg13g2_o21ai_1
XFILLER_23_829 VPWR VGND sg13g2_decap_4
XFILLER_35_667 VPWR VGND sg13g2_decap_4
XFILLER_16_892 VPWR VGND sg13g2_decap_8
XFILLER_34_177 VPWR VGND sg13g2_fill_1
X_2953_ net538 VGND VPWR _0144_ sdr_i.DP_4.matrix\[63\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1904_ net272 net284 _0072_ VPWR VGND sg13g2_and2_1
X_2884_ net246 _0147_ VPWR VGND sg13g2_buf_1
XFILLER_30_383 VPWR VGND sg13g2_decap_8
XFILLER_31_884 VPWR VGND sg13g2_decap_8
X_1835_ VGND VPWR _0379_ net13 _0377_ _0374_ sg13g2_a21oi_2
X_1766_ VGND VPWR _1187_ net453 _1333_ net512 sg13g2_a21oi_1
XFILLER_7_590 VPWR VGND sg13g2_decap_8
X_1697_ _1098_ net457 _1267_ VPWR VGND sg13g2_nor2_1
X_2318_ net392 net384 _0739_ VPWR VGND sg13g2_nor2_2
X_2249_ _0551_ _0672_ _0673_ VPWR VGND sg13g2_nor2_2
XFILLER_39_995 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_25_155 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_21_372 VPWR VGND sg13g2_decap_8
XFILLER_22_884 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_decap_8
Xoutput9 net9 uio_oe[5] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_oe[7] VPWR VGND sg13g2_buf_1
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_0_232 VPWR VGND sg13g2_decap_8
XFILLER_49_748 VPWR VGND sg13g2_decap_8
XFILLER_48_258 VPWR VGND sg13g2_decap_8
XFILLER_36_409 VPWR VGND sg13g2_fill_2
XFILLER_17_612 VPWR VGND sg13g2_fill_2
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_44_497 VPWR VGND sg13g2_fill_2
XFILLER_44_486 VPWR VGND sg13g2_decap_8
XFILLER_16_177 VPWR VGND sg13g2_fill_2
XFILLER_16_199 VPWR VGND sg13g2_fill_1
XFILLER_9_833 VPWR VGND sg13g2_fill_1
XFILLER_9_877 VPWR VGND sg13g2_decap_8
X_1620_ VPWR _1191_ net697 VGND sg13g2_inv_1
X_1551_ VPWR _1122_ net368 VGND sg13g2_inv_1
XFILLER_4_582 VPWR VGND sg13g2_fill_1
XFILLER_4_571 VPWR VGND sg13g2_decap_8
X_3221_ net199 VGND VPWR net319 ppwm_i.u_ppwm.u_ex.state_q\[1\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3152_ net529 VGND VPWR _0058_ sdr_i.mac1.products_ff\[68\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_39_203 VPWR VGND sg13g2_decap_4
X_2103_ _0531_ net511 net389 VPWR VGND sg13g2_nand2_1
X_3083_ net106 VGND VPWR net620 ppwm_i.u_ppwm.u_mem.memory\[59\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_39_269 VPWR VGND sg13g2_decap_8
X_2034_ _0481_ _0482_ _0170_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_954 VPWR VGND sg13g2_decap_8
X_2936_ net538 VGND VPWR _0127_ sdr_i.DP_3.matrix\[64\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2867_ net280 _0130_ VPWR VGND sg13g2_buf_1
X_1818_ _0367_ _0366_ _1312_ VPWR VGND sg13g2_nand2b_1
Xhold310 ppwm_i.u_ppwm.u_mem.state_q\[2\] VPWR VGND net690 sg13g2_dlygate4sd3_1
X_2798_ _1082_ VPWR _1083_ VGND ppwm_i.u_ppwm.u_pwm.counter\[2\] _1246_ sg13g2_o21ai_1
Xhold321 _0296_ VPWR VGND net701 sg13g2_dlygate4sd3_1
X_1749_ _1316_ net438 _1139_ net442 _1146_ VPWR VGND sg13g2_a22oi_1
Xhold332 ppwm_i.u_ppwm.polarity VPWR VGND net712 sg13g2_dlygate4sd3_1
Xhold343 _0441_ VPWR VGND net723 sg13g2_dlygate4sd3_1
Xhold387 _0512_ VPWR VGND net767 sg13g2_dlygate4sd3_1
Xhold365 _0028_ VPWR VGND net745 sg13g2_dlygate4sd3_1
Xhold354 sdr_i.mac1.products_ff\[0\] VPWR VGND net734 sg13g2_dlygate4sd3_1
Xhold376 _0037_ VPWR VGND net756 sg13g2_dlygate4sd3_1
X_3419_ net549 net6 VPWR VGND sg13g2_buf_1
Xhold398 sdr_i.mac1.products_ff\[51\] VPWR VGND net778 sg13g2_dlygate4sd3_1
XFILLER_39_792 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_27_954 VPWR VGND sg13g2_decap_8
XFILLER_42_902 VPWR VGND sg13g2_decap_8
X_3082__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_26_453 VPWR VGND sg13g2_decap_8
XFILLER_42_979 VPWR VGND sg13g2_decap_8
X_3046__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_42_43 VPWR VGND sg13g2_decap_8
XFILLER_41_478 VPWR VGND sg13g2_fill_2
XFILLER_9_118 VPWR VGND sg13g2_fill_1
XFILLER_3_37 VPWR VGND sg13g2_fill_2
XFILLER_1_552 VPWR VGND sg13g2_decap_8
XFILLER_49_512 VPWR VGND sg13g2_fill_2
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_18_932 VPWR VGND sg13g2_decap_8
XFILLER_33_902 VPWR VGND sg13g2_decap_8
XFILLER_33_979 VPWR VGND sg13g2_decap_8
XFILLER_34_1001 VPWR VGND sg13g2_decap_8
XFILLER_41_990 VPWR VGND sg13g2_decap_8
X_2721_ VGND VPWR net475 _1123_ _0300_ _1039_ sg13g2_a21oi_1
XFILLER_13_681 VPWR VGND sg13g2_fill_1
XFILLER_9_663 VPWR VGND sg13g2_decap_8
XFILLER_12_191 VPWR VGND sg13g2_decap_8
X_2652_ net430 VPWR _1005_ VGND net488 net366 sg13g2_o21ai_1
X_1603_ VPWR _1174_ net714 VGND sg13g2_inv_1
X_2583_ VGND VPWR net484 _1192_ _0231_ _0970_ sg13g2_a21oi_1
X_1534_ VPWR _1105_ net645 VGND sg13g2_inv_1
XFILLER_4_390 VPWR VGND sg13g2_fill_2
X_3204_ net533 VGND VPWR _0070_ sdr_i.mac2.products_ff\[136\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3135_ net164 VGND VPWR _0326_ ppwm_i.u_ppwm.u_mem.memory\[111\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3066_ net174 VGND VPWR net683 ppwm_i.u_ppwm.u_mem.memory\[42\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_42_209 VPWR VGND sg13g2_decap_8
X_2017_ _1254_ _1255_ _0469_ _0472_ VPWR VGND sg13g2_nor3_2
XFILLER_23_423 VPWR VGND sg13g2_fill_1
XFILLER_24_924 VPWR VGND sg13g2_decap_8
X_2919_ net521 VGND VPWR _0110_ sdr_i.DP_2.matrix\[72\] clknet_leaf_3_clk sg13g2_dfrbpq_1
Xhold162 ppwm_i.u_ppwm.u_mem.memory\[100\] VPWR VGND net362 sg13g2_dlygate4sd3_1
Xhold151 _0193_ VPWR VGND net351 sg13g2_dlygate4sd3_1
Xhold140 _1069_ VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold184 _0272_ VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold195 _0282_ VPWR VGND net575 sg13g2_dlygate4sd3_1
Xhold173 _0413_ VPWR VGND net553 sg13g2_dlygate4sd3_1
XFILLER_37_32 VPWR VGND sg13g2_fill_1
XFILLER_15_913 VPWR VGND sg13g2_decap_8
XFILLER_14_401 VPWR VGND sg13g2_decap_8
XFILLER_41_220 VPWR VGND sg13g2_decap_4
XFILLER_42_776 VPWR VGND sg13g2_decap_8
XFILLER_30_916 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_393 VPWR VGND sg13g2_fill_2
XFILLER_49_386 VPWR VGND sg13g2_decap_8
XFILLER_37_526 VPWR VGND sg13g2_decap_8
XFILLER_18_784 VPWR VGND sg13g2_decap_4
XFILLER_45_592 VPWR VGND sg13g2_fill_2
XFILLER_21_905 VPWR VGND sg13g2_decap_8
XFILLER_33_776 VPWR VGND sg13g2_decap_8
X_2704_ net417 VPWR _1031_ VGND net478 net652 sg13g2_o21ai_1
X_2635_ VGND VPWR net491 _1166_ _0257_ _0996_ sg13g2_a21oi_1
X_2566_ net432 VPWR _0962_ VGND net495 ppwm_i.u_ppwm.u_mem.memory\[8\] sg13g2_o21ai_1
X_2497_ net423 VPWR _0907_ VGND net818 net374 sg13g2_o21ai_1
X_3118_ net72 VGND VPWR net598 ppwm_i.u_ppwm.u_mem.memory\[94\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
Xtiny_wrapper_16 VPWR VGND uio_out[0] sg13g2_tielo
Xtiny_wrapper_27 VPWR VGND uo_out[7] sg13g2_tielo
X_3049_ net52 VGND VPWR _0240_ ppwm_i.u_ppwm.u_mem.memory\[25\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_12_905 VPWR VGND sg13g2_decap_8
XFILLER_11_415 VPWR VGND sg13g2_fill_2
XFILLER_23_253 VPWR VGND sg13g2_decap_4
XFILLER_24_798 VPWR VGND sg13g2_fill_1
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_23_275 VPWR VGND sg13g2_fill_1
XFILLER_11_459 VPWR VGND sg13g2_decap_4
XFILLER_23_67 VPWR VGND sg13g2_fill_2
XFILLER_23_78 VPWR VGND sg13g2_fill_2
XFILLER_20_982 VPWR VGND sg13g2_decap_8
XFILLER_2_157 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_fill_1
Xfanout450 net452 net450 VPWR VGND sg13g2_buf_8
Xfanout483 net486 net483 VPWR VGND sg13g2_buf_8
Xfanout461 _1233_ net461 VPWR VGND sg13g2_buf_1
Xfanout472 net501 net472 VPWR VGND sg13g2_buf_8
XFILLER_24_1022 VPWR VGND sg13g2_decap_8
Xfanout494 net496 net494 VPWR VGND sg13g2_buf_1
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_9_36 VPWR VGND sg13g2_decap_8
XFILLER_9_69 VPWR VGND sg13g2_fill_1
XFILLER_7_920 VPWR VGND sg13g2_decap_8
XFILLER_11_993 VPWR VGND sg13g2_decap_8
XFILLER_10_481 VPWR VGND sg13g2_fill_1
XFILLER_7_997 VPWR VGND sg13g2_decap_8
XFILLER_6_496 VPWR VGND sg13g2_decap_8
X_2420_ _0836_ _0763_ _0725_ VPWR VGND sg13g2_nand2b_1
X_2351_ _0771_ ppwm_i.u_ppwm.global_counter\[14\] net403 VPWR VGND sg13g2_nand2_1
X_2282_ VGND VPWR _0687_ _0704_ _0705_ _0685_ sg13g2_a21oi_1
XFILLER_38_868 VPWR VGND sg13g2_decap_8
XFILLER_37_389 VPWR VGND sg13g2_fill_1
X_1997_ _1261_ _0461_ _0462_ VPWR VGND sg13g2_nor2_1
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
X_2618_ net430 VPWR _0988_ VGND net489 net675 sg13g2_o21ai_1
X_2549_ VPWR VGND _0953_ net459 _0950_ _1210_ _0214_ _0861_ sg13g2_a221oi_1
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_29_857 VPWR VGND sg13g2_decap_8
XFILLER_11_212 VPWR VGND sg13g2_fill_1
XFILLER_8_706 VPWR VGND sg13g2_decap_8
XFILLER_4_923 VPWR VGND sg13g2_decap_8
XFILLER_3_433 VPWR VGND sg13g2_fill_2
XFILLER_3_455 VPWR VGND sg13g2_decap_8
XFILLER_46_142 VPWR VGND sg13g2_fill_1
XFILLER_47_698 VPWR VGND sg13g2_decap_8
XFILLER_46_164 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_34_337 VPWR VGND sg13g2_decap_8
X_3023__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_30_510 VPWR VGND sg13g2_fill_1
X_1920_ sdr_i.mac2.sum_lvl2_ff\[1\] sdr_i.mac2.sum_lvl2_ff\[5\] _0421_ VPWR VGND sg13g2_xor2_1
X_1851_ _0390_ net312 net263 VPWR VGND sg13g2_nand2_1
XFILLER_30_554 VPWR VGND sg13g2_decap_8
X_1782_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[90\] net447 _1349_ net460 sg13g2_a21oi_1
XFILLER_6_271 VPWR VGND sg13g2_fill_1
XFILLER_41_2 VPWR VGND sg13g2_fill_1
X_2403_ VPWR VGND _0666_ _0692_ _0739_ _0350_ _0820_ _0723_ sg13g2_a221oi_1
X_2334_ _1225_ net391 _0754_ VPWR VGND sg13g2_nor2_1
XFILLER_29_109 VPWR VGND sg13g2_fill_2
X_2265_ net377 _0687_ _0678_ _0689_ VPWR VGND sg13g2_nand3_1
X_2196_ VPWR VGND _0621_ _1312_ _0620_ _1210_ _0622_ ppwm_i.u_ppwm.global_counter\[9\]
+ sg13g2_a221oi_1
XFILLER_37_120 VPWR VGND sg13g2_decap_8
XFILLER_25_304 VPWR VGND sg13g2_fill_1
XFILLER_37_164 VPWR VGND sg13g2_fill_2
XFILLER_38_687 VPWR VGND sg13g2_fill_1
XFILLER_37_197 VPWR VGND sg13g2_fill_1
XFILLER_41_808 VPWR VGND sg13g2_decap_8
XFILLER_25_359 VPWR VGND sg13g2_decap_8
XFILLER_34_882 VPWR VGND sg13g2_decap_8
XFILLER_4_208 VPWR VGND sg13g2_fill_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
Xhold22 sdr_i.DP_4.matrix\[10\] VPWR VGND net222 sg13g2_dlygate4sd3_1
Xhold11 sdr_i.mac2.sum_lvl1_ff\[32\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold55 _0032_ VPWR VGND net255 sg13g2_dlygate4sd3_1
Xhold44 sdr_i.DP_1.matrix\[46\] VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold33 sdr_i.DP_2.matrix\[64\] VPWR VGND net233 sg13g2_dlygate4sd3_1
Xhold88 sdr_i.DP_3.matrix\[0\] VPWR VGND net288 sg13g2_dlygate4sd3_1
XFILLER_21_1003 VPWR VGND sg13g2_decap_8
Xhold99 sdr_i.DP_3.matrix\[36\] VPWR VGND net299 sg13g2_dlygate4sd3_1
Xhold77 sdr_i.DP_4.matrix\[36\] VPWR VGND net277 sg13g2_dlygate4sd3_1
Xhold66 _0036_ VPWR VGND net266 sg13g2_dlygate4sd3_1
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_602 VPWR VGND sg13g2_decap_4
XFILLER_16_304 VPWR VGND sg13g2_decap_4
XFILLER_17_816 VPWR VGND sg13g2_fill_1
XFILLER_44_657 VPWR VGND sg13g2_decap_8
XFILLER_28_197 VPWR VGND sg13g2_fill_1
XFILLER_44_668 VPWR VGND sg13g2_fill_1
XFILLER_43_145 VPWR VGND sg13g2_decap_8
XFILLER_40_885 VPWR VGND sg13g2_decap_8
XFILLER_12_565 VPWR VGND sg13g2_decap_8
XFILLER_8_558 VPWR VGND sg13g2_fill_1
XFILLER_39_429 VPWR VGND sg13g2_fill_1
X_2050_ _0493_ _1242_ net410 VPWR VGND sg13g2_nand2_1
XFILLER_48_996 VPWR VGND sg13g2_decap_8
XFILLER_19_142 VPWR VGND sg13g2_fill_1
XFILLER_35_613 VPWR VGND sg13g2_decap_8
XFILLER_47_484 VPWR VGND sg13g2_decap_8
XFILLER_35_657 VPWR VGND sg13g2_fill_1
XFILLER_15_370 VPWR VGND sg13g2_fill_1
X_2952_ net537 VGND VPWR _0143_ sdr_i.DP_4.matrix\[55\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1903_ net316 net315 _0070_ VPWR VGND sg13g2_and2_1
XFILLER_31_863 VPWR VGND sg13g2_decap_8
X_2883_ net315 _0146_ VPWR VGND sg13g2_buf_1
X_1834_ _0379_ net548 _0378_ VPWR VGND sg13g2_nand2_1
X_1765_ ppwm_i.u_ppwm.u_mem.memory\[1\] net514 net517 _1332_ VPWR VGND sg13g2_nor3_1
X_1696_ net457 ppwm_i.rst_n VPWR VGND sg13g2_inv_4
X_2317_ _0736_ _0735_ _0737_ _0738_ VPWR VGND sg13g2_a21o_1
X_2248_ _0672_ net394 _0547_ VPWR VGND sg13g2_nand2_2
XFILLER_39_974 VPWR VGND sg13g2_decap_8
XFILLER_26_613 VPWR VGND sg13g2_fill_1
XFILLER_38_451 VPWR VGND sg13g2_decap_8
X_2179_ VGND VPWR _0586_ _0604_ _0605_ _0585_ sg13g2_a21oi_1
XFILLER_26_624 VPWR VGND sg13g2_decap_8
XFILLER_14_819 VPWR VGND sg13g2_decap_8
XFILLER_15_13 VPWR VGND sg13g2_decap_8
XFILLER_25_134 VPWR VGND sg13g2_decap_8
XFILLER_40_115 VPWR VGND sg13g2_decap_8
XFILLER_25_189 VPWR VGND sg13g2_decap_8
XFILLER_21_351 VPWR VGND sg13g2_fill_1
XFILLER_31_56 VPWR VGND sg13g2_decap_4
XFILLER_5_539 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_211 VPWR VGND sg13g2_fill_2
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_decap_8
XFILLER_48_237 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_16_101 VPWR VGND sg13g2_decap_8
XFILLER_29_495 VPWR VGND sg13g2_fill_1
XFILLER_16_145 VPWR VGND sg13g2_decap_4
XFILLER_32_616 VPWR VGND sg13g2_decap_8
XFILLER_12_351 VPWR VGND sg13g2_fill_2
XFILLER_12_362 VPWR VGND sg13g2_fill_1
XFILLER_13_885 VPWR VGND sg13g2_decap_8
XFILLER_40_693 VPWR VGND sg13g2_decap_4
XFILLER_9_856 VPWR VGND sg13g2_decap_8
XFILLER_8_399 VPWR VGND sg13g2_decap_8
X_1550_ VPWR _1121_ net354 VGND sg13g2_inv_1
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
X_3134__29 VPWR VGND net29 sg13g2_tiehi
X_3220_ net198 VGND VPWR net760 ppwm_i.u_ppwm.u_ex.state_q\[0\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3151_ net535 VGND VPWR _0043_ sdr_i.mac1.products_ff\[52\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2102_ VGND VPWR _0522_ _0524_ _0530_ _0523_ sg13g2_a21oi_1
X_3082_ net110 VGND VPWR _0273_ ppwm_i.u_ppwm.u_mem.memory\[58\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_48_793 VPWR VGND sg13g2_decap_8
XFILLER_47_281 VPWR VGND sg13g2_fill_1
XFILLER_36_933 VPWR VGND sg13g2_decap_8
X_2033_ VGND VPWR _1246_ net409 _0482_ net456 sg13g2_a21oi_1
XFILLER_35_454 VPWR VGND sg13g2_decap_4
XFILLER_16_690 VPWR VGND sg13g2_decap_8
X_2935_ net538 VGND VPWR _0126_ sdr_i.DP_3.matrix\[63\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2866_ net238 _0129_ VPWR VGND sg13g2_buf_1
X_1817_ _1339_ _0351_ _0365_ _0366_ VPWR VGND sg13g2_nor3_1
Xhold300 ppwm_i.u_ppwm.u_mem.memory\[97\] VPWR VGND net680 sg13g2_dlygate4sd3_1
Xhold311 ppwm_i.u_ppwm.u_mem.memory\[26\] VPWR VGND net691 sg13g2_dlygate4sd3_1
X_2797_ _1081_ VPWR _1082_ VGND _1240_ ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] sg13g2_o21ai_1
Xhold322 ppwm_i.u_ppwm.u_mem.memory\[41\] VPWR VGND net702 sg13g2_dlygate4sd3_1
XFILLER_2_509 VPWR VGND sg13g2_decap_4
X_1748_ VPWR VGND _1118_ _1313_ net442 _1104_ _1315_ net450 sg13g2_a221oi_1
Xhold333 _0194_ VPWR VGND net713 sg13g2_dlygate4sd3_1
Xhold344 _0012_ VPWR VGND net724 sg13g2_dlygate4sd3_1
Xhold377 sdr_i.mac2.products_ff\[17\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold366 sdr_i.mac1.sum_lvl1_ff\[24\] VPWR VGND net746 sg13g2_dlygate4sd3_1
Xhold355 _0016_ VPWR VGND net735 sg13g2_dlygate4sd3_1
X_1679_ VPWR _1250_ ppwm_i.u_ppwm.data_o VGND sg13g2_inv_1
X_3418_ net549 net5 VPWR VGND sg13g2_buf_1
Xhold399 _0018_ VPWR VGND net779 sg13g2_dlygate4sd3_1
Xhold388 ppwm_i.u_ppwm.u_ex.state_q\[2\] VPWR VGND net768 sg13g2_dlygate4sd3_1
XFILLER_27_933 VPWR VGND sg13g2_decap_8
XFILLER_38_281 VPWR VGND sg13g2_fill_1
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_42_958 VPWR VGND sg13g2_decap_8
XFILLER_41_457 VPWR VGND sg13g2_decap_8
XFILLER_10_811 VPWR VGND sg13g2_decap_4
XFILLER_42_77 VPWR VGND sg13g2_decap_8
X_3061__28 VPWR VGND net28 sg13g2_tiehi
XFILLER_10_888 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_fill_2
XFILLER_18_911 VPWR VGND sg13g2_decap_8
XFILLER_37_719 VPWR VGND sg13g2_decap_8
XFILLER_18_988 VPWR VGND sg13g2_decap_8
XFILLER_29_292 VPWR VGND sg13g2_decap_8
XFILLER_17_465 VPWR VGND sg13g2_decap_8
XFILLER_17_487 VPWR VGND sg13g2_decap_8
XFILLER_32_446 VPWR VGND sg13g2_decap_8
XFILLER_33_958 VPWR VGND sg13g2_decap_8
XFILLER_13_660 VPWR VGND sg13g2_fill_2
XFILLER_12_170 VPWR VGND sg13g2_decap_8
X_2720_ net418 VPWR _1039_ VGND net476 net358 sg13g2_o21ai_1
X_2651_ VGND VPWR net487 _1158_ _0265_ _1004_ sg13g2_a21oi_1
XFILLER_8_185 VPWR VGND sg13g2_decap_8
X_1602_ VPWR _1173_ net584 VGND sg13g2_inv_1
X_2582_ net427 VPWR _0970_ VGND net484 ppwm_i.u_ppwm.u_mem.memory\[16\] sg13g2_o21ai_1
XFILLER_5_881 VPWR VGND sg13g2_decap_8
X_1533_ VPWR _1104_ net749 VGND sg13g2_inv_1
X_3203_ net538 VGND VPWR _0069_ sdr_i.mac2.products_ff\[120\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3134_ net29 VGND VPWR net583 ppwm_i.u_ppwm.u_mem.memory\[110\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_27_207 VPWR VGND sg13g2_decap_8
X_3065_ net178 VGND VPWR _0256_ ppwm_i.u_ppwm.u_mem.memory\[41\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_2
X_2016_ _0163_ net572 _0469_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_903 VPWR VGND sg13g2_decap_8
XFILLER_36_741 VPWR VGND sg13g2_decap_8
XFILLER_23_413 VPWR VGND sg13g2_fill_2
XFILLER_23_446 VPWR VGND sg13g2_fill_2
XFILLER_23_457 VPWR VGND sg13g2_decap_8
X_2918_ net528 VGND VPWR _0109_ sdr_i.DP_2.matrix\[64\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_12_25 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_30_clk clknet_3_5__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_2849_ net288 _0112_ VPWR VGND sg13g2_buf_1
Xhold152 ppwm_i.u_ppwm.u_mem.memory\[17\] VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold130 ppwm_i.u_ppwm.u_mem.bit_count\[5\] VPWR VGND net330 sg13g2_dlygate4sd3_1
Xhold141 _0328_ VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold185 ppwm_i.u_ppwm.u_pwm.counter\[5\] VPWR VGND net565 sg13g2_dlygate4sd3_1
Xhold163 _0314_ VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold174 _0029_ VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold196 ppwm_i.u_ppwm.u_mem.memory\[30\] VPWR VGND net576 sg13g2_dlygate4sd3_1
XFILLER_46_505 VPWR VGND sg13g2_decap_4
XFILLER_18_229 VPWR VGND sg13g2_decap_8
XFILLER_37_55 VPWR VGND sg13g2_decap_8
XFILLER_42_722 VPWR VGND sg13g2_fill_1
XFILLER_42_700 VPWR VGND sg13g2_fill_2
XFILLER_15_969 VPWR VGND sg13g2_decap_8
XFILLER_14_468 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_21_clk clknet_3_6__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
XFILLER_5_111 VPWR VGND sg13g2_fill_1
XFILLER_6_689 VPWR VGND sg13g2_decap_8
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_fill_2
XFILLER_33_711 VPWR VGND sg13g2_decap_8
XFILLER_32_232 VPWR VGND sg13g2_fill_1
XFILLER_20_405 VPWR VGND sg13g2_decap_4
XFILLER_32_243 VPWR VGND sg13g2_fill_1
XFILLER_14_991 VPWR VGND sg13g2_decap_8
XFILLER_20_438 VPWR VGND sg13g2_decap_4
XFILLER_9_461 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_12_clk clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_2703_ VGND VPWR net466 _1132_ _0291_ _1030_ sg13g2_a21oi_1
X_2634_ net428 VPWR _0996_ VGND net491 net682 sg13g2_o21ai_1
X_3033__83 VPWR VGND net83 sg13g2_tiehi
X_2565_ VGND VPWR net494 _1201_ _0222_ _0961_ sg13g2_a21oi_1
X_2496_ _0770_ _0904_ _0905_ _0906_ VPWR VGND sg13g2_nor3_1
X_3117_ net80 VGND VPWR net641 ppwm_i.u_ppwm.u_mem.memory\[93\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_43_508 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_17 VPWR VGND uio_out[1] sg13g2_tielo
X_3048_ net53 VGND VPWR net587 ppwm_i.u_ppwm.u_mem.memory\[24\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_23_232 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_7_409 VPWR VGND sg13g2_decap_8
XFILLER_20_961 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 net441 net440 VPWR VGND sg13g2_buf_8
XFILLER_24_1001 VPWR VGND sg13g2_decap_8
Xfanout473 net476 net473 VPWR VGND sg13g2_buf_8
Xfanout462 net463 net462 VPWR VGND sg13g2_buf_8
Xfanout484 net486 net484 VPWR VGND sg13g2_buf_1
Xfanout451 net452 net451 VPWR VGND sg13g2_buf_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_46_302 VPWR VGND sg13g2_fill_2
Xfanout495 net496 net495 VPWR VGND sg13g2_buf_8
XFILLER_19_549 VPWR VGND sg13g2_fill_1
XFILLER_34_508 VPWR VGND sg13g2_decap_8
XFILLER_14_210 VPWR VGND sg13g2_decap_8
XFILLER_11_972 VPWR VGND sg13g2_decap_8
XFILLER_7_976 VPWR VGND sg13g2_decap_8
XFILLER_9_1017 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
X_2350_ _0769_ VPWR _0770_ VGND _0761_ _0765_ sg13g2_o21ai_1
XFILLER_2_670 VPWR VGND sg13g2_decap_4
X_2281_ _0704_ net507 net386 VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_1_clk clknet_3_1__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_49_184 VPWR VGND sg13g2_decap_8
XFILLER_38_847 VPWR VGND sg13g2_decap_8
XFILLER_37_346 VPWR VGND sg13g2_fill_2
XFILLER_25_519 VPWR VGND sg13g2_fill_2
XFILLER_33_541 VPWR VGND sg13g2_fill_2
XFILLER_33_563 VPWR VGND sg13g2_decap_8
XFILLER_21_725 VPWR VGND sg13g2_fill_2
XFILLER_33_596 VPWR VGND sg13g2_decap_4
XFILLER_20_257 VPWR VGND sg13g2_decap_8
X_1996_ _0153_ net333 _0459_ VPWR VGND sg13g2_xnor2_1
X_3000__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
X_2617_ VGND VPWR net489 _1175_ _0248_ _0987_ sg13g2_a21oi_1
X_2548_ VPWR VGND _0671_ _0861_ _0952_ _0691_ _0953_ _0850_ sg13g2_a221oi_1
XFILLER_0_618 VPWR VGND sg13g2_decap_8
X_2479_ _0879_ _0888_ _0877_ _0890_ VPWR VGND sg13g2_nand3_1
XFILLER_18_13 VPWR VGND sg13g2_decap_4
XFILLER_29_836 VPWR VGND sg13g2_decap_8
X_3088__86 VPWR VGND net86 sg13g2_tiehi
XFILLER_28_379 VPWR VGND sg13g2_decap_8
XFILLER_12_769 VPWR VGND sg13g2_fill_2
XFILLER_11_279 VPWR VGND sg13g2_fill_2
Xclkload0 clkload0/Y clknet_3_6__leaf_clk VPWR VGND sg13g2_inv_2
XFILLER_4_902 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_fill_1
XFILLER_4_979 VPWR VGND sg13g2_decap_8
XFILLER_34_316 VPWR VGND sg13g2_decap_8
XFILLER_15_530 VPWR VGND sg13g2_decap_8
X_3127__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_43_894 VPWR VGND sg13g2_decap_8
X_1850_ _0389_ _0388_ _0057_ VPWR VGND sg13g2_xor2_1
XFILLER_30_533 VPWR VGND sg13g2_decap_8
X_1781_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[76\] net510 net438 ppwm_i.u_ppwm.u_mem.memory\[62\]
+ _1348_ net447 sg13g2_a221oi_1
XFILLER_7_740 VPWR VGND sg13g2_decap_8
XFILLER_7_795 VPWR VGND sg13g2_fill_1
X_2402_ _0819_ _0763_ _0698_ VPWR VGND sg13g2_nand2b_1
X_2333_ _0753_ _0752_ _0198_ VPWR VGND sg13g2_nor2b_1
X_2264_ net800 net371 _0688_ VPWR VGND sg13g2_nor2_1
XFILLER_38_600 VPWR VGND sg13g2_fill_2
X_2195_ _0621_ _1260_ ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] _1259_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_633 VPWR VGND sg13g2_decap_8
XFILLER_38_655 VPWR VGND sg13g2_fill_2
XFILLER_37_154 VPWR VGND sg13g2_fill_2
XFILLER_38_666 VPWR VGND sg13g2_fill_2
XFILLER_25_338 VPWR VGND sg13g2_fill_2
XFILLER_34_861 VPWR VGND sg13g2_decap_8
X_1979_ _0452_ net279 net248 VPWR VGND sg13g2_nand2_1
XFILLER_1_905 VPWR VGND sg13g2_decap_8
XFILLER_49_909 VPWR VGND sg13g2_decap_8
Xhold23 sdr_i.DP_3.matrix\[1\] VPWR VGND net223 sg13g2_dlygate4sd3_1
XFILLER_0_459 VPWR VGND sg13g2_decap_8
Xhold12 sdr_i.mac2.products_ff\[137\] VPWR VGND net212 sg13g2_dlygate4sd3_1
Xhold34 sdr_i.DP_4.matrix\[19\] VPWR VGND net234 sg13g2_dlygate4sd3_1
Xhold45 sdr_i.DP_3.matrix\[19\] VPWR VGND net245 sg13g2_dlygate4sd3_1
XFILLER_29_56 VPWR VGND sg13g2_decap_4
Xhold56 sdr_i.DP_3.matrix\[37\] VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold78 sdr_i.DP_3.matrix\[27\] VPWR VGND net278 sg13g2_dlygate4sd3_1
Xhold67 sdr_i.mac1.sum_lvl1_ff\[16\] VPWR VGND net267 sg13g2_dlygate4sd3_1
Xhold89 sdr_i.DP_1.matrix\[63\] VPWR VGND net289 sg13g2_dlygate4sd3_1
XFILLER_29_644 VPWR VGND sg13g2_decap_8
XFILLER_43_113 VPWR VGND sg13g2_fill_2
XFILLER_45_99 VPWR VGND sg13g2_fill_2
XFILLER_45_88 VPWR VGND sg13g2_decap_8
XFILLER_43_135 VPWR VGND sg13g2_fill_1
XFILLER_25_894 VPWR VGND sg13g2_decap_8
XFILLER_40_864 VPWR VGND sg13g2_decap_8
XFILLER_8_537 VPWR VGND sg13g2_fill_2
XFILLER_8_526 VPWR VGND sg13g2_fill_1
XFILLER_4_721 VPWR VGND sg13g2_fill_1
XFILLER_10_91 VPWR VGND sg13g2_fill_1
XFILLER_48_975 VPWR VGND sg13g2_decap_8
XFILLER_43_680 VPWR VGND sg13g2_decap_8
XFILLER_15_360 VPWR VGND sg13g2_decap_8
X_2951_ net535 VGND VPWR _0142_ sdr_i.DP_4.matrix\[54\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_15_382 VPWR VGND sg13g2_fill_2
X_3140__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_31_842 VPWR VGND sg13g2_decap_8
X_1902_ net271 net302 _0068_ VPWR VGND sg13g2_and2_1
X_2882_ net253 _0145_ VPWR VGND sg13g2_buf_1
X_1833_ VGND VPWR _0378_ _0377_ _0374_ sg13g2_or2_1
X_1764_ _1331_ _1329_ _1330_ _1328_ _1326_ VPWR VGND sg13g2_a22oi_1
X_1695_ _1266_ net2 _1248_ VPWR VGND sg13g2_nand2_1
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
X_2316_ net378 VPWR _0737_ VGND _0735_ _0736_ sg13g2_o21ai_1
XFILLER_39_953 VPWR VGND sg13g2_decap_8
X_2247_ _0671_ net395 net394 _0365_ VPWR VGND sg13g2_and3_2
X_2178_ _0587_ VPWR _0604_ VGND _0601_ _0603_ sg13g2_o21ai_1
X_3058__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_13_308 VPWR VGND sg13g2_fill_2
XFILLER_22_831 VPWR VGND sg13g2_fill_1
XFILLER_31_35 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_706 VPWR VGND sg13g2_decap_8
XFILLER_0_278 VPWR VGND sg13g2_decap_8
XFILLER_1_779 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_31_127 VPWR VGND sg13g2_fill_1
XFILLER_13_864 VPWR VGND sg13g2_decap_8
XFILLER_8_345 VPWR VGND sg13g2_fill_2
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_3150_ net536 VGND VPWR _0042_ sdr_i.mac1.products_ff\[51\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_3081_ net114 VGND VPWR net564 ppwm_i.u_ppwm.u_mem.memory\[57\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2101_ VGND VPWR _0525_ _0529_ _0190_ net458 sg13g2_a21oi_1
XFILLER_48_772 VPWR VGND sg13g2_decap_8
X_2032_ net794 net409 _0481_ VPWR VGND sg13g2_nor2_1
XFILLER_36_912 VPWR VGND sg13g2_decap_8
XFILLER_47_260 VPWR VGND sg13g2_fill_1
XFILLER_36_989 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_4
X_3222__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_31_672 VPWR VGND sg13g2_decap_4
X_2934_ net535 VGND VPWR _0125_ sdr_i.DP_3.matrix\[55\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2865_ net316 _0128_ VPWR VGND sg13g2_buf_1
XFILLER_30_182 VPWR VGND sg13g2_fill_2
XFILLER_11_1014 VPWR VGND sg13g2_decap_8
X_1816_ _0358_ _0357_ _0364_ _0365_ VPWR VGND sg13g2_a21o_2
Xhold301 ppwm_i.u_ppwm.u_mem.memory\[84\] VPWR VGND net681 sg13g2_dlygate4sd3_1
X_2796_ _1080_ VPWR _1081_ VGND ppwm_i.u_ppwm.u_pwm.counter\[0\] _1247_ sg13g2_o21ai_1
Xhold334 ppwm_i.u_ppwm.u_mem.memory\[35\] VPWR VGND net714 sg13g2_dlygate4sd3_1
X_1747_ VGND VPWR _1111_ net438 _1314_ net460 sg13g2_a21oi_1
Xhold323 ppwm_i.u_ppwm.u_mem.memory\[47\] VPWR VGND net703 sg13g2_dlygate4sd3_1
Xhold312 ppwm_i.u_ppwm.u_mem.memory\[7\] VPWR VGND net692 sg13g2_dlygate4sd3_1
Xhold345 ppwm_i.u_ppwm.u_pwm.cmp_value\[9\] VPWR VGND net725 sg13g2_dlygate4sd3_1
Xhold378 _0033_ VPWR VGND net758 sg13g2_dlygate4sd3_1
Xhold367 _0026_ VPWR VGND net747 sg13g2_dlygate4sd3_1
Xhold356 sdr_i.mac1.sum_lvl1_ff\[1\] VPWR VGND net736 sg13g2_dlygate4sd3_1
X_1678_ VPWR _1249_ net326 VGND sg13g2_inv_1
X_3417_ net548 net4 VPWR VGND sg13g2_buf_1
Xhold389 ppwm_i.u_ppwm.u_pwm.counter\[0\] VPWR VGND net769 sg13g2_dlygate4sd3_1
XFILLER_27_912 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_fill_1
XFILLER_27_989 VPWR VGND sg13g2_decap_8
XFILLER_42_937 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_10_867 VPWR VGND sg13g2_decap_8
XFILLER_6_849 VPWR VGND sg13g2_decap_8
XFILLER_27_1010 VPWR VGND sg13g2_decap_8
XFILLER_1_587 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_45_742 VPWR VGND sg13g2_decap_8
XFILLER_44_241 VPWR VGND sg13g2_fill_1
XFILLER_18_967 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_8
XFILLER_33_937 VPWR VGND sg13g2_decap_8
XFILLER_9_610 VPWR VGND sg13g2_decap_8
XFILLER_8_120 VPWR VGND sg13g2_decap_8
X_2650_ net428 VPWR _1004_ VGND net491 ppwm_i.u_ppwm.u_mem.memory\[50\] sg13g2_o21ai_1
XFILLER_8_164 VPWR VGND sg13g2_decap_8
X_1601_ VPWR _1172_ net606 VGND sg13g2_inv_1
XFILLER_9_698 VPWR VGND sg13g2_decap_8
XFILLER_5_860 VPWR VGND sg13g2_decap_8
X_2581_ VGND VPWR net489 _1193_ _0230_ _0969_ sg13g2_a21oi_1
X_1532_ VPWR _1103_ ppwm_i.u_ppwm.u_mem.memory\[106\] VGND sg13g2_inv_1
X_3202_ net538 VGND VPWR _0068_ sdr_i.mac2.products_ff\[119\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
X_3133_ net45 VGND VPWR net605 ppwm_i.u_ppwm.u_mem.memory\[109\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3115__96 VPWR VGND net96 sg13g2_tiehi
X_3064_ net181 VGND VPWR _0255_ ppwm_i.u_ppwm.u_mem.memory\[40\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2015_ _1255_ _0469_ _0471_ VPWR VGND sg13g2_nor2_1
XFILLER_35_263 VPWR VGND sg13g2_fill_2
XFILLER_36_786 VPWR VGND sg13g2_decap_8
XFILLER_24_959 VPWR VGND sg13g2_decap_8
X_2917_ net530 VGND VPWR _0108_ sdr_i.DP_2.matrix\[63\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2848_ net224 _0111_ VPWR VGND sg13g2_buf_1
XFILLER_3_819 VPWR VGND sg13g2_decap_8
X_2779_ _1070_ net339 ppwm_i.u_ppwm.u_mem.bit_count\[0\] net472 VPWR VGND sg13g2_and3_1
Xhold120 ppwm_i.u_ppwm.global_counter\[6\] VPWR VGND net320 sg13g2_dlygate4sd3_1
Xhold153 _0231_ VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold142 ppwm_i.u_ppwm.u_mem.memory\[3\] VPWR VGND net342 sg13g2_dlygate4sd3_1
Xhold131 _1076_ VPWR VGND net331 sg13g2_dlygate4sd3_1
Xhold186 _0506_ VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold175 ppwm_i.u_ppwm.u_mem.memory\[99\] VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold164 ppwm_i.u_ppwm.u_mem.memory\[79\] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold197 _0244_ VPWR VGND net577 sg13g2_dlygate4sd3_1
X_3010__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_18_208 VPWR VGND sg13g2_decap_8
XFILLER_27_753 VPWR VGND sg13g2_fill_1
XFILLER_37_89 VPWR VGND sg13g2_fill_2
XFILLER_15_948 VPWR VGND sg13g2_decap_8
XFILLER_18_1009 VPWR VGND sg13g2_decap_8
XFILLER_23_992 VPWR VGND sg13g2_decap_8
XFILLER_6_668 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_49_366 VPWR VGND sg13g2_decap_4
XFILLER_45_594 VPWR VGND sg13g2_fill_1
XFILLER_17_285 VPWR VGND sg13g2_fill_2
XFILLER_14_970 VPWR VGND sg13g2_decap_8
X_2702_ net412 VPWR _1030_ VGND net466 net677 sg13g2_o21ai_1
XFILLER_13_491 VPWR VGND sg13g2_decap_8
X_2633_ VGND VPWR net491 _1167_ _0256_ _0995_ sg13g2_a21oi_1
X_2564_ net432 VPWR _0961_ VGND net494 net692 sg13g2_o21ai_1
X_2495_ net374 VPWR _0905_ VGND _0901_ _0902_ sg13g2_o21ai_1
X_3116_ net88 VGND VPWR _0307_ ppwm_i.u_ppwm.u_mem.memory\[92\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_28_528 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_18 VPWR VGND uio_out[2] sg13g2_tielo
X_3047_ net55 VGND VPWR net600 ppwm_i.u_ppwm.u_mem.memory\[23\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_24_789 VPWR VGND sg13g2_decap_8
XFILLER_11_417 VPWR VGND sg13g2_fill_1
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_23_288 VPWR VGND sg13g2_fill_1
XFILLER_20_940 VPWR VGND sg13g2_decap_8
XFILLER_3_649 VPWR VGND sg13g2_fill_2
Xfanout430 net434 net430 VPWR VGND sg13g2_buf_8
Xfanout441 _1283_ net441 VPWR VGND sg13g2_buf_8
Xfanout474 net476 net474 VPWR VGND sg13g2_buf_8
Xfanout463 net464 net463 VPWR VGND sg13g2_buf_8
Xfanout452 _1276_ net452 VPWR VGND sg13g2_buf_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
Xfanout485 net486 net485 VPWR VGND sg13g2_buf_8
Xfanout496 net500 net496 VPWR VGND sg13g2_buf_8
XFILLER_46_358 VPWR VGND sg13g2_fill_1
XFILLER_0_29 VPWR VGND sg13g2_decap_8
XFILLER_15_723 VPWR VGND sg13g2_decap_4
XFILLER_14_266 VPWR VGND sg13g2_decap_8
XFILLER_14_277 VPWR VGND sg13g2_fill_1
XFILLER_11_951 VPWR VGND sg13g2_decap_8
XFILLER_31_1017 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_955 VPWR VGND sg13g2_decap_8
XFILLER_6_476 VPWR VGND sg13g2_fill_1
X_2280_ _1228_ _0341_ _0347_ _0703_ VPWR VGND sg13g2_nor3_1
XFILLER_49_163 VPWR VGND sg13g2_decap_8
XFILLER_49_152 VPWR VGND sg13g2_fill_2
XFILLER_37_314 VPWR VGND sg13g2_decap_4
XFILLER_38_826 VPWR VGND sg13g2_decap_8
XFILLER_18_561 VPWR VGND sg13g2_decap_4
XFILLER_46_892 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_4
XFILLER_21_737 VPWR VGND sg13g2_decap_8
X_1995_ ppwm_i.u_ppwm.global_counter\[4\] ppwm_i.u_ppwm.global_counter\[3\] net333
+ _0461_ VPWR VGND _0458_ sg13g2_nand4_1
X_2616_ net431 VPWR _0987_ VGND net484 ppwm_i.u_ppwm.u_mem.memory\[33\] sg13g2_o21ai_1
X_2547_ VGND VPWR _1220_ net381 _0952_ _0951_ sg13g2_a21oi_1
X_2478_ _0879_ _0877_ _0888_ _0889_ VPWR VGND sg13g2_a21o_1
XFILLER_29_815 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_fill_2
XFILLER_28_358 VPWR VGND sg13g2_decap_8
X_3009__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_34_35 VPWR VGND sg13g2_decap_4
XFILLER_36_391 VPWR VGND sg13g2_decap_8
XFILLER_24_575 VPWR VGND sg13g2_decap_4
XFILLER_24_586 VPWR VGND sg13g2_decap_4
XFILLER_34_79 VPWR VGND sg13g2_fill_2
XFILLER_20_770 VPWR VGND sg13g2_decap_4
Xclkload1 clknet_3_7__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_958 VPWR VGND sg13g2_decap_8
XFILLER_47_667 VPWR VGND sg13g2_fill_2
XFILLER_35_829 VPWR VGND sg13g2_decap_8
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_fill_2
XFILLER_15_586 VPWR VGND sg13g2_decap_8
XFILLER_42_383 VPWR VGND sg13g2_decap_8
X_1780_ _1347_ net442 ppwm_i.u_ppwm.u_mem.memory\[69\] net450 ppwm_i.u_ppwm.u_mem.memory\[83\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_30_589 VPWR VGND sg13g2_decap_4
XFILLER_6_251 VPWR VGND sg13g2_fill_1
X_2401_ VGND VPWR _0814_ _0816_ _0818_ _0685_ sg13g2_a21oi_1
XFILLER_3_980 VPWR VGND sg13g2_decap_8
X_2332_ net435 VPWR _0753_ VGND net506 net373 sg13g2_o21ai_1
X_2263_ _0687_ ppwm_i.u_ppwm.pwm_value\[0\] net396 VPWR VGND sg13g2_nand2_1
X_2194_ _0619_ VPWR _0620_ VGND _0606_ _0618_ sg13g2_o21ai_1
XFILLER_26_818 VPWR VGND sg13g2_decap_8
XFILLER_38_678 VPWR VGND sg13g2_decap_8
XFILLER_25_317 VPWR VGND sg13g2_fill_2
XFILLER_34_840 VPWR VGND sg13g2_decap_8
XFILLER_14_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_567 VPWR VGND sg13g2_fill_1
X_1978_ _0451_ _0450_ _0047_ VPWR VGND sg13g2_xor2_1
XFILLER_0_416 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_fill_1
Xhold13 sdr_i.mac2.products_ff\[51\] VPWR VGND net213 sg13g2_dlygate4sd3_1
XFILLER_29_13 VPWR VGND sg13g2_decap_8
Xhold24 sdr_i.DP_2.matrix\[73\] VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold46 sdr_i.DP_4.matrix\[73\] VPWR VGND net246 sg13g2_dlygate4sd3_1
Xhold35 sdr_i.DP_1.matrix\[28\] VPWR VGND net235 sg13g2_dlygate4sd3_1
Xhold79 sdr_i.DP_1.matrix\[45\] VPWR VGND net279 sg13g2_dlygate4sd3_1
Xhold68 _0025_ VPWR VGND net268 sg13g2_dlygate4sd3_1
Xhold57 sdr_i.mac2.products_ff\[119\] VPWR VGND net257 sg13g2_dlygate4sd3_1
XFILLER_29_678 VPWR VGND sg13g2_decap_8
XFILLER_45_67 VPWR VGND sg13g2_decap_8
XFILLER_25_873 VPWR VGND sg13g2_decap_8
XFILLER_40_843 VPWR VGND sg13g2_decap_8
XFILLER_12_523 VPWR VGND sg13g2_fill_1
XFILLER_3_276 VPWR VGND sg13g2_fill_1
XFILLER_3_265 VPWR VGND sg13g2_decap_8
XFILLER_0_983 VPWR VGND sg13g2_decap_8
XFILLER_48_954 VPWR VGND sg13g2_decap_8
XFILLER_47_431 VPWR VGND sg13g2_fill_1
XFILLER_13_8 VPWR VGND sg13g2_fill_1
XFILLER_19_90 VPWR VGND sg13g2_fill_2
XFILLER_35_648 VPWR VGND sg13g2_fill_1
XFILLER_16_851 VPWR VGND sg13g2_decap_4
XFILLER_43_670 VPWR VGND sg13g2_fill_2
XFILLER_31_821 VPWR VGND sg13g2_decap_8
X_2950_ net542 VGND VPWR _0141_ sdr_i.DP_4.matrix\[46\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_37_1012 VPWR VGND sg13g2_decap_8
X_1901_ net309 net300 _0066_ VPWR VGND sg13g2_and2_1
X_2881_ net302 _0144_ VPWR VGND sg13g2_buf_1
X_1832_ _0377_ sdr_i.mac1.total_sum\[1\] sdr_i.mac2.total_sum\[1\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_397 VPWR VGND sg13g2_fill_2
XFILLER_31_898 VPWR VGND sg13g2_decap_8
X_1763_ VPWR VGND _1145_ net510 net443 _1131_ _1330_ net451 sg13g2_a221oi_1
X_1694_ VPWR _1265_ ppwm_i.u_ppwm.global_counter\[2\] VGND sg13g2_inv_1
XFILLER_44_1005 VPWR VGND sg13g2_decap_8
X_2315_ VGND VPWR _0713_ _0717_ _0736_ _0715_ sg13g2_a21oi_1
XFILLER_39_932 VPWR VGND sg13g2_decap_8
X_2246_ ppwm_i.u_ppwm.global_counter\[10\] ppwm_i.u_ppwm.global_counter\[0\] net398
+ _0670_ VPWR VGND sg13g2_mux2_1
XFILLER_26_604 VPWR VGND sg13g2_fill_2
X_2177_ _0602_ VPWR _0603_ VGND _1221_ ppwm_i.u_ppwm.global_counter\[8\] sg13g2_o21ai_1
XFILLER_38_497 VPWR VGND sg13g2_fill_1
XFILLER_41_629 VPWR VGND sg13g2_decap_8
XFILLER_33_180 VPWR VGND sg13g2_decap_8
XFILLER_21_386 VPWR VGND sg13g2_decap_8
XFILLER_22_898 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
Xoutput14 net14 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_246 VPWR VGND sg13g2_fill_1
XFILLER_0_213 VPWR VGND sg13g2_fill_1
XFILLER_1_758 VPWR VGND sg13g2_decap_8
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_44_401 VPWR VGND sg13g2_decap_8
XFILLER_29_486 VPWR VGND sg13g2_fill_1
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_44_456 VPWR VGND sg13g2_decap_8
XFILLER_44_445 VPWR VGND sg13g2_decap_8
XFILLER_40_662 VPWR VGND sg13g2_decap_8
XFILLER_12_331 VPWR VGND sg13g2_fill_2
XFILLER_12_386 VPWR VGND sg13g2_decap_4
XFILLER_4_552 VPWR VGND sg13g2_decap_8
XFILLER_21_80 VPWR VGND sg13g2_decap_4
XFILLER_4_596 VPWR VGND sg13g2_fill_2
X_3080_ net117 VGND VPWR net633 ppwm_i.u_ppwm.u_mem.memory\[56\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_0_780 VPWR VGND sg13g2_decap_8
X_2100_ _0529_ _0526_ _0528_ VPWR VGND sg13g2_nand2b_1
XFILLER_48_751 VPWR VGND sg13g2_decap_8
X_2031_ net457 _0479_ _0480_ _0169_ VPWR VGND sg13g2_nor3_1
XFILLER_47_272 VPWR VGND sg13g2_decap_8
XFILLER_36_968 VPWR VGND sg13g2_decap_8
XFILLER_23_629 VPWR VGND sg13g2_decap_8
X_2933_ net535 VGND VPWR _0124_ sdr_i.DP_3.matrix\[54\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_31_640 VPWR VGND sg13g2_fill_1
X_2864_ net250 _0127_ VPWR VGND sg13g2_buf_1
X_1815_ VPWR VGND _0363_ net509 _0361_ _0359_ _0364_ _0360_ sg13g2_a221oi_1
X_2795_ _1080_ ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] ppwm_i.u_ppwm.u_pwm.counter\[1\]
+ VPWR VGND sg13g2_nand2b_1
Xhold302 ppwm_i.u_ppwm.u_mem.memory\[42\] VPWR VGND net682 sg13g2_dlygate4sd3_1
XFILLER_7_71 VPWR VGND sg13g2_fill_2
XFILLER_7_60 VPWR VGND sg13g2_decap_8
X_1746_ ppwm_i.u_ppwm.u_mem.memory\[84\] net515 net518 _1313_ VPWR VGND sg13g2_nor3_1
Xhold324 ppwm_i.u_ppwm.u_mem.memory\[73\] VPWR VGND net704 sg13g2_dlygate4sd3_1
Xhold313 _0222_ VPWR VGND net693 sg13g2_dlygate4sd3_1
Xhold335 ppwm_i.u_ppwm.mem_write_done VPWR VGND net715 sg13g2_dlygate4sd3_1
Xhold346 ppwm_i.u_ppwm.u_mem.memory\[53\] VPWR VGND net726 sg13g2_dlygate4sd3_1
Xhold357 _0431_ VPWR VGND net737 sg13g2_dlygate4sd3_1
X_1677_ VPWR _1248_ net548 VGND sg13g2_inv_1
Xhold368 ppwm_i.u_ppwm.u_mem.bit_count\[4\] VPWR VGND net748 sg13g2_dlygate4sd3_1
Xhold379 ppwm_i.u_ppwm.u_ex.state_q\[0\] VPWR VGND net759 sg13g2_dlygate4sd3_1
X_3118__72 VPWR VGND net72 sg13g2_tiehi
X_2229_ net396 net395 net390 _0653_ VGND VPWR _0651_ sg13g2_nor4_2
XFILLER_38_250 VPWR VGND sg13g2_fill_1
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_27_968 VPWR VGND sg13g2_decap_8
XFILLER_42_916 VPWR VGND sg13g2_decap_8
XFILLER_41_415 VPWR VGND sg13g2_decap_8
XFILLER_14_607 VPWR VGND sg13g2_fill_2
XFILLER_14_629 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_4
XFILLER_41_437 VPWR VGND sg13g2_decap_4
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_42_13 VPWR VGND sg13g2_decap_4
XFILLER_42_57 VPWR VGND sg13g2_fill_1
XFILLER_22_684 VPWR VGND sg13g2_fill_1
XFILLER_6_828 VPWR VGND sg13g2_decap_8
XFILLER_21_183 VPWR VGND sg13g2_fill_2
XFILLER_1_566 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_fill_1
XFILLER_45_710 VPWR VGND sg13g2_decap_8
XFILLER_18_946 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
XFILLER_33_916 VPWR VGND sg13g2_decap_8
XFILLER_26_990 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_fill_1
XFILLER_32_459 VPWR VGND sg13g2_decap_4
XFILLER_34_1015 VPWR VGND sg13g2_decap_8
XFILLER_40_481 VPWR VGND sg13g2_decap_8
X_3060__30 VPWR VGND net30 sg13g2_tiehi
X_1600_ VPWR _1171_ net643 VGND sg13g2_inv_1
X_2580_ net431 VPWR _0969_ VGND net489 net588 sg13g2_o21ai_1
X_1531_ VPWR _1102_ net612 VGND sg13g2_inv_1
X_3201_ net537 VGND VPWR _0045_ sdr_i.mac2.products_ff\[103\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3132_ net60 VGND VPWR _0323_ ppwm_i.u_ppwm.u_mem.memory\[108\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_3063_ net185 VGND VPWR _0254_ ppwm_i.u_ppwm.u_mem.memory\[39\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2014_ _0469_ _0470_ _0162_ VPWR VGND sg13g2_and2_1
XFILLER_24_938 VPWR VGND sg13g2_decap_8
XFILLER_35_242 VPWR VGND sg13g2_decap_8
XFILLER_23_415 VPWR VGND sg13g2_fill_1
X_2916_ net528 VGND VPWR _0107_ sdr_i.DP_2.matrix\[55\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_32_982 VPWR VGND sg13g2_decap_8
X_2981__184 VPWR VGND net184 sg13g2_tiehi
X_2847_ net284 _0110_ VPWR VGND sg13g2_buf_1
Xhold110 sdr_i.DP_2.matrix\[54\] VPWR VGND net310 sg13g2_dlygate4sd3_1
X_2778_ VGND VPWR ppwm_i.u_ppwm.u_mem.bit_count\[0\] net472 _1069_ net339 sg13g2_a21oi_1
Xhold121 _0154_ VPWR VGND net321 sg13g2_dlygate4sd3_1
X_1729_ VGND VPWR _1296_ _1294_ _1288_ sg13g2_or2_1
Xhold143 ppwm_i.u_ppwm.u_mem.memory\[1\] VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold132 _0332_ VPWR VGND net332 sg13g2_dlygate4sd3_1
Xhold176 _0313_ VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold165 _0293_ VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold154 ppwm_i.u_ppwm.u_mem.memory\[88\] VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold198 ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] VPWR VGND net578 sg13g2_dlygate4sd3_1
Xhold187 _0188_ VPWR VGND net567 sg13g2_dlygate4sd3_1
XFILLER_37_13 VPWR VGND sg13g2_decap_8
XFILLER_39_570 VPWR VGND sg13g2_fill_2
XFILLER_26_231 VPWR VGND sg13g2_decap_8
XFILLER_15_927 VPWR VGND sg13g2_decap_8
XFILLER_26_242 VPWR VGND sg13g2_fill_1
XFILLER_26_297 VPWR VGND sg13g2_decap_8
XFILLER_41_267 VPWR VGND sg13g2_fill_2
XFILLER_23_971 VPWR VGND sg13g2_decap_8
XFILLER_6_603 VPWR VGND sg13g2_decap_4
XFILLER_10_654 VPWR VGND sg13g2_fill_2
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_49_323 VPWR VGND sg13g2_fill_2
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_17_242 VPWR VGND sg13g2_decap_8
XFILLER_17_264 VPWR VGND sg13g2_decap_8
XFILLER_45_584 VPWR VGND sg13g2_fill_2
XFILLER_32_223 VPWR VGND sg13g2_decap_8
XFILLER_33_746 VPWR VGND sg13g2_decap_8
XFILLER_21_919 VPWR VGND sg13g2_decap_8
XFILLER_33_757 VPWR VGND sg13g2_fill_1
XFILLER_32_278 VPWR VGND sg13g2_decap_8
X_2701_ VGND VPWR net465 _1133_ _0290_ _1029_ sg13g2_a21oi_1
X_2632_ net428 VPWR _0995_ VGND net487 net702 sg13g2_o21ai_1
X_2563_ VGND VPWR net494 _1202_ _0221_ _0960_ sg13g2_a21oi_1
X_2494_ VGND VPWR _1225_ net382 _0904_ _0903_ sg13g2_a21oi_1
XFILLER_4_94 VPWR VGND sg13g2_decap_8
X_3115_ net96 VGND VPWR net569 ppwm_i.u_ppwm.u_mem.memory\[91\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_28_507 VPWR VGND sg13g2_decap_8
X_3046_ net57 VGND VPWR net618 ppwm_i.u_ppwm.u_mem.memory\[22\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
Xtiny_wrapper_19 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_36_562 VPWR VGND sg13g2_decap_8
XFILLER_36_584 VPWR VGND sg13g2_decap_4
XFILLER_12_919 VPWR VGND sg13g2_decap_8
XFILLER_20_996 VPWR VGND sg13g2_decap_8
Xfanout420 net424 net420 VPWR VGND sg13g2_buf_8
Xfanout431 net433 net431 VPWR VGND sg13g2_buf_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
Xfanout464 net470 net464 VPWR VGND sg13g2_buf_8
Xfanout475 net476 net475 VPWR VGND sg13g2_buf_1
Xfanout453 net454 net453 VPWR VGND sg13g2_buf_8
Xfanout442 _1282_ net442 VPWR VGND sg13g2_buf_8
XFILLER_46_304 VPWR VGND sg13g2_fill_1
Xfanout486 net501 net486 VPWR VGND sg13g2_buf_8
XFILLER_19_518 VPWR VGND sg13g2_decap_8
XFILLER_19_529 VPWR VGND sg13g2_fill_2
Xfanout497 net498 net497 VPWR VGND sg13g2_buf_8
XFILLER_27_540 VPWR VGND sg13g2_fill_2
XFILLER_27_562 VPWR VGND sg13g2_fill_1
XFILLER_42_565 VPWR VGND sg13g2_fill_2
XFILLER_14_245 VPWR VGND sg13g2_decap_8
XFILLER_15_757 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_4
XFILLER_11_930 VPWR VGND sg13g2_decap_8
XFILLER_7_934 VPWR VGND sg13g2_decap_8
XFILLER_6_444 VPWR VGND sg13g2_fill_2
XFILLER_6_466 VPWR VGND sg13g2_fill_1
XFILLER_6_455 VPWR VGND sg13g2_decap_8
X_3136__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_49_131 VPWR VGND sg13g2_decap_8
XFILLER_1_171 VPWR VGND sg13g2_fill_1
XFILLER_38_805 VPWR VGND sg13g2_decap_8
XFILLER_46_871 VPWR VGND sg13g2_decap_8
XFILLER_33_510 VPWR VGND sg13g2_decap_8
X_1994_ _0459_ _0460_ _0152_ VPWR VGND sg13g2_and2_1
X_2615_ VGND VPWR net483 _1176_ _0247_ _0986_ sg13g2_a21oi_1
X_2546_ net381 _0852_ _0951_ VPWR VGND sg13g2_nor2_1
X_2477_ _0888_ _0886_ _0887_ VPWR VGND sg13g2_nand2_1
XFILLER_43_318 VPWR VGND sg13g2_fill_2
X_3029_ net91 VGND VPWR net629 ppwm_i.u_ppwm.u_mem.memory\[5\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
XFILLER_37_893 VPWR VGND sg13g2_decap_8
XFILLER_34_14 VPWR VGND sg13g2_decap_8
Xclkload2 VPWR clkload2/Y clknet_leaf_46_clk VGND sg13g2_inv_1
XFILLER_4_937 VPWR VGND sg13g2_decap_8
XFILLER_19_315 VPWR VGND sg13g2_fill_1
XFILLER_47_679 VPWR VGND sg13g2_fill_2
XFILLER_35_808 VPWR VGND sg13g2_decap_8
XFILLER_46_178 VPWR VGND sg13g2_decap_8
XFILLER_43_852 VPWR VGND sg13g2_decap_8
XFILLER_30_568 VPWR VGND sg13g2_decap_8
XFILLER_11_793 VPWR VGND sg13g2_decap_8
XFILLER_10_281 VPWR VGND sg13g2_decap_8
XFILLER_7_753 VPWR VGND sg13g2_fill_2
X_2400_ _0817_ _0815_ _0814_ VPWR VGND sg13g2_nand2b_1
X_2331_ _0738_ _0748_ net373 _0752_ VPWR VGND _0751_ sg13g2_nand4_1
X_2262_ VPWR VGND _1309_ _1229_ _1306_ net508 _0686_ _1302_ sg13g2_a221oi_1
XFILLER_38_602 VPWR VGND sg13g2_fill_1
X_2193_ _0619_ _1211_ ppwm_i.u_ppwm.global_counter\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_37_134 VPWR VGND sg13g2_decap_8
XFILLER_37_145 VPWR VGND sg13g2_fill_1
XFILLER_38_657 VPWR VGND sg13g2_fill_1
XFILLER_34_896 VPWR VGND sg13g2_decap_8
X_1977_ _0451_ net277 net256 VPWR VGND sg13g2_nand2_1
X_2529_ _0934_ _0935_ _0212_ VPWR VGND sg13g2_nor2_1
Xhold14 _0034_ VPWR VGND net214 sg13g2_dlygate4sd3_1
XFILLER_0_439 VPWR VGND sg13g2_decap_8
Xhold47 sdr_i.DP_4.matrix\[1\] VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold36 sdr_i.DP_3.matrix\[28\] VPWR VGND net236 sg13g2_dlygate4sd3_1
Xhold25 sdr_i.DP_2.matrix\[55\] VPWR VGND net225 sg13g2_dlygate4sd3_1
XFILLER_21_1017 VPWR VGND sg13g2_decap_8
Xhold58 _0038_ VPWR VGND net258 sg13g2_dlygate4sd3_1
Xhold69 sdr_i.mac2.sum_lvl1_ff\[24\] VPWR VGND net269 sg13g2_dlygate4sd3_1
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_45_46 VPWR VGND sg13g2_fill_1
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_44_627 VPWR VGND sg13g2_fill_2
XFILLER_43_159 VPWR VGND sg13g2_decap_8
XFILLER_40_822 VPWR VGND sg13g2_decap_8
XFILLER_8_506 VPWR VGND sg13g2_fill_2
XFILLER_12_579 VPWR VGND sg13g2_decap_4
XFILLER_40_899 VPWR VGND sg13g2_decap_8
XFILLER_8_539 VPWR VGND sg13g2_fill_1
XFILLER_3_200 VPWR VGND sg13g2_fill_1
XFILLER_10_82 VPWR VGND sg13g2_decap_8
XFILLER_3_288 VPWR VGND sg13g2_decap_8
XFILLER_0_962 VPWR VGND sg13g2_decap_8
XFILLER_48_933 VPWR VGND sg13g2_decap_8
XFILLER_19_101 VPWR VGND sg13g2_fill_1
XFILLER_34_115 VPWR VGND sg13g2_decap_8
XFILLER_28_690 VPWR VGND sg13g2_decap_8
XFILLER_16_885 VPWR VGND sg13g2_decap_8
XFILLER_31_800 VPWR VGND sg13g2_decap_8
X_1900_ net278 net301 _0064_ VPWR VGND sg13g2_and2_1
XFILLER_42_170 VPWR VGND sg13g2_decap_4
XFILLER_15_384 VPWR VGND sg13g2_fill_1
X_2880_ net227 _0143_ VPWR VGND sg13g2_buf_1
X_1831_ _0376_ sdr_i.mac1.total_sum\[1\] sdr_i.mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_30_332 VPWR VGND sg13g2_fill_2
XFILLER_31_877 VPWR VGND sg13g2_decap_8
X_1762_ _1329_ net439 _1138_ net447 _1152_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_583 VPWR VGND sg13g2_decap_8
X_1693_ _1264_ net789 VPWR VGND sg13g2_inv_2
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_911 VPWR VGND sg13g2_decap_8
X_2314_ _0735_ _0733_ _0734_ VPWR VGND sg13g2_nand2_1
X_2245_ _0669_ _0659_ _0668_ _0658_ net379 VPWR VGND sg13g2_a22oi_1
X_2176_ _0602_ net503 ppwm_i.u_ppwm.global_counter\[7\] VPWR VGND sg13g2_nand2b_1
XFILLER_39_988 VPWR VGND sg13g2_decap_8
XFILLER_25_148 VPWR VGND sg13g2_decap_8
XFILLER_40_129 VPWR VGND sg13g2_decap_4
XFILLER_34_693 VPWR VGND sg13g2_decap_8
XFILLER_21_343 VPWR VGND sg13g2_fill_2
XFILLER_22_877 VPWR VGND sg13g2_decap_8
XFILLER_21_365 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_0_225 VPWR VGND sg13g2_decap_8
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_48_207 VPWR VGND sg13g2_fill_2
XFILLER_0_258 VPWR VGND sg13g2_decap_4
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_44_435 VPWR VGND sg13g2_decap_4
XFILLER_25_693 VPWR VGND sg13g2_fill_2
XFILLER_9_826 VPWR VGND sg13g2_decap_8
X_3020__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_8_336 VPWR VGND sg13g2_fill_1
XFILLER_8_325 VPWR VGND sg13g2_fill_2
XFILLER_13_899 VPWR VGND sg13g2_decap_8
XFILLER_4_531 VPWR VGND sg13g2_decap_8
XFILLER_48_730 VPWR VGND sg13g2_decap_8
X_2030_ net578 net409 _0480_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_947 VPWR VGND sg13g2_decap_8
XFILLER_35_435 VPWR VGND sg13g2_decap_8
XFILLER_44_991 VPWR VGND sg13g2_decap_8
X_2932_ net543 VGND VPWR _0123_ sdr_i.DP_3.matrix\[46\] clknet_leaf_10_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_42_clk clknet_3_1__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
XFILLER_31_663 VPWR VGND sg13g2_fill_1
X_2863_ net271 _0126_ VPWR VGND sg13g2_buf_1
X_1814_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[44\] _0362_ net440 ppwm_i.u_ppwm.u_mem.memory\[37\]
+ _0363_ net444 sg13g2_a221oi_1
X_2794_ net457 _1078_ net695 _0333_ VPWR VGND sg13g2_nor3_1
XFILLER_30_184 VPWR VGND sg13g2_fill_1
XFILLER_8_881 VPWR VGND sg13g2_decap_8
X_1745_ _1312_ net404 _1311_ VPWR VGND sg13g2_nand2_2
Xhold303 _0257_ VPWR VGND net683 sg13g2_dlygate4sd3_1
Xhold325 ppwm_i.u_ppwm.u_mem.memory\[19\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xhold314 ppwm_i.u_ppwm.u_mem.bit_count\[6\] VPWR VGND net694 sg13g2_dlygate4sd3_1
Xhold347 ppwm_i.u_ppwm.u_mem.memory\[91\] VPWR VGND net727 sg13g2_dlygate4sd3_1
Xhold358 _0024_ VPWR VGND net738 sg13g2_dlygate4sd3_1
Xhold369 ppwm_i.u_ppwm.u_mem.memory\[105\] VPWR VGND net749 sg13g2_dlygate4sd3_1
Xhold336 ppwm_i.u_ppwm.u_mem.bit_count\[2\] VPWR VGND net716 sg13g2_dlygate4sd3_1
X_1676_ VPWR _1247_ net322 VGND sg13g2_inv_1
XFILLER_39_785 VPWR VGND sg13g2_decap_8
X_2228_ _1325_ net394 _0365_ _0652_ VPWR VGND sg13g2_nor3_1
XFILLER_26_446 VPWR VGND sg13g2_decap_8
XFILLER_27_947 VPWR VGND sg13g2_decap_8
X_2159_ _0585_ net398 _1311_ VPWR VGND sg13g2_nand2_2
Xclkbuf_leaf_33_clk clknet_3_5__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_10_836 VPWR VGND sg13g2_fill_2
XFILLER_22_663 VPWR VGND sg13g2_fill_2
XFILLER_22_696 VPWR VGND sg13g2_fill_1
XFILLER_18_925 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_fill_2
XFILLER_32_405 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_40_460 VPWR VGND sg13g2_fill_1
XFILLER_13_674 VPWR VGND sg13g2_decap_8
XFILLER_13_696 VPWR VGND sg13g2_decap_8
XFILLER_12_184 VPWR VGND sg13g2_decap_8
XFILLER_8_155 VPWR VGND sg13g2_fill_1
XFILLER_8_199 VPWR VGND sg13g2_fill_2
XFILLER_4_350 VPWR VGND sg13g2_fill_1
X_1530_ VPWR _1101_ net616 VGND sg13g2_inv_1
XFILLER_5_895 VPWR VGND sg13g2_decap_8
XFILLER_4_383 VPWR VGND sg13g2_decap_8
X_3200_ net537 VGND VPWR _0044_ sdr_i.mac2.products_ff\[102\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3131_ net76 VGND VPWR _0322_ ppwm_i.u_ppwm.u_mem.memory\[107\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_3062_ net189 VGND VPWR _0253_ ppwm_i.u_ppwm.u_mem.memory\[38\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2013_ _0467_ net776 net813 _0470_ VPWR VGND sg13g2_a21o_1
XFILLER_24_917 VPWR VGND sg13g2_decap_8
XFILLER_35_232 VPWR VGND sg13g2_fill_1
XFILLER_17_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_3_3__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_32_961 VPWR VGND sg13g2_decap_8
X_2915_ net528 VGND VPWR _0106_ sdr_i.DP_2.matrix\[54\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_2846_ net233 _0109_ VPWR VGND sg13g2_buf_1
XFILLER_12_39 VPWR VGND sg13g2_fill_2
X_2777_ _1067_ _1068_ _0327_ VPWR VGND sg13g2_nor2_1
Xhold100 sdr_i.DP_4.matrix\[45\] VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold111 sdr_i.DP_2.matrix\[45\] VPWR VGND net311 sg13g2_dlygate4sd3_1
X_1728_ _1288_ _1294_ _1295_ VPWR VGND sg13g2_nor2_2
Xhold144 _0215_ VPWR VGND net344 sg13g2_dlygate4sd3_1
Xhold122 ppwm_i.u_ppwm.u_pwm.cmp_value\[0\] VPWR VGND net322 sg13g2_dlygate4sd3_1
Xhold133 ppwm_i.u_ppwm.global_counter\[5\] VPWR VGND net333 sg13g2_dlygate4sd3_1
Xhold166 ppwm_i.u_ppwm.u_mem.memory\[51\] VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold155 _0302_ VPWR VGND net355 sg13g2_dlygate4sd3_1
X_1659_ VPWR _1230_ net712 VGND sg13g2_inv_1
Xhold177 ppwm_i.u_ppwm.global_counter\[10\] VPWR VGND net557 sg13g2_dlygate4sd3_1
Xhold188 ppwm_i.u_ppwm.u_mem.memory\[92\] VPWR VGND net568 sg13g2_dlygate4sd3_1
Xhold199 _0169_ VPWR VGND net579 sg13g2_dlygate4sd3_1
XFILLER_46_519 VPWR VGND sg13g2_decap_4
XFILLER_39_582 VPWR VGND sg13g2_fill_2
XFILLER_15_906 VPWR VGND sg13g2_decap_8
XFILLER_27_788 VPWR VGND sg13g2_decap_4
XFILLER_41_224 VPWR VGND sg13g2_fill_2
XFILLER_41_213 VPWR VGND sg13g2_decap_8
XFILLER_23_950 VPWR VGND sg13g2_decap_8
XFILLER_30_909 VPWR VGND sg13g2_decap_8
XFILLER_22_493 VPWR VGND sg13g2_decap_8
X_3019__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_5_158 VPWR VGND sg13g2_decap_4
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_49_302 VPWR VGND sg13g2_decap_4
XFILLER_1_364 VPWR VGND sg13g2_fill_1
XFILLER_49_357 VPWR VGND sg13g2_decap_4
XFILLER_49_379 VPWR VGND sg13g2_decap_8
XFILLER_37_519 VPWR VGND sg13g2_decap_8
XFILLER_45_530 VPWR VGND sg13g2_decap_4
XFILLER_27_80 VPWR VGND sg13g2_decap_8
XFILLER_17_287 VPWR VGND sg13g2_fill_1
XFILLER_27_91 VPWR VGND sg13g2_fill_1
XFILLER_43_90 VPWR VGND sg13g2_decap_8
XFILLER_41_780 VPWR VGND sg13g2_decap_8
X_2700_ net413 VPWR _1029_ VGND net462 net607 sg13g2_o21ai_1
XFILLER_13_471 VPWR VGND sg13g2_decap_8
XFILLER_40_290 VPWR VGND sg13g2_decap_8
XFILLER_9_475 VPWR VGND sg13g2_fill_2
X_2631_ VGND VPWR net487 _1168_ _0255_ _0994_ sg13g2_a21oi_1
X_2562_ net432 VPWR _0960_ VGND net494 net628 sg13g2_o21ai_1
XFILLER_5_681 VPWR VGND sg13g2_fill_1
XFILLER_4_191 VPWR VGND sg13g2_decap_4
X_2493_ net380 VPWR _0903_ VGND net382 _0772_ sg13g2_o21ai_1
Xclkbuf_leaf_4_clk clknet_3_0__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_3114_ net104 VGND VPWR _0305_ ppwm_i.u_ppwm.u_mem.memory\[90\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_3045_ net59 VGND VPWR net622 ppwm_i.u_ppwm.u_mem.memory\[21\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_36_541 VPWR VGND sg13g2_decap_8
XFILLER_23_202 VPWR VGND sg13g2_fill_2
XFILLER_24_736 VPWR VGND sg13g2_decap_4
XFILLER_23_246 VPWR VGND sg13g2_decap_8
XFILLER_17_1022 VPWR VGND sg13g2_decap_8
XFILLER_23_268 VPWR VGND sg13g2_decap_8
XFILLER_20_975 VPWR VGND sg13g2_decap_8
XFILLER_31_290 VPWR VGND sg13g2_decap_8
X_2829_ net272 _0092_ VPWR VGND sg13g2_buf_1
XFILLER_3_629 VPWR VGND sg13g2_decap_8
Xfanout410 net411 net410 VPWR VGND sg13g2_buf_8
Xfanout432 net433 net432 VPWR VGND sg13g2_buf_8
Xfanout421 net422 net421 VPWR VGND sg13g2_buf_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
Xfanout465 net467 net465 VPWR VGND sg13g2_buf_8
Xfanout443 _1282_ net443 VPWR VGND sg13g2_buf_2
Xfanout454 _1276_ net454 VPWR VGND sg13g2_buf_2
XFILLER_24_1015 VPWR VGND sg13g2_decap_8
Xfanout487 net488 net487 VPWR VGND sg13g2_buf_8
Xfanout476 net480 net476 VPWR VGND sg13g2_buf_8
Xfanout498 net500 net498 VPWR VGND sg13g2_buf_8
XFILLER_42_511 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_4
XFILLER_7_913 VPWR VGND sg13g2_decap_8
XFILLER_11_986 VPWR VGND sg13g2_decap_8
X_3030__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_49_110 VPWR VGND sg13g2_decap_8
XFILLER_49_198 VPWR VGND sg13g2_decap_8
XFILLER_46_850 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_33_555 VPWR VGND sg13g2_fill_2
XFILLER_21_706 VPWR VGND sg13g2_decap_4
XFILLER_20_227 VPWR VGND sg13g2_fill_1
X_1993_ _0458_ net789 net806 _0460_ VPWR VGND sg13g2_a21o_1
XFILLER_9_294 VPWR VGND sg13g2_decap_8
X_2614_ net427 VPWR _0986_ VGND net483 net345 sg13g2_o21ai_1
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
X_2545_ _0949_ VPWR _0950_ VGND _0947_ _0948_ sg13g2_o21ai_1
X_2476_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] net407 net405 _0887_ VPWR VGND sg13g2_or3_1
XFILLER_28_305 VPWR VGND sg13g2_fill_2
XFILLER_18_38 VPWR VGND sg13g2_fill_2
XFILLER_44_809 VPWR VGND sg13g2_decap_8
X_3028_ net93 VGND VPWR net685 ppwm_i.u_ppwm.u_mem.memory\[4\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_37_872 VPWR VGND sg13g2_decap_8
XFILLER_12_728 VPWR VGND sg13g2_fill_2
XFILLER_24_599 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_leaf_8_clk VGND sg13g2_inv_1
XFILLER_4_916 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_647 VPWR VGND sg13g2_fill_2
XFILLER_46_102 VPWR VGND sg13g2_decap_8
XFILLER_47_669 VPWR VGND sg13g2_fill_1
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_43_831 VPWR VGND sg13g2_decap_8
XFILLER_15_555 VPWR VGND sg13g2_fill_2
X_3062__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_11_761 VPWR VGND sg13g2_decap_8
XFILLER_24_70 VPWR VGND sg13g2_decap_4
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_10_260 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
X_2330_ _0751_ _0750_ net376 net375 net816 VPWR VGND sg13g2_a22oi_1
XFILLER_2_470 VPWR VGND sg13g2_fill_1
X_2261_ _0685_ net395 VPWR VGND _0651_ sg13g2_nand2b_2
X_3110__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_27_4 VPWR VGND sg13g2_decap_4
X_2192_ VPWR VGND _0616_ _0617_ _0615_ _1212_ _0618_ ppwm_i.u_ppwm.global_counter\[7\]
+ sg13g2_a221oi_1
XFILLER_37_113 VPWR VGND sg13g2_decap_8
XFILLER_38_647 VPWR VGND sg13g2_fill_2
XFILLER_19_850 VPWR VGND sg13g2_fill_1
XFILLER_25_319 VPWR VGND sg13g2_fill_1
XFILLER_34_875 VPWR VGND sg13g2_decap_8
XFILLER_21_514 VPWR VGND sg13g2_decap_8
XFILLER_21_547 VPWR VGND sg13g2_decap_8
X_1976_ _0450_ net299 net251 VPWR VGND sg13g2_nand2_1
X_2528_ net423 VPWR _0935_ VGND net817 _0860_ sg13g2_o21ai_1
XFILLER_1_919 VPWR VGND sg13g2_decap_8
Xhold15 sdr_i.mac1.sum_lvl1_ff\[0\] VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold37 sdr_i.DP_2.matrix\[10\] VPWR VGND net237 sg13g2_dlygate4sd3_1
Xhold26 sdr_i.DP_2.matrix\[28\] VPWR VGND net226 sg13g2_dlygate4sd3_1
X_2459_ net380 VPWR _0872_ VGND net383 _0709_ sg13g2_o21ai_1
Xhold48 sdr_i.DP_2.matrix\[46\] VPWR VGND net248 sg13g2_dlygate4sd3_1
Xhold59 sdr_i.mac2.sum_lvl3_ff\[0\] VPWR VGND net259 sg13g2_dlygate4sd3_1
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_37_691 VPWR VGND sg13g2_decap_4
XFILLER_40_801 VPWR VGND sg13g2_decap_8
XFILLER_40_878 VPWR VGND sg13g2_decap_8
XFILLER_12_558 VPWR VGND sg13g2_decap_8
XFILLER_20_591 VPWR VGND sg13g2_decap_4
XFILLER_3_223 VPWR VGND sg13g2_fill_1
XFILLER_0_941 VPWR VGND sg13g2_decap_8
XFILLER_48_912 VPWR VGND sg13g2_decap_8
XFILLER_47_400 VPWR VGND sg13g2_fill_2
XFILLER_48_989 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_fill_1
XFILLER_47_444 VPWR VGND sg13g2_decap_4
XFILLER_19_135 VPWR VGND sg13g2_decap_8
XFILLER_47_477 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_decap_8
XFILLER_35_639 VPWR VGND sg13g2_fill_1
XFILLER_16_831 VPWR VGND sg13g2_decap_4
XFILLER_15_341 VPWR VGND sg13g2_decap_4
XFILLER_42_182 VPWR VGND sg13g2_decap_8
XFILLER_30_322 VPWR VGND sg13g2_decap_4
X_1830_ _0375_ VPWR net12 VGND net548 _1250_ sg13g2_o21ai_1
XFILLER_31_856 VPWR VGND sg13g2_decap_8
X_1761_ VPWR VGND _1110_ _1327_ net439 _1117_ _1328_ net443 sg13g2_a221oi_1
X_1692_ VPWR _1263_ ppwm_i.u_ppwm.global_counter\[4\] VGND sg13g2_inv_1
X_2313_ net506 net408 net405 _0734_ VPWR VGND sg13g2_or3_1
X_2244_ _0663_ _0667_ _0668_ VPWR VGND sg13g2_nor2_1
X_2175_ VPWR VGND _1223_ _0600_ ppwm_i.u_ppwm.global_counter\[6\] _1222_ _0601_ ppwm_i.u_ppwm.global_counter\[7\]
+ sg13g2_a221oi_1
XFILLER_39_967 VPWR VGND sg13g2_decap_8
XFILLER_38_444 VPWR VGND sg13g2_decap_8
XFILLER_25_127 VPWR VGND sg13g2_decap_8
XFILLER_40_108 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_fill_1
XFILLER_22_845 VPWR VGND sg13g2_fill_2
XFILLER_22_856 VPWR VGND sg13g2_fill_1
XFILLER_31_49 VPWR VGND sg13g2_fill_2
X_1959_ sdr_i.mac2.sum_lvl1_ff\[16\] net269 _0011_ VPWR VGND sg13g2_xor2_1
XFILLER_1_716 VPWR VGND sg13g2_decap_8
X_2991__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_0_204 VPWR VGND sg13g2_decap_8
XFILLER_45_926 VPWR VGND sg13g2_decap_8
XFILLER_29_466 VPWR VGND sg13g2_fill_2
XFILLER_16_149 VPWR VGND sg13g2_fill_1
XFILLER_12_300 VPWR VGND sg13g2_fill_2
XFILLER_25_672 VPWR VGND sg13g2_decap_8
XFILLER_40_631 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_fill_1
XFILLER_13_878 VPWR VGND sg13g2_decap_8
XFILLER_40_697 VPWR VGND sg13g2_fill_2
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_40_675 VPWR VGND sg13g2_decap_8
XFILLER_9_849 VPWR VGND sg13g2_decap_8
XFILLER_4_521 VPWR VGND sg13g2_fill_1
XFILLER_48_786 VPWR VGND sg13g2_decap_8
XFILLER_36_926 VPWR VGND sg13g2_decap_8
XFILLER_35_447 VPWR VGND sg13g2_decap_8
XFILLER_44_970 VPWR VGND sg13g2_decap_8
X_2931_ net542 VGND VPWR _0122_ sdr_i.DP_3.matrix\[45\] clknet_leaf_8_clk sg13g2_dfrbpq_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_686 VPWR VGND sg13g2_fill_1
X_2862_ net242 _0125_ VPWR VGND sg13g2_buf_1
X_1813_ _0362_ ppwm_i.u_ppwm.u_mem.memory\[51\] net516 net519 VPWR VGND sg13g2_and3_1
X_2793_ VGND VPWR net694 _1066_ _1079_ _1077_ sg13g2_a21oi_1
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_1744_ net397 _1311_ VPWR VGND sg13g2_inv_4
Xhold326 ppwm_i.u_ppwm.u_mem.memory\[80\] VPWR VGND net706 sg13g2_dlygate4sd3_1
Xhold304 ppwm_i.u_ppwm.u_mem.memory\[5\] VPWR VGND net684 sg13g2_dlygate4sd3_1
Xhold315 _1079_ VPWR VGND net695 sg13g2_dlygate4sd3_1
Xhold348 ppwm_i.u_ppwm.u_mem.memory\[59\] VPWR VGND net728 sg13g2_dlygate4sd3_1
Xhold337 _1071_ VPWR VGND net717 sg13g2_dlygate4sd3_1
Xhold359 sdr_i.mac2.products_ff\[102\] VPWR VGND net739 sg13g2_dlygate4sd3_1
X_1675_ VPWR _1246_ ppwm_i.u_ppwm.u_pwm.cmp_value\[2\] VGND sg13g2_inv_1
XFILLER_39_720 VPWR VGND sg13g2_decap_8
X_2227_ VGND VPWR _0651_ _0365_ net394 sg13g2_or2_1
XFILLER_27_926 VPWR VGND sg13g2_decap_8
XFILLER_38_241 VPWR VGND sg13g2_fill_1
X_2158_ _0584_ _1252_ ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] _1251_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_274 VPWR VGND sg13g2_decap_8
X_2089_ net401 _0518_ _0519_ VPWR VGND sg13g2_nor2_1
XFILLER_10_826 VPWR VGND sg13g2_fill_1
XFILLER_21_141 VPWR VGND sg13g2_decap_8
XFILLER_5_329 VPWR VGND sg13g2_fill_2
XFILLER_1_524 VPWR VGND sg13g2_fill_1
XFILLER_27_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_18_904 VPWR VGND sg13g2_decap_8
XFILLER_29_285 VPWR VGND sg13g2_decap_8
XFILLER_44_277 VPWR VGND sg13g2_decap_4
XFILLER_32_439 VPWR VGND sg13g2_decap_8
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_9_635 VPWR VGND sg13g2_fill_1
XFILLER_12_163 VPWR VGND sg13g2_decap_8
XFILLER_8_134 VPWR VGND sg13g2_decap_4
XFILLER_8_178 VPWR VGND sg13g2_decap_8
XFILLER_5_874 VPWR VGND sg13g2_decap_8
XFILLER_4_362 VPWR VGND sg13g2_decap_8
X_3130_ net92 VGND VPWR net613 ppwm_i.u_ppwm.u_mem.memory\[106\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_0_590 VPWR VGND sg13g2_decap_8
X_3061_ net28 VGND VPWR net644 ppwm_i.u_ppwm.u_mem.memory\[37\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_2
XFILLER_36_734 VPWR VGND sg13g2_decap_8
X_2012_ net776 _0467_ net813 _0469_ VPWR VGND sg13g2_nand3_1
XFILLER_23_439 VPWR VGND sg13g2_decap_8
XFILLER_32_940 VPWR VGND sg13g2_decap_8
X_2914_ net532 VGND VPWR _0105_ sdr_i.DP_2.matrix\[46\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_2845_ net286 _0108_ VPWR VGND sg13g2_buf_1
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_472 VPWR VGND sg13g2_decap_8
XFILLER_31_483 VPWR VGND sg13g2_fill_1
Xhold101 sdr_i.DP_4.matrix\[27\] VPWR VGND net301 sg13g2_dlygate4sd3_1
X_2776_ _1068_ net751 net471 VPWR VGND sg13g2_xnor2_1
Xhold112 sdr_i.DP_2.matrix\[36\] VPWR VGND net312 sg13g2_dlygate4sd3_1
X_1727_ VPWR VGND _1293_ net509 _1292_ _1290_ _1294_ _1291_ sg13g2_a221oi_1
Xhold123 _0168_ VPWR VGND net323 sg13g2_dlygate4sd3_1
Xhold134 _0153_ VPWR VGND net334 sg13g2_dlygate4sd3_1
Xhold167 _0265_ VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold156 ppwm_i.u_ppwm.u_mem.memory\[44\] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold145 ppwm_i.u_ppwm.u_mem.memory\[32\] VPWR VGND net345 sg13g2_dlygate4sd3_1
X_1658_ ppwm_i.u_ppwm.pwm_value\[0\] _1229_ VPWR VGND sg13g2_inv_4
Xhold189 _0306_ VPWR VGND net569 sg13g2_dlygate4sd3_1
Xhold178 _0158_ VPWR VGND net558 sg13g2_dlygate4sd3_1
X_1589_ VPWR _1160_ net638 VGND sg13g2_inv_1
XFILLER_46_509 VPWR VGND sg13g2_fill_2
XFILLER_39_550 VPWR VGND sg13g2_fill_1
XFILLER_37_48 VPWR VGND sg13g2_decap_8
XFILLER_39_594 VPWR VGND sg13g2_decap_8
XFILLER_39_572 VPWR VGND sg13g2_fill_1
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_211 VPWR VGND sg13g2_decap_8
XFILLER_42_715 VPWR VGND sg13g2_fill_2
XFILLER_14_417 VPWR VGND sg13g2_fill_1
XFILLER_22_472 VPWR VGND sg13g2_decap_8
X_3027__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_6_627 VPWR VGND sg13g2_decap_8
XFILLER_10_656 VPWR VGND sg13g2_fill_1
X_3042__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_17_211 VPWR VGND sg13g2_decap_4
XFILLER_18_734 VPWR VGND sg13g2_fill_1
XFILLER_45_586 VPWR VGND sg13g2_fill_1
XFILLER_14_984 VPWR VGND sg13g2_decap_8
XFILLER_20_409 VPWR VGND sg13g2_fill_2
XFILLER_9_443 VPWR VGND sg13g2_fill_2
X_2630_ net430 VPWR _0994_ VGND net488 net699 sg13g2_o21ai_1
X_2561_ VGND VPWR net499 _1203_ _0220_ _0959_ sg13g2_a21oi_1
X_2492_ net378 VPWR _0902_ VGND _0896_ _0900_ sg13g2_o21ai_1
XFILLER_4_63 VPWR VGND sg13g2_decap_4
X_3113_ net112 VGND VPWR net615 ppwm_i.u_ppwm.u_mem.memory\[89\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_49_881 VPWR VGND sg13g2_decap_8
X_3044_ net61 VGND VPWR _0235_ ppwm_i.u_ppwm.u_mem.memory\[20\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
XFILLER_36_520 VPWR VGND sg13g2_decap_8
XFILLER_48_391 VPWR VGND sg13g2_fill_2
XFILLER_17_1001 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_20_954 VPWR VGND sg13g2_decap_8
X_2828_ net221 _0091_ VPWR VGND sg13g2_buf_1
X_2759_ VGND VPWR net468 _1104_ _0319_ _1058_ sg13g2_a21oi_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout411 _0477_ net411 VPWR VGND sg13g2_buf_8
Xfanout400 _1296_ net400 VPWR VGND sg13g2_buf_8
Xfanout422 net423 net422 VPWR VGND sg13g2_buf_8
Xfanout455 net459 net455 VPWR VGND sg13g2_buf_8
Xfanout466 net467 net466 VPWR VGND sg13g2_buf_8
Xfanout444 net446 net444 VPWR VGND sg13g2_buf_8
Xfanout433 net434 net433 VPWR VGND sg13g2_buf_8
Xfanout488 net490 net488 VPWR VGND sg13g2_buf_2
Xfanout477 net478 net477 VPWR VGND sg13g2_buf_8
Xfanout499 net500 net499 VPWR VGND sg13g2_buf_8
XFILLER_39_380 VPWR VGND sg13g2_decap_8
XFILLER_10_453 VPWR VGND sg13g2_fill_2
XFILLER_11_965 VPWR VGND sg13g2_decap_8
XFILLER_22_280 VPWR VGND sg13g2_decap_8
XFILLER_13_72 VPWR VGND sg13g2_decap_8
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_2_685 VPWR VGND sg13g2_fill_1
XFILLER_2_674 VPWR VGND sg13g2_fill_2
XFILLER_29_8 VPWR VGND sg13g2_fill_1
XFILLER_49_177 VPWR VGND sg13g2_decap_8
XFILLER_37_339 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_4
X_3100__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_45_394 VPWR VGND sg13g2_decap_8
XFILLER_33_534 VPWR VGND sg13g2_fill_2
XFILLER_33_589 VPWR VGND sg13g2_decap_8
XFILLER_14_781 VPWR VGND sg13g2_fill_2
X_1992_ net789 _0458_ net806 _0459_ VPWR VGND sg13g2_nand3_1
XFILLER_13_280 VPWR VGND sg13g2_fill_1
Xclkload10 clkload10/Y clknet_leaf_24_clk VPWR VGND sg13g2_inv_2
X_2613_ VGND VPWR net483 _1177_ _0246_ _0985_ sg13g2_a21oi_1
X_2544_ VGND VPWR _0947_ _0948_ _0949_ _0685_ sg13g2_a21oi_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] VPWR _0886_ VGND net407 net405 sg13g2_o21ai_1
XFILLER_18_17 VPWR VGND sg13g2_fill_2
XFILLER_29_829 VPWR VGND sg13g2_decap_8
XFILLER_18_28 VPWR VGND sg13g2_fill_2
XFILLER_37_851 VPWR VGND sg13g2_decap_8
X_3027_ net95 VGND VPWR _0218_ ppwm_i.u_ppwm.u_mem.memory\[3\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_34_49 VPWR VGND sg13g2_decap_4
Xclkload4 VPWR clkload4/Y clknet_leaf_37_clk VGND sg13g2_inv_1
XFILLER_3_427 VPWR VGND sg13g2_fill_2
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_4
XFILLER_43_810 VPWR VGND sg13g2_decap_8
XFILLER_15_512 VPWR VGND sg13g2_fill_2
XFILLER_28_862 VPWR VGND sg13g2_decap_8
X_3087__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_15_523 VPWR VGND sg13g2_decap_8
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_15_567 VPWR VGND sg13g2_fill_1
XFILLER_7_733 VPWR VGND sg13g2_decap_8
XFILLER_6_210 VPWR VGND sg13g2_decap_8
XFILLER_3_994 VPWR VGND sg13g2_decap_8
X_2260_ _0651_ net395 _0684_ VPWR VGND sg13g2_nor2b_2
X_2191_ net502 _1261_ _0617_ VPWR VGND sg13g2_nor2_1
XFILLER_38_615 VPWR VGND sg13g2_fill_2
XFILLER_38_626 VPWR VGND sg13g2_decap_8
XFILLER_1_64 VPWR VGND sg13g2_decap_8
XFILLER_45_180 VPWR VGND sg13g2_fill_1
XFILLER_19_895 VPWR VGND sg13g2_decap_8
XFILLER_33_320 VPWR VGND sg13g2_fill_2
XFILLER_34_854 VPWR VGND sg13g2_decap_8
XFILLER_33_364 VPWR VGND sg13g2_fill_1
XFILLER_33_397 VPWR VGND sg13g2_decap_8
X_1975_ _0449_ _0448_ _0045_ VPWR VGND sg13g2_xor2_1
XFILLER_14_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_18 VPWR VGND sg13g2_decap_4
X_2527_ VPWR VGND net380 _0933_ _0932_ _0929_ _0934_ _0930_ sg13g2_a221oi_1
X_2458_ VGND VPWR _0863_ _0869_ _0871_ _0870_ sg13g2_a21oi_1
Xhold16 _0023_ VPWR VGND net216 sg13g2_dlygate4sd3_1
Xhold38 sdr_i.DP_3.matrix\[73\] VPWR VGND net238 sg13g2_dlygate4sd3_1
Xhold27 sdr_i.DP_4.matrix\[55\] VPWR VGND net227 sg13g2_dlygate4sd3_1
X_2389_ _0807_ _0806_ _0659_ _0768_ net379 VPWR VGND sg13g2_a22oi_1
Xhold49 sdr_i.DP_2.matrix\[37\] VPWR VGND net249 sg13g2_dlygate4sd3_1
XFILLER_28_103 VPWR VGND sg13g2_decap_8
XFILLER_29_615 VPWR VGND sg13g2_fill_2
XFILLER_29_637 VPWR VGND sg13g2_decap_8
XFILLER_29_659 VPWR VGND sg13g2_fill_1
XFILLER_43_128 VPWR VGND sg13g2_decap_8
XFILLER_25_887 VPWR VGND sg13g2_decap_8
XFILLER_40_857 VPWR VGND sg13g2_decap_8
XFILLER_10_40 VPWR VGND sg13g2_decap_8
XFILLER_0_920 VPWR VGND sg13g2_decap_8
XFILLER_0_997 VPWR VGND sg13g2_decap_8
XFILLER_48_968 VPWR VGND sg13g2_decap_8
XFILLER_16_821 VPWR VGND sg13g2_decap_4
XFILLER_31_835 VPWR VGND sg13g2_decap_8
XFILLER_37_1026 VPWR VGND sg13g2_fill_2
X_1760_ ppwm_i.u_ppwm.u_mem.memory\[85\] net515 net518 _1327_ VPWR VGND sg13g2_nor3_1
XFILLER_7_552 VPWR VGND sg13g2_decap_8
X_1691_ VPWR _1262_ ppwm_i.u_ppwm.global_counter\[5\] VGND sg13g2_inv_1
XFILLER_44_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_791 VPWR VGND sg13g2_decap_8
X_2312_ net506 VPWR _0733_ VGND net408 net405 sg13g2_o21ai_1
XFILLER_39_946 VPWR VGND sg13g2_decap_8
X_2243_ net388 _0664_ _0665_ _0667_ VPWR VGND sg13g2_nor3_1
X_2174_ _0600_ _0598_ _0599_ _1261_ net504 VPWR VGND sg13g2_a22oi_1
XFILLER_15_29 VPWR VGND sg13g2_fill_2
XFILLER_33_150 VPWR VGND sg13g2_decap_8
X_3006__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_33_194 VPWR VGND sg13g2_fill_2
XFILLER_31_28 VPWR VGND sg13g2_decap_8
X_1958_ _0440_ net269 sdr_i.mac2.sum_lvl1_ff\[16\] VPWR VGND sg13g2_nand2_1
X_1889_ net295 net312 _0058_ VPWR VGND sg13g2_and2_1
XFILLER_48_209 VPWR VGND sg13g2_fill_1
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_44_415 VPWR VGND sg13g2_decap_8
XFILLER_16_128 VPWR VGND sg13g2_decap_4
XFILLER_40_610 VPWR VGND sg13g2_decap_8
XFILLER_24_161 VPWR VGND sg13g2_decap_4
XFILLER_25_695 VPWR VGND sg13g2_fill_1
XFILLER_31_109 VPWR VGND sg13g2_decap_8
XFILLER_4_588 VPWR VGND sg13g2_decap_4
XFILLER_0_794 VPWR VGND sg13g2_decap_8
XFILLER_48_765 VPWR VGND sg13g2_decap_8
XFILLER_35_404 VPWR VGND sg13g2_fill_2
XFILLER_36_905 VPWR VGND sg13g2_decap_8
XFILLER_29_990 VPWR VGND sg13g2_decap_8
XFILLER_16_640 VPWR VGND sg13g2_decap_8
XFILLER_16_662 VPWR VGND sg13g2_fill_1
XFILLER_22_109 VPWR VGND sg13g2_decap_8
X_2930_ net536 VGND VPWR _0121_ sdr_i.DP_3.matrix\[37\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_31_632 VPWR VGND sg13g2_fill_1
XFILLER_30_164 VPWR VGND sg13g2_fill_2
X_2861_ net282 _0124_ VPWR VGND sg13g2_buf_1
XFILLER_7_30 VPWR VGND sg13g2_decap_8
X_1812_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[30\] net449 _0361_ net461 sg13g2_a21oi_1
X_2792_ net694 _1077_ _1078_ VPWR VGND sg13g2_and2_1
XFILLER_30_175 VPWR VGND sg13g2_decap_8
XFILLER_31_698 VPWR VGND sg13g2_decap_8
XFILLER_11_1007 VPWR VGND sg13g2_decap_8
X_1743_ _1310_ _1306_ _1309_ _1302_ net508 VPWR VGND sg13g2_a22oi_1
Xhold305 _0219_ VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold316 _0333_ VPWR VGND net696 sg13g2_dlygate4sd3_1
X_1674_ VPWR _1245_ ppwm_i.u_ppwm.u_pwm.cmp_value\[3\] VGND sg13g2_inv_1
Xhold349 sdr_i.mac2.products_ff\[34\] VPWR VGND net729 sg13g2_dlygate4sd3_1
Xhold338 _0329_ VPWR VGND net718 sg13g2_dlygate4sd3_1
Xhold327 ppwm_i.u_ppwm.u_pwm.counter\[1\] VPWR VGND net707 sg13g2_dlygate4sd3_1
XFILLER_30_0 VPWR VGND sg13g2_decap_4
X_3133__45 VPWR VGND net45 sg13g2_tiehi
X_2226_ VGND VPWR _1230_ _0649_ _0194_ _0650_ sg13g2_a21oi_1
XFILLER_38_220 VPWR VGND sg13g2_decap_8
XFILLER_27_905 VPWR VGND sg13g2_decap_8
X_2157_ _0569_ VPWR _0583_ VGND _0581_ _0582_ sg13g2_o21ai_1
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_26_415 VPWR VGND sg13g2_fill_2
X_2088_ _0517_ VPWR _0518_ VGND ppwm_i.u_ppwm.u_ex.cmp_flag_q net394 sg13g2_o21ai_1
X_3039__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_22_621 VPWR VGND sg13g2_decap_8
XFILLER_10_838 VPWR VGND sg13g2_fill_1
XFILLER_27_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
XFILLER_44_212 VPWR VGND sg13g2_fill_1
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_16_72 VPWR VGND sg13g2_fill_2
XFILLER_16_94 VPWR VGND sg13g2_decap_8
XFILLER_9_603 VPWR VGND sg13g2_decap_8
XFILLER_12_153 VPWR VGND sg13g2_fill_1
XFILLER_8_113 VPWR VGND sg13g2_decap_8
XFILLER_13_687 VPWR VGND sg13g2_fill_1
XFILLER_5_853 VPWR VGND sg13g2_decap_8
X_3060_ net30 VGND VPWR _0251_ ppwm_i.u_ppwm.u_mem.memory\[36\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2011_ _0161_ _1256_ _0467_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_256 VPWR VGND sg13g2_decap_8
XFILLER_36_779 VPWR VGND sg13g2_decap_8
XFILLER_23_429 VPWR VGND sg13g2_decap_4
X_2913_ net532 VGND VPWR _0104_ sdr_i.DP_2.matrix\[45\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_2844_ net225 _0107_ VPWR VGND sg13g2_buf_1
XFILLER_32_996 VPWR VGND sg13g2_decap_8
X_2775_ _1067_ net421 _1066_ VPWR VGND sg13g2_nand2_2
Xhold135 ppwm_i.u_ppwm.global_counter\[9\] VPWR VGND net335 sg13g2_dlygate4sd3_1
X_1726_ VPWR VGND _1171_ net460 net446 _1157_ _1293_ net454 sg13g2_a221oi_1
Xhold113 sdr_i.mac1.products_ff\[34\] VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold124 ppwm_i.u_ppwm.u_mem.state_q\[0\] VPWR VGND net324 sg13g2_dlygate4sd3_1
Xhold102 sdr_i.DP_4.matrix\[63\] VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold157 _0258_ VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold146 _0246_ VPWR VGND net346 sg13g2_dlygate4sd3_1
Xhold168 ppwm_i.u_ppwm.u_mem.memory\[87\] VPWR VGND net368 sg13g2_dlygate4sd3_1
X_1657_ _1228_ net507 VPWR VGND sg13g2_inv_2
X_1588_ VPWR _1159_ net639 VGND sg13g2_inv_1
Xhold179 ppwm_i.u_ppwm.u_mem.memory\[72\] VPWR VGND net559 sg13g2_dlygate4sd3_1
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
X_3189_ net545 VGND VPWR _0057_ sdr_i.mac2.products_ff\[1\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2209_ _0635_ _1212_ net503 VPWR VGND sg13g2_nand2_1
XFILLER_39_584 VPWR VGND sg13g2_fill_1
XFILLER_42_727 VPWR VGND sg13g2_decap_4
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_311 VPWR VGND sg13g2_fill_2
XFILLER_1_355 VPWR VGND sg13g2_decap_4
XFILLER_40_1011 VPWR VGND sg13g2_decap_8
XFILLER_17_256 VPWR VGND sg13g2_decap_4
XFILLER_17_278 VPWR VGND sg13g2_decap_8
XFILLER_26_790 VPWR VGND sg13g2_fill_2
XFILLER_14_963 VPWR VGND sg13g2_decap_8
XFILLER_9_411 VPWR VGND sg13g2_fill_1
XFILLER_13_484 VPWR VGND sg13g2_decap_8
X_2560_ net433 VPWR _0959_ VGND net499 ppwm_i.u_ppwm.u_mem.memory\[5\] sg13g2_o21ai_1
XFILLER_5_672 VPWR VGND sg13g2_decap_8
X_2491_ _0896_ _0900_ _0901_ VPWR VGND sg13g2_and2_1
X_3113__112 VPWR VGND net112 sg13g2_tiehi
XFILLER_49_860 VPWR VGND sg13g2_decap_8
X_3112_ net119 VGND VPWR _0303_ ppwm_i.u_ppwm.u_mem.memory\[88\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_3043_ net63 VGND VPWR net624 ppwm_i.u_ppwm.u_mem.memory\[19\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_23_204 VPWR VGND sg13g2_fill_1
XFILLER_36_576 VPWR VGND sg13g2_decap_4
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_20_933 VPWR VGND sg13g2_decap_8
XFILLER_32_793 VPWR VGND sg13g2_decap_8
X_2827_ net289 _0090_ VPWR VGND sg13g2_buf_1
X_2758_ net415 VPWR _1058_ VGND net468 net645 sg13g2_o21ai_1
X_1709_ net514 net517 _1276_ VPWR VGND sg13g2_and2_1
X_2689_ VGND VPWR net462 _1139_ _0284_ _1023_ sg13g2_a21oi_1
Xfanout423 net424 net423 VPWR VGND sg13g2_buf_8
Xfanout412 net415 net412 VPWR VGND sg13g2_buf_8
Xfanout401 _1295_ net401 VPWR VGND sg13g2_buf_8
Xfanout456 net459 net456 VPWR VGND sg13g2_buf_1
Xfanout445 net446 net445 VPWR VGND sg13g2_buf_1
Xfanout434 ppwm_i.rst_n net434 VPWR VGND sg13g2_buf_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
Xfanout478 net479 net478 VPWR VGND sg13g2_buf_8
Xfanout467 net470 net467 VPWR VGND sg13g2_buf_2
Xfanout489 net490 net489 VPWR VGND sg13g2_buf_8
XFILLER_46_318 VPWR VGND sg13g2_decap_8
XFILLER_15_705 VPWR VGND sg13g2_decap_4
XFILLER_15_716 VPWR VGND sg13g2_decap_8
XFILLER_15_727 VPWR VGND sg13g2_fill_2
XFILLER_27_576 VPWR VGND sg13g2_decap_4
XFILLER_14_259 VPWR VGND sg13g2_decap_8
XFILLER_11_944 VPWR VGND sg13g2_decap_8
XFILLER_13_40 VPWR VGND sg13g2_fill_1
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_49_145 VPWR VGND sg13g2_decap_8
XFILLER_38_819 VPWR VGND sg13g2_decap_8
XFILLER_37_307 VPWR VGND sg13g2_decap_8
XFILLER_37_329 VPWR VGND sg13g2_fill_1
XFILLER_18_532 VPWR VGND sg13g2_decap_8
XFILLER_46_885 VPWR VGND sg13g2_decap_8
XFILLER_18_554 VPWR VGND sg13g2_decap_8
XFILLER_18_565 VPWR VGND sg13g2_fill_2
XFILLER_14_760 VPWR VGND sg13g2_decap_8
XFILLER_14_771 VPWR VGND sg13g2_fill_2
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_20_218 VPWR VGND sg13g2_fill_1
X_1991_ _0151_ _1264_ _0458_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_590 VPWR VGND sg13g2_decap_8
X_2612_ net426 VPWR _0985_ VGND net483 ppwm_i.u_ppwm.u_mem.memory\[31\] sg13g2_o21ai_1
Xclkload11 clknet_leaf_28_clk clkload11/Y VPWR VGND sg13g2_inv_4
X_2543_ _0948_ net805 net392 VPWR VGND sg13g2_xnor2_1
X_2474_ VPWR VGND _0885_ net458 _0881_ _1217_ _0207_ net370 sg13g2_a221oi_1
XFILLER_29_808 VPWR VGND sg13g2_decap_8
XFILLER_28_307 VPWR VGND sg13g2_fill_1
XFILLER_37_830 VPWR VGND sg13g2_decap_8
X_3026_ net97 VGND VPWR _0217_ ppwm_i.u_ppwm.u_mem.memory\[2\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_24_524 VPWR VGND sg13g2_decap_4
XFILLER_24_546 VPWR VGND sg13g2_fill_1
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_24_579 VPWR VGND sg13g2_fill_2
XFILLER_34_39 VPWR VGND sg13g2_fill_1
Xclkload5 VPWR clkload5/Y clknet_leaf_38_clk VGND sg13g2_inv_1
XFILLER_20_763 VPWR VGND sg13g2_decap_8
XFILLER_20_774 VPWR VGND sg13g2_fill_2
XFILLER_30_1021 VPWR VGND sg13g2_decap_8
X_3016__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_15_579 VPWR VGND sg13g2_decap_8
XFILLER_23_590 VPWR VGND sg13g2_decap_8
X_3142__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_11_785 VPWR VGND sg13g2_decap_4
XFILLER_6_299 VPWR VGND sg13g2_decap_8
XFILLER_3_973 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
X_2190_ _0616_ _1262_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] _1261_ net502 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_18_362 VPWR VGND sg13g2_decap_4
XFILLER_46_682 VPWR VGND sg13g2_decap_8
XFILLER_34_833 VPWR VGND sg13g2_decap_8
XFILLER_14_1005 VPWR VGND sg13g2_decap_8
X_1974_ _0449_ net282 net227 VPWR VGND sg13g2_nand2_1
X_2526_ _0933_ _0821_ _0860_ VPWR VGND sg13g2_nand2_1
XFILLER_0_409 VPWR VGND sg13g2_decap_8
X_2457_ net377 VPWR _0870_ VGND _0863_ _0869_ sg13g2_o21ai_1
Xhold28 sdr_i.DP_4.matrix\[28\] VPWR VGND net228 sg13g2_dlygate4sd3_1
Xhold17 sdr_i.mac1.products_ff\[17\] VPWR VGND net217 sg13g2_dlygate4sd3_1
XFILLER_29_39 VPWR VGND sg13g2_decap_4
X_2388_ net384 _0785_ _0806_ VPWR VGND sg13g2_and2_1
XFILLER_29_627 VPWR VGND sg13g2_decap_4
Xhold39 sdr_i.DP_4.matrix\[46\] VPWR VGND net239 sg13g2_dlygate4sd3_1
XFILLER_25_822 VPWR VGND sg13g2_decap_8
X_3009_ net130 VGND VPWR net829 ppwm_i.u_ppwm.pwm_value\[5\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_25_866 VPWR VGND sg13g2_decap_8
XFILLER_40_836 VPWR VGND sg13g2_decap_8
XFILLER_12_516 VPWR VGND sg13g2_decap_8
XFILLER_4_748 VPWR VGND sg13g2_fill_1
XFILLER_3_258 VPWR VGND sg13g2_decap_8
X_3172__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_0_976 VPWR VGND sg13g2_decap_8
XFILLER_48_947 VPWR VGND sg13g2_decap_8
XFILLER_19_83 VPWR VGND sg13g2_decap_8
XFILLER_19_115 VPWR VGND sg13g2_decap_4
XFILLER_15_321 VPWR VGND sg13g2_fill_1
XFILLER_16_855 VPWR VGND sg13g2_fill_2
XFILLER_37_1005 VPWR VGND sg13g2_decap_8
XFILLER_15_376 VPWR VGND sg13g2_fill_1
XFILLER_16_899 VPWR VGND sg13g2_decap_8
XFILLER_31_814 VPWR VGND sg13g2_decap_8
XFILLER_7_531 VPWR VGND sg13g2_decap_8
X_3220__198 VPWR VGND net198 sg13g2_tiehi
X_1690_ _1261_ net320 VPWR VGND sg13g2_inv_2
XFILLER_7_597 VPWR VGND sg13g2_decap_8
X_2977__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_3_770 VPWR VGND sg13g2_fill_2
X_2311_ _0732_ _0731_ _0197_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_925 VPWR VGND sg13g2_decap_8
X_2242_ _0664_ _0665_ _0666_ VPWR VGND sg13g2_nor2_1
X_2173_ _0599_ _1224_ ppwm_i.u_ppwm.global_counter\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_47_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_45_clk clknet_3_1__leaf_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
XFILLER_34_652 VPWR VGND sg13g2_decap_8
XFILLER_33_173 VPWR VGND sg13g2_decap_8
XFILLER_21_379 VPWR VGND sg13g2_decap_8
X_1957_ _0039_ _0438_ _0439_ VPWR VGND sg13g2_xnor2_1
X_1888_ net288 net280 _0056_ VPWR VGND sg13g2_and2_1
X_2509_ net390 VPWR _0917_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] ppwm_i.u_ppwm.u_ex.reg_value_q\[4\]
+ sg13g2_o21ai_1
XFILLER_0_239 VPWR VGND sg13g2_decap_8
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
XFILLER_29_468 VPWR VGND sg13g2_fill_1
XFILLER_38_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_36_clk clknet_3_4__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_13_803 VPWR VGND sg13g2_fill_1
XFILLER_12_324 VPWR VGND sg13g2_fill_2
XFILLER_12_379 VPWR VGND sg13g2_decap_8
XFILLER_21_891 VPWR VGND sg13g2_decap_8
XFILLER_21_73 VPWR VGND sg13g2_decap_8
XFILLER_4_545 VPWR VGND sg13g2_decap_8
XFILLER_21_84 VPWR VGND sg13g2_fill_2
XFILLER_4_578 VPWR VGND sg13g2_decap_4
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
XFILLER_0_773 VPWR VGND sg13g2_decap_8
XFILLER_48_744 VPWR VGND sg13g2_decap_8
XFILLER_47_265 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_27_clk clknet_3_7__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_43_482 VPWR VGND sg13g2_decap_8
X_2860_ net243 _0123_ VPWR VGND sg13g2_buf_1
X_1811_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[9\] net513 net445 ppwm_i.u_ppwm.u_mem.memory\[23\]
+ _0360_ net454 sg13g2_a221oi_1
XFILLER_30_132 VPWR VGND sg13g2_decap_8
XFILLER_7_20 VPWR VGND sg13g2_fill_1
XFILLER_12_891 VPWR VGND sg13g2_decap_8
X_2791_ _1067_ net331 _1077_ _0332_ VPWR VGND sg13g2_nor3_1
XFILLER_7_53 VPWR VGND sg13g2_decap_8
X_1742_ VGND VPWR net509 _1309_ _1308_ _1307_ sg13g2_a21oi_2
XFILLER_30_198 VPWR VGND sg13g2_fill_2
X_1673_ VPWR _1244_ net796 VGND sg13g2_inv_1
XFILLER_8_895 VPWR VGND sg13g2_decap_8
XFILLER_7_372 VPWR VGND sg13g2_fill_2
XFILLER_7_361 VPWR VGND sg13g2_decap_8
Xhold317 ppwm_i.u_ppwm.u_mem.memory\[18\] VPWR VGND net697 sg13g2_dlygate4sd3_1
Xhold306 ppwm_i.u_ppwm.u_mem.memory\[12\] VPWR VGND net686 sg13g2_dlygate4sd3_1
Xhold339 ppwm_i.u_ppwm.global_counter\[12\] VPWR VGND net719 sg13g2_dlygate4sd3_1
Xhold328 _0498_ VPWR VGND net708 sg13g2_dlygate4sd3_1
X_2225_ net419 VPWR _0650_ VGND net401 _0649_ sg13g2_o21ai_1
X_2156_ _1212_ ppwm_i.u_ppwm.global_counter\[17\] _0582_ VPWR VGND sg13g2_nor2_1
XFILLER_39_799 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_3__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_42_909 VPWR VGND sg13g2_decap_8
XFILLER_19_490 VPWR VGND sg13g2_decap_8
X_2087_ net395 _0365_ _0517_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_21_110 VPWR VGND sg13g2_decap_8
X_3054__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_21_176 VPWR VGND sg13g2_decap_8
X_2989_ net169 VGND VPWR _0180_ ppwm_i.u_ppwm.u_pwm.counter\[2\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
XFILLER_1_559 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_4
XFILLER_29_210 VPWR VGND sg13g2_fill_1
XFILLER_18_939 VPWR VGND sg13g2_decap_8
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_decap_4
XFILLER_33_909 VPWR VGND sg13g2_decap_8
XFILLER_13_600 VPWR VGND sg13g2_decap_8
XFILLER_26_983 VPWR VGND sg13g2_decap_8
XFILLER_41_920 VPWR VGND sg13g2_decap_8
XFILLER_34_1008 VPWR VGND sg13g2_decap_8
XFILLER_41_997 VPWR VGND sg13g2_decap_8
XFILLER_12_198 VPWR VGND sg13g2_decap_8
XFILLER_5_832 VPWR VGND sg13g2_decap_8
XFILLER_4_320 VPWR VGND sg13g2_decap_8
XFILLER_48_541 VPWR VGND sg13g2_fill_2
X_2010_ _0467_ net720 _0160_ VPWR VGND sg13g2_nor2_1
X_2912_ net529 VGND VPWR _0103_ sdr_i.DP_2.matrix\[37\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_16_482 VPWR VGND sg13g2_fill_1
XFILLER_17_994 VPWR VGND sg13g2_decap_8
XFILLER_32_975 VPWR VGND sg13g2_decap_8
X_2843_ net310 _0106_ VPWR VGND sg13g2_buf_1
XFILLER_31_496 VPWR VGND sg13g2_decap_8
X_2774_ _1066_ net324 net471 VPWR VGND sg13g2_nand2b_1
XFILLER_8_681 VPWR VGND sg13g2_decap_8
X_1725_ _1292_ net441 _1164_ net448 _1178_ VPWR VGND sg13g2_a22oi_1
Xhold103 sdr_i.DP_1.matrix\[54\] VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold114 _0017_ VPWR VGND net314 sg13g2_dlygate4sd3_1
Xhold125 _0005_ VPWR VGND net325 sg13g2_dlygate4sd3_1
Xhold136 _0157_ VPWR VGND net336 sg13g2_dlygate4sd3_1
Xhold147 ppwm_i.u_ppwm.u_mem.memory\[65\] VPWR VGND net347 sg13g2_dlygate4sd3_1
Xhold158 ppwm_i.u_ppwm.u_mem.memory\[85\] VPWR VGND net358 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_6__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_1656_ _1227_ ppwm_i.u_ppwm.pwm_value\[2\] VPWR VGND sg13g2_inv_2
X_1587_ VPWR _1158_ net366 VGND sg13g2_inv_1
Xhold169 _0301_ VPWR VGND net369 sg13g2_dlygate4sd3_1
X_3188_ net544 VGND VPWR _0056_ sdr_i.mac2.products_ff\[0\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2208_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] _0633_ _1223_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\]
+ _0634_ _1222_ sg13g2_a221oi_1
XFILLER_39_563 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_3121__49 VPWR VGND net49 sg13g2_tiehi
X_2139_ _0564_ VPWR _0565_ VGND net504 _1254_ sg13g2_o21ai_1
XFILLER_42_717 VPWR VGND sg13g2_fill_1
XFILLER_14_408 VPWR VGND sg13g2_decap_4
XFILLER_23_964 VPWR VGND sg13g2_decap_8
XFILLER_10_625 VPWR VGND sg13g2_decap_4
XFILLER_10_669 VPWR VGND sg13g2_decap_4
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_49_316 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_decap_4
X_3065__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_14_942 VPWR VGND sg13g2_decap_8
XFILLER_32_216 VPWR VGND sg13g2_decap_8
XFILLER_41_794 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_fill_1
X_2490_ _0897_ _0875_ _0898_ _0900_ VPWR VGND sg13g2_a21o_2
X_3072__149 VPWR VGND net149 sg13g2_tiehi
X_3111_ net127 VGND VPWR net355 ppwm_i.u_ppwm.u_mem.memory\[87\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_3042_ net65 VGND VPWR _0233_ ppwm_i.u_ppwm.u_mem.memory\[18\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_48_393 VPWR VGND sg13g2_fill_1
XFILLER_36_588 VPWR VGND sg13g2_fill_2
XFILLER_20_912 VPWR VGND sg13g2_decap_8
X_2826_ net264 _0089_ VPWR VGND sg13g2_buf_1
XFILLER_31_282 VPWR VGND sg13g2_decap_4
XFILLER_20_989 VPWR VGND sg13g2_decap_8
X_2757_ VGND VPWR net464 _1105_ _0318_ _1057_ sg13g2_a21oi_1
X_2688_ net413 VPWR _1023_ VGND net462 net637 sg13g2_o21ai_1
X_1708_ _1275_ VPWR _0005_ VGND _1271_ _1272_ sg13g2_o21ai_1
X_1639_ _1210_ net805 VPWR VGND sg13g2_inv_2
Xfanout402 net403 net402 VPWR VGND sg13g2_buf_8
Xfanout413 net415 net413 VPWR VGND sg13g2_buf_8
Xfanout446 _1282_ net446 VPWR VGND sg13g2_buf_1
Xfanout424 ppwm_i.rst_n net424 VPWR VGND sg13g2_buf_8
Xfanout457 net459 net457 VPWR VGND sg13g2_buf_8
Xfanout435 net437 net435 VPWR VGND sg13g2_buf_8
Xfanout479 net480 net479 VPWR VGND sg13g2_buf_8
Xfanout468 net470 net468 VPWR VGND sg13g2_buf_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_27_533 VPWR VGND sg13g2_decap_8
XFILLER_42_536 VPWR VGND sg13g2_decap_8
XFILLER_10_400 VPWR VGND sg13g2_decap_8
XFILLER_11_923 VPWR VGND sg13g2_decap_8
XFILLER_23_772 VPWR VGND sg13g2_fill_2
XFILLER_13_30 VPWR VGND sg13g2_decap_4
XFILLER_7_927 VPWR VGND sg13g2_decap_8
XFILLER_13_52 VPWR VGND sg13g2_decap_4
XFILLER_6_437 VPWR VGND sg13g2_decap_8
XFILLER_2_610 VPWR VGND sg13g2_decap_8
XFILLER_1_142 VPWR VGND sg13g2_fill_2
XFILLER_49_124 VPWR VGND sg13g2_decap_8
XFILLER_46_864 VPWR VGND sg13g2_decap_8
XFILLER_33_503 VPWR VGND sg13g2_decap_8
XFILLER_33_536 VPWR VGND sg13g2_fill_1
X_1990_ _0150_ net710 _0456_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_242 VPWR VGND sg13g2_decap_8
X_2611_ VGND VPWR net484 _1178_ _0245_ _0984_ sg13g2_a21oi_1
Xclkload12 clkload12/Y clknet_leaf_29_clk VPWR VGND sg13g2_inv_2
X_2542_ _0940_ VPWR _0947_ VGND _0939_ _0941_ sg13g2_o21ai_1
XFILLER_6_982 VPWR VGND sg13g2_decap_8
X_2473_ _0885_ _0726_ net374 _0884_ VPWR VGND sg13g2_and3_1
XFILLER_28_319 VPWR VGND sg13g2_fill_1
XFILLER_49_691 VPWR VGND sg13g2_decap_4
X_3025_ net99 VGND VPWR net338 ppwm_i.u_ppwm.u_mem.memory\[1\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_37_886 VPWR VGND sg13g2_decap_8
XFILLER_20_742 VPWR VGND sg13g2_decap_8
Xclkload6 clkload6/Y clknet_leaf_30_clk VPWR VGND sg13g2_inv_2
XFILLER_30_1000 VPWR VGND sg13g2_decap_8
X_2809_ _1094_ _1242_ net839 _1241_ ppwm_i.u_ppwm.u_pwm.counter\[9\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_429 VPWR VGND sg13g2_fill_1
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_43_845 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_11_742 VPWR VGND sg13g2_decap_8
XFILLER_11_775 VPWR VGND sg13g2_decap_4
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_10_274 VPWR VGND sg13g2_decap_8
XFILLER_40_72 VPWR VGND sg13g2_fill_2
XFILLER_40_94 VPWR VGND sg13g2_decap_8
XFILLER_3_952 VPWR VGND sg13g2_decap_8
XFILLER_38_617 VPWR VGND sg13g2_fill_1
XFILLER_37_127 VPWR VGND sg13g2_decap_8
XFILLER_18_341 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_fill_2
XFILLER_34_812 VPWR VGND sg13g2_decap_8
XFILLER_34_889 VPWR VGND sg13g2_decap_8
X_1973_ _0448_ net283 net242 VPWR VGND sg13g2_nand2_1
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_2525_ VGND VPWR _1222_ net382 _0932_ _0931_ sg13g2_a21oi_1
X_2456_ _0869_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] net389 VPWR VGND sg13g2_xnor2_1
Xhold18 _0015_ VPWR VGND net218 sg13g2_dlygate4sd3_1
Xhold29 sdr_i.DP_1.matrix\[1\] VPWR VGND net229 sg13g2_dlygate4sd3_1
XFILLER_29_617 VPWR VGND sg13g2_fill_1
X_2387_ _0803_ _0804_ _0691_ _0805_ VPWR VGND sg13g2_nand3_1
XFILLER_45_28 VPWR VGND sg13g2_decap_8
X_3008_ net132 VGND VPWR _0199_ ppwm_i.u_ppwm.pwm_value\[4\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_3126__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_40_815 VPWR VGND sg13g2_decap_8
XFILLER_20_572 VPWR VGND sg13g2_decap_4
XFILLER_10_75 VPWR VGND sg13g2_decap_8
XFILLER_0_955 VPWR VGND sg13g2_decap_8
XFILLER_48_926 VPWR VGND sg13g2_decap_8
XFILLER_19_62 VPWR VGND sg13g2_decap_8
XFILLER_28_683 VPWR VGND sg13g2_decap_8
XFILLER_34_108 VPWR VGND sg13g2_decap_8
XFILLER_42_163 VPWR VGND sg13g2_decap_8
XFILLER_35_94 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_594 VPWR VGND sg13g2_decap_8
X_2310_ net435 VPWR _0732_ VGND net794 net373 sg13g2_o21ai_1
X_2241_ _1226_ net403 _0665_ VPWR VGND sg13g2_nor2_1
XFILLER_39_904 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_38_425 VPWR VGND sg13g2_decap_8
X_2172_ _0597_ VPWR _0598_ VGND _0594_ _0596_ sg13g2_o21ai_1
XFILLER_20_1010 VPWR VGND sg13g2_decap_8
XFILLER_38_458 VPWR VGND sg13g2_fill_2
XFILLER_34_620 VPWR VGND sg13g2_decap_4
XFILLER_34_686 VPWR VGND sg13g2_fill_2
X_1956_ sdr_i.mac2.products_ff\[120\] sdr_i.mac2.products_ff\[103\] _0439_ VPWR VGND
+ sg13g2_xor2_1
XFILLER_30_881 VPWR VGND sg13g2_decap_8
X_1887_ _0016_ _0406_ _0407_ VPWR VGND sg13g2_xnor2_1
X_2508_ _0916_ net502 net393 VPWR VGND sg13g2_xnor2_1
XFILLER_0_218 VPWR VGND sg13g2_decap_8
X_2439_ _0854_ net373 _0853_ VPWR VGND sg13g2_nand2_1
XFILLER_29_436 VPWR VGND sg13g2_decap_8
XFILLER_44_439 VPWR VGND sg13g2_fill_2
XFILLER_16_108 VPWR VGND sg13g2_decap_8
XFILLER_25_653 VPWR VGND sg13g2_fill_1
XFILLER_40_601 VPWR VGND sg13g2_decap_4
XFILLER_25_686 VPWR VGND sg13g2_decap_8
XFILLER_40_645 VPWR VGND sg13g2_fill_2
XFILLER_24_174 VPWR VGND sg13g2_fill_1
XFILLER_12_347 VPWR VGND sg13g2_decap_4
XFILLER_12_358 VPWR VGND sg13g2_decap_4
XFILLER_21_870 VPWR VGND sg13g2_decap_8
XFILLER_4_502 VPWR VGND sg13g2_decap_8
XFILLER_0_752 VPWR VGND sg13g2_decap_8
XFILLER_48_723 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_fill_1
XFILLER_47_299 VPWR VGND sg13g2_decap_8
XFILLER_44_984 VPWR VGND sg13g2_decap_8
XFILLER_43_461 VPWR VGND sg13g2_decap_8
XFILLER_15_152 VPWR VGND sg13g2_decap_8
XFILLER_16_653 VPWR VGND sg13g2_fill_1
XFILLER_43_494 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_fill_2
X_1810_ _0359_ net441 ppwm_i.u_ppwm.u_mem.memory\[16\] net448 ppwm_i.u_ppwm.u_mem.memory\[2\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_12_870 VPWR VGND sg13g2_decap_8
X_2790_ _1077_ net330 ppwm_i.u_ppwm.u_mem.bit_count\[4\] _1073_ VPWR VGND sg13g2_and3_1
XFILLER_8_874 VPWR VGND sg13g2_decap_8
XFILLER_11_391 VPWR VGND sg13g2_decap_8
X_1741_ VPWR VGND _1198_ net512 net444 _1205_ _1308_ net448 sg13g2_a221oi_1
X_1672_ VPWR _1243_ net791 VGND sg13g2_inv_1
Xhold307 ppwm_i.u_ppwm.u_mem.memory\[89\] VPWR VGND net687 sg13g2_dlygate4sd3_1
XFILLER_7_395 VPWR VGND sg13g2_decap_8
Xhold318 ppwm_i.u_ppwm.u_mem.memory\[39\] VPWR VGND net698 sg13g2_dlygate4sd3_1
Xhold329 _0179_ VPWR VGND net709 sg13g2_dlygate4sd3_1
X_2224_ net396 _0366_ ppwm_i.u_ppwm.u_ex.state_q\[2\] _0649_ VPWR VGND sg13g2_nand3_1
X_2155_ VPWR VGND _0579_ _0580_ _0578_ _1213_ _0581_ ppwm_i.u_ppwm.global_counter\[16\]
+ sg13g2_a221oi_1
XFILLER_39_778 VPWR VGND sg13g2_decap_8
XFILLER_16_0 VPWR VGND sg13g2_fill_2
X_2086_ net566 _0515_ _0516_ _0188_ VPWR VGND sg13g2_nor3_1
XFILLER_26_439 VPWR VGND sg13g2_decap_8
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_21_155 VPWR VGND sg13g2_decap_8
XFILLER_22_689 VPWR VGND sg13g2_decap_8
X_2988_ net171 VGND VPWR net709 ppwm_i.u_ppwm.u_pwm.counter\[1\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
X_1939_ net215 sdr_i.mac1.sum_lvl1_ff\[8\] _0023_ VPWR VGND sg13g2_xor2_1
XFILLER_18_918 VPWR VGND sg13g2_decap_8
XFILLER_29_255 VPWR VGND sg13g2_fill_2
XFILLER_29_299 VPWR VGND sg13g2_fill_2
XFILLER_26_962 VPWR VGND sg13g2_decap_8
XFILLER_12_111 VPWR VGND sg13g2_fill_1
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_40_453 VPWR VGND sg13g2_fill_2
XFILLER_40_442 VPWR VGND sg13g2_decap_8
XFILLER_13_667 VPWR VGND sg13g2_decap_8
XFILLER_12_177 VPWR VGND sg13g2_decap_8
XFILLER_5_811 VPWR VGND sg13g2_decap_8
XFILLER_5_888 VPWR VGND sg13g2_decap_8
XFILLER_4_376 VPWR VGND sg13g2_decap_8
XFILLER_17_973 VPWR VGND sg13g2_decap_8
XFILLER_44_781 VPWR VGND sg13g2_decap_8
X_2911_ net529 VGND VPWR _0102_ sdr_i.DP_2.matrix\[36\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_16_461 VPWR VGND sg13g2_decap_8
XFILLER_16_494 VPWR VGND sg13g2_decap_8
XFILLER_32_954 VPWR VGND sg13g2_decap_8
X_2842_ net248 _0105_ VPWR VGND sg13g2_buf_1
X_2773_ VGND VPWR _1098_ net471 _0326_ _1065_ sg13g2_a21oi_1
X_1724_ VPWR VGND _1199_ _1289_ net444 _1185_ _1291_ net453 sg13g2_a221oi_1
Xhold115 sdr_i.DP_4.matrix\[72\] VPWR VGND net315 sg13g2_dlygate4sd3_1
Xhold104 sdr_i.DP_1.matrix\[27\] VPWR VGND net304 sg13g2_dlygate4sd3_1
Xhold126 ppwm_i.u_ppwm.period_start VPWR VGND net326 sg13g2_dlygate4sd3_1
Xhold148 _0279_ VPWR VGND net348 sg13g2_dlygate4sd3_1
Xhold159 _0299_ VPWR VGND net359 sg13g2_dlygate4sd3_1
Xhold137 ppwm_i.u_ppwm.u_mem.memory\[2\] VPWR VGND net337 sg13g2_dlygate4sd3_1
X_1655_ _1226_ net506 VPWR VGND sg13g2_inv_2
X_1586_ VPWR _1157_ net657 VGND sg13g2_inv_1
X_2207_ VPWR VGND _0631_ _0632_ _0630_ _1214_ _0633_ ppwm_i.u_ppwm.pwm_value\[5\]
+ sg13g2_a221oi_1
XFILLER_39_531 VPWR VGND sg13g2_decap_8
X_3187_ net525 VGND VPWR net554 sdr_i.total_sum1\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2138_ _0564_ _1222_ ppwm_i.u_ppwm.global_counter\[17\] VPWR VGND sg13g2_nand2_1
XFILLER_26_225 VPWR VGND sg13g2_fill_2
X_2069_ _0504_ _0505_ _0182_ VPWR VGND sg13g2_nor2_1
XFILLER_23_943 VPWR VGND sg13g2_decap_8
XFILLER_34_291 VPWR VGND sg13g2_decap_4
XFILLER_22_486 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
XFILLER_49_306 VPWR VGND sg13g2_fill_1
XFILLER_45_534 VPWR VGND sg13g2_fill_2
XFILLER_14_921 VPWR VGND sg13g2_decap_8
XFILLER_32_206 VPWR VGND sg13g2_fill_1
XFILLER_43_83 VPWR VGND sg13g2_decap_8
XFILLER_41_773 VPWR VGND sg13g2_decap_8
XFILLER_13_464 VPWR VGND sg13g2_decap_8
XFILLER_14_998 VPWR VGND sg13g2_decap_8
XFILLER_40_272 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_4
XFILLER_4_184 VPWR VGND sg13g2_decap_8
XFILLER_4_22 VPWR VGND sg13g2_fill_2
XFILLER_4_195 VPWR VGND sg13g2_fill_2
X_3110_ net135 VGND VPWR net369 ppwm_i.u_ppwm.u_mem.memory\[86\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
XFILLER_1_891 VPWR VGND sg13g2_decap_8
XFILLER_49_895 VPWR VGND sg13g2_decap_8
X_3041_ net67 VGND VPWR _0232_ ppwm_i.u_ppwm.u_mem.memory\[17\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_36_534 VPWR VGND sg13g2_decap_8
XFILLER_17_781 VPWR VGND sg13g2_fill_2
XFILLER_17_792 VPWR VGND sg13g2_decap_8
XFILLER_17_1015 VPWR VGND sg13g2_decap_8
XFILLER_23_239 VPWR VGND sg13g2_decap_8
X_2825_ net303 _0088_ VPWR VGND sg13g2_buf_1
XFILLER_20_968 VPWR VGND sg13g2_decap_8
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_2756_ net414 VPWR _1057_ VGND net464 net594 sg13g2_o21ai_1
X_2687_ VGND VPWR net463 _1140_ _0283_ _1022_ sg13g2_a21oi_1
X_1707_ _1275_ net324 _1267_ VPWR VGND sg13g2_nand2_1
X_1638_ VPWR _1209_ ppwm_i.u_ppwm.u_mem.memory\[0\] VGND sg13g2_inv_1
Xfanout414 net415 net414 VPWR VGND sg13g2_buf_8
Xfanout403 net404 net403 VPWR VGND sg13g2_buf_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
Xfanout436 net437 net436 VPWR VGND sg13g2_buf_8
Xfanout447 net449 net447 VPWR VGND sg13g2_buf_8
X_1569_ VPWR _1140_ net637 VGND sg13g2_inv_1
Xfanout425 net426 net425 VPWR VGND sg13g2_buf_8
XFILLER_24_1008 VPWR VGND sg13g2_decap_8
Xfanout469 net470 net469 VPWR VGND sg13g2_buf_1
Xfanout458 net459 net458 VPWR VGND sg13g2_buf_8
XFILLER_39_394 VPWR VGND sg13g2_fill_1
XFILLER_42_504 VPWR VGND sg13g2_decap_8
XFILLER_14_217 VPWR VGND sg13g2_fill_1
XFILLER_11_902 VPWR VGND sg13g2_decap_8
XFILLER_7_906 VPWR VGND sg13g2_decap_8
XFILLER_13_20 VPWR VGND sg13g2_fill_1
XFILLER_22_294 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_11_979 VPWR VGND sg13g2_decap_8
XFILLER_13_86 VPWR VGND sg13g2_decap_8
XFILLER_8_2 VPWR VGND sg13g2_fill_1
XFILLER_49_103 VPWR VGND sg13g2_decap_8
XFILLER_46_843 VPWR VGND sg13g2_decap_8
XFILLER_18_512 VPWR VGND sg13g2_decap_8
XFILLER_18_523 VPWR VGND sg13g2_fill_1
XFILLER_33_548 VPWR VGND sg13g2_decap_8
XFILLER_41_570 VPWR VGND sg13g2_fill_1
XFILLER_13_250 VPWR VGND sg13g2_fill_1
X_2610_ net425 VPWR _0984_ VGND net484 ppwm_i.u_ppwm.u_mem.memory\[30\] sg13g2_o21ai_1
X_2541_ VPWR VGND _0946_ net459 _0943_ _1211_ _0213_ net370 sg13g2_a221oi_1
XFILLER_6_961 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
X_2472_ VGND VPWR net380 _0883_ _0884_ _0727_ sg13g2_a21oi_1
XFILLER_49_670 VPWR VGND sg13g2_decap_8
X_3024_ net101 VGND VPWR net344 ppwm_i.u_ppwm.u_mem.memory\[0\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_2987__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_37_865 VPWR VGND sg13g2_decap_8
XFILLER_20_721 VPWR VGND sg13g2_decap_4
Xclkload7 VPWR clkload7/Y clknet_leaf_32_clk VGND sg13g2_inv_1
X_2808_ _1092_ VPWR _1093_ VGND _1089_ _1091_ sg13g2_o21ai_1
XFILLER_4_909 VPWR VGND sg13g2_decap_8
X_2739_ VGND VPWR net468 _1114_ _0309_ _1048_ sg13g2_a21oi_1
XFILLER_47_607 VPWR VGND sg13g2_decap_4
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_43_824 VPWR VGND sg13g2_decap_8
XFILLER_15_548 VPWR VGND sg13g2_decap_8
XFILLER_27_397 VPWR VGND sg13g2_decap_8
XFILLER_11_721 VPWR VGND sg13g2_fill_2
XFILLER_24_74 VPWR VGND sg13g2_fill_2
XFILLER_10_253 VPWR VGND sg13g2_fill_2
XFILLER_11_754 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_3_931 VPWR VGND sg13g2_decap_8
XFILLER_49_82 VPWR VGND sg13g2_decap_8
XFILLER_2_485 VPWR VGND sg13g2_fill_2
XFILLER_27_8 VPWR VGND sg13g2_fill_1
XFILLER_19_821 VPWR VGND sg13g2_fill_1
XFILLER_18_320 VPWR VGND sg13g2_fill_2
XFILLER_45_172 VPWR VGND sg13g2_decap_4
XFILLER_33_334 VPWR VGND sg13g2_fill_2
XFILLER_34_868 VPWR VGND sg13g2_decap_8
X_1972_ net602 VPWR _0006_ VGND _0416_ _0418_ sg13g2_o21ai_1
X_2524_ net381 _0822_ _0931_ VPWR VGND sg13g2_nor2_1
X_2455_ _1218_ _0341_ _0347_ _0868_ VPWR VGND sg13g2_nor3_1
Xhold19 sdr_i.DP_3.matrix\[10\] VPWR VGND net219 sg13g2_dlygate4sd3_1
X_2386_ _0763_ VPWR _0804_ VGND _0663_ _0667_ sg13g2_o21ai_1
XFILLER_43_109 VPWR VGND sg13g2_decap_4
X_3007_ net134 VGND VPWR _0198_ ppwm_i.u_ppwm.pwm_value\[3\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_37_684 VPWR VGND sg13g2_decap_8
XFILLER_37_695 VPWR VGND sg13g2_fill_1
XFILLER_20_595 VPWR VGND sg13g2_fill_1
XFILLER_0_934 VPWR VGND sg13g2_decap_8
XFILLER_48_905 VPWR VGND sg13g2_decap_8
XFILLER_47_437 VPWR VGND sg13g2_decap_8
XFILLER_47_415 VPWR VGND sg13g2_decap_8
XFILLER_19_128 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_fill_2
XFILLER_28_640 VPWR VGND sg13g2_decap_8
XFILLER_16_835 VPWR VGND sg13g2_fill_1
XFILLER_43_654 VPWR VGND sg13g2_fill_2
XFILLER_43_643 VPWR VGND sg13g2_fill_1
XFILLER_15_334 VPWR VGND sg13g2_decap_8
XFILLER_15_345 VPWR VGND sg13g2_fill_1
XFILLER_27_172 VPWR VGND sg13g2_fill_1
XFILLER_30_326 VPWR VGND sg13g2_fill_1
XFILLER_31_849 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_fill_1
XFILLER_11_584 VPWR VGND sg13g2_fill_2
X_2240_ _1216_ net398 _0664_ VPWR VGND sg13g2_nor2_1
XFILLER_38_437 VPWR VGND sg13g2_decap_8
X_2171_ _0597_ _1263_ ppwm_i.u_ppwm.pwm_value\[4\] _1262_ ppwm_i.u_ppwm.pwm_value\[5\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_18_161 VPWR VGND sg13g2_decap_4
XFILLER_19_662 VPWR VGND sg13g2_decap_4
XFILLER_19_695 VPWR VGND sg13g2_fill_1
XFILLER_22_827 VPWR VGND sg13g2_decap_4
XFILLER_33_164 VPWR VGND sg13g2_fill_1
X_1955_ net257 sdr_i.mac2.products_ff\[102\] _0038_ VPWR VGND sg13g2_xor2_1
XFILLER_30_860 VPWR VGND sg13g2_decap_8
X_1886_ sdr_i.mac1.products_ff\[18\] sdr_i.mac1.products_ff\[1\] _0407_ VPWR VGND
+ sg13g2_xor2_1
X_2507_ _1213_ net393 _0915_ VPWR VGND sg13g2_nor2_1
X_2438_ _0853_ _0852_ _0673_ _0676_ net805 VPWR VGND sg13g2_a22oi_1
X_2369_ _0659_ _0787_ _0788_ VPWR VGND sg13g2_and2_1
XFILLER_29_426 VPWR VGND sg13g2_fill_1
XFILLER_45_919 VPWR VGND sg13g2_decap_8
XFILLER_25_632 VPWR VGND sg13g2_decap_8
XFILLER_37_492 VPWR VGND sg13g2_decap_8
XFILLER_25_665 VPWR VGND sg13g2_decap_8
XFILLER_40_624 VPWR VGND sg13g2_decap_8
XFILLER_12_315 VPWR VGND sg13g2_decap_4
XFILLER_12_326 VPWR VGND sg13g2_fill_1
XFILLER_0_731 VPWR VGND sg13g2_decap_8
XFILLER_48_779 VPWR VGND sg13g2_decap_8
XFILLER_47_256 VPWR VGND sg13g2_decap_4
XFILLER_36_919 VPWR VGND sg13g2_decap_8
XFILLER_46_50 VPWR VGND sg13g2_fill_2
X_3068__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_28_481 VPWR VGND sg13g2_decap_8
XFILLER_44_963 VPWR VGND sg13g2_decap_8
XFILLER_15_131 VPWR VGND sg13g2_decap_8
XFILLER_8_853 VPWR VGND sg13g2_decap_8
XFILLER_7_341 VPWR VGND sg13g2_fill_2
X_1740_ _1307_ net440 _1191_ net453 _1184_ VPWR VGND sg13g2_a22oi_1
X_1671_ VPWR _1242_ net802 VGND sg13g2_inv_1
X_3075__137 VPWR VGND net137 sg13g2_tiehi
Xhold308 ppwm_i.u_ppwm.u_mem.memory\[33\] VPWR VGND net688 sg13g2_dlygate4sd3_1
Xhold319 ppwm_i.u_ppwm.u_mem.memory\[40\] VPWR VGND net699 sg13g2_dlygate4sd3_1
XFILLER_39_713 VPWR VGND sg13g2_fill_2
X_2223_ VGND VPWR net350 _0648_ _0193_ net458 sg13g2_a21oi_1
X_2154_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] ppwm_i.u_ppwm.global_counter\[17\] _0580_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_27_919 VPWR VGND sg13g2_decap_8
XFILLER_38_234 VPWR VGND sg13g2_decap_8
X_2085_ ppwm_i.u_ppwm.u_pwm.counter\[6\] ppwm_i.u_ppwm.u_pwm.counter\[1\] ppwm_i.u_ppwm.u_pwm.counter\[7\]
+ _0516_ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[0\] sg13g2_nand4_1
XFILLER_35_941 VPWR VGND sg13g2_decap_8
XFILLER_34_440 VPWR VGND sg13g2_decap_8
XFILLER_22_635 VPWR VGND sg13g2_fill_1
XFILLER_10_819 VPWR VGND sg13g2_decap_8
X_2987_ net173 VGND VPWR _0178_ ppwm_i.u_ppwm.u_pwm.counter\[0\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
X_1938_ _0430_ sdr_i.mac1.sum_lvl1_ff\[8\] net215 VPWR VGND sg13g2_nand2_1
X_1869_ _0402_ net284 net232 VPWR VGND sg13g2_nand2_1
XFILLER_27_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_201 VPWR VGND sg13g2_decap_8
XFILLER_44_237 VPWR VGND sg13g2_decap_4
XFILLER_26_941 VPWR VGND sg13g2_decap_8
XFILLER_13_635 VPWR VGND sg13g2_decap_4
XFILLER_25_484 VPWR VGND sg13g2_decap_8
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_40_421 VPWR VGND sg13g2_decap_8
XFILLER_9_617 VPWR VGND sg13g2_fill_1
XFILLER_8_127 VPWR VGND sg13g2_decap_8
XFILLER_10_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_867 VPWR VGND sg13g2_decap_8
XFILLER_4_355 VPWR VGND sg13g2_decap_8
XFILLER_0_583 VPWR VGND sg13g2_decap_8
XFILLER_48_543 VPWR VGND sg13g2_fill_1
XFILLER_17_952 VPWR VGND sg13g2_decap_8
X_2910_ net535 VGND VPWR _0101_ sdr_i.DP_2.matrix\[28\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_32_933 VPWR VGND sg13g2_decap_8
XFILLER_31_443 VPWR VGND sg13g2_decap_4
X_2841_ net311 _0104_ VPWR VGND sg13g2_buf_1
X_3036__77 VPWR VGND net77 sg13g2_tiehi
X_2772_ net414 VPWR _1065_ VGND net582 net471 sg13g2_o21ai_1
X_1723_ VGND VPWR _1192_ net441 _1290_ net512 sg13g2_a21oi_1
XFILLER_8_694 VPWR VGND sg13g2_fill_2
Xhold105 sdr_i.mac1.sum_lvl2_ff\[0\] VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold116 sdr_i.DP_3.matrix\[72\] VPWR VGND net316 sg13g2_dlygate4sd3_1
Xhold138 _0216_ VPWR VGND net338 sg13g2_dlygate4sd3_1
Xhold149 ppwm_i.u_ppwm.u_ex.cmp_flag_q VPWR VGND net349 sg13g2_dlygate4sd3_1
Xhold127 _0148_ VPWR VGND net327 sg13g2_dlygate4sd3_1
X_1654_ net505 _1225_ VPWR VGND sg13g2_inv_4
X_1585_ VPWR _1156_ ppwm_i.u_ppwm.u_mem.memory\[53\] VGND sg13g2_inv_1
XFILLER_39_510 VPWR VGND sg13g2_decap_8
X_2206_ ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] _1223_ _0632_ VPWR VGND sg13g2_nor2_1
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
X_3186_ net525 VGND VPWR net775 sdr_i.mac1.total_sum\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_26_204 VPWR VGND sg13g2_decap_8
X_2137_ VPWR VGND _0561_ _0562_ _0560_ net504 _0563_ _1254_ sg13g2_a221oi_1
XFILLER_27_749 VPWR VGND sg13g2_decap_4
X_2068_ net422 VPWR _0505_ VGND net785 _0502_ sg13g2_o21ai_1
XFILLER_23_922 VPWR VGND sg13g2_decap_8
XFILLER_22_421 VPWR VGND sg13g2_decap_8
XFILLER_22_465 VPWR VGND sg13g2_decap_8
XFILLER_23_999 VPWR VGND sg13g2_decap_8
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
X_2997__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_40_1025 VPWR VGND sg13g2_decap_4
XFILLER_17_204 VPWR VGND sg13g2_decap_8
XFILLER_45_557 VPWR VGND sg13g2_fill_1
XFILLER_14_900 VPWR VGND sg13g2_decap_8
XFILLER_41_752 VPWR VGND sg13g2_decap_4
XFILLER_14_977 VPWR VGND sg13g2_decap_8
XFILLER_9_436 VPWR VGND sg13g2_decap_8
XFILLER_13_498 VPWR VGND sg13g2_fill_2
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_1_870 VPWR VGND sg13g2_decap_8
XFILLER_49_874 VPWR VGND sg13g2_decap_8
X_3040_ net69 VGND VPWR net353 ppwm_i.u_ppwm.u_mem.memory\[16\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_48_384 VPWR VGND sg13g2_decap_8
XFILLER_36_513 VPWR VGND sg13g2_decap_8
X_2824_ net244 _0087_ VPWR VGND sg13g2_buf_1
XFILLER_20_947 VPWR VGND sg13g2_decap_8
X_2755_ VGND VPWR net472 _1106_ _0317_ _1056_ sg13g2_a21oi_1
X_2686_ net413 VPWR _1022_ VGND net463 net574 sg13g2_o21ai_1
X_1706_ _0004_ _1273_ _1274_ VPWR VGND sg13g2_nand2_1
X_1637_ VPWR _1208_ net343 VGND sg13g2_inv_1
Xfanout404 _1295_ net404 VPWR VGND sg13g2_buf_2
X_1568_ VPWR _1139_ net667 VGND sg13g2_inv_1
Xfanout426 net427 net426 VPWR VGND sg13g2_buf_8
Xfanout448 net449 net448 VPWR VGND sg13g2_buf_8
Xfanout415 net420 net415 VPWR VGND sg13g2_buf_8
Xfanout437 ppwm_i.rst_n net437 VPWR VGND sg13g2_buf_8
Xfanout459 _1266_ net459 VPWR VGND sg13g2_buf_8
X_3169_ net530 VGND VPWR net763 sdr_i.mac1.sum_lvl1_ff\[25\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_23_752 VPWR VGND sg13g2_fill_1
XFILLER_23_774 VPWR VGND sg13g2_fill_1
XFILLER_11_958 VPWR VGND sg13g2_decap_8
XFILLER_22_273 VPWR VGND sg13g2_decap_8
XFILLER_13_65 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_decap_8
XFILLER_45_354 VPWR VGND sg13g2_fill_1
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_46_899 VPWR VGND sg13g2_decap_8
XFILLER_6_940 VPWR VGND sg13g2_decap_8
X_2540_ _0946_ _0838_ _0860_ _0945_ VPWR VGND sg13g2_and3_1
X_2471_ VGND VPWR _1227_ net383 _0883_ _0882_ sg13g2_a21oi_1
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
X_3023_ net103 VGND VPWR _0214_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
XFILLER_37_844 VPWR VGND sg13g2_decap_8
XFILLER_36_354 VPWR VGND sg13g2_decap_4
XFILLER_36_398 VPWR VGND sg13g2_decap_8
Xclkload8 VPWR clkload8/Y clknet_leaf_19_clk VGND sg13g2_inv_1
X_2807_ _1092_ ppwm_i.u_ppwm.u_pwm.cmp_value\[7\] _1237_ ppwm_i.u_ppwm.u_pwm.cmp_value\[8\]
+ _1236_ VPWR VGND sg13g2_a22oi_1
X_2738_ net419 VPWR _1048_ VGND net474 ppwm_i.u_ppwm.u_mem.memory\[94\] sg13g2_o21ai_1
X_2669_ VGND VPWR net466 _1149_ _0274_ _1013_ sg13g2_a21oi_1
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
XFILLER_43_803 VPWR VGND sg13g2_decap_8
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_42_302 VPWR VGND sg13g2_decap_8
XFILLER_15_505 VPWR VGND sg13g2_decap_8
XFILLER_11_700 VPWR VGND sg13g2_decap_8
XFILLER_10_232 VPWR VGND sg13g2_decap_8
XFILLER_40_30 VPWR VGND sg13g2_decap_8
XFILLER_6_269 VPWR VGND sg13g2_fill_2
XFILLER_3_910 VPWR VGND sg13g2_decap_8
XFILLER_3_987 VPWR VGND sg13g2_decap_8
XFILLER_18_310 VPWR VGND sg13g2_fill_1
XFILLER_46_652 VPWR VGND sg13g2_fill_1
XFILLER_46_674 VPWR VGND sg13g2_fill_1
XFILLER_45_151 VPWR VGND sg13g2_decap_8
XFILLER_18_376 VPWR VGND sg13g2_decap_8
XFILLER_19_888 VPWR VGND sg13g2_decap_8
XFILLER_33_302 VPWR VGND sg13g2_fill_1
XFILLER_46_696 VPWR VGND sg13g2_decap_4
XFILLER_34_847 VPWR VGND sg13g2_decap_8
XFILLER_21_508 VPWR VGND sg13g2_fill_1
X_1971_ _0447_ _0446_ _0043_ VPWR VGND sg13g2_xor2_1
XFILLER_14_1019 VPWR VGND sg13g2_decap_8
X_2523_ VGND VPWR _0926_ _0928_ _0930_ _0685_ sg13g2_a21oi_1
X_2454_ _1218_ VPWR _0867_ VGND _0341_ _0347_ sg13g2_o21ai_1
X_2385_ _0764_ VPWR _0803_ VGND _0657_ _0724_ sg13g2_o21ai_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_29_608 VPWR VGND sg13g2_decap_8
Xinput1 ena net1 VPWR VGND sg13g2_buf_2
XFILLER_37_652 VPWR VGND sg13g2_decap_8
X_3006_ net136 VGND VPWR _0197_ ppwm_i.u_ppwm.pwm_value\[2\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_36_184 VPWR VGND sg13g2_fill_2
XFILLER_36_195 VPWR VGND sg13g2_decap_8
XFILLER_0_913 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_39_clk clknet_3_4__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_16_825 VPWR VGND sg13g2_fill_2
XFILLER_43_622 VPWR VGND sg13g2_decap_8
XFILLER_35_41 VPWR VGND sg13g2_decap_4
XFILLER_43_666 VPWR VGND sg13g2_decap_4
XFILLER_37_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_828 VPWR VGND sg13g2_decap_8
X_3090__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_7_545 VPWR VGND sg13g2_decap_8
XFILLER_3_784 VPWR VGND sg13g2_decap_8
XFILLER_39_939 VPWR VGND sg13g2_decap_8
X_2170_ _0595_ VPWR _0596_ VGND net505 _1263_ sg13g2_o21ai_1
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_46_460 VPWR VGND sg13g2_decap_8
XFILLER_18_140 VPWR VGND sg13g2_decap_8
XFILLER_19_685 VPWR VGND sg13g2_decap_4
XFILLER_46_471 VPWR VGND sg13g2_fill_1
XFILLER_33_143 VPWR VGND sg13g2_decap_8
XFILLER_33_187 VPWR VGND sg13g2_decap_8
XFILLER_34_688 VPWR VGND sg13g2_fill_1
XFILLER_21_349 VPWR VGND sg13g2_fill_2
X_1954_ _0438_ net739 net257 VPWR VGND sg13g2_nand2_1
X_1885_ net285 net274 _0054_ VPWR VGND sg13g2_and2_1
X_2506_ VPWR VGND _0914_ net459 _0911_ _1214_ _0210_ net370 sg13g2_a221oi_1
X_2437_ _0851_ VPWR _0852_ VGND _1259_ net402 sg13g2_o21ai_1
X_2368_ _0766_ _0785_ net386 _0787_ VPWR VGND sg13g2_mux2_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_405 VPWR VGND sg13g2_fill_2
X_2299_ VPWR VGND net386 _0720_ _0695_ _0350_ _0721_ _0655_ sg13g2_a221oi_1
XFILLER_44_408 VPWR VGND sg13g2_decap_8
XFILLER_38_994 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_fill_1
XFILLER_40_647 VPWR VGND sg13g2_fill_1
XFILLER_4_559 VPWR VGND sg13g2_decap_8
XFILLER_0_710 VPWR VGND sg13g2_decap_8
XFILLER_0_787 VPWR VGND sg13g2_decap_8
XFILLER_48_758 VPWR VGND sg13g2_decap_8
XFILLER_47_279 VPWR VGND sg13g2_fill_2
XFILLER_28_460 VPWR VGND sg13g2_decap_8
XFILLER_29_983 VPWR VGND sg13g2_decap_8
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_16_633 VPWR VGND sg13g2_decap_8
XFILLER_43_430 VPWR VGND sg13g2_decap_4
X_3048__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_31_625 VPWR VGND sg13g2_decap_8
X_1670_ VPWR _1241_ net725 VGND sg13g2_inv_1
XFILLER_7_67 VPWR VGND sg13g2_decap_4
Xhold309 _0247_ VPWR VGND net689 sg13g2_dlygate4sd3_1
XFILLER_3_592 VPWR VGND sg13g2_fill_2
XFILLER_30_4 VPWR VGND sg13g2_fill_1
XFILLER_39_736 VPWR VGND sg13g2_fill_2
X_2222_ _0645_ _0623_ _0647_ _0648_ VPWR VGND sg13g2_a21o_1
X_2153_ _0579_ _1255_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] _1254_ net502 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_39_747 VPWR VGND sg13g2_fill_2
XFILLER_38_213 VPWR VGND sg13g2_decap_8
XFILLER_38_246 VPWR VGND sg13g2_decap_4
XFILLER_47_791 VPWR VGND sg13g2_decap_8
X_2084_ ppwm_i.u_ppwm.u_pwm.counter\[8\] net423 ppwm_i.u_ppwm.u_pwm.counter\[9\] _0515_
+ VPWR VGND sg13g2_nand3_1
XFILLER_35_920 VPWR VGND sg13g2_decap_8
XFILLER_22_614 VPWR VGND sg13g2_decap_8
XFILLER_34_485 VPWR VGND sg13g2_decap_4
XFILLER_35_997 VPWR VGND sg13g2_decap_8
X_2986_ net175 VGND VPWR _0177_ ppwm_i.u_ppwm.u_pwm.cmp_value\[9\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_1937_ _0022_ _0428_ net762 VPWR VGND sg13g2_xnor2_1
X_1868_ _0401_ _0400_ _0071_ VPWR VGND sg13g2_xor2_1
X_1799_ _0341_ _0347_ _0348_ VPWR VGND sg13g2_nor2_1
X_3132__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_26_920 VPWR VGND sg13g2_decap_8
XFILLER_38_791 VPWR VGND sg13g2_decap_8
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_13_614 VPWR VGND sg13g2_fill_2
XFILLER_16_65 VPWR VGND sg13g2_decap_8
XFILLER_16_87 VPWR VGND sg13g2_decap_8
XFILLER_26_997 VPWR VGND sg13g2_decap_8
XFILLER_12_135 VPWR VGND sg13g2_fill_2
XFILLER_40_466 VPWR VGND sg13g2_decap_4
XFILLER_8_106 VPWR VGND sg13g2_decap_8
XFILLER_12_146 VPWR VGND sg13g2_decap_8
XFILLER_32_31 VPWR VGND sg13g2_fill_1
XFILLER_40_488 VPWR VGND sg13g2_decap_4
XFILLER_10_1000 VPWR VGND sg13g2_decap_8
XFILLER_5_846 VPWR VGND sg13g2_decap_8
XFILLER_0_562 VPWR VGND sg13g2_decap_8
XFILLER_17_931 VPWR VGND sg13g2_decap_8
XFILLER_29_780 VPWR VGND sg13g2_decap_8
XFILLER_35_249 VPWR VGND sg13g2_decap_8
XFILLER_32_912 VPWR VGND sg13g2_decap_8
XFILLER_43_293 VPWR VGND sg13g2_decap_8
X_2840_ net249 _0103_ VPWR VGND sg13g2_buf_1
XFILLER_32_989 VPWR VGND sg13g2_decap_8
X_2771_ VGND VPWR _1097_ net471 _0325_ _1064_ sg13g2_a21oi_1
X_3051__48 VPWR VGND net48 sg13g2_tiehi
X_1722_ ppwm_i.u_ppwm.u_mem.memory\[3\] net516 net519 _1289_ VPWR VGND sg13g2_nor3_1
X_1653_ ppwm_i.u_ppwm.pwm_value\[5\] _1224_ VPWR VGND sg13g2_inv_4
Xhold106 _0027_ VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold117 ppwm_i.u_ppwm.u_ex.state_q\[1\] VPWR VGND net317 sg13g2_dlygate4sd3_1
Xhold128 ppwm_i.u_ppwm.global_counter\[19\] VPWR VGND net328 sg13g2_dlygate4sd3_1
Xhold139 ppwm_i.u_ppwm.u_mem.bit_count\[1\] VPWR VGND net339 sg13g2_dlygate4sd3_1
X_1584_ VPWR _1155_ net669 VGND sg13g2_inv_1
X_2205_ _0631_ _1225_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] _1224_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\]
+ VPWR VGND sg13g2_a22oi_1
X_3185_ net525 VGND VPWR net262 sdr_i.mac1.total_sum\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2136_ _1224_ ppwm_i.u_ppwm.global_counter\[15\] _0562_ VPWR VGND sg13g2_nor2_1
X_2067_ net785 _0502_ _0504_ VPWR VGND sg13g2_and2_1
XFILLER_26_238 VPWR VGND sg13g2_decap_4
XFILLER_23_901 VPWR VGND sg13g2_decap_8
XFILLER_35_794 VPWR VGND sg13g2_decap_8
XFILLER_23_978 VPWR VGND sg13g2_decap_8
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
X_2969_ net435 VGND VPWR net721 ppwm_i.u_ppwm.global_counter\[12\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_5_109 VPWR VGND sg13g2_fill_2
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_1_348 VPWR VGND sg13g2_decap_8
XFILLER_40_1004 VPWR VGND sg13g2_decap_8
XFILLER_45_503 VPWR VGND sg13g2_fill_2
XFILLER_45_525 VPWR VGND sg13g2_fill_1
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_17_249 VPWR VGND sg13g2_decap_8
XFILLER_25_260 VPWR VGND sg13g2_fill_1
XFILLER_14_956 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_fill_2
XFILLER_5_665 VPWR VGND sg13g2_decap_8
XFILLER_4_24 VPWR VGND sg13g2_fill_1
XFILLER_0_381 VPWR VGND sg13g2_decap_8
XFILLER_49_853 VPWR VGND sg13g2_decap_8
XFILLER_36_569 VPWR VGND sg13g2_decap_8
XFILLER_17_783 VPWR VGND sg13g2_fill_1
XFILLER_20_926 VPWR VGND sg13g2_decap_8
X_2823_ net279 _0086_ VPWR VGND sg13g2_buf_1
XFILLER_32_786 VPWR VGND sg13g2_decap_8
X_2754_ net415 VPWR _1056_ VGND net472 ppwm_i.u_ppwm.u_mem.memory\[102\] sg13g2_o21ai_1
XFILLER_9_982 VPWR VGND sg13g2_decap_8
X_1705_ net715 net421 _1098_ _1274_ VPWR VGND sg13g2_nand3_1
X_2685_ VGND VPWR net467 _1141_ _0282_ _1021_ sg13g2_a21oi_1
X_1636_ VPWR _1207_ net337 VGND sg13g2_inv_1
X_1567_ VPWR _1138_ ppwm_i.u_ppwm.u_mem.memory\[71\] VGND sg13g2_inv_1
Xfanout405 net406 net405 VPWR VGND sg13g2_buf_2
Xfanout416 net418 net416 VPWR VGND sg13g2_buf_8
Xfanout427 net434 net427 VPWR VGND sg13g2_buf_8
Xfanout438 _1283_ net438 VPWR VGND sg13g2_buf_8
Xfanout449 _1280_ net449 VPWR VGND sg13g2_buf_8
X_3168_ net529 VGND VPWR net231 sdr_i.mac1.sum_lvl1_ff\[24\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_15_709 VPWR VGND sg13g2_fill_1
X_2119_ _0546_ _0542_ _0545_ _1232_ net508 VPWR VGND sg13g2_a22oi_1
X_3099_ net43 VGND VPWR _0290_ ppwm_i.u_ppwm.u_mem.memory\[75\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3064__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_22_230 VPWR VGND sg13g2_decap_4
XFILLER_10_414 VPWR VGND sg13g2_fill_2
XFILLER_11_937 VPWR VGND sg13g2_decap_8
XFILLER_10_469 VPWR VGND sg13g2_fill_1
XFILLER_2_624 VPWR VGND sg13g2_decap_4
XFILLER_49_138 VPWR VGND sg13g2_decap_8
XFILLER_46_801 VPWR VGND sg13g2_decap_8
XFILLER_46_878 VPWR VGND sg13g2_decap_8
XFILLER_45_377 VPWR VGND sg13g2_decap_4
XFILLER_33_517 VPWR VGND sg13g2_decap_8
XFILLER_14_753 VPWR VGND sg13g2_decap_8
XFILLER_41_583 VPWR VGND sg13g2_decap_8
XFILLER_9_201 VPWR VGND sg13g2_fill_2
XFILLER_9_278 VPWR VGND sg13g2_fill_2
XFILLER_6_996 VPWR VGND sg13g2_decap_8
XFILLER_5_462 VPWR VGND sg13g2_decap_8
X_2470_ net383 _0729_ _0882_ VPWR VGND sg13g2_nor2_1
X_3022_ net105 VGND VPWR net810 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
XFILLER_36_300 VPWR VGND sg13g2_decap_4
XFILLER_37_823 VPWR VGND sg13g2_decap_8
XFILLER_24_517 VPWR VGND sg13g2_decap_8
XFILLER_24_528 VPWR VGND sg13g2_fill_2
XFILLER_24_539 VPWR VGND sg13g2_decap_8
XFILLER_20_756 VPWR VGND sg13g2_decap_8
Xclkload9 clkload9/Y clknet_leaf_22_clk VPWR VGND sg13g2_inv_8
X_2806_ _1090_ VPWR _1091_ VGND _1238_ ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] sg13g2_o21ai_1
XFILLER_30_1014 VPWR VGND sg13g2_decap_8
X_2737_ VGND VPWR net474 _1115_ _0308_ _1047_ sg13g2_a21oi_1
X_2668_ net416 VPWR _1013_ VGND net474 ppwm_i.u_ppwm.u_mem.memory\[59\] sg13g2_o21ai_1
X_1619_ VPWR _1190_ net705 VGND sg13g2_inv_1
X_2599_ VGND VPWR net497 _1184_ _0239_ _0978_ sg13g2_a21oi_1
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_27_333 VPWR VGND sg13g2_fill_1
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_42_325 VPWR VGND sg13g2_fill_2
XFILLER_24_32 VPWR VGND sg13g2_fill_2
XFILLER_23_561 VPWR VGND sg13g2_decap_8
XFILLER_40_20 VPWR VGND sg13g2_fill_1
XFILLER_10_255 VPWR VGND sg13g2_fill_1
XFILLER_3_966 VPWR VGND sg13g2_decap_8
XFILLER_2_454 VPWR VGND sg13g2_fill_1
XFILLER_49_51 VPWR VGND sg13g2_decap_8
XFILLER_49_40 VPWR VGND sg13g2_decap_8
XFILLER_19_812 VPWR VGND sg13g2_decap_8
XFILLER_18_355 VPWR VGND sg13g2_decap_8
XFILLER_34_826 VPWR VGND sg13g2_decap_8
XFILLER_33_314 VPWR VGND sg13g2_fill_1
X_1970_ _0447_ net275 net235 VPWR VGND sg13g2_nand2_1
XFILLER_42_881 VPWR VGND sg13g2_decap_8
XFILLER_14_561 VPWR VGND sg13g2_fill_2
X_3078__125 VPWR VGND net125 sg13g2_tiehi
X_2522_ _0929_ _0927_ _0926_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_292 VPWR VGND sg13g2_decap_4
X_2453_ VPWR VGND _0669_ net458 _0866_ _1219_ _0205_ net370 sg13g2_a221oi_1
X_2384_ VGND VPWR _0796_ _0800_ _0802_ _0801_ sg13g2_a21oi_1
Xinput2 rst_n net2 VPWR VGND sg13g2_buf_2
XFILLER_28_119 VPWR VGND sg13g2_decap_8
XFILLER_49_491 VPWR VGND sg13g2_fill_1
XFILLER_49_480 VPWR VGND sg13g2_decap_8
X_3005_ net138 VGND VPWR net832 ppwm_i.u_ppwm.pwm_value\[1\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_25_859 VPWR VGND sg13g2_decap_8
XFILLER_12_509 VPWR VGND sg13g2_decap_8
XFILLER_40_829 VPWR VGND sg13g2_decap_8
XFILLER_33_881 VPWR VGND sg13g2_decap_8
XFILLER_20_520 VPWR VGND sg13g2_fill_2
XFILLER_20_542 VPWR VGND sg13g2_fill_2
XFILLER_10_89 VPWR VGND sg13g2_fill_2
XFILLER_0_969 VPWR VGND sg13g2_decap_8
XFILLER_19_76 VPWR VGND sg13g2_decap_8
XFILLER_15_314 VPWR VGND sg13g2_fill_2
XFILLER_28_697 VPWR VGND sg13g2_decap_8
XFILLER_43_656 VPWR VGND sg13g2_fill_1
XFILLER_31_807 VPWR VGND sg13g2_decap_8
XFILLER_23_380 VPWR VGND sg13g2_decap_4
XFILLER_7_524 VPWR VGND sg13g2_decap_8
XFILLER_7_502 VPWR VGND sg13g2_decap_8
XFILLER_3_763 VPWR VGND sg13g2_decap_8
XFILLER_2_251 VPWR VGND sg13g2_decap_8
XFILLER_39_918 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_18_130 VPWR VGND sg13g2_fill_1
XFILLER_20_1024 VPWR VGND sg13g2_decap_4
XFILLER_34_634 VPWR VGND sg13g2_fill_2
XFILLER_22_807 VPWR VGND sg13g2_fill_2
XFILLER_33_122 VPWR VGND sg13g2_decap_8
XFILLER_34_645 VPWR VGND sg13g2_decap_8
X_1953_ _0035_ _0436_ _0437_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_892 VPWR VGND sg13g2_decap_8
XFILLER_21_339 VPWR VGND sg13g2_decap_4
X_1884_ net217 sdr_i.mac1.products_ff\[0\] _0015_ VPWR VGND sg13g2_xor2_1
XFILLER_30_895 VPWR VGND sg13g2_decap_8
X_2505_ _0914_ _0789_ net374 _0913_ VPWR VGND sg13g2_and3_1
X_2436_ _0851_ ppwm_i.u_ppwm.global_counter\[19\] net402 VPWR VGND sg13g2_nand2_1
X_2367_ net386 _0766_ _0786_ VPWR VGND sg13g2_nor2_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_2298_ _0720_ net392 _0691_ VPWR VGND sg13g2_nand2_1
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_25_612 VPWR VGND sg13g2_fill_2
XFILLER_21_884 VPWR VGND sg13g2_decap_8
XFILLER_4_516 VPWR VGND sg13g2_fill_2
XFILLER_4_538 VPWR VGND sg13g2_decap_8
XFILLER_21_66 VPWR VGND sg13g2_decap_8
XFILLER_21_99 VPWR VGND sg13g2_fill_2
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_48_737 VPWR VGND sg13g2_decap_8
XFILLER_0_766 VPWR VGND sg13g2_decap_8
XFILLER_29_962 VPWR VGND sg13g2_decap_8
XFILLER_46_74 VPWR VGND sg13g2_fill_1
XFILLER_44_921 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_fill_2
X_3109__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_44_998 VPWR VGND sg13g2_decap_8
XFILLER_43_475 VPWR VGND sg13g2_decap_8
XFILLER_15_166 VPWR VGND sg13g2_fill_2
XFILLER_12_840 VPWR VGND sg13g2_decap_4
XFILLER_8_811 VPWR VGND sg13g2_fill_1
XFILLER_8_800 VPWR VGND sg13g2_fill_1
XFILLER_7_46 VPWR VGND sg13g2_decap_8
XFILLER_7_13 VPWR VGND sg13g2_decap_8
XFILLER_12_884 VPWR VGND sg13g2_decap_8
XFILLER_8_888 VPWR VGND sg13g2_decap_8
X_2221_ _0647_ _0549_ _0646_ VPWR VGND sg13g2_nand2_1
XFILLER_39_715 VPWR VGND sg13g2_fill_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
X_2152_ _0577_ VPWR _0578_ VGND _0574_ _0576_ sg13g2_o21ai_1
X_2083_ net455 net753 _0187_ VPWR VGND sg13g2_nor2_1
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_19_483 VPWR VGND sg13g2_decap_8
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_22_604 VPWR VGND sg13g2_decap_4
X_2985_ net177 VGND VPWR _0176_ ppwm_i.u_ppwm.u_pwm.cmp_value\[8\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_1936_ net761 sdr_i.mac1.products_ff\[120\] _0429_ VPWR VGND sg13g2_xor2_1
XFILLER_30_681 VPWR VGND sg13g2_fill_1
X_1867_ _0401_ net316 net246 VPWR VGND sg13g2_nand2_1
X_1798_ VPWR VGND _0346_ net509 _0345_ _0342_ _0347_ _0343_ sg13g2_a221oi_1
X_2419_ _0833_ _0834_ net377 _0835_ VPWR VGND sg13g2_nand3_1
X_3117__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_44_217 VPWR VGND sg13g2_decap_8
XFILLER_38_770 VPWR VGND sg13g2_decap_8
XFILLER_26_976 VPWR VGND sg13g2_decap_8
XFILLER_41_913 VPWR VGND sg13g2_decap_8
XFILLER_40_401 VPWR VGND sg13g2_decap_8
XFILLER_40_412 VPWR VGND sg13g2_fill_1
XFILLER_21_670 VPWR VGND sg13g2_fill_1
XFILLER_32_43 VPWR VGND sg13g2_fill_2
XFILLER_20_191 VPWR VGND sg13g2_fill_2
XFILLER_5_825 VPWR VGND sg13g2_decap_8
XFILLER_4_313 VPWR VGND sg13g2_decap_8
XFILLER_4_302 VPWR VGND sg13g2_fill_2
XFILLER_4_346 VPWR VGND sg13g2_decap_4
XFILLER_0_541 VPWR VGND sg13g2_decap_8
XFILLER_17_910 VPWR VGND sg13g2_decap_8
XFILLER_35_228 VPWR VGND sg13g2_decap_4
XFILLER_16_420 VPWR VGND sg13g2_decap_4
XFILLER_16_453 VPWR VGND sg13g2_fill_2
XFILLER_17_987 VPWR VGND sg13g2_decap_8
XFILLER_44_795 VPWR VGND sg13g2_decap_8
XFILLER_32_968 VPWR VGND sg13g2_decap_8
XFILLER_40_990 VPWR VGND sg13g2_decap_8
X_2770_ net414 VPWR _1064_ VGND net471 ppwm_i.u_ppwm.u_mem.memory\[110\] sg13g2_o21ai_1
XFILLER_8_674 VPWR VGND sg13g2_decap_8
XFILLER_11_180 VPWR VGND sg13g2_decap_4
X_1721_ VPWR VGND _1287_ _1231_ _1286_ _1284_ _1288_ _1285_ sg13g2_a221oi_1
X_1652_ _1223_ net504 VPWR VGND sg13g2_inv_2
XFILLER_8_696 VPWR VGND sg13g2_fill_1
Xhold107 sdr_i.mac1.products_ff\[85\] VPWR VGND net307 sg13g2_dlygate4sd3_1
Xhold129 _0167_ VPWR VGND net329 sg13g2_dlygate4sd3_1
Xhold118 _0372_ VPWR VGND net318 sg13g2_dlygate4sd3_1
X_1583_ VPWR _1154_ ppwm_i.u_ppwm.u_mem.memory\[55\] VGND sg13g2_inv_1
X_3184_ net524 VGND VPWR net205 sdr_i.mac1.sum_lvl3_ff\[3\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2204_ _0629_ VPWR _0630_ VGND _0626_ _0628_ sg13g2_o21ai_1
X_2135_ _0561_ ppwm_i.u_ppwm.global_counter\[14\] _1225_ ppwm_i.u_ppwm.global_counter\[15\]
+ _1224_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
XFILLER_19_291 VPWR VGND sg13g2_decap_8
X_2066_ _0502_ _0503_ _0181_ VPWR VGND sg13g2_nor2_1
XFILLER_23_957 VPWR VGND sg13g2_decap_8
XFILLER_34_272 VPWR VGND sg13g2_decap_8
X_2968_ net435 VGND VPWR _0159_ ppwm_i.u_ppwm.global_counter\[11\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
X_1919_ net297 sdr_i.mac2.sum_lvl2_ff\[4\] _0009_ VPWR VGND sg13g2_xor2_1
X_2899_ net528 VGND VPWR _0090_ sdr_i.DP_1.matrix\[63\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_45_548 VPWR VGND sg13g2_fill_2
XFILLER_27_87 VPWR VGND sg13g2_decap_4
XFILLER_26_751 VPWR VGND sg13g2_fill_1
XFILLER_13_412 VPWR VGND sg13g2_decap_8
XFILLER_14_935 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
X_3106__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_13_445 VPWR VGND sg13g2_fill_2
XFILLER_43_97 VPWR VGND sg13g2_fill_2
XFILLER_41_787 VPWR VGND sg13g2_decap_8
XFILLER_13_478 VPWR VGND sg13g2_fill_1
XFILLER_40_297 VPWR VGND sg13g2_decap_4
X_3002__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_4_121 VPWR VGND sg13g2_decap_8
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
XFILLER_36_548 VPWR VGND sg13g2_fill_1
XFILLER_44_581 VPWR VGND sg13g2_decap_8
XFILLER_20_905 VPWR VGND sg13g2_decap_8
X_2822_ net263 _0085_ VPWR VGND sg13g2_buf_1
XFILLER_13_990 VPWR VGND sg13g2_decap_8
XFILLER_31_275 VPWR VGND sg13g2_decap_8
XFILLER_9_961 VPWR VGND sg13g2_decap_8
X_2753_ VGND VPWR net474 _1107_ _0316_ _1055_ sg13g2_a21oi_1
XFILLER_31_297 VPWR VGND sg13g2_decap_8
X_1704_ net421 _1271_ net471 _1273_ VPWR VGND sg13g2_nand3_1
X_2684_ net412 VPWR _1021_ VGND net465 ppwm_i.u_ppwm.u_mem.memory\[67\] sg13g2_o21ai_1
XFILLER_8_493 VPWR VGND sg13g2_fill_2
X_1635_ VPWR _1206_ net342 VGND sg13g2_inv_1
X_1566_ VPWR _1137_ net559 VGND sg13g2_inv_1
Xfanout417 net418 net417 VPWR VGND sg13g2_buf_8
Xfanout428 net434 net428 VPWR VGND sg13g2_buf_8
Xfanout439 _1283_ net439 VPWR VGND sg13g2_buf_8
Xfanout406 _1352_ net406 VPWR VGND sg13g2_buf_1
XFILLER_39_320 VPWR VGND sg13g2_fill_2
X_3167_ net531 VGND VPWR net742 sdr_i.mac1.sum_lvl1_ff\[17\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_27_504 VPWR VGND sg13g2_decap_8
X_3098_ net47 VGND VPWR net608 ppwm_i.u_ppwm.u_mem.memory\[74\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3102__31 VPWR VGND net31 sg13g2_tiehi
X_2118_ net768 _0544_ _0545_ VPWR VGND sg13g2_and2_1
X_2049_ net455 _0491_ _0492_ _0175_ VPWR VGND sg13g2_nor3_1
XFILLER_11_916 VPWR VGND sg13g2_decap_8
XFILLER_23_765 VPWR VGND sg13g2_decap_8
XFILLER_13_45 VPWR VGND sg13g2_decap_8
XFILLER_2_603 VPWR VGND sg13g2_decap_8
Xhold460 _1094_ VPWR VGND net840 sg13g2_dlygate4sd3_1
XFILLER_1_135 VPWR VGND sg13g2_decap_8
XFILLER_49_117 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_46_857 VPWR VGND sg13g2_decap_8
XFILLER_14_732 VPWR VGND sg13g2_decap_4
XFILLER_41_540 VPWR VGND sg13g2_fill_2
XFILLER_14_798 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_10_993 VPWR VGND sg13g2_decap_8
XFILLER_6_975 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_fill_1
XFILLER_49_684 VPWR VGND sg13g2_decap_8
X_3021_ net107 VGND VPWR _0212_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
XFILLER_37_802 VPWR VGND sg13g2_decap_8
XFILLER_49_695 VPWR VGND sg13g2_fill_2
XFILLER_37_879 VPWR VGND sg13g2_decap_8
XFILLER_17_592 VPWR VGND sg13g2_decap_8
XFILLER_32_562 VPWR VGND sg13g2_fill_2
X_2805_ _1090_ ppwm_i.u_ppwm.u_pwm.counter\[7\] ppwm_i.u_ppwm.u_pwm.cmp_value\[7\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_20_735 VPWR VGND sg13g2_decap_8
XFILLER_32_595 VPWR VGND sg13g2_decap_4
XFILLER_20_779 VPWR VGND sg13g2_decap_8
X_2736_ net417 VPWR _1047_ VGND net479 ppwm_i.u_ppwm.u_mem.memory\[93\] sg13g2_o21ai_1
X_2667_ VGND VPWR net479 _1150_ _0273_ _1012_ sg13g2_a21oi_1
X_1618_ VPWR _1189_ net623 VGND sg13g2_inv_1
X_2598_ net431 VPWR _0978_ VGND net497 ppwm_i.u_ppwm.u_mem.memory\[24\] sg13g2_o21ai_1
X_1549_ VPWR _1120_ net687 VGND sg13g2_inv_1
XFILLER_28_813 VPWR VGND sg13g2_decap_8
X_3219_ net544 VGND VPWR net724 sdr_i.mac2.sum_lvl2_ff\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_43_838 VPWR VGND sg13g2_decap_8
XFILLER_23_540 VPWR VGND sg13g2_fill_1
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_267 VPWR VGND sg13g2_decap_8
XFILLER_11_768 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_fill_2
XFILLER_40_87 VPWR VGND sg13g2_decap_8
XFILLER_40_65 VPWR VGND sg13g2_decap_8
XFILLER_3_945 VPWR VGND sg13g2_decap_8
XFILLER_2_411 VPWR VGND sg13g2_decap_8
XFILLER_46_1011 VPWR VGND sg13g2_decap_8
Xhold290 _0269_ VPWR VGND net670 sg13g2_dlygate4sd3_1
XFILLER_49_96 VPWR VGND sg13g2_decap_8
XFILLER_18_334 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_34_805 VPWR VGND sg13g2_decap_8
XFILLER_42_860 VPWR VGND sg13g2_decap_8
X_3093__66 VPWR VGND net66 sg13g2_tiehi
X_2521_ VPWR _0928_ _0927_ VGND sg13g2_inv_1
XFILLER_6_761 VPWR VGND sg13g2_decap_4
X_2452_ net374 _0865_ _0866_ VPWR VGND sg13g2_and2_1
X_2383_ net377 VPWR _0801_ VGND _0796_ _0800_ sg13g2_o21ai_1
Xinput3 ui_in[0] net3 VPWR VGND sg13g2_buf_1
X_3004_ net140 VGND VPWR net801 ppwm_i.u_ppwm.pwm_value\[0\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_18_890 VPWR VGND sg13g2_decap_8
XFILLER_36_186 VPWR VGND sg13g2_fill_1
XFILLER_40_808 VPWR VGND sg13g2_decap_8
XFILLER_33_860 VPWR VGND sg13g2_decap_8
XFILLER_20_576 VPWR VGND sg13g2_fill_2
X_2719_ VGND VPWR net467 _1124_ _0299_ _1038_ sg13g2_a21oi_1
XFILLER_10_13 VPWR VGND sg13g2_decap_4
XFILLER_3_219 VPWR VGND sg13g2_decap_4
XFILLER_0_948 VPWR VGND sg13g2_decap_8
XFILLER_48_919 VPWR VGND sg13g2_decap_8
XFILLER_19_55 VPWR VGND sg13g2_decap_8
XFILLER_28_632 VPWR VGND sg13g2_fill_2
XFILLER_28_654 VPWR VGND sg13g2_fill_1
XFILLER_15_304 VPWR VGND sg13g2_fill_1
XFILLER_35_54 VPWR VGND sg13g2_decap_4
XFILLER_24_882 VPWR VGND sg13g2_decap_8
XFILLER_30_318 VPWR VGND sg13g2_fill_1
XFILLER_35_87 VPWR VGND sg13g2_decap_8
XFILLER_2_230 VPWR VGND sg13g2_decap_8
XFILLER_38_418 VPWR VGND sg13g2_decap_8
XFILLER_20_1003 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_34_613 VPWR VGND sg13g2_decap_8
XFILLER_34_624 VPWR VGND sg13g2_fill_2
X_2984__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_15_871 VPWR VGND sg13g2_decap_8
XFILLER_34_679 VPWR VGND sg13g2_decap_8
X_1952_ sdr_i.mac2.products_ff\[52\] sdr_i.mac2.products_ff\[35\] _0437_ VPWR VGND
+ sg13g2_xor2_1
XFILLER_14_370 VPWR VGND sg13g2_fill_2
X_1883_ _0406_ net734 net217 VPWR VGND sg13g2_nand2_1
XFILLER_30_874 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_2504_ _0912_ VPWR _0913_ VGND net382 _0791_ sg13g2_o21ai_1
X_2435_ _0849_ VPWR _0850_ VGND _0786_ _0848_ sg13g2_o21ai_1
X_2366_ _0784_ VPWR _0785_ VGND _1220_ net404 sg13g2_o21ai_1
XFILLER_29_407 VPWR VGND sg13g2_fill_1
X_2297_ VGND VPWR _0719_ _0718_ _0685_ sg13g2_or2_1
XFILLER_37_451 VPWR VGND sg13g2_decap_8
XFILLER_38_952 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_fill_2
XFILLER_25_646 VPWR VGND sg13g2_decap_8
XFILLER_25_679 VPWR VGND sg13g2_decap_8
XFILLER_36_1010 VPWR VGND sg13g2_decap_8
XFILLER_40_638 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XFILLER_20_351 VPWR VGND sg13g2_fill_1
XFILLER_21_863 VPWR VGND sg13g2_decap_8
XFILLER_0_745 VPWR VGND sg13g2_decap_8
XFILLER_48_716 VPWR VGND sg13g2_decap_8
XFILLER_47_215 VPWR VGND sg13g2_fill_2
XFILLER_29_941 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_16_602 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_fill_2
XFILLER_44_977 VPWR VGND sg13g2_decap_8
XFILLER_28_495 VPWR VGND sg13g2_decap_4
XFILLER_15_145 VPWR VGND sg13g2_decap_8
XFILLER_30_104 VPWR VGND sg13g2_fill_1
XFILLER_31_638 VPWR VGND sg13g2_fill_2
XFILLER_11_340 VPWR VGND sg13g2_fill_1
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_7_388 VPWR VGND sg13g2_decap_8
XFILLER_3_550 VPWR VGND sg13g2_decap_8
X_2220_ net396 VPWR _0646_ VGND net401 net389 sg13g2_o21ai_1
X_3012__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_39_705 VPWR VGND sg13g2_decap_4
XFILLER_39_749 VPWR VGND sg13g2_fill_1
XFILLER_39_738 VPWR VGND sg13g2_fill_1
X_2151_ _0577_ ppwm_i.u_ppwm.global_counter\[14\] _1215_ ppwm_i.u_ppwm.global_counter\[15\]
+ _1214_ VPWR VGND sg13g2_a22oi_1
X_2082_ _0514_ net752 _0513_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_462 VPWR VGND sg13g2_decap_8
X_3141__84 VPWR VGND net84 sg13g2_tiehi
XFILLER_35_955 VPWR VGND sg13g2_decap_8
XFILLER_34_454 VPWR VGND sg13g2_decap_4
X_2984_ net179 VGND VPWR net581 ppwm_i.u_ppwm.u_pwm.cmp_value\[7\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_1935_ net230 sdr_i.mac1.products_ff\[119\] _0021_ VPWR VGND sg13g2_xor2_1
XFILLER_21_148 VPWR VGND sg13g2_decap_8
X_1866_ _0400_ net315 net238 VPWR VGND sg13g2_nand2_1
X_1797_ VGND VPWR _1183_ net453 _0346_ net512 sg13g2_a21oi_1
X_2418_ _0834_ _0832_ _0830_ VPWR VGND sg13g2_nand2b_1
X_2349_ _0769_ _0768_ _0659_ _0725_ net379 VPWR VGND sg13g2_a22oi_1
XFILLER_25_443 VPWR VGND sg13g2_decap_4
XFILLER_26_955 VPWR VGND sg13g2_decap_8
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_5_804 VPWR VGND sg13g2_decap_8
XFILLER_4_369 VPWR VGND sg13g2_decap_4
XFILLER_0_520 VPWR VGND sg13g2_decap_8
XFILLER_0_597 VPWR VGND sg13g2_decap_8
XFILLER_17_966 VPWR VGND sg13g2_decap_8
XFILLER_44_774 VPWR VGND sg13g2_decap_8
XFILLER_43_251 VPWR VGND sg13g2_decap_8
XFILLER_43_262 VPWR VGND sg13g2_fill_1
XFILLER_16_487 VPWR VGND sg13g2_decap_8
XFILLER_32_947 VPWR VGND sg13g2_decap_8
XFILLER_31_479 VPWR VGND sg13g2_decap_4
X_1720_ VPWR VGND _1150_ net510 net447 _1129_ _1287_ net451 sg13g2_a221oi_1
X_1651_ _1222_ net503 VPWR VGND sg13g2_inv_2
Xhold108 _0019_ VPWR VGND net308 sg13g2_dlygate4sd3_1
Xhold119 _0001_ VPWR VGND net319 sg13g2_dlygate4sd3_1
X_1582_ _1153_ net673 VPWR VGND sg13g2_inv_2
XFILLER_4_881 VPWR VGND sg13g2_decap_8
XFILLER_3_380 VPWR VGND sg13g2_decap_8
XFILLER_39_524 VPWR VGND sg13g2_decap_8
X_3183_ net526 VGND VPWR net210 sdr_i.mac1.sum_lvl3_ff\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2203_ _0629_ net506 _1216_ ppwm_i.u_ppwm.pwm_value\[4\] _1215_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_546 VPWR VGND sg13g2_decap_4
X_2134_ _0558_ VPWR _0560_ VGND _0553_ _0559_ sg13g2_o21ai_1
XFILLER_26_218 VPWR VGND sg13g2_decap_8
X_2065_ net422 VPWR _0503_ VGND net786 _0500_ sg13g2_o21ai_1
XFILLER_23_936 VPWR VGND sg13g2_decap_8
XFILLER_34_284 VPWR VGND sg13g2_decap_8
XFILLER_22_479 VPWR VGND sg13g2_decap_8
X_2967_ net435 VGND VPWR net558 ppwm_i.u_ppwm.global_counter\[10\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
X_2898_ net529 VGND VPWR _0089_ sdr_i.DP_1.matrix\[55\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_1918_ _0420_ net764 net297 VPWR VGND sg13g2_nand2_1
X_1849_ _0389_ net288 net247 VPWR VGND sg13g2_nand2_1
X_3050__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_27_33 VPWR VGND sg13g2_fill_1
XFILLER_14_914 VPWR VGND sg13g2_decap_8
XFILLER_41_733 VPWR VGND sg13g2_fill_2
XFILLER_41_766 VPWR VGND sg13g2_decap_8
XFILLER_40_243 VPWR VGND sg13g2_fill_2
XFILLER_13_435 VPWR VGND sg13g2_fill_2
XFILLER_13_457 VPWR VGND sg13g2_decap_8
XFILLER_43_76 VPWR VGND sg13g2_decap_8
XFILLER_40_265 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_3_3__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_612 VPWR VGND sg13g2_fill_2
XFILLER_4_155 VPWR VGND sg13g2_fill_2
XFILLER_4_15 VPWR VGND sg13g2_decap_8
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_36_527 VPWR VGND sg13g2_fill_2
XFILLER_16_284 VPWR VGND sg13g2_decap_4
XFILLER_17_1008 VPWR VGND sg13g2_decap_8
X_2821_ net295 _0084_ VPWR VGND sg13g2_buf_1
XFILLER_9_940 VPWR VGND sg13g2_decap_8
X_2752_ net419 VPWR _1055_ VGND net474 ppwm_i.u_ppwm.u_mem.memory\[101\] sg13g2_o21ai_1
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_1703_ _1272_ net471 net421 VPWR VGND sg13g2_nand2_1
X_2683_ VGND VPWR net466 _1142_ _0281_ _1020_ sg13g2_a21oi_1
X_1634_ VPWR _1205_ net656 VGND sg13g2_inv_1
X_1565_ VPWR _1136_ net704 VGND sg13g2_inv_1
Xfanout418 net420 net418 VPWR VGND sg13g2_buf_8
Xfanout429 net430 net429 VPWR VGND sg13g2_buf_1
Xfanout407 net408 net407 VPWR VGND sg13g2_buf_8
X_3166_ net531 VGND VPWR net308 sdr_i.mac1.sum_lvl1_ff\[16\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_39_387 VPWR VGND sg13g2_fill_2
X_3097_ net51 VGND VPWR net631 ppwm_i.u_ppwm.u_mem.memory\[73\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_2117_ _0518_ VPWR _0544_ VGND _1277_ _0543_ sg13g2_o21ai_1
X_2048_ net580 net411 _0492_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_733 VPWR VGND sg13g2_fill_2
XFILLER_35_593 VPWR VGND sg13g2_fill_2
XFILLER_22_243 VPWR VGND sg13g2_fill_1
XFILLER_10_416 VPWR VGND sg13g2_fill_1
XFILLER_13_13 VPWR VGND sg13g2_decap_8
XFILLER_22_287 VPWR VGND sg13g2_decap_8
XFILLER_13_79 VPWR VGND sg13g2_decap_8
Xhold461 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] VPWR VGND net841 sg13g2_dlygate4sd3_1
Xhold450 ppwm_i.u_ppwm.pwm_value\[6\] VPWR VGND net830 sg13g2_dlygate4sd3_1
X_3071__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_18_505 VPWR VGND sg13g2_decap_8
XFILLER_46_836 VPWR VGND sg13g2_decap_8
XFILLER_14_700 VPWR VGND sg13g2_decap_4
XFILLER_26_571 VPWR VGND sg13g2_fill_2
XFILLER_13_243 VPWR VGND sg13g2_decap_8
XFILLER_41_563 VPWR VGND sg13g2_decap_8
XFILLER_10_972 VPWR VGND sg13g2_decap_8
XFILLER_6_954 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_fill_1
XFILLER_49_663 VPWR VGND sg13g2_decap_8
X_3020_ net109 VGND VPWR net837 ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_48_173 VPWR VGND sg13g2_fill_2
XFILLER_36_335 VPWR VGND sg13g2_decap_8
XFILLER_37_858 VPWR VGND sg13g2_decap_8
XFILLER_45_891 VPWR VGND sg13g2_decap_8
XFILLER_20_714 VPWR VGND sg13g2_decap_8
X_2804_ VPWR VGND _1239_ _1088_ ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] _1238_ _1089_ ppwm_i.u_ppwm.u_pwm.cmp_value\[6\]
+ sg13g2_a221oi_1
X_2735_ VGND VPWR net478 _1116_ _0307_ _1046_ sg13g2_a21oi_1
X_2994__159 VPWR VGND net159 sg13g2_tiehi
X_2666_ net417 VPWR _1012_ VGND net479 net563 sg13g2_o21ai_1
X_1617_ VPWR _1188_ net733 VGND sg13g2_inv_1
X_2597_ VGND VPWR net489 _1185_ _0238_ _0977_ sg13g2_a21oi_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_1548_ VPWR _1119_ net614 VGND sg13g2_inv_1
XFILLER_27_302 VPWR VGND sg13g2_decap_8
X_3218_ net536 VGND VPWR net270 sdr_i.mac2.sum_lvl2_ff\[4\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3149_ net526 VGND VPWR _0041_ sdr_i.mac1.products_ff\[35\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_27_313 VPWR VGND sg13g2_fill_1
XFILLER_43_817 VPWR VGND sg13g2_decap_8
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_42_327 VPWR VGND sg13g2_fill_1
XFILLER_42_316 VPWR VGND sg13g2_fill_2
XFILLER_36_891 VPWR VGND sg13g2_decap_8
XFILLER_24_34 VPWR VGND sg13g2_fill_1
XFILLER_10_246 VPWR VGND sg13g2_decap_8
XFILLER_6_217 VPWR VGND sg13g2_decap_8
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_3_924 VPWR VGND sg13g2_decap_8
Xhold280 ppwm_i.u_ppwm.u_mem.memory\[62\] VPWR VGND net660 sg13g2_dlygate4sd3_1
Xhold291 ppwm_i.u_ppwm.u_mem.memory\[67\] VPWR VGND net671 sg13g2_dlygate4sd3_1
XFILLER_46_600 VPWR VGND sg13g2_decap_4
XFILLER_46_611 VPWR VGND sg13g2_fill_1
XFILLER_45_165 VPWR VGND sg13g2_decap_8
XFILLER_27_891 VPWR VGND sg13g2_decap_8
XFILLER_33_327 VPWR VGND sg13g2_decap_8
X_2520_ _0927_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] net393 VPWR VGND sg13g2_xnor2_1
XFILLER_6_795 VPWR VGND sg13g2_decap_4
X_2451_ VPWR VGND net377 _0675_ _0864_ net380 _0865_ _0858_ sg13g2_a221oi_1
X_2382_ _0799_ _0758_ _0798_ _0800_ VPWR VGND sg13g2_a21o_1
X_3003_ net142 VGND VPWR net713 ppwm_i.u_ppwm.polarity clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_36_143 VPWR VGND sg13g2_fill_2
XFILLER_37_666 VPWR VGND sg13g2_decap_8
XFILLER_24_305 VPWR VGND sg13g2_fill_2
XFILLER_24_349 VPWR VGND sg13g2_fill_1
XFILLER_20_544 VPWR VGND sg13g2_fill_1
X_2718_ net412 VPWR _1038_ VGND net466 ppwm_i.u_ppwm.u_mem.memory\[84\] sg13g2_o21ai_1
XFILLER_3_209 VPWR VGND sg13g2_fill_1
XFILLER_10_47 VPWR VGND sg13g2_fill_1
X_2649_ VGND VPWR net491 _1159_ _0264_ _1003_ sg13g2_a21oi_1
XFILLER_0_927 VPWR VGND sg13g2_decap_8
XFILLER_15_327 VPWR VGND sg13g2_decap_8
XFILLER_27_165 VPWR VGND sg13g2_decap_8
XFILLER_43_636 VPWR VGND sg13g2_decap_8
XFILLER_42_113 VPWR VGND sg13g2_decap_4
XFILLER_24_861 VPWR VGND sg13g2_decap_8
XFILLER_13_1011 VPWR VGND sg13g2_decap_8
XFILLER_7_559 VPWR VGND sg13g2_fill_2
XFILLER_3_710 VPWR VGND sg13g2_fill_2
XFILLER_3_754 VPWR VGND sg13g2_decap_4
XFILLER_3_798 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_18_8 VPWR VGND sg13g2_fill_1
XFILLER_46_485 VPWR VGND sg13g2_decap_8
XFILLER_18_154 VPWR VGND sg13g2_decap_8
XFILLER_18_165 VPWR VGND sg13g2_fill_1
XFILLER_18_198 VPWR VGND sg13g2_fill_1
XFILLER_22_809 VPWR VGND sg13g2_fill_1
XFILLER_34_636 VPWR VGND sg13g2_fill_1
XFILLER_15_850 VPWR VGND sg13g2_decap_8
XFILLER_15_861 VPWR VGND sg13g2_fill_1
X_3125__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_33_157 VPWR VGND sg13g2_decap_8
XFILLER_42_691 VPWR VGND sg13g2_fill_1
X_1951_ net213 sdr_i.mac2.products_ff\[34\] _0034_ VPWR VGND sg13g2_xor2_1
X_1882_ net289 net286 _0052_ VPWR VGND sg13g2_and2_1
XFILLER_30_853 VPWR VGND sg13g2_decap_8
X_2503_ VGND VPWR _1224_ net382 _0912_ _0672_ sg13g2_a21oi_1
X_2434_ _0849_ _0746_ _0763_ VPWR VGND sg13g2_nand2_1
X_2365_ _0784_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] net404 VPWR VGND sg13g2_nand2_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_2296_ _0718_ _0713_ _0717_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_931 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_25_625 VPWR VGND sg13g2_decap_8
XFILLER_37_485 VPWR VGND sg13g2_decap_8
XFILLER_25_658 VPWR VGND sg13g2_decap_8
XFILLER_40_617 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_fill_1
XFILLER_21_13 VPWR VGND sg13g2_decap_4
XFILLER_0_724 VPWR VGND sg13g2_decap_8
XFILLER_29_920 VPWR VGND sg13g2_decap_8
XFILLER_47_249 VPWR VGND sg13g2_decap_8
XFILLER_46_32 VPWR VGND sg13g2_fill_2
XFILLER_46_21 VPWR VGND sg13g2_fill_2
XFILLER_46_65 VPWR VGND sg13g2_fill_1
XFILLER_28_474 VPWR VGND sg13g2_decap_8
XFILLER_29_997 VPWR VGND sg13g2_decap_8
XFILLER_44_956 VPWR VGND sg13g2_decap_8
XFILLER_15_124 VPWR VGND sg13g2_decap_8
XFILLER_16_647 VPWR VGND sg13g2_fill_1
X_2983__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_8_846 VPWR VGND sg13g2_decap_8
X_2150_ _0575_ VPWR _0576_ VGND _1215_ ppwm_i.u_ppwm.global_counter\[14\] sg13g2_o21ai_1
XFILLER_38_227 VPWR VGND sg13g2_decap_8
X_2081_ net455 net767 _0513_ _0186_ VPWR VGND sg13g2_nor3_1
XFILLER_34_433 VPWR VGND sg13g2_decap_8
XFILLER_35_934 VPWR VGND sg13g2_decap_8
X_2983_ net180 VGND VPWR net665 ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
XFILLER_22_628 VPWR VGND sg13g2_decap_8
X_1934_ _0428_ sdr_i.mac1.products_ff\[119\] net230 VPWR VGND sg13g2_nand2_1
X_1865_ _0399_ _0398_ _0069_ VPWR VGND sg13g2_xor2_1
X_1796_ VPWR VGND _1190_ _0344_ net441 _1197_ _0345_ net445 sg13g2_a221oi_1
X_2417_ _0833_ _0830_ _0832_ VPWR VGND sg13g2_nand2b_1
X_2348_ VGND VPWR net384 _0744_ _0768_ _0767_ sg13g2_a21oi_1
X_2279_ _1228_ VPWR _0702_ VGND _0341_ _0347_ sg13g2_o21ai_1
X_3067__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_26_934 VPWR VGND sg13g2_decap_8
XFILLER_25_466 VPWR VGND sg13g2_fill_1
XFILLER_41_948 VPWR VGND sg13g2_decap_8
XFILLER_13_639 VPWR VGND sg13g2_fill_1
X_3045__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_20_193 VPWR VGND sg13g2_fill_1
XFILLER_4_304 VPWR VGND sg13g2_fill_1
XFILLER_10_1014 VPWR VGND sg13g2_decap_8
X_3074__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_0_510 VPWR VGND sg13g2_decap_8
XFILLER_0_576 VPWR VGND sg13g2_decap_8
XFILLER_16_433 VPWR VGND sg13g2_fill_1
XFILLER_17_945 VPWR VGND sg13g2_decap_8
XFILLER_29_794 VPWR VGND sg13g2_decap_8
XFILLER_16_455 VPWR VGND sg13g2_fill_1
XFILLER_32_926 VPWR VGND sg13g2_decap_8
XFILLER_8_643 VPWR VGND sg13g2_fill_2
X_1650_ _1221_ ppwm_i.u_ppwm.pwm_value\[8\] VPWR VGND sg13g2_inv_2
X_1581_ VPWR _1152_ net632 VGND sg13g2_inv_1
Xhold109 sdr_i.DP_3.matrix\[45\] VPWR VGND net309 sg13g2_dlygate4sd3_1
XFILLER_4_860 VPWR VGND sg13g2_decap_8
XFILLER_3_392 VPWR VGND sg13g2_fill_1
X_3182_ net533 VGND VPWR net745 sdr_i.mac1.sum_lvl3_ff\[1\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_2202_ _0628_ _0625_ _0627_ ppwm_i.u_ppwm.pwm_value\[2\] _1217_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_2 VPWR VGND sg13g2_fill_1
X_2133_ VPWR VGND ppwm_i.u_ppwm.pwm_value\[2\] _0557_ _1257_ net506 _0559_ _1256_
+ sg13g2_a221oi_1
XFILLER_35_742 VPWR VGND sg13g2_decap_8
X_2064_ net786 _0500_ _0502_ VPWR VGND sg13g2_and2_1
XFILLER_23_915 VPWR VGND sg13g2_decap_8
XFILLER_22_458 VPWR VGND sg13g2_decap_8
X_2966_ net437 VGND VPWR net336 ppwm_i.u_ppwm.global_counter\[9\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
X_2897_ net528 VGND VPWR _0088_ sdr_i.DP_1.matrix\[54\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_1917_ _0008_ _0416_ _0419_ VPWR VGND sg13g2_xnor2_1
X_1848_ _0388_ net280 net223 VPWR VGND sg13g2_nand2_1
X_1779_ VPWR VGND _1345_ net509 _1343_ _1340_ _1346_ _1342_ sg13g2_a221oi_1
XFILLER_40_1018 VPWR VGND sg13g2_decap_8
XFILLER_26_742 VPWR VGND sg13g2_decap_4
XFILLER_26_775 VPWR VGND sg13g2_fill_2
XFILLER_41_756 VPWR VGND sg13g2_fill_1
XFILLER_41_745 VPWR VGND sg13g2_decap_8
XFILLER_43_99 VPWR VGND sg13g2_fill_1
XFILLER_9_429 VPWR VGND sg13g2_decap_8
XFILLER_5_657 VPWR VGND sg13g2_decap_4
XFILLER_4_101 VPWR VGND sg13g2_fill_2
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_679 VPWR VGND sg13g2_fill_2
XFILLER_1_863 VPWR VGND sg13g2_decap_8
XFILLER_0_351 VPWR VGND sg13g2_decap_8
XFILLER_49_867 VPWR VGND sg13g2_decap_8
XFILLER_0_395 VPWR VGND sg13g2_decap_8
XFILLER_16_241 VPWR VGND sg13g2_decap_8
XFILLER_17_764 VPWR VGND sg13g2_decap_4
XFILLER_32_734 VPWR VGND sg13g2_decap_4
X_2820_ net235 _0083_ VPWR VGND sg13g2_buf_1
XFILLER_31_255 VPWR VGND sg13g2_decap_4
X_2751_ VGND VPWR net475 _1108_ _0315_ _1054_ sg13g2_a21oi_1
X_2682_ net418 VPWR _1020_ VGND net473 net659 sg13g2_o21ai_1
XFILLER_9_996 VPWR VGND sg13g2_decap_8
X_1702_ net748 _1269_ _1270_ _1271_ VPWR VGND sg13g2_nor3_1
X_1633_ VPWR _1204_ net684 VGND sg13g2_inv_1
X_1564_ VPWR _1135_ net630 VGND sg13g2_inv_1
Xfanout408 _1346_ net408 VPWR VGND sg13g2_buf_2
Xfanout419 net420 net419 VPWR VGND sg13g2_buf_8
XFILLER_39_300 VPWR VGND sg13g2_decap_8
XFILLER_39_344 VPWR VGND sg13g2_decap_4
X_3165_ net526 VGND VPWR net779 sdr_i.mac1.sum_lvl1_ff\[9\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_39_399 VPWR VGND sg13g2_decap_4
X_3096_ net54 VGND VPWR _0287_ ppwm_i.u_ppwm.u_mem.memory\[72\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_2116_ VGND VPWR net511 net451 _0543_ net508 sg13g2_a21oi_1
X_2047_ net503 net410 _0491_ VPWR VGND sg13g2_nor2_1
XFILLER_35_572 VPWR VGND sg13g2_decap_8
X_2949_ net542 VGND VPWR _0140_ sdr_i.DP_4.matrix\[45\] clknet_leaf_10_clk sg13g2_dfrbpq_1
Xhold440 ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] VPWR VGND net820 sg13g2_dlygate4sd3_1
Xhold451 ppwm_i.u_ppwm.pwm_value\[1\] VPWR VGND net831 sg13g2_dlygate4sd3_1
XFILLER_46_815 VPWR VGND sg13g2_decap_8
XFILLER_18_539 VPWR VGND sg13g2_decap_8
XFILLER_41_542 VPWR VGND sg13g2_fill_1
XFILLER_14_767 VPWR VGND sg13g2_decap_4
XFILLER_41_597 VPWR VGND sg13g2_fill_2
XFILLER_10_951 VPWR VGND sg13g2_decap_8
XFILLER_6_933 VPWR VGND sg13g2_decap_8
XFILLER_5_432 VPWR VGND sg13g2_fill_1
XFILLER_5_476 VPWR VGND sg13g2_decap_4
XFILLER_49_642 VPWR VGND sg13g2_decap_8
XFILLER_0_170 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_837 VPWR VGND sg13g2_decap_8
X_3096__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_36_358 VPWR VGND sg13g2_fill_1
XFILLER_45_870 VPWR VGND sg13g2_decap_8
XFILLER_20_704 VPWR VGND sg13g2_fill_1
XFILLER_32_564 VPWR VGND sg13g2_fill_1
X_2803_ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[4\] _1087_ _1244_ net520 _1088_ _1243_
+ sg13g2_a221oi_1
XFILLER_9_771 VPWR VGND sg13g2_decap_8
X_2734_ net416 VPWR _1046_ VGND net478 net568 sg13g2_o21ai_1
XFILLER_9_793 VPWR VGND sg13g2_fill_1
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_2665_ VGND VPWR net485 _1151_ _0272_ _1011_ sg13g2_a21oi_1
X_1616_ VPWR _1187_ net621 VGND sg13g2_inv_1
X_2596_ net431 VPWR _0977_ VGND net490 ppwm_i.u_ppwm.u_mem.memory\[23\] sg13g2_o21ai_1
X_1547_ VPWR _1118_ net727 VGND sg13g2_inv_1
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
X_3217_ net544 VGND VPWR net732 sdr_i.mac2.sum_lvl2_ff\[1\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3148_ net526 VGND VPWR _0040_ sdr_i.mac1.products_ff\[34\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_39_196 VPWR VGND sg13g2_decap_8
X_3079_ net121 VGND VPWR net674 ppwm_i.u_ppwm.u_mem.memory\[55\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_2
XFILLER_36_870 VPWR VGND sg13g2_decap_8
XFILLER_42_339 VPWR VGND sg13g2_fill_1
XFILLER_23_531 VPWR VGND sg13g2_decap_8
XFILLER_23_575 VPWR VGND sg13g2_fill_2
XFILLER_11_726 VPWR VGND sg13g2_fill_2
XFILLER_23_597 VPWR VGND sg13g2_decap_8
XFILLER_3_903 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_4
Xhold270 ppwm_i.u_ppwm.u_mem.memory\[63\] VPWR VGND net650 sg13g2_dlygate4sd3_1
Xhold292 ppwm_i.u_ppwm.u_mem.memory\[93\] VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold281 ppwm_i.u_ppwm.u_mem.bit_count\[3\] VPWR VGND net661 sg13g2_dlygate4sd3_1
XFILLER_19_848 VPWR VGND sg13g2_fill_2
XFILLER_45_144 VPWR VGND sg13g2_decap_8
XFILLER_46_689 VPWR VGND sg13g2_decap_8
XFILLER_18_369 VPWR VGND sg13g2_decap_8
XFILLER_27_870 VPWR VGND sg13g2_decap_8
XFILLER_42_895 VPWR VGND sg13g2_decap_8
XFILLER_41_383 VPWR VGND sg13g2_decap_4
X_2450_ _0864_ _1219_ net397 VPWR VGND sg13g2_xnor2_1
XFILLER_46_5 VPWR VGND sg13g2_decap_8
X_2381_ _0755_ _0778_ _0799_ VPWR VGND sg13g2_and2_1
XFILLER_2_991 VPWR VGND sg13g2_decap_8
XFILLER_49_450 VPWR VGND sg13g2_decap_8
X_3002_ net144 VGND VPWR net351 ppwm_i.u_ppwm.u_ex.cmp_flag_q clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_37_612 VPWR VGND sg13g2_fill_2
XFILLER_25_829 VPWR VGND sg13g2_fill_2
XFILLER_36_177 VPWR VGND sg13g2_decap_8
X_3022__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_33_895 VPWR VGND sg13g2_decap_8
XFILLER_20_556 VPWR VGND sg13g2_fill_2
X_2717_ VGND VPWR net463 _1125_ _0298_ _1037_ sg13g2_a21oi_1
X_2648_ net428 VPWR _1003_ VGND net492 net638 sg13g2_o21ai_1
XFILLER_0_906 VPWR VGND sg13g2_decap_8
X_2579_ VGND VPWR net495 _1194_ _0229_ _0968_ sg13g2_a21oi_1
XFILLER_27_100 VPWR VGND sg13g2_fill_2
XFILLER_43_615 VPWR VGND sg13g2_decap_8
XFILLER_35_34 VPWR VGND sg13g2_decap_8
XFILLER_24_840 VPWR VGND sg13g2_decap_8
XFILLER_23_350 VPWR VGND sg13g2_decap_8
XFILLER_30_309 VPWR VGND sg13g2_decap_4
XFILLER_7_538 VPWR VGND sg13g2_decap_8
XFILLER_3_777 VPWR VGND sg13g2_decap_8
XFILLER_2_265 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_46_453 VPWR VGND sg13g2_decap_8
XFILLER_19_689 VPWR VGND sg13g2_fill_2
XFILLER_18_188 VPWR VGND sg13g2_fill_1
XFILLER_33_136 VPWR VGND sg13g2_decap_8
XFILLER_34_659 VPWR VGND sg13g2_decap_8
X_1950_ _0436_ net729 net213 VPWR VGND sg13g2_nand2_1
XFILLER_14_372 VPWR VGND sg13g2_fill_1
XFILLER_30_832 VPWR VGND sg13g2_decap_8
X_1881_ net303 net310 _0050_ VPWR VGND sg13g2_and2_1
XFILLER_14_394 VPWR VGND sg13g2_decap_8
X_2502_ _0909_ _0910_ net378 _0911_ VPWR VGND sg13g2_nand3_1
X_2433_ _0764_ VPWR _0848_ VGND net384 _0697_ sg13g2_o21ai_1
X_2364_ VPWR VGND _0655_ _0692_ _0739_ _0350_ _0783_ _0661_ sg13g2_a221oi_1
X_2295_ _0714_ _0716_ _0717_ VPWR VGND sg13g2_and2_1
XFILLER_38_910 VPWR VGND sg13g2_decap_8
XFILLER_37_420 VPWR VGND sg13g2_decap_8
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_33_670 VPWR VGND sg13g2_fill_2
XFILLER_21_843 VPWR VGND sg13g2_fill_2
XFILLER_21_898 VPWR VGND sg13g2_decap_8
XFILLER_0_703 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_217 VPWR VGND sg13g2_fill_1
XFILLER_29_976 VPWR VGND sg13g2_decap_8
XFILLER_44_935 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_fill_1
XFILLER_43_445 VPWR VGND sg13g2_fill_1
XFILLER_31_618 VPWR VGND sg13g2_decap_8
XFILLER_7_302 VPWR VGND sg13g2_fill_2
XFILLER_12_898 VPWR VGND sg13g2_decap_8
XFILLER_7_368 VPWR VGND sg13g2_decap_4
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_38_206 VPWR VGND sg13g2_decap_8
X_2080_ net766 _0511_ _0513_ VPWR VGND sg13g2_and2_1
XFILLER_4_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_46_250 VPWR VGND sg13g2_decap_4
XFILLER_35_913 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_decap_8
XFILLER_34_412 VPWR VGND sg13g2_decap_8
X_2982_ net182 VGND VPWR _0173_ ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
XFILLER_21_117 VPWR VGND sg13g2_fill_2
XFILLER_34_478 VPWR VGND sg13g2_decap_8
XFILLER_34_489 VPWR VGND sg13g2_fill_2
X_1933_ _0020_ _0426_ _0427_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_191 VPWR VGND sg13g2_fill_1
X_1864_ _0399_ net271 net253 VPWR VGND sg13g2_nand2_1
X_1795_ ppwm_i.u_ppwm.u_mem.memory\[5\] net516 net519 _0344_ VPWR VGND sg13g2_nor3_1
X_2416_ _0832_ ppwm_i.u_ppwm.pwm_value\[8\] net391 VPWR VGND sg13g2_xnor2_1
X_2347_ net384 _0766_ _0767_ VPWR VGND sg13g2_nor2_1
X_2278_ VPWR VGND net379 _0696_ _0700_ _0659_ _0701_ _0698_ sg13g2_a221oi_1
XFILLER_26_913 VPWR VGND sg13g2_decap_8
XFILLER_38_751 VPWR VGND sg13g2_fill_2
XFILLER_38_784 VPWR VGND sg13g2_decap_8
XFILLER_37_272 VPWR VGND sg13g2_decap_8
XFILLER_13_607 VPWR VGND sg13g2_decap_8
XFILLER_16_58 VPWR VGND sg13g2_decap_8
XFILLER_41_927 VPWR VGND sg13g2_decap_8
XFILLER_12_128 VPWR VGND sg13g2_decap_8
XFILLER_21_651 VPWR VGND sg13g2_decap_8
XFILLER_5_839 VPWR VGND sg13g2_decap_8
XFILLER_4_327 VPWR VGND sg13g2_decap_8
XFILLER_0_555 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_4
XFILLER_29_762 VPWR VGND sg13g2_fill_2
XFILLER_29_773 VPWR VGND sg13g2_decap_8
XFILLER_17_924 VPWR VGND sg13g2_decap_8
XFILLER_32_905 VPWR VGND sg13g2_decap_8
XFILLER_16_478 VPWR VGND sg13g2_decap_4
XFILLER_31_459 VPWR VGND sg13g2_decap_8
XFILLER_8_688 VPWR VGND sg13g2_fill_2
X_1580_ VPWR _1151_ net563 VGND sg13g2_inv_1
XFILLER_26_1011 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_fill_2
X_3181_ net526 VGND VPWR net306 sdr_i.mac1.sum_lvl3_ff\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2201_ _0627_ _1228_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _1227_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2132_ _0558_ net505 ppwm_i.u_ppwm.global_counter\[14\] VPWR VGND sg13g2_nand2b_1
X_2063_ _0500_ _0501_ _0180_ VPWR VGND sg13g2_nor2_1
XFILLER_34_220 VPWR VGND sg13g2_decap_8
XFILLER_35_787 VPWR VGND sg13g2_decap_8
XFILLER_16_990 VPWR VGND sg13g2_decap_8
X_2965_ net436 VGND VPWR _0156_ ppwm_i.u_ppwm.global_counter\[8\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_31_982 VPWR VGND sg13g2_decap_8
X_2896_ net531 VGND VPWR _0087_ sdr_i.DP_1.matrix\[46\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_1916_ net782 net601 _0419_ VPWR VGND sg13g2_xor2_1
XFILLER_30_470 VPWR VGND sg13g2_decap_8
XFILLER_30_492 VPWR VGND sg13g2_decap_4
XFILLER_8_92 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_4
X_1847_ _0387_ _0386_ _0055_ VPWR VGND sg13g2_xor2_1
XFILLER_2_809 VPWR VGND sg13g2_decap_8
X_1778_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[48\] _1344_ net440 ppwm_i.u_ppwm.u_mem.memory\[41\]
+ _1345_ net444 sg13g2_a221oi_1
XFILLER_45_518 VPWR VGND sg13g2_fill_2
XFILLER_27_13 VPWR VGND sg13g2_decap_8
X_3120__56 VPWR VGND net56 sg13g2_tiehi
XFILLER_41_713 VPWR VGND sg13g2_fill_2
XFILLER_41_702 VPWR VGND sg13g2_decap_8
XFILLER_14_949 VPWR VGND sg13g2_decap_8
XFILLER_25_253 VPWR VGND sg13g2_decap_8
XFILLER_25_275 VPWR VGND sg13g2_fill_2
XFILLER_41_735 VPWR VGND sg13g2_fill_1
XFILLER_40_223 VPWR VGND sg13g2_fill_2
XFILLER_40_212 VPWR VGND sg13g2_decap_8
XFILLER_13_437 VPWR VGND sg13g2_fill_1
XFILLER_25_297 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_fill_1
XFILLER_22_982 VPWR VGND sg13g2_decap_8
XFILLER_5_614 VPWR VGND sg13g2_fill_1
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
XFILLER_0_330 VPWR VGND sg13g2_decap_8
XFILLER_1_842 VPWR VGND sg13g2_decap_8
XFILLER_49_846 VPWR VGND sg13g2_decap_8
XFILLER_0_374 VPWR VGND sg13g2_decap_8
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_581 VPWR VGND sg13g2_decap_8
XFILLER_17_743 VPWR VGND sg13g2_fill_1
XFILLER_44_562 VPWR VGND sg13g2_decap_4
XFILLER_44_595 VPWR VGND sg13g2_decap_8
XFILLER_16_297 VPWR VGND sg13g2_decap_8
XFILLER_31_234 VPWR VGND sg13g2_decap_4
XFILLER_20_919 VPWR VGND sg13g2_decap_8
XFILLER_32_779 VPWR VGND sg13g2_decap_8
XFILLER_12_470 VPWR VGND sg13g2_decap_4
XFILLER_12_481 VPWR VGND sg13g2_fill_1
X_2750_ net419 VPWR _1054_ VGND net475 net362 sg13g2_o21ai_1
XFILLER_8_463 VPWR VGND sg13g2_decap_4
X_2681_ VGND VPWR net478 _1143_ _0280_ _1019_ sg13g2_a21oi_1
XFILLER_9_975 VPWR VGND sg13g2_decap_8
X_1701_ net716 net339 net661 _1270_ VPWR VGND net751 sg13g2_nand4_1
X_1632_ VPWR _1203_ net628 VGND sg13g2_inv_1
X_3032__85 VPWR VGND net85 sg13g2_tiehi
X_1563_ VPWR _1134_ net607 VGND sg13g2_inv_1
Xfanout409 net411 net409 VPWR VGND sg13g2_buf_8
X_3164_ net526 VGND VPWR net314 sdr_i.mac1.sum_lvl1_ff\[8\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_27_518 VPWR VGND sg13g2_decap_4
X_3095_ net58 VGND VPWR net560 ppwm_i.u_ppwm.u_mem.memory\[71\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_2115_ _0541_ VPWR _0542_ VGND _0539_ _0540_ sg13g2_o21ai_1
X_2046_ net456 _0489_ _0490_ _0174_ VPWR VGND sg13g2_nor3_1
XFILLER_35_551 VPWR VGND sg13g2_fill_1
XFILLER_22_223 VPWR VGND sg13g2_decap_8
XFILLER_10_407 VPWR VGND sg13g2_decap_8
X_2948_ net536 VGND VPWR _0139_ sdr_i.DP_4.matrix\[37\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2879_ net283 _0142_ VPWR VGND sg13g2_buf_1
Xhold430 _0213_ VPWR VGND net810 sg13g2_dlygate4sd3_1
XFILLER_2_617 VPWR VGND sg13g2_decap_8
XFILLER_2_628 VPWR VGND sg13g2_fill_2
XFILLER_2_639 VPWR VGND sg13g2_fill_1
Xhold452 _0196_ VPWR VGND net832 sg13g2_dlygate4sd3_1
Xhold441 ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] VPWR VGND net821 sg13g2_dlygate4sd3_1
XFILLER_38_34 VPWR VGND sg13g2_fill_2
XFILLER_45_326 VPWR VGND sg13g2_fill_2
XFILLER_45_315 VPWR VGND sg13g2_decap_4
XFILLER_39_890 VPWR VGND sg13g2_decap_8
XFILLER_26_573 VPWR VGND sg13g2_fill_1
XFILLER_14_746 VPWR VGND sg13g2_decap_8
XFILLER_41_576 VPWR VGND sg13g2_fill_2
XFILLER_9_216 VPWR VGND sg13g2_fill_2
XFILLER_9_249 VPWR VGND sg13g2_fill_2
XFILLER_10_930 VPWR VGND sg13g2_decap_8
XFILLER_13_278 VPWR VGND sg13g2_fill_2
XFILLER_6_912 VPWR VGND sg13g2_decap_8
XFILLER_6_989 VPWR VGND sg13g2_decap_8
XFILLER_49_621 VPWR VGND sg13g2_decap_8
XFILLER_37_816 VPWR VGND sg13g2_decap_8
XFILLER_36_304 VPWR VGND sg13g2_fill_1
X_2802_ VGND VPWR _1083_ _1084_ _1087_ _1086_ sg13g2_a21oi_1
XFILLER_20_749 VPWR VGND sg13g2_decap_8
X_2733_ VGND VPWR net473 _1117_ _0306_ _1045_ sg13g2_a21oi_1
XFILLER_30_1007 VPWR VGND sg13g2_decap_8
XFILLER_8_260 VPWR VGND sg13g2_decap_4
X_2664_ net426 VPWR _1011_ VGND net485 ppwm_i.u_ppwm.u_mem.memory\[57\] sg13g2_o21ai_1
X_1615_ VPWR _1186_ net617 VGND sg13g2_inv_1
X_2595_ VGND VPWR net495 _1186_ _0237_ _0976_ sg13g2_a21oi_1
X_1546_ VPWR _1117_ net568 VGND sg13g2_inv_1
XFILLER_5_71 VPWR VGND sg13g2_decap_8
X_3135__164 VPWR VGND net164 sg13g2_tiehi
X_3216_ net544 VGND VPWR net292 sdr_i.mac2.sum_lvl2_ff\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3147_ net523 VGND VPWR _0055_ sdr_i.mac1.products_ff\[18\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_28_827 VPWR VGND sg13g2_decap_8
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_42_318 VPWR VGND sg13g2_fill_1
X_3078_ net125 VGND VPWR net670 ppwm_i.u_ppwm.u_mem.memory\[54\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2029_ net507 net409 _0479_ VPWR VGND sg13g2_nor2_1
XFILLER_23_554 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_10_204 VPWR VGND sg13g2_fill_1
XFILLER_40_13 VPWR VGND sg13g2_decap_8
XFILLER_3_959 VPWR VGND sg13g2_decap_8
Xhold271 _0278_ VPWR VGND net651 sg13g2_dlygate4sd3_1
Xhold260 ppwm_i.u_ppwm.u_mem.memory\[94\] VPWR VGND net640 sg13g2_dlygate4sd3_1
XFILLER_49_33 VPWR VGND sg13g2_decap_8
XFILLER_46_1025 VPWR VGND sg13g2_decap_4
Xhold293 ppwm_i.u_ppwm.u_mem.memory\[56\] VPWR VGND net673 sg13g2_dlygate4sd3_1
Xhold282 _1074_ VPWR VGND net662 sg13g2_dlygate4sd3_1
XFILLER_19_805 VPWR VGND sg13g2_decap_8
XFILLER_46_624 VPWR VGND sg13g2_decap_4
XFILLER_18_326 VPWR VGND sg13g2_fill_2
XFILLER_46_646 VPWR VGND sg13g2_fill_2
XFILLER_18_348 VPWR VGND sg13g2_decap_8
XFILLER_33_307 VPWR VGND sg13g2_decap_8
XFILLER_34_819 VPWR VGND sg13g2_decap_8
XFILLER_14_521 VPWR VGND sg13g2_decap_4
XFILLER_26_370 VPWR VGND sg13g2_decap_8
XFILLER_26_381 VPWR VGND sg13g2_fill_1
XFILLER_42_874 VPWR VGND sg13g2_decap_8
XFILLER_14_543 VPWR VGND sg13g2_fill_2
X_2993__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_5_296 VPWR VGND sg13g2_fill_1
XFILLER_5_285 VPWR VGND sg13g2_decap_8
XFILLER_30_90 VPWR VGND sg13g2_decap_8
X_2380_ VGND VPWR _1224_ _1225_ _0798_ net392 sg13g2_a21oi_1
XFILLER_2_970 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
X_3001_ net146 VGND VPWR _0192_ ppwm_i.u_ppwm.pc\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_37_635 VPWR VGND sg13g2_decap_4
XFILLER_24_307 VPWR VGND sg13g2_fill_1
XFILLER_36_167 VPWR VGND sg13g2_fill_1
XFILLER_17_370 VPWR VGND sg13g2_decap_4
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_32_340 VPWR VGND sg13g2_fill_1
XFILLER_33_874 VPWR VGND sg13g2_decap_8
XFILLER_20_513 VPWR VGND sg13g2_decap_8
XFILLER_20_535 VPWR VGND sg13g2_decap_8
X_2716_ net413 VPWR _1037_ VGND net463 net678 sg13g2_o21ai_1
X_2647_ VGND VPWR net492 _1160_ _0263_ _1002_ sg13g2_a21oi_1
X_3139__37 VPWR VGND net37 sg13g2_tiehi
X_2578_ net432 VPWR _0968_ VGND net495 ppwm_i.u_ppwm.u_mem.memory\[14\] sg13g2_o21ai_1
X_1529_ VPWR _1100_ net627 VGND sg13g2_inv_1
XFILLER_19_69 VPWR VGND sg13g2_decap_8
XFILLER_28_602 VPWR VGND sg13g2_decap_8
XFILLER_28_613 VPWR VGND sg13g2_fill_2
XFILLER_35_13 VPWR VGND sg13g2_decap_4
XFILLER_36_690 VPWR VGND sg13g2_decap_4
XFILLER_11_513 VPWR VGND sg13g2_decap_4
XFILLER_11_524 VPWR VGND sg13g2_fill_2
XFILLER_23_373 VPWR VGND sg13g2_decap_8
XFILLER_23_384 VPWR VGND sg13g2_fill_2
XFILLER_24_896 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_712 VPWR VGND sg13g2_fill_1
XFILLER_3_745 VPWR VGND sg13g2_fill_1
XFILLER_2_244 VPWR VGND sg13g2_decap_8
XFILLER_2_299 VPWR VGND sg13g2_fill_1
XFILLER_19_624 VPWR VGND sg13g2_fill_1
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_18_101 VPWR VGND sg13g2_fill_2
XFILLER_18_112 VPWR VGND sg13g2_decap_8
XFILLER_19_646 VPWR VGND sg13g2_decap_8
XFILLER_20_1017 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_33_115 VPWR VGND sg13g2_decap_8
XFILLER_15_885 VPWR VGND sg13g2_decap_8
XFILLER_30_811 VPWR VGND sg13g2_decap_8
X_1880_ net279 net311 _0048_ VPWR VGND sg13g2_and2_1
XFILLER_14_384 VPWR VGND sg13g2_decap_4
XFILLER_30_888 VPWR VGND sg13g2_decap_8
X_2501_ _0895_ _0901_ _0908_ _0910_ VPWR VGND sg13g2_or3_1
X_2432_ _0845_ _0846_ net377 _0847_ VPWR VGND sg13g2_nand3_1
X_2363_ _0782_ _0763_ _0700_ VPWR VGND sg13g2_nand2b_1
X_2294_ ppwm_i.u_ppwm.pwm_value\[2\] VPWR _0716_ VGND net407 net405 sg13g2_o21ai_1
XFILLER_38_966 VPWR VGND sg13g2_decap_8
X_3057__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_33_682 VPWR VGND sg13g2_fill_1
XFILLER_36_1024 VPWR VGND sg13g2_decap_4
XFILLER_21_877 VPWR VGND sg13g2_decap_8
XFILLER_4_509 VPWR VGND sg13g2_decap_8
XFILLER_21_59 VPWR VGND sg13g2_decap_8
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_759 VPWR VGND sg13g2_decap_8
XFILLER_46_34 VPWR VGND sg13g2_fill_1
XFILLER_46_12 VPWR VGND sg13g2_fill_1
XFILLER_29_955 VPWR VGND sg13g2_decap_8
XFILLER_44_914 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_16_627 VPWR VGND sg13g2_fill_1
XFILLER_43_468 VPWR VGND sg13g2_decap_8
XFILLER_15_159 VPWR VGND sg13g2_decap_8
XFILLER_12_800 VPWR VGND sg13g2_decap_8
XFILLER_12_833 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_fill_1
XFILLER_12_877 VPWR VGND sg13g2_decap_8
XFILLER_11_398 VPWR VGND sg13g2_decap_4
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_decap_8
XFILLER_22_608 VPWR VGND sg13g2_fill_1
XFILLER_35_969 VPWR VGND sg13g2_decap_8
X_2981_ net184 VGND VPWR _0172_ ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_41_clk clknet_3_4__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_1932_ sdr_i.mac1.products_ff\[86\] sdr_i.mac1.products_ff\[69\] _0427_ VPWR VGND
+ sg13g2_xor2_1
XFILLER_30_674 VPWR VGND sg13g2_decap_8
X_1863_ _0398_ net302 net250 VPWR VGND sg13g2_nand2_1
X_1794_ VPWR VGND _1169_ net461 net444 _1155_ _0343_ net453 sg13g2_a221oi_1
XFILLER_7_892 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_2415_ _0831_ net814 _0336_ VPWR VGND sg13g2_nand2_1
X_2346_ ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] ppwm_i.u_ppwm.pwm_value\[8\] net399 _0766_
+ VPWR VGND sg13g2_mux2_1
X_2277_ VGND VPWR net386 _0666_ _0700_ _0699_ sg13g2_a21oi_1
XFILLER_38_730 VPWR VGND sg13g2_decap_8
XFILLER_38_763 VPWR VGND sg13g2_decap_8
XFILLER_41_906 VPWR VGND sg13g2_decap_8
XFILLER_26_969 VPWR VGND sg13g2_decap_8
XFILLER_34_980 VPWR VGND sg13g2_decap_8
XFILLER_40_449 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_32_clk clknet_3_5__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_32_36 VPWR VGND sg13g2_decap_8
XFILLER_20_162 VPWR VGND sg13g2_fill_2
XFILLER_5_818 VPWR VGND sg13g2_decap_8
XFILLER_4_339 VPWR VGND sg13g2_fill_2
XFILLER_0_534 VPWR VGND sg13g2_decap_8
XFILLER_17_903 VPWR VGND sg13g2_decap_8
XFILLER_29_752 VPWR VGND sg13g2_fill_1
XFILLER_44_711 VPWR VGND sg13g2_decap_8
XFILLER_16_424 VPWR VGND sg13g2_fill_1
XFILLER_43_232 VPWR VGND sg13g2_decap_8
X_3081__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_16_446 VPWR VGND sg13g2_decap_8
XFILLER_44_788 VPWR VGND sg13g2_decap_8
XFILLER_16_468 VPWR VGND sg13g2_fill_2
X_3029__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_40_983 VPWR VGND sg13g2_decap_8
XFILLER_11_173 VPWR VGND sg13g2_decap_8
X_3044__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_8_667 VPWR VGND sg13g2_decap_8
XFILLER_4_895 VPWR VGND sg13g2_decap_8
X_2200_ _1216_ net506 _0626_ VPWR VGND sg13g2_nor2_1
X_3180_ net522 VGND VPWR net206 sdr_i.mac1.sum_lvl2_ff\[9\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_39_538 VPWR VGND sg13g2_fill_2
X_2131_ VPWR VGND _0556_ _0555_ _0554_ _1227_ _0557_ ppwm_i.u_ppwm.global_counter\[12\]
+ sg13g2_a221oi_1
X_2062_ net422 VPWR _0501_ VGND net784 _0499_ sg13g2_o21ai_1
XFILLER_47_582 VPWR VGND sg13g2_decap_8
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_35_700 VPWR VGND sg13g2_decap_4
XFILLER_34_265 VPWR VGND sg13g2_decap_8
X_2964_ net436 VGND VPWR net655 ppwm_i.u_ppwm.global_counter\[7\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
X_1915_ net601 sdr_i.mac2.sum_lvl3_ff\[1\] _0418_ VPWR VGND sg13g2_nor2_1
XFILLER_31_961 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_3_3__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_2895_ net531 VGND VPWR _0086_ sdr_i.DP_1.matrix\[45\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_1846_ _0387_ net285 net237 VPWR VGND sg13g2_nand2_1
X_1777_ _1344_ ppwm_i.u_ppwm.u_mem.memory\[55\] net514 net517 VPWR VGND sg13g2_and3_1
X_2329_ _0749_ VPWR _0750_ VGND _1264_ net403 sg13g2_o21ai_1
XFILLER_25_210 VPWR VGND sg13g2_decap_8
XFILLER_25_232 VPWR VGND sg13g2_decap_8
XFILLER_38_593 VPWR VGND sg13g2_decap_8
XFILLER_13_405 VPWR VGND sg13g2_decap_8
XFILLER_14_928 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_22_961 VPWR VGND sg13g2_decap_8
XFILLER_40_279 VPWR VGND sg13g2_fill_2
XFILLER_4_114 VPWR VGND sg13g2_decap_8
XFILLER_1_821 VPWR VGND sg13g2_decap_8
XFILLER_49_825 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_17_722 VPWR VGND sg13g2_decap_4
XFILLER_29_560 VPWR VGND sg13g2_decap_4
XFILLER_17_733 VPWR VGND sg13g2_fill_1
XFILLER_17_755 VPWR VGND sg13g2_decap_4
XFILLER_44_552 VPWR VGND sg13g2_decap_4
XFILLER_31_202 VPWR VGND sg13g2_decap_8
XFILLER_31_268 VPWR VGND sg13g2_decap_8
XFILLER_40_780 VPWR VGND sg13g2_decap_8
XFILLER_9_954 VPWR VGND sg13g2_decap_8
XFILLER_13_983 VPWR VGND sg13g2_decap_8
X_2680_ net417 VPWR _1019_ VGND net477 net347 sg13g2_o21ai_1
X_1700_ _1269_ net694 net330 VPWR VGND sg13g2_nand2_1
X_1631_ VPWR _1202_ net692 VGND sg13g2_inv_1
X_1562_ VPWR _1133_ net677 VGND sg13g2_inv_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ net526 VGND VPWR net735 sdr_i.mac1.sum_lvl1_ff\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2114_ VGND VPWR _0539_ _0540_ _0541_ _0518_ sg13g2_a21oi_1
XFILLER_48_891 VPWR VGND sg13g2_decap_8
X_3094_ net62 VGND VPWR net668 ppwm_i.u_ppwm.u_mem.memory\[70\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_2045_ net664 net410 _0490_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_202 VPWR VGND sg13g2_decap_8
XFILLER_11_909 VPWR VGND sg13g2_decap_8
XFILLER_13_38 VPWR VGND sg13g2_fill_2
X_2947_ net536 VGND VPWR _0138_ sdr_i.DP_4.matrix\[36\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2878_ net239 _0141_ VPWR VGND sg13g2_buf_1
X_1829_ _0373_ _0374_ net548 _0375_ VPWR VGND sg13g2_nand3_1
Xhold420 ppwm_i.u_ppwm.pwm_value\[0\] VPWR VGND net800 sg13g2_dlygate4sd3_1
Xhold453 ppwm_i.u_ppwm.pwm_value\[7\] VPWR VGND net833 sg13g2_dlygate4sd3_1
XFILLER_1_106 VPWR VGND sg13g2_fill_2
Xhold431 ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] VPWR VGND net811 sg13g2_dlygate4sd3_1
Xhold442 ppwm_i.u_ppwm.global_counter\[1\] VPWR VGND net822 sg13g2_dlygate4sd3_1
XFILLER_18_519 VPWR VGND sg13g2_decap_4
XFILLER_41_533 VPWR VGND sg13g2_decap_8
XFILLER_14_725 VPWR VGND sg13g2_decap_8
XFILLER_16_1011 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_22_780 VPWR VGND sg13g2_fill_1
XFILLER_21_290 VPWR VGND sg13g2_fill_1
XFILLER_5_412 VPWR VGND sg13g2_fill_1
XFILLER_10_986 VPWR VGND sg13g2_decap_8
XFILLER_6_968 VPWR VGND sg13g2_decap_8
XFILLER_48_110 VPWR VGND sg13g2_fill_1
XFILLER_49_677 VPWR VGND sg13g2_decap_8
XFILLER_17_585 VPWR VGND sg13g2_decap_8
XFILLER_32_555 VPWR VGND sg13g2_decap_8
X_2801_ _1085_ VPWR _1086_ VGND ppwm_i.u_ppwm.u_pwm.counter\[3\] _1245_ sg13g2_o21ai_1
XFILLER_20_728 VPWR VGND sg13g2_decap_8
XFILLER_32_588 VPWR VGND sg13g2_decap_8
X_2732_ net416 VPWR _1045_ VGND net473 ppwm_i.u_ppwm.u_mem.memory\[91\] sg13g2_o21ai_1
X_2663_ VGND VPWR net485 _1152_ _0271_ _1010_ sg13g2_a21oi_1
X_2594_ net429 VPWR _0976_ VGND net493 ppwm_i.u_ppwm.u_mem.memory\[22\] sg13g2_o21ai_1
X_1614_ VPWR _1185_ net599 VGND sg13g2_inv_1
X_1545_ VPWR _1116_ net672 VGND sg13g2_inv_1
XFILLER_5_50 VPWR VGND sg13g2_decap_8
X_3215_ net536 VGND VPWR net212 sdr_i.mac2.sum_lvl1_ff\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_806 VPWR VGND sg13g2_decap_8
X_3146_ net523 VGND VPWR _0054_ sdr_i.mac1.products_ff\[17\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3077_ net129 VGND VPWR _0268_ ppwm_i.u_ppwm.u_mem.memory\[53\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2028_ VGND VPWR _1247_ net409 _0168_ _0478_ sg13g2_a21oi_1
XFILLER_11_717 VPWR VGND sg13g2_decap_4
XFILLER_3_938 VPWR VGND sg13g2_decap_8
XFILLER_2_404 VPWR VGND sg13g2_decap_8
XFILLER_49_12 VPWR VGND sg13g2_decap_8
XFILLER_46_1004 VPWR VGND sg13g2_decap_8
Xhold250 ppwm_i.u_ppwm.u_mem.memory\[74\] VPWR VGND net630 sg13g2_dlygate4sd3_1
Xhold261 _0308_ VPWR VGND net641 sg13g2_dlygate4sd3_1
Xhold294 _0270_ VPWR VGND net674 sg13g2_dlygate4sd3_1
Xhold272 ppwm_i.u_ppwm.u_mem.memory\[77\] VPWR VGND net652 sg13g2_dlygate4sd3_1
Xhold283 _0330_ VPWR VGND net663 sg13g2_dlygate4sd3_1
XFILLER_49_89 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_45_135 VPWR VGND sg13g2_decap_4
XFILLER_45_124 VPWR VGND sg13g2_fill_2
XFILLER_42_853 VPWR VGND sg13g2_decap_8
X_3008__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_14_70 VPWR VGND sg13g2_fill_1
XFILLER_6_710 VPWR VGND sg13g2_decap_8
XFILLER_6_754 VPWR VGND sg13g2_decap_8
XFILLER_6_776 VPWR VGND sg13g2_fill_2
XFILLER_5_264 VPWR VGND sg13g2_fill_2
XFILLER_1_481 VPWR VGND sg13g2_fill_1
X_3000_ net148 VGND VPWR _0191_ ppwm_i.u_ppwm.pc\[2\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_37_614 VPWR VGND sg13g2_fill_1
XFILLER_18_883 VPWR VGND sg13g2_decap_8
XFILLER_33_853 VPWR VGND sg13g2_decap_8
X_3092__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_32_352 VPWR VGND sg13g2_decap_8
XFILLER_20_558 VPWR VGND sg13g2_fill_1
X_2715_ VGND VPWR net462 _1126_ _0297_ _1036_ sg13g2_a21oi_1
XFILLER_10_17 VPWR VGND sg13g2_fill_2
X_2646_ net428 VPWR _1002_ VGND net492 net570 sg13g2_o21ai_1
X_2577_ VGND VPWR net495 _1195_ _0228_ _0967_ sg13g2_a21oi_1
X_1528_ VPWR _1099_ net604 VGND sg13g2_inv_1
XFILLER_28_647 VPWR VGND sg13g2_decap_8
X_3129_ net108 VGND VPWR net750 ppwm_i.u_ppwm.u_mem.memory\[105\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_24_820 VPWR VGND sg13g2_decap_8
XFILLER_35_58 VPWR VGND sg13g2_fill_2
XFILLER_24_875 VPWR VGND sg13g2_decap_8
XFILLER_13_1025 VPWR VGND sg13g2_decap_4
XFILLER_46_400 VPWR VGND sg13g2_decap_4
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_34_606 VPWR VGND sg13g2_decap_8
XFILLER_15_831 VPWR VGND sg13g2_decap_8
XFILLER_14_363 VPWR VGND sg13g2_decap_8
XFILLER_30_867 VPWR VGND sg13g2_decap_8
X_2500_ _0908_ VPWR _0909_ VGND _0895_ _0901_ sg13g2_o21ai_1
X_2431_ _0834_ _0831_ _0844_ _0846_ VPWR VGND sg13g2_a21o_1
XFILLER_6_595 VPWR VGND sg13g2_fill_2
X_2362_ _0779_ _0780_ net377 _0781_ VPWR VGND sg13g2_nand3_1
X_2293_ _1227_ net393 _0715_ VPWR VGND sg13g2_nor2_1
XFILLER_49_282 VPWR VGND sg13g2_decap_8
XFILLER_38_945 VPWR VGND sg13g2_decap_8
XFILLER_37_444 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_25_639 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_decap_4
XFILLER_36_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_300 VPWR VGND sg13g2_decap_8
X_2629_ VGND VPWR net481 _1169_ _0254_ _0993_ sg13g2_a21oi_1
XFILLER_0_738 VPWR VGND sg13g2_decap_8
XFILLER_28_400 VPWR VGND sg13g2_decap_8
XFILLER_29_934 VPWR VGND sg13g2_decap_8
XFILLER_46_46 VPWR VGND sg13g2_decap_4
XFILLER_28_488 VPWR VGND sg13g2_decap_8
XFILLER_15_138 VPWR VGND sg13g2_decap_8
XFILLER_12_812 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_fill_2
XFILLER_11_355 VPWR VGND sg13g2_fill_2
XFILLER_23_193 VPWR VGND sg13g2_fill_1
XFILLER_7_337 VPWR VGND sg13g2_decap_4
XFILLER_7_326 VPWR VGND sg13g2_fill_2
XFILLER_39_709 VPWR VGND sg13g2_fill_1
Xfanout390 _0336_ net390 VPWR VGND sg13g2_buf_8
XFILLER_19_400 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_35_948 VPWR VGND sg13g2_decap_8
XFILLER_34_447 VPWR VGND sg13g2_decap_8
XFILLER_34_458 VPWR VGND sg13g2_fill_2
XFILLER_34_469 VPWR VGND sg13g2_fill_1
X_2980_ net186 VGND VPWR net772 ppwm_i.u_ppwm.u_pwm.cmp_value\[3\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_43_992 VPWR VGND sg13g2_decap_8
X_1931_ net307 sdr_i.mac1.products_ff\[68\] _0019_ VPWR VGND sg13g2_xor2_1
X_1862_ _0397_ _0396_ _0067_ VPWR VGND sg13g2_xor2_1
X_1793_ _0342_ net441 _1162_ net448 _1176_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_871 VPWR VGND sg13g2_decap_8
X_2414_ VGND VPWR _0758_ _0827_ _0830_ _0829_ sg13g2_a21oi_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_29_208 VPWR VGND sg13g2_fill_2
X_2345_ _0762_ VPWR _0765_ VGND _0658_ _0764_ sg13g2_o21ai_1
X_2276_ net386 _0656_ _0699_ VPWR VGND sg13g2_nor2_1
XFILLER_38_753 VPWR VGND sg13g2_fill_1
XFILLER_26_948 VPWR VGND sg13g2_decap_8
XFILLER_25_436 VPWR VGND sg13g2_decap_8
XFILLER_25_447 VPWR VGND sg13g2_fill_2
XFILLER_40_428 VPWR VGND sg13g2_decap_4
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
X_3123__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_29_742 VPWR VGND sg13g2_fill_2
XFILLER_16_403 VPWR VGND sg13g2_decap_4
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_17_959 VPWR VGND sg13g2_decap_8
XFILLER_25_992 VPWR VGND sg13g2_decap_8
XFILLER_40_962 VPWR VGND sg13g2_decap_8
XFILLER_12_653 VPWR VGND sg13g2_decap_4
XFILLER_12_697 VPWR VGND sg13g2_fill_1
XFILLER_4_874 VPWR VGND sg13g2_decap_8
XFILLER_3_362 VPWR VGND sg13g2_decap_4
XFILLER_39_517 VPWR VGND sg13g2_decap_8
X_2130_ _0556_ ppwm_i.u_ppwm.pwm_value\[0\] ppwm_i.u_ppwm.global_counter\[10\] VPWR
+ VGND sg13g2_nand2b_1
X_2061_ net784 _0499_ _0500_ VPWR VGND sg13g2_and2_1
XFILLER_47_572 VPWR VGND sg13g2_fill_1
XFILLER_23_929 VPWR VGND sg13g2_decap_8
X_2963_ net436 VGND VPWR net321 ppwm_i.u_ppwm.global_counter\[6\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_22_428 VPWR VGND sg13g2_fill_2
X_1914_ _0417_ net601 sdr_i.mac2.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_31_940 VPWR VGND sg13g2_decap_8
X_2894_ net529 VGND VPWR _0085_ sdr_i.DP_1.matrix\[37\] clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
X_1845_ _0386_ net274 net220 VPWR VGND sg13g2_nand2_1
X_1776_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[34\] net448 _1343_ net461 sg13g2_a21oi_1
X_2328_ _0749_ ppwm_i.u_ppwm.global_counter\[13\] net403 VPWR VGND sg13g2_nand2_1
X_2259_ VGND VPWR _0682_ _0683_ net375 _0585_ sg13g2_a21oi_2
XFILLER_14_907 VPWR VGND sg13g2_decap_8
XFILLER_41_726 VPWR VGND sg13g2_decap_8
XFILLER_13_428 VPWR VGND sg13g2_decap_8
XFILLER_25_277 VPWR VGND sg13g2_fill_1
XFILLER_40_236 VPWR VGND sg13g2_decap_8
XFILLER_22_940 VPWR VGND sg13g2_decap_8
X_2980__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_1_800 VPWR VGND sg13g2_decap_8
XFILLER_0_321 VPWR VGND sg13g2_decap_4
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_1_877 VPWR VGND sg13g2_decap_8
XFILLER_0_365 VPWR VGND sg13g2_decap_4
XFILLER_44_531 VPWR VGND sg13g2_fill_2
XFILLER_16_255 VPWR VGND sg13g2_fill_2
XFILLER_13_962 VPWR VGND sg13g2_decap_8
XFILLER_9_933 VPWR VGND sg13g2_decap_8
XFILLER_33_91 VPWR VGND sg13g2_decap_8
X_1630_ VPWR _1201_ ppwm_i.u_ppwm.u_mem.memory\[8\] VGND sg13g2_inv_1
X_1561_ VPWR _1132_ net652 VGND sg13g2_inv_1
X_3231_ net525 VGND VPWR net603 sdr_i.mac2.total_sum\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3162_ net533 VGND VPWR net218 sdr_i.mac1.sum_lvl1_ff\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3099__43 VPWR VGND net43 sg13g2_tiehi
X_2113_ _0531_ VPWR _0540_ VGND _0530_ _0532_ sg13g2_o21ai_1
XFILLER_48_870 VPWR VGND sg13g2_decap_8
X_3093_ net66 VGND VPWR _0284_ ppwm_i.u_ppwm.u_mem.memory\[69\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_2044_ net504 net411 _0489_ VPWR VGND sg13g2_nor2_1
XFILLER_23_748 VPWR VGND sg13g2_decap_4
XFILLER_35_586 VPWR VGND sg13g2_decap_8
XFILLER_22_258 VPWR VGND sg13g2_decap_8
X_2946_ net540 VGND VPWR _0137_ sdr_i.DP_4.matrix\[28\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2877_ net300 _0140_ VPWR VGND sg13g2_buf_1
X_1828_ _0374_ sdr_i.mac1.total_sum\[0\] sdr_i.mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
Xhold410 _0151_ VPWR VGND net790 sg13g2_dlygate4sd3_1
Xhold454 _0202_ VPWR VGND net834 sg13g2_dlygate4sd3_1
X_1759_ VGND VPWR _1103_ net451 _1326_ net460 sg13g2_a21oi_1
Xhold421 _0195_ VPWR VGND net801 sg13g2_dlygate4sd3_1
Xhold432 ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] VPWR VGND net812 sg13g2_dlygate4sd3_1
Xhold443 _0457_ VPWR VGND net823 sg13g2_dlygate4sd3_1
XFILLER_38_36 VPWR VGND sg13g2_fill_1
XFILLER_38_69 VPWR VGND sg13g2_decap_4
XFILLER_46_829 VPWR VGND sg13g2_decap_8
XFILLER_45_339 VPWR VGND sg13g2_fill_1
XFILLER_26_564 VPWR VGND sg13g2_decap_8
XFILLER_41_512 VPWR VGND sg13g2_fill_2
XFILLER_26_586 VPWR VGND sg13g2_fill_2
XFILLER_41_556 VPWR VGND sg13g2_decap_8
XFILLER_13_236 VPWR VGND sg13g2_decap_8
XFILLER_9_218 VPWR VGND sg13g2_fill_1
XFILLER_10_965 VPWR VGND sg13g2_decap_8
XFILLER_6_947 VPWR VGND sg13g2_decap_8
XFILLER_49_656 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_542 VPWR VGND sg13g2_fill_2
XFILLER_45_884 VPWR VGND sg13g2_decap_8
XFILLER_32_501 VPWR VGND sg13g2_decap_4
X_2800_ _1085_ ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] ppwm_i.u_ppwm.u_pwm.counter\[4\]
+ VPWR VGND sg13g2_nand2b_1
X_2731_ VGND VPWR net465 _1118_ _0305_ _1044_ sg13g2_a21oi_1
XFILLER_12_280 VPWR VGND sg13g2_decap_4
XFILLER_13_792 VPWR VGND sg13g2_decap_8
X_2662_ net426 VPWR _1010_ VGND net485 ppwm_i.u_ppwm.u_mem.memory\[56\] sg13g2_o21ai_1
X_2593_ VGND VPWR net493 _1187_ _0236_ _0975_ sg13g2_a21oi_1
X_1613_ VPWR _1184_ net586 VGND sg13g2_inv_1
X_1544_ VPWR _1115_ net640 VGND sg13g2_inv_1
X_3214_ net532 VGND VPWR net202 sdr_i.mac2.sum_lvl1_ff\[32\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3145_ net523 VGND VPWR _0075_ sdr_i.mac1.products_ff\[1\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3076_ net133 VGND VPWR net658 ppwm_i.u_ppwm.u_mem.memory\[52\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_42_309 VPWR VGND sg13g2_decap_8
X_2027_ net421 VPWR _0478_ VGND ppwm_i.u_ppwm.pwm_value\[0\] net409 sg13g2_o21ai_1
XFILLER_39_1023 VPWR VGND sg13g2_decap_4
XFILLER_36_884 VPWR VGND sg13g2_decap_8
XFILLER_11_707 VPWR VGND sg13g2_fill_2
XFILLER_10_239 VPWR VGND sg13g2_decap_8
X_2929_ net537 VGND VPWR _0120_ sdr_i.DP_3.matrix\[36\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_40_37 VPWR VGND sg13g2_fill_1
XFILLER_3_917 VPWR VGND sg13g2_decap_8
Xhold240 _0274_ VPWR VGND net620 sg13g2_dlygate4sd3_1
Xhold251 _0288_ VPWR VGND net631 sg13g2_dlygate4sd3_1
Xhold262 ppwm_i.u_ppwm.u_mem.memory\[10\] VPWR VGND net642 sg13g2_dlygate4sd3_1
Xhold284 ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold273 _0292_ VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold295 ppwm_i.u_ppwm.u_mem.memory\[34\] VPWR VGND net675 sg13g2_dlygate4sd3_1
XFILLER_18_328 VPWR VGND sg13g2_fill_1
XFILLER_45_158 VPWR VGND sg13g2_decap_8
XFILLER_42_832 VPWR VGND sg13g2_decap_8
XFILLER_27_884 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_fill_1
XFILLER_6_788 VPWR VGND sg13g2_decap_8
XFILLER_6_799 VPWR VGND sg13g2_fill_2
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_464 VPWR VGND sg13g2_decap_4
XFILLER_39_90 VPWR VGND sg13g2_decap_8
XFILLER_37_659 VPWR VGND sg13g2_decap_8
XFILLER_33_832 VPWR VGND sg13g2_decap_8
XFILLER_45_692 VPWR VGND sg13g2_fill_1
XFILLER_44_191 VPWR VGND sg13g2_fill_1
X_2714_ net413 VPWR _1036_ VGND net462 ppwm_i.u_ppwm.u_mem.memory\[82\] sg13g2_o21ai_1
XFILLER_9_582 VPWR VGND sg13g2_decap_8
X_2645_ VGND VPWR net492 _1161_ _0262_ _1001_ sg13g2_a21oi_1
X_2576_ net432 VPWR _0967_ VGND net499 net609 sg13g2_o21ai_1
X_1527_ VPWR _1098_ net3 VGND sg13g2_inv_1
XFILLER_19_27 VPWR VGND sg13g2_fill_1
X_3128_ net123 VGND VPWR _0319_ ppwm_i.u_ppwm.u_mem.memory\[104\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_43_629 VPWR VGND sg13g2_decap_8
XFILLER_42_117 VPWR VGND sg13g2_fill_2
X_3059_ net32 VGND VPWR net585 ppwm_i.u_ppwm.u_mem.memory\[35\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_23_331 VPWR VGND sg13g2_decap_8
XFILLER_24_854 VPWR VGND sg13g2_decap_8
XFILLER_13_1004 VPWR VGND sg13g2_decap_8
XFILLER_3_703 VPWR VGND sg13g2_decap_8
XFILLER_3_758 VPWR VGND sg13g2_fill_1
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_46_423 VPWR VGND sg13g2_decap_8
X_3084__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_46_467 VPWR VGND sg13g2_decap_4
XFILLER_18_147 VPWR VGND sg13g2_decap_8
XFILLER_46_478 VPWR VGND sg13g2_decap_8
XFILLER_15_810 VPWR VGND sg13g2_fill_1
XFILLER_27_670 VPWR VGND sg13g2_decap_8
XFILLER_27_681 VPWR VGND sg13g2_fill_1
XFILLER_14_331 VPWR VGND sg13g2_fill_1
XFILLER_42_684 VPWR VGND sg13g2_decap_8
XFILLER_41_172 VPWR VGND sg13g2_decap_4
XFILLER_41_161 VPWR VGND sg13g2_fill_2
XFILLER_30_846 VPWR VGND sg13g2_decap_8
X_2430_ _0834_ _0844_ _0831_ _0845_ VPWR VGND sg13g2_nand3_1
XFILLER_29_1011 VPWR VGND sg13g2_decap_8
X_2361_ _0780_ _0778_ _0777_ VPWR VGND sg13g2_nand2b_1
X_3171__196 VPWR VGND net196 sg13g2_tiehi
X_2292_ ppwm_i.u_ppwm.pwm_value\[2\] net407 net405 _0714_ VPWR VGND sg13g2_or3_1
XFILLER_2_30 VPWR VGND sg13g2_decap_8
XFILLER_38_924 VPWR VGND sg13g2_decap_8
XFILLER_49_261 VPWR VGND sg13g2_decap_8
XFILLER_46_990 VPWR VGND sg13g2_decap_8
XFILLER_25_618 VPWR VGND sg13g2_decap_8
XFILLER_37_478 VPWR VGND sg13g2_decap_8
XFILLER_33_640 VPWR VGND sg13g2_fill_1
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_21_17 VPWR VGND sg13g2_fill_2
X_2628_ net425 VPWR _0993_ VGND net481 net698 sg13g2_o21ai_1
XFILLER_0_717 VPWR VGND sg13g2_decap_8
X_2559_ VGND VPWR net498 _1204_ _0219_ _0958_ sg13g2_a21oi_1
XFILLER_29_913 VPWR VGND sg13g2_decap_8
XFILLER_28_467 VPWR VGND sg13g2_decap_8
XFILLER_44_949 VPWR VGND sg13g2_decap_8
XFILLER_8_806 VPWR VGND sg13g2_fill_1
XFILLER_8_839 VPWR VGND sg13g2_decap_8
XFILLER_11_61 VPWR VGND sg13g2_decap_8
Xfanout391 net392 net391 VPWR VGND sg13g2_buf_8
Xfanout380 _0671_ net380 VPWR VGND sg13g2_buf_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_35_927 VPWR VGND sg13g2_decap_8
XFILLER_34_426 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_42_470 VPWR VGND sg13g2_fill_1
X_1930_ _0426_ net741 net307 VPWR VGND sg13g2_nand2_1
XFILLER_30_654 VPWR VGND sg13g2_fill_1
X_1861_ _0397_ net309 net239 VPWR VGND sg13g2_nand2_1
XFILLER_7_850 VPWR VGND sg13g2_decap_8
X_1792_ VPWR VGND _0340_ _1231_ _0339_ _0337_ _0341_ _0338_ sg13g2_a221oi_1
XFILLER_6_382 VPWR VGND sg13g2_decap_4
X_2413_ _0829_ _0797_ _0828_ VPWR VGND sg13g2_nand2_1
X_2344_ _0764_ _0351_ _0740_ VPWR VGND sg13g2_nand2_2
XFILLER_28_0 VPWR VGND sg13g2_fill_1
X_2275_ _0662_ _0697_ net387 _0698_ VPWR VGND sg13g2_mux2_1
XFILLER_26_927 VPWR VGND sg13g2_decap_8
XFILLER_38_798 VPWR VGND sg13g2_decap_8
XFILLER_25_459 VPWR VGND sg13g2_decap_8
XFILLER_33_481 VPWR VGND sg13g2_decap_8
XFILLER_21_665 VPWR VGND sg13g2_fill_2
XFILLER_21_676 VPWR VGND sg13g2_fill_2
XFILLER_10_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_503 VPWR VGND sg13g2_decap_8
XFILLER_0_569 VPWR VGND sg13g2_decap_8
XFILLER_17_938 VPWR VGND sg13g2_decap_8
XFILLER_29_787 VPWR VGND sg13g2_decap_8
XFILLER_25_971 VPWR VGND sg13g2_decap_8
XFILLER_32_919 VPWR VGND sg13g2_decap_8
XFILLER_43_289 VPWR VGND sg13g2_fill_1
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_40_941 VPWR VGND sg13g2_decap_8
XFILLER_12_632 VPWR VGND sg13g2_fill_2
XFILLER_4_853 VPWR VGND sg13g2_decap_8
XFILLER_26_1025 VPWR VGND sg13g2_decap_4
X_2060_ net455 net708 _0499_ _0179_ VPWR VGND sg13g2_nor3_1
XFILLER_19_242 VPWR VGND sg13g2_decap_8
XFILLER_35_724 VPWR VGND sg13g2_decap_4
XFILLER_34_234 VPWR VGND sg13g2_decap_4
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_35_757 VPWR VGND sg13g2_fill_2
XFILLER_23_908 VPWR VGND sg13g2_decap_8
X_2962_ net435 VGND VPWR net334 ppwm_i.u_ppwm.global_counter\[5\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_1913_ net259 sdr_i.mac2.sum_lvl3_ff\[2\] _0007_ VPWR VGND sg13g2_xor2_1
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
X_2893_ net529 VGND VPWR _0084_ sdr_i.DP_1.matrix\[36\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_31_996 VPWR VGND sg13g2_decap_8
X_1844_ _0385_ _0384_ _0053_ VPWR VGND sg13g2_xor2_1
X_1775_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[20\] _1341_ net440 ppwm_i.u_ppwm.u_mem.memory\[6\]
+ _1342_ net449 sg13g2_a221oi_1
X_2327_ VPWR VGND _0691_ _0747_ _0742_ net379 _0748_ _0698_ sg13g2_a221oi_1
X_2258_ _0682_ ppwm_i.u_ppwm.u_ex.state_q\[2\] _0681_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_49 VPWR VGND sg13g2_decap_4
XFILLER_38_573 VPWR VGND sg13g2_fill_2
XFILLER_26_735 VPWR VGND sg13g2_decap_8
X_2189_ _0614_ VPWR _0615_ VGND _0611_ _0613_ sg13g2_o21ai_1
XFILLER_22_996 VPWR VGND sg13g2_decap_8
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_0_300 VPWR VGND sg13g2_decap_8
XFILLER_0_344 VPWR VGND sg13g2_decap_8
XFILLER_1_856 VPWR VGND sg13g2_decap_8
XFILLER_0_388 VPWR VGND sg13g2_decap_8
XFILLER_48_348 VPWR VGND sg13g2_decap_4
XFILLER_29_595 VPWR VGND sg13g2_fill_2
XFILLER_16_234 VPWR VGND sg13g2_decap_8
XFILLER_17_768 VPWR VGND sg13g2_fill_1
XFILLER_32_705 VPWR VGND sg13g2_decap_4
XFILLER_32_727 VPWR VGND sg13g2_decap_8
XFILLER_32_738 VPWR VGND sg13g2_fill_2
XFILLER_32_749 VPWR VGND sg13g2_fill_2
XFILLER_9_912 VPWR VGND sg13g2_decap_8
XFILLER_13_941 VPWR VGND sg13g2_decap_8
XFILLER_31_248 VPWR VGND sg13g2_decap_8
XFILLER_9_989 VPWR VGND sg13g2_decap_8
XFILLER_8_499 VPWR VGND sg13g2_decap_8
X_1560_ VPWR _1131_ ppwm_i.u_ppwm.u_mem.memory\[78\] VGND sg13g2_inv_1
X_3018__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_3_193 VPWR VGND sg13g2_decap_8
X_3230_ net525 VGND VPWR net783 sdr_i.mac2.total_sum\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3161_ net522 VGND VPWR _0073_ sdr_i.mac1.products_ff\[137\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_39_337 VPWR VGND sg13g2_decap_8
X_2112_ net408 _0538_ _0539_ VPWR VGND sg13g2_nor2_1
X_3092_ net70 VGND VPWR _0283_ ppwm_i.u_ppwm.u_mem.memory\[68\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_3129__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_47_370 VPWR VGND sg13g2_fill_2
X_2043_ net455 net792 _0173_ VPWR VGND sg13g2_nor2_1
X_2945_ net539 VGND VPWR _0136_ sdr_i.DP_4.matrix\[27\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2876_ net251 _0139_ VPWR VGND sg13g2_buf_1
XFILLER_31_793 VPWR VGND sg13g2_decap_8
X_1827_ VGND VPWR _0373_ sdr_i.mac2.total_sum\[0\] sdr_i.mac1.total_sum\[0\] sg13g2_or2_1
Xhold400 ppwm_i.u_ppwm.global_counter\[16\] VPWR VGND net780 sg13g2_dlygate4sd3_1
Xhold411 ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] VPWR VGND net791 sg13g2_dlygate4sd3_1
Xhold422 ppwm_i.u_ppwm.u_pwm.cmp_value\[8\] VPWR VGND net802 sg13g2_dlygate4sd3_1
X_1758_ _1324_ _1231_ _1318_ _1325_ VPWR VGND sg13g2_a21o_2
Xhold444 _0149_ VPWR VGND net824 sg13g2_dlygate4sd3_1
Xhold433 ppwm_i.u_ppwm.global_counter\[14\] VPWR VGND net813 sg13g2_dlygate4sd3_1
X_1689_ VPWR _1260_ ppwm_i.u_ppwm.global_counter\[8\] VGND sg13g2_inv_1
Xhold455 ppwm_i.u_ppwm.pc\[3\] VPWR VGND net835 sg13g2_dlygate4sd3_1
XFILLER_46_808 VPWR VGND sg13g2_decap_8
XFILLER_10_944 VPWR VGND sg13g2_decap_8
XFILLER_6_926 VPWR VGND sg13g2_decap_8
XFILLER_5_469 VPWR VGND sg13g2_decap_8
XFILLER_0_130 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_48_101 VPWR VGND sg13g2_decap_8
XFILLER_0_152 VPWR VGND sg13g2_decap_8
XFILLER_49_635 VPWR VGND sg13g2_decap_8
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_45_863 VPWR VGND sg13g2_decap_8
XFILLER_44_362 VPWR VGND sg13g2_decap_8
XFILLER_13_771 VPWR VGND sg13g2_fill_2
X_2730_ net415 VPWR _1044_ VGND net465 net614 sg13g2_o21ai_1
X_2661_ VGND VPWR net485 _1153_ _0270_ _1009_ sg13g2_a21oi_1
X_1612_ _1183_ net691 VPWR VGND sg13g2_inv_2
X_2592_ net428 VPWR _0975_ VGND net493 ppwm_i.u_ppwm.u_mem.memory\[21\] sg13g2_o21ai_1
X_1543_ VPWR _1114_ net597 VGND sg13g2_inv_1
X_3213_ net541 VGND VPWR net740 sdr_i.mac2.sum_lvl1_ff\[25\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_39_123 VPWR VGND sg13g2_fill_2
X_3144_ net523 VGND VPWR _0074_ sdr_i.mac1.products_ff\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3075_ net137 VGND VPWR _0266_ ppwm_i.u_ppwm.u_mem.memory\[51\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_39_189 VPWR VGND sg13g2_decap_8
X_2026_ _1236_ _0475_ _1234_ _0477_ VPWR VGND _0476_ sg13g2_nand4_1
XFILLER_39_1002 VPWR VGND sg13g2_decap_8
XFILLER_36_863 VPWR VGND sg13g2_decap_8
XFILLER_23_524 VPWR VGND sg13g2_decap_8
XFILLER_23_568 VPWR VGND sg13g2_decap_8
X_2928_ net539 VGND VPWR _0119_ sdr_i.DP_3.matrix\[28\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2859_ net309 _0122_ VPWR VGND sg13g2_buf_1
Xhold252 ppwm_i.u_ppwm.u_mem.memory\[57\] VPWR VGND net632 sg13g2_dlygate4sd3_1
Xhold241 ppwm_i.u_ppwm.u_mem.memory\[22\] VPWR VGND net621 sg13g2_dlygate4sd3_1
Xhold230 _0227_ VPWR VGND net610 sg13g2_dlygate4sd3_1
Xhold274 ppwm_i.u_ppwm.global_counter\[7\] VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold285 _0174_ VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold263 ppwm_i.u_ppwm.u_mem.memory\[38\] VPWR VGND net643 sg13g2_dlygate4sd3_1
Xhold296 _0248_ VPWR VGND net676 sg13g2_dlygate4sd3_1
XFILLER_49_69 VPWR VGND sg13g2_decap_4
XFILLER_49_58 VPWR VGND sg13g2_fill_2
XFILLER_19_819 VPWR VGND sg13g2_fill_2
XFILLER_27_863 VPWR VGND sg13g2_decap_8
XFILLER_42_811 VPWR VGND sg13g2_decap_8
XFILLER_26_351 VPWR VGND sg13g2_decap_8
XFILLER_42_888 VPWR VGND sg13g2_decap_8
XFILLER_41_376 VPWR VGND sg13g2_decap_8
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_49_421 VPWR VGND sg13g2_decap_8
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_49_443 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_4
XFILLER_18_863 VPWR VGND sg13g2_fill_2
XFILLER_33_811 VPWR VGND sg13g2_decap_8
XFILLER_33_888 VPWR VGND sg13g2_decap_8
XFILLER_20_549 VPWR VGND sg13g2_decap_8
X_2713_ VGND VPWR net463 _1127_ _0296_ _1035_ sg13g2_a21oi_1
X_2644_ net428 VPWR _1001_ VGND net492 ppwm_i.u_ppwm.u_mem.memory\[47\] sg13g2_o21ai_1
X_2575_ VGND VPWR net499 _1196_ _0227_ _0966_ sg13g2_a21oi_1
X_1526_ VPWR _1097_ net582 VGND sg13g2_inv_1
X_3127_ net139 VGND VPWR _0318_ ppwm_i.u_ppwm.u_mem.memory\[103\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_43_608 VPWR VGND sg13g2_decap_8
X_3058_ net34 VGND VPWR _0249_ ppwm_i.u_ppwm.u_mem.memory\[34\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2009_ VGND VPWR ppwm_i.u_ppwm.global_counter\[11\] _0466_ _0468_ net719 sg13g2_a21oi_1
XFILLER_35_192 VPWR VGND sg13g2_fill_2
XFILLER_23_343 VPWR VGND sg13g2_decap_8
XFILLER_7_509 VPWR VGND sg13g2_fill_2
XFILLER_2_258 VPWR VGND sg13g2_decap_8
Xfanout540 net541 net540 VPWR VGND sg13g2_buf_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_19_638 VPWR VGND sg13g2_decap_4
XFILLER_46_446 VPWR VGND sg13g2_decap_8
XFILLER_46_435 VPWR VGND sg13g2_fill_1
XFILLER_18_126 VPWR VGND sg13g2_decap_4
XFILLER_15_844 VPWR VGND sg13g2_fill_1
XFILLER_33_129 VPWR VGND sg13g2_decap_8
XFILLER_42_663 VPWR VGND sg13g2_decap_4
XFILLER_42_696 VPWR VGND sg13g2_decap_4
XFILLER_41_151 VPWR VGND sg13g2_fill_2
XFILLER_15_899 VPWR VGND sg13g2_decap_8
XFILLER_30_825 VPWR VGND sg13g2_decap_8
XFILLER_6_597 VPWR VGND sg13g2_fill_1
X_2360_ _0779_ _0777_ _0778_ VPWR VGND sg13g2_nand2b_1
XFILLER_2_781 VPWR VGND sg13g2_decap_8
X_2291_ _0702_ _0686_ _0703_ _0713_ VPWR VGND sg13g2_a21o_2
XFILLER_49_240 VPWR VGND sg13g2_decap_8
XFILLER_2_20 VPWR VGND sg13g2_fill_1
XFILLER_38_903 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_decap_8
XFILLER_18_671 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_44_clk clknet_3_1__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_33_663 VPWR VGND sg13g2_decap_8
XFILLER_32_151 VPWR VGND sg13g2_fill_2
XFILLER_9_380 VPWR VGND sg13g2_decap_4
X_2627_ VGND VPWR net482 _1170_ _0253_ _0992_ sg13g2_a21oi_1
X_2558_ net433 VPWR _0958_ VGND net498 net656 sg13g2_o21ai_1
X_2489_ VGND VPWR _0875_ _0897_ _0899_ _0898_ sg13g2_a21oi_1
XFILLER_29_969 VPWR VGND sg13g2_decap_8
XFILLER_44_928 VPWR VGND sg13g2_decap_8
XFILLER_37_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_35_clk clknet_3_5__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_11_357 VPWR VGND sg13g2_fill_1
XFILLER_20_891 VPWR VGND sg13g2_decap_8
XFILLER_3_501 VPWR VGND sg13g2_decap_8
X_2990__167 VPWR VGND net167 sg13g2_tiehi
Xfanout392 _0335_ net392 VPWR VGND sg13g2_buf_8
Xfanout370 _0861_ net370 VPWR VGND sg13g2_buf_8
Xfanout381 net382 net381 VPWR VGND sg13g2_buf_8
XFILLER_4_1014 VPWR VGND sg13g2_decap_8
XFILLER_46_232 VPWR VGND sg13g2_fill_2
XFILLER_35_906 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_46_254 VPWR VGND sg13g2_fill_2
XFILLER_46_243 VPWR VGND sg13g2_decap_8
XFILLER_34_405 VPWR VGND sg13g2_decap_8
XFILLER_43_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_7__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_14_162 VPWR VGND sg13g2_fill_1
XFILLER_14_184 VPWR VGND sg13g2_decap_8
X_1860_ _0396_ net300 net243 VPWR VGND sg13g2_nand2_1
X_1791_ VPWR VGND _1141_ net510 net442 _1127_ _0340_ net450 sg13g2_a221oi_1
XFILLER_6_350 VPWR VGND sg13g2_decap_8
X_2412_ _0336_ VPWR _0828_ VGND net503 net504 sg13g2_o21ai_1
X_2343_ _0350_ _0739_ _0763_ VPWR VGND sg13g2_nor2_2
X_2274_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] ppwm_i.u_ppwm.pwm_value\[5\] net399 _0697_
+ VPWR VGND sg13g2_mux2_1
XFILLER_26_906 VPWR VGND sg13g2_decap_8
XFILLER_38_744 VPWR VGND sg13g2_decap_8
XFILLER_25_416 VPWR VGND sg13g2_fill_1
XFILLER_37_265 VPWR VGND sg13g2_decap_8
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_16_29 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_17_clk clknet_3_3__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_40_408 VPWR VGND sg13g2_decap_4
XFILLER_34_994 VPWR VGND sg13g2_decap_8
XFILLER_21_644 VPWR VGND sg13g2_decap_8
X_1989_ net326 net710 ppwm_i.u_ppwm.global_counter\[1\] ppwm_i.u_ppwm.global_counter\[0\]
+ _0458_ VPWR VGND sg13g2_and4_1
XFILLER_48_508 VPWR VGND sg13g2_fill_1
XFILLER_0_548 VPWR VGND sg13g2_decap_8
XFILLER_28_232 VPWR VGND sg13g2_decap_8
XFILLER_17_917 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_43_246 VPWR VGND sg13g2_fill_1
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_25_950 VPWR VGND sg13g2_decap_8
XFILLER_43_279 VPWR VGND sg13g2_fill_2
XFILLER_40_920 VPWR VGND sg13g2_decap_8
XFILLER_40_997 VPWR VGND sg13g2_decap_8
XFILLER_7_169 VPWR VGND sg13g2_decap_4
XFILLER_4_832 VPWR VGND sg13g2_decap_8
XFILLER_26_1004 VPWR VGND sg13g2_decap_8
XFILLER_21_8 VPWR VGND sg13g2_fill_1
XFILLER_19_232 VPWR VGND sg13g2_fill_1
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_34_213 VPWR VGND sg13g2_decap_8
XFILLER_16_983 VPWR VGND sg13g2_decap_8
XFILLER_34_279 VPWR VGND sg13g2_fill_1
X_2961_ net435 VGND VPWR _0152_ ppwm_i.u_ppwm.global_counter\[4\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_1912_ _0416_ sdr_i.mac2.sum_lvl3_ff\[2\] net259 VPWR VGND sg13g2_nand2_1
XFILLER_8_30 VPWR VGND sg13g2_decap_4
X_2892_ net535 VGND VPWR _0083_ sdr_i.DP_1.matrix\[28\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_30_463 VPWR VGND sg13g2_decap_8
XFILLER_31_975 VPWR VGND sg13g2_decap_8
XFILLER_8_85 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_fill_2
X_1843_ _0385_ net289 net233 VPWR VGND sg13g2_nand2_1
XFILLER_30_496 VPWR VGND sg13g2_fill_1
X_1774_ _1341_ ppwm_i.u_ppwm.u_mem.memory\[27\] net514 net517 VPWR VGND sg13g2_and3_1
Xclkbuf_leaf_6_clk clknet_3_0__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
X_2326_ _0659_ _0746_ _0747_ VPWR VGND sg13g2_and2_1
X_2257_ _0681_ _0680_ net398 _0679_ net380 VPWR VGND sg13g2_a22oi_1
XFILLER_26_703 VPWR VGND sg13g2_fill_2
XFILLER_26_714 VPWR VGND sg13g2_fill_2
X_2188_ _0614_ ppwm_i.u_ppwm.global_counter\[4\] _1215_ ppwm_i.u_ppwm.global_counter\[5\]
+ _1214_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_246 VPWR VGND sg13g2_decap_8
XFILLER_40_205 VPWR VGND sg13g2_decap_8
XFILLER_34_791 VPWR VGND sg13g2_decap_8
XFILLER_22_975 VPWR VGND sg13g2_decap_8
X_3026__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_21_496 VPWR VGND sg13g2_decap_8
X_3041__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_4_128 VPWR VGND sg13g2_fill_1
XFILLER_1_835 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_decap_8
XFILLER_29_530 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_fill_1
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_588 VPWR VGND sg13g2_decap_8
XFILLER_13_920 VPWR VGND sg13g2_decap_8
XFILLER_25_780 VPWR VGND sg13g2_fill_2
XFILLER_31_216 VPWR VGND sg13g2_decap_8
XFILLER_31_227 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_fill_2
XFILLER_12_452 VPWR VGND sg13g2_fill_2
XFILLER_40_794 VPWR VGND sg13g2_decap_8
XFILLER_9_968 VPWR VGND sg13g2_decap_8
XFILLER_12_474 VPWR VGND sg13g2_fill_2
XFILLER_13_997 VPWR VGND sg13g2_decap_8
XFILLER_8_489 VPWR VGND sg13g2_decap_4
XFILLER_8_467 VPWR VGND sg13g2_fill_2
XFILLER_8_456 VPWR VGND sg13g2_decap_8
XFILLER_4_684 VPWR VGND sg13g2_fill_1
X_3160_ net522 VGND VPWR _0072_ sdr_i.mac1.products_ff\[136\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3091_ net74 VGND VPWR net575 ppwm_i.u_ppwm.u_mem.memory\[67\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_12_4 VPWR VGND sg13g2_decap_8
Xhold1 sdr_i.mac1.products_ff\[136\] VPWR VGND net201 sg13g2_dlygate4sd3_1
X_2111_ _1231_ net406 _0538_ VPWR VGND sg13g2_nor2_1
X_2042_ _0487_ VPWR _0488_ VGND ppwm_i.u_ppwm.pwm_value\[5\] net410 sg13g2_o21ai_1
XFILLER_22_216 VPWR VGND sg13g2_decap_8
XFILLER_35_599 VPWR VGND sg13g2_decap_8
XFILLER_22_249 VPWR VGND sg13g2_decap_4
X_2944_ net539 VGND VPWR _0135_ sdr_i.DP_4.matrix\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_31_772 VPWR VGND sg13g2_decap_8
X_2875_ net277 _0138_ VPWR VGND sg13g2_buf_1
X_1826_ net318 VPWR _0001_ VGND _1279_ _0367_ sg13g2_o21ai_1
Xhold401 _0164_ VPWR VGND net781 sg13g2_dlygate4sd3_1
Xhold434 ppwm_i.u_ppwm.pwm_value\[8\] VPWR VGND net814 sg13g2_dlygate4sd3_1
Xhold423 _0494_ VPWR VGND net803 sg13g2_dlygate4sd3_1
Xhold412 _0488_ VPWR VGND net792 sg13g2_dlygate4sd3_1
X_1757_ _1324_ _1322_ _1323_ _1321_ _1319_ VPWR VGND sg13g2_a22oi_1
Xhold445 ppwm_i.u_ppwm.pc\[1\] VPWR VGND net825 sg13g2_dlygate4sd3_1
X_1688_ _1259_ net335 VPWR VGND sg13g2_inv_2
Xhold456 ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] VPWR VGND net836 sg13g2_dlygate4sd3_1
X_2309_ _0719_ _0726_ net373 _0731_ VPWR VGND _0730_ sg13g2_nand4_1
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_45_319 VPWR VGND sg13g2_fill_2
XFILLER_39_883 VPWR VGND sg13g2_decap_8
XFILLER_26_544 VPWR VGND sg13g2_decap_4
XFILLER_41_514 VPWR VGND sg13g2_fill_1
XFILLER_16_1025 VPWR VGND sg13g2_decap_4
XFILLER_10_923 VPWR VGND sg13g2_decap_8
XFILLER_22_794 VPWR VGND sg13g2_fill_1
XFILLER_6_905 VPWR VGND sg13g2_decap_8
XFILLER_5_426 VPWR VGND sg13g2_fill_2
XFILLER_49_614 VPWR VGND sg13g2_decap_8
XFILLER_0_197 VPWR VGND sg13g2_decap_8
XFILLER_0_186 VPWR VGND sg13g2_fill_2
XFILLER_37_809 VPWR VGND sg13g2_decap_8
XFILLER_28_82 VPWR VGND sg13g2_decap_8
XFILLER_45_842 VPWR VGND sg13g2_decap_8
XFILLER_44_341 VPWR VGND sg13g2_decap_8
XFILLER_17_544 VPWR VGND sg13g2_fill_1
XFILLER_8_264 VPWR VGND sg13g2_fill_2
XFILLER_8_253 VPWR VGND sg13g2_decap_8
X_2660_ net426 VPWR _1009_ VGND net485 ppwm_i.u_ppwm.u_mem.memory\[55\] sg13g2_o21ai_1
XFILLER_8_286 VPWR VGND sg13g2_decap_8
XFILLER_8_275 VPWR VGND sg13g2_fill_2
X_1611_ VPWR _1182_ net550 VGND sg13g2_inv_1
X_2591_ VGND VPWR net493 _1188_ _0235_ _0974_ sg13g2_a21oi_1
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_1542_ VPWR _1113_ net635 VGND sg13g2_inv_1
X_3212_ net541 VGND VPWR net258 sdr_i.mac2.sum_lvl1_ff\[24\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3143_ net194 VGND VPWR _0334_ ppwm_i.u_ppwm.data_o clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_39_168 VPWR VGND sg13g2_decap_8
X_3074_ net141 VGND VPWR net367 ppwm_i.u_ppwm.u_mem.memory\[50\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2025_ ppwm_i.u_ppwm.u_pwm.counter\[7\] ppwm_i.u_ppwm.u_pwm.counter\[6\] net520 ppwm_i.u_ppwm.u_pwm.counter\[4\]
+ _0476_ VPWR VGND sg13g2_nor4_1
XFILLER_36_842 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
X_2927_ net540 VGND VPWR _0118_ sdr_i.DP_3.matrix\[27\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2858_ net256 _0121_ VPWR VGND sg13g2_buf_1
X_1809_ VGND VPWR _0352_ _0353_ _0358_ _1231_ sg13g2_a21oi_1
Xhold220 _0238_ VPWR VGND net600 sg13g2_dlygate4sd3_1
X_2789_ VGND VPWR ppwm_i.u_ppwm.u_mem.bit_count\[4\] _1073_ _1076_ net330 sg13g2_a21oi_1
Xhold253 _0271_ VPWR VGND net633 sg13g2_dlygate4sd3_1
XFILLER_2_418 VPWR VGND sg13g2_decap_4
Xhold231 ppwm_i.u_ppwm.u_mem.memory\[45\] VPWR VGND net611 sg13g2_dlygate4sd3_1
Xhold242 _0236_ VPWR VGND net622 sg13g2_dlygate4sd3_1
XFILLER_49_26 VPWR VGND sg13g2_decap_8
XFILLER_46_1018 VPWR VGND sg13g2_decap_8
Xhold275 _0155_ VPWR VGND net655 sg13g2_dlygate4sd3_1
Xhold264 _0252_ VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold286 ppwm_i.u_ppwm.u_mem.memory\[14\] VPWR VGND net666 sg13g2_dlygate4sd3_1
Xhold297 ppwm_i.u_ppwm.u_mem.memory\[76\] VPWR VGND net677 sg13g2_dlygate4sd3_1
XFILLER_46_639 VPWR VGND sg13g2_decap_8
XFILLER_46_628 VPWR VGND sg13g2_fill_1
XFILLER_39_680 VPWR VGND sg13g2_fill_1
XFILLER_27_842 VPWR VGND sg13g2_decap_8
XFILLER_14_525 VPWR VGND sg13g2_fill_1
XFILLER_42_867 VPWR VGND sg13g2_decap_8
XFILLER_22_580 VPWR VGND sg13g2_fill_1
XFILLER_10_742 VPWR VGND sg13g2_fill_2
XFILLER_10_764 VPWR VGND sg13g2_decap_4
XFILLER_5_256 VPWR VGND sg13g2_decap_4
XFILLER_30_83 VPWR VGND sg13g2_decap_8
XFILLER_49_400 VPWR VGND sg13g2_decap_8
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_37_628 VPWR VGND sg13g2_decap_8
XFILLER_37_639 VPWR VGND sg13g2_fill_2
XFILLER_18_831 VPWR VGND sg13g2_decap_8
XFILLER_17_363 VPWR VGND sg13g2_decap_8
XFILLER_18_897 VPWR VGND sg13g2_decap_8
XFILLER_17_374 VPWR VGND sg13g2_fill_1
XFILLER_20_506 VPWR VGND sg13g2_fill_2
XFILLER_33_867 VPWR VGND sg13g2_decap_8
X_2712_ net413 VPWR _1035_ VGND net462 net700 sg13g2_o21ai_1
X_2643_ VGND VPWR net483 _1162_ _0261_ _1000_ sg13g2_a21oi_1
X_2574_ net433 VPWR _0966_ VGND net499 ppwm_i.u_ppwm.u_mem.memory\[12\] sg13g2_o21ai_1
X_3126_ net156 VGND VPWR net595 ppwm_i.u_ppwm.u_mem.memory\[102\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_28_628 VPWR VGND sg13g2_decap_4
X_3057_ net36 VGND VPWR net676 ppwm_i.u_ppwm.u_mem.memory\[33\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_35_17 VPWR VGND sg13g2_fill_2
XFILLER_35_28 VPWR VGND sg13g2_fill_2
XFILLER_36_661 VPWR VGND sg13g2_fill_1
XFILLER_24_834 VPWR VGND sg13g2_fill_2
X_2008_ _0467_ net719 net787 _0466_ VPWR VGND sg13g2_and3_2
XFILLER_36_683 VPWR VGND sg13g2_decap_8
XFILLER_11_506 VPWR VGND sg13g2_decap_8
XFILLER_24_889 VPWR VGND sg13g2_decap_8
XFILLER_11_517 VPWR VGND sg13g2_fill_2
XFILLER_3_749 VPWR VGND sg13g2_fill_2
XFILLER_2_215 VPWR VGND sg13g2_fill_2
XFILLER_2_237 VPWR VGND sg13g2_decap_8
Xfanout530 net534 net530 VPWR VGND sg13g2_buf_8
Xfanout541 net547 net541 VPWR VGND sg13g2_buf_8
XFILLER_19_606 VPWR VGND sg13g2_fill_2
XFILLER_19_617 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_14_322 VPWR VGND sg13g2_decap_8
XFILLER_15_878 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_fill_2
XFILLER_30_804 VPWR VGND sg13g2_decap_8
XFILLER_14_388 VPWR VGND sg13g2_fill_2
XFILLER_25_83 VPWR VGND sg13g2_fill_2
XFILLER_6_510 VPWR VGND sg13g2_decap_8
XFILLER_10_583 VPWR VGND sg13g2_fill_1
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
X_2290_ _0712_ _0711_ _0196_ VPWR VGND sg13g2_nor2b_1
XFILLER_1_281 VPWR VGND sg13g2_fill_2
XFILLER_49_296 VPWR VGND sg13g2_fill_2
XFILLER_37_458 VPWR VGND sg13g2_decap_8
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_18_650 VPWR VGND sg13g2_decap_8
XFILLER_45_480 VPWR VGND sg13g2_decap_8
XFILLER_17_193 VPWR VGND sg13g2_fill_2
XFILLER_36_1017 VPWR VGND sg13g2_decap_8
XFILLER_21_826 VPWR VGND sg13g2_decap_4
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_347 VPWR VGND sg13g2_decap_4
X_2626_ net425 VPWR _0992_ VGND net482 net643 sg13g2_o21ai_1
X_2557_ VGND VPWR net497 _1205_ _0218_ _0957_ sg13g2_a21oi_1
X_2488_ _0898_ _0877_ _0886_ VPWR VGND sg13g2_nand2_1
XFILLER_28_414 VPWR VGND sg13g2_fill_1
XFILLER_29_948 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
X_3109_ net143 VGND VPWR _0300_ ppwm_i.u_ppwm.u_mem.memory\[85\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_2
XFILLER_16_609 VPWR VGND sg13g2_decap_4
XFILLER_37_970 VPWR VGND sg13g2_decap_8
XFILLER_12_826 VPWR VGND sg13g2_decap_8
XFILLER_11_336 VPWR VGND sg13g2_decap_4
X_3005__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_11_85 VPWR VGND sg13g2_decap_4
XFILLER_3_557 VPWR VGND sg13g2_fill_1
XFILLER_47_712 VPWR VGND sg13g2_decap_4
Xfanout393 _0335_ net393 VPWR VGND sg13g2_buf_8
Xfanout371 net373 net371 VPWR VGND sg13g2_buf_8
Xfanout382 _0639_ net382 VPWR VGND sg13g2_buf_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_36_71 VPWR VGND sg13g2_decap_8
X_1790_ _0339_ net438 _1134_ net447 _1148_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_881 VPWR VGND sg13g2_decap_8
XFILLER_7_885 VPWR VGND sg13g2_decap_8
X_2411_ _0755_ _0778_ _0796_ _0815_ _0827_ VPWR VGND sg13g2_and4_1
X_2342_ _0762_ _0350_ _0666_ VPWR VGND sg13g2_nand2_1
XFILLER_42_1021 VPWR VGND sg13g2_decap_8
X_2273_ _0351_ _0692_ _0695_ _0696_ VPWR VGND sg13g2_nor3_1
XFILLER_38_723 VPWR VGND sg13g2_decap_8
X_3108__151 VPWR VGND net151 sg13g2_tiehi
X_3038__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_21_612 VPWR VGND sg13g2_decap_8
XFILLER_34_973 VPWR VGND sg13g2_decap_8
XFILLER_20_155 VPWR VGND sg13g2_decap_8
XFILLER_21_678 VPWR VGND sg13g2_fill_1
X_1988_ _0456_ net823 _0149_ VPWR VGND sg13g2_and2_1
X_2609_ VGND VPWR net487 _1179_ _0244_ _0983_ sg13g2_a21oi_1
XFILLER_0_527 VPWR VGND sg13g2_fill_2
XFILLER_44_704 VPWR VGND sg13g2_decap_8
XFILLER_44_737 VPWR VGND sg13g2_fill_2
XFILLER_16_439 VPWR VGND sg13g2_decap_8
XFILLER_43_258 VPWR VGND sg13g2_decap_4
XFILLER_12_612 VPWR VGND sg13g2_fill_1
XFILLER_11_111 VPWR VGND sg13g2_decap_4
XFILLER_12_634 VPWR VGND sg13g2_fill_1
XFILLER_40_976 VPWR VGND sg13g2_decap_8
XFILLER_8_627 VPWR VGND sg13g2_fill_2
XFILLER_7_104 VPWR VGND sg13g2_decap_8
XFILLER_4_811 VPWR VGND sg13g2_decap_8
XFILLER_22_62 VPWR VGND sg13g2_decap_4
XFILLER_4_888 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_35_704 VPWR VGND sg13g2_fill_2
XFILLER_16_962 VPWR VGND sg13g2_decap_8
X_2960_ net435 VGND VPWR net790 ppwm_i.u_ppwm.global_counter\[3\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_1911_ net276 net287 _0074_ VPWR VGND sg13g2_and2_1
X_2891_ net535 VGND VPWR _0082_ sdr_i.DP_1.matrix\[27\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_30_431 VPWR VGND sg13g2_decap_8
XFILLER_31_954 VPWR VGND sg13g2_decap_8
X_1842_ _0384_ net286 net221 VPWR VGND sg13g2_nand2_1
X_1773_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[13\] net445 _1340_ net513 sg13g2_a21oi_1
XFILLER_7_682 VPWR VGND sg13g2_fill_2
XFILLER_33_0 VPWR VGND sg13g2_decap_8
X_2325_ VGND VPWR net387 _0744_ _0746_ _0745_ sg13g2_a21oi_1
X_2256_ VGND VPWR net395 _1338_ _0680_ _0365_ sg13g2_a21oi_1
XFILLER_38_553 VPWR VGND sg13g2_fill_1
XFILLER_25_203 VPWR VGND sg13g2_decap_8
X_2187_ _0612_ VPWR _0613_ VGND _1215_ ppwm_i.u_ppwm.global_counter\[4\] sg13g2_o21ai_1
XFILLER_25_225 VPWR VGND sg13g2_decap_8
XFILLER_22_954 VPWR VGND sg13g2_decap_8
XFILLER_21_442 VPWR VGND sg13g2_decap_8
XFILLER_21_453 VPWR VGND sg13g2_fill_2
XFILLER_4_107 VPWR VGND sg13g2_decap_8
XFILLER_1_814 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_fill_2
XFILLER_17_715 VPWR VGND sg13g2_decap_8
XFILLER_17_726 VPWR VGND sg13g2_fill_2
XFILLER_29_597 VPWR VGND sg13g2_fill_1
XFILLER_44_556 VPWR VGND sg13g2_fill_1
XFILLER_17_51 VPWR VGND sg13g2_decap_8
XFILLER_17_62 VPWR VGND sg13g2_fill_1
XFILLER_17_748 VPWR VGND sg13g2_decap_8
XFILLER_40_773 VPWR VGND sg13g2_decap_8
XFILLER_13_976 VPWR VGND sg13g2_decap_8
XFILLER_33_50 VPWR VGND sg13g2_fill_2
XFILLER_33_61 VPWR VGND sg13g2_fill_2
XFILLER_9_947 VPWR VGND sg13g2_decap_8
XFILLER_33_72 VPWR VGND sg13g2_fill_2
X_3090_ net78 VGND VPWR _0281_ ppwm_i.u_ppwm.u_mem.memory\[66\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xhold2 sdr_i.mac2.products_ff\[136\] VPWR VGND net202 sg13g2_dlygate4sd3_1
X_2110_ VGND VPWR _0534_ _0537_ _0191_ net458 sg13g2_a21oi_1
X_2041_ _0487_ _1243_ net410 VPWR VGND sg13g2_nand2_1
XFILLER_48_884 VPWR VGND sg13g2_decap_8
XFILLER_47_372 VPWR VGND sg13g2_fill_1
XFILLER_35_523 VPWR VGND sg13g2_fill_2
X_2943_ net539 VGND VPWR _0134_ sdr_i.DP_4.matrix\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_15_280 VPWR VGND sg13g2_fill_2
X_3105__176 VPWR VGND net176 sg13g2_tiehi
X_2874_ net228 _0137_ VPWR VGND sg13g2_buf_1
X_1825_ net317 net414 _1249_ _0372_ VPWR VGND sg13g2_nand3_1
X_1756_ VPWR VGND _1195_ net512 net440 _1202_ _1323_ net445 sg13g2_a221oi_1
Xhold402 sdr_i.mac2.sum_lvl3_ff\[1\] VPWR VGND net782 sg13g2_dlygate4sd3_1
Xhold424 ppwm_i.u_ppwm.global_counter\[18\] VPWR VGND net804 sg13g2_dlygate4sd3_1
Xhold435 _0203_ VPWR VGND net815 sg13g2_dlygate4sd3_1
Xhold413 ppwm_i.u_ppwm.pwm_value\[9\] VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold457 _0211_ VPWR VGND net837 sg13g2_dlygate4sd3_1
Xhold446 ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] VPWR VGND net826 sg13g2_dlygate4sd3_1
X_1687_ _1258_ net787 VPWR VGND sg13g2_inv_2
X_2308_ VPWR VGND net376 _0727_ _0729_ net820 _0730_ net375 sg13g2_a221oi_1
XFILLER_39_862 VPWR VGND sg13g2_decap_8
XFILLER_38_372 VPWR VGND sg13g2_decap_8
X_2239_ net384 _0662_ _0663_ VPWR VGND sg13g2_nor2_1
XFILLER_38_383 VPWR VGND sg13g2_fill_2
XFILLER_14_718 VPWR VGND sg13g2_decap_8
XFILLER_10_902 VPWR VGND sg13g2_decap_8
XFILLER_16_1004 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_fill_2
XFILLER_21_250 VPWR VGND sg13g2_fill_1
XFILLER_10_979 VPWR VGND sg13g2_decap_8
XFILLER_5_405 VPWR VGND sg13g2_decap_8
XFILLER_1_655 VPWR VGND sg13g2_fill_2
XFILLER_1_688 VPWR VGND sg13g2_fill_1
XFILLER_48_169 VPWR VGND sg13g2_decap_4
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_17_501 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_fill_1
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_13_773 VPWR VGND sg13g2_fill_1
X_1610_ VPWR _1181_ net596 VGND sg13g2_inv_1
X_2590_ net432 VPWR _0974_ VGND net493 net623 sg13g2_o21ai_1
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_1541_ VPWR _1112_ net680 VGND sg13g2_inv_1
XFILLER_5_65 VPWR VGND sg13g2_fill_1
XFILLER_4_482 VPWR VGND sg13g2_fill_2
X_3211_ net542 VGND VPWR net756 sdr_i.mac2.sum_lvl1_ff\[17\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3142_ net193 VGND VPWR net696 ppwm_i.u_ppwm.u_mem.bit_count\[6\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_39_125 VPWR VGND sg13g2_fill_1
X_3073_ net145 VGND VPWR _0264_ ppwm_i.u_ppwm.u_mem.memory\[49\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_27_309 VPWR VGND sg13g2_decap_4
XFILLER_36_821 VPWR VGND sg13g2_decap_8
XFILLER_47_191 VPWR VGND sg13g2_fill_2
X_2024_ ppwm_i.u_ppwm.u_pwm.counter\[3\] ppwm_i.u_ppwm.u_pwm.counter\[2\] ppwm_i.u_ppwm.u_pwm.counter\[1\]
+ ppwm_i.u_ppwm.u_pwm.counter\[0\] _0475_ VPWR VGND sg13g2_nor4_1
XFILLER_36_898 VPWR VGND sg13g2_decap_8
XFILLER_35_375 VPWR VGND sg13g2_fill_2
X_2926_ net538 VGND VPWR _0117_ sdr_i.DP_3.matrix\[19\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2857_ net299 _0120_ VPWR VGND sg13g2_buf_1
XFILLER_31_592 VPWR VGND sg13g2_decap_4
X_1808_ _0355_ _0356_ _0354_ _0357_ VPWR VGND sg13g2_nand3_1
Xhold210 ppwm_i.u_ppwm.u_mem.memory\[61\] VPWR VGND net590 sg13g2_dlygate4sd3_1
X_2788_ _1067_ _1075_ _0331_ VPWR VGND sg13g2_nor2_1
X_1739_ _1303_ _1304_ net512 _1306_ VPWR VGND _1305_ sg13g2_nand4_1
Xhold232 ppwm_i.u_ppwm.u_mem.memory\[107\] VPWR VGND net612 sg13g2_dlygate4sd3_1
Xhold243 ppwm_i.u_ppwm.u_mem.memory\[20\] VPWR VGND net623 sg13g2_dlygate4sd3_1
Xhold221 sdr_i.mac2.sum_lvl3_ff\[3\] VPWR VGND net601 sg13g2_dlygate4sd3_1
Xhold287 ppwm_i.u_ppwm.u_mem.memory\[70\] VPWR VGND net667 sg13g2_dlygate4sd3_1
Xhold265 ppwm_i.u_ppwm.u_mem.memory\[104\] VPWR VGND net645 sg13g2_dlygate4sd3_1
Xhold254 ppwm_i.u_ppwm.u_mem.memory\[86\] VPWR VGND net634 sg13g2_dlygate4sd3_1
Xhold276 ppwm_i.u_ppwm.u_mem.memory\[4\] VPWR VGND net656 sg13g2_dlygate4sd3_1
Xhold298 ppwm_i.u_ppwm.u_mem.memory\[83\] VPWR VGND net678 sg13g2_dlygate4sd3_1
XFILLER_45_117 VPWR VGND sg13g2_decap_8
XFILLER_27_821 VPWR VGND sg13g2_decap_8
XFILLER_26_331 VPWR VGND sg13g2_decap_8
XFILLER_14_504 VPWR VGND sg13g2_fill_1
XFILLER_42_846 VPWR VGND sg13g2_decap_8
XFILLER_27_898 VPWR VGND sg13g2_decap_8
XFILLER_14_30 VPWR VGND sg13g2_fill_2
XFILLER_14_41 VPWR VGND sg13g2_fill_2
XFILLER_22_570 VPWR VGND sg13g2_decap_4
XFILLER_6_703 VPWR VGND sg13g2_decap_8
XFILLER_6_769 VPWR VGND sg13g2_decap_8
XFILLER_6_747 VPWR VGND sg13g2_decap_8
XFILLER_2_942 VPWR VGND sg13g2_decap_8
X_3015__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_17_331 VPWR VGND sg13g2_decap_8
XFILLER_45_651 VPWR VGND sg13g2_fill_1
XFILLER_18_876 VPWR VGND sg13g2_decap_8
XFILLER_33_846 VPWR VGND sg13g2_decap_8
XFILLER_32_345 VPWR VGND sg13g2_decap_8
X_2711_ VGND VPWR net469 _1128_ _0295_ _1034_ sg13g2_a21oi_1
XFILLER_9_596 VPWR VGND sg13g2_decap_8
X_2642_ net425 VPWR _1000_ VGND net483 net592 sg13g2_o21ai_1
X_2573_ VGND VPWR net499 _1197_ _0226_ _0965_ sg13g2_a21oi_1
X_3125_ net172 VGND VPWR net626 ppwm_i.u_ppwm.u_mem.memory\[101\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_3056_ net38 VGND VPWR net689 ppwm_i.u_ppwm.u_mem.memory\[32\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_24_813 VPWR VGND sg13g2_decap_8
X_2007_ _0159_ _1258_ _0466_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_161 VPWR VGND sg13g2_fill_2
XFILLER_24_868 VPWR VGND sg13g2_decap_8
XFILLER_13_1018 VPWR VGND sg13g2_decap_8
X_2909_ net535 VGND VPWR _0100_ sdr_i.DP_2.matrix\[27\] clknet_leaf_11_clk sg13g2_dfrbpq_1
Xfanout520 net565 net520 VPWR VGND sg13g2_buf_8
Xfanout531 net534 net531 VPWR VGND sg13g2_buf_8
Xfanout542 net543 net542 VPWR VGND sg13g2_buf_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_46_404 VPWR VGND sg13g2_fill_2
XFILLER_27_651 VPWR VGND sg13g2_decap_4
XFILLER_14_301 VPWR VGND sg13g2_decap_8
XFILLER_15_824 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_41_131 VPWR VGND sg13g2_decap_8
XFILLER_14_356 VPWR VGND sg13g2_decap_8
XFILLER_15_857 VPWR VGND sg13g2_decap_4
XFILLER_10_562 VPWR VGND sg13g2_decap_8
XFILLER_6_588 VPWR VGND sg13g2_decap_8
XFILLER_29_1025 VPWR VGND sg13g2_decap_4
XFILLER_37_7 VPWR VGND sg13g2_fill_2
XFILLER_2_44 VPWR VGND sg13g2_decap_8
XFILLER_49_275 VPWR VGND sg13g2_decap_8
XFILLER_38_938 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_fill_1
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XFILLER_33_621 VPWR VGND sg13g2_decap_8
XFILLER_32_153 VPWR VGND sg13g2_fill_1
X_2625_ VGND VPWR net482 _1171_ _0252_ _0991_ sg13g2_a21oi_1
X_2556_ net431 VPWR _0957_ VGND net497 net342 sg13g2_o21ai_1
X_2487_ _0876_ _0877_ _0886_ _0887_ _0897_ VPWR VGND sg13g2_and4_1
XFILLER_29_927 VPWR VGND sg13g2_decap_8
XFILLER_46_39 VPWR VGND sg13g2_decap_8
XFILLER_46_17 VPWR VGND sg13g2_decap_4
X_3108_ net151 VGND VPWR net359 ppwm_i.u_ppwm.u_mem.memory\[84\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
X_3039_ net71 VGND VPWR _0230_ ppwm_i.u_ppwm.u_mem.memory\[15\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_24_610 VPWR VGND sg13g2_fill_2
XFILLER_36_481 VPWR VGND sg13g2_fill_2
XFILLER_24_643 VPWR VGND sg13g2_decap_4
XFILLER_23_142 VPWR VGND sg13g2_fill_1
XFILLER_24_676 VPWR VGND sg13g2_fill_2
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_11_75 VPWR VGND sg13g2_fill_2
Xfanout372 net373 net372 VPWR VGND sg13g2_buf_1
Xfanout383 _0639_ net383 VPWR VGND sg13g2_buf_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
Xfanout394 _1338_ net394 VPWR VGND sg13g2_buf_8
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_15_632 VPWR VGND sg13g2_decap_8
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_42_484 VPWR VGND sg13g2_fill_1
XFILLER_15_698 VPWR VGND sg13g2_decap_8
XFILLER_30_624 VPWR VGND sg13g2_fill_1
X_2999__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_7_864 VPWR VGND sg13g2_decap_8
X_2410_ _0825_ _0826_ _0202_ VPWR VGND sg13g2_nor2_1
X_2341_ _0691_ VPWR _0761_ VGND _0694_ _0740_ sg13g2_o21ai_1
XFILLER_42_1000 VPWR VGND sg13g2_decap_8
X_2272_ VPWR _0695_ _0694_ VGND sg13g2_inv_1
XFILLER_37_234 VPWR VGND sg13g2_fill_2
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_34_952 VPWR VGND sg13g2_decap_8
X_3053__44 VPWR VGND net44 sg13g2_tiehi
X_1987_ ppwm_i.u_ppwm.global_counter\[0\] net326 net822 _0457_ VPWR VGND sg13g2_a21o_1
XFILLER_9_190 VPWR VGND sg13g2_decap_8
X_2608_ net430 VPWR _0983_ VGND net487 ppwm_i.u_ppwm.u_mem.memory\[29\] sg13g2_o21ai_1
X_2539_ _0944_ VPWR _0945_ VGND net381 _0840_ sg13g2_o21ai_1
XFILLER_16_407 VPWR VGND sg13g2_fill_2
XFILLER_16_429 VPWR VGND sg13g2_decap_4
XFILLER_25_985 VPWR VGND sg13g2_decap_8
XFILLER_40_955 VPWR VGND sg13g2_decap_8
XFILLER_12_657 VPWR VGND sg13g2_fill_1
XFILLER_8_639 VPWR VGND sg13g2_decap_4
XFILLER_7_138 VPWR VGND sg13g2_decap_4
XFILLER_22_41 VPWR VGND sg13g2_decap_8
XFILLER_4_867 VPWR VGND sg13g2_decap_8
XFILLER_3_366 VPWR VGND sg13g2_fill_2
XFILLER_3_355 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_fill_2
XFILLER_47_521 VPWR VGND sg13g2_fill_2
XFILLER_19_256 VPWR VGND sg13g2_fill_2
XFILLER_47_93 VPWR VGND sg13g2_decap_8
XFILLER_16_941 VPWR VGND sg13g2_decap_8
XFILLER_15_462 VPWR VGND sg13g2_decap_4
XFILLER_43_782 VPWR VGND sg13g2_decap_8
XFILLER_42_281 VPWR VGND sg13g2_decap_8
X_1910_ _0031_ _0412_ _0415_ VPWR VGND sg13g2_xnor2_1
X_2890_ net525 VGND VPWR _0081_ sdr_i.DP_1.matrix\[19\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_31_933 VPWR VGND sg13g2_decap_8
X_1841_ VGND VPWR _1248_ net15 _0383_ _0380_ sg13g2_a21oi_2
X_1772_ _1339_ _1325_ net394 VPWR VGND sg13g2_nand2_1
X_2324_ net387 _0722_ _0745_ VPWR VGND sg13g2_nor2_1
X_2255_ net385 VPWR _0679_ VGND net401 net397 sg13g2_o21ai_1
XFILLER_38_510 VPWR VGND sg13g2_fill_1
X_2186_ _0612_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _1264_ VPWR VGND sg13g2_nand2_1
XFILLER_19_790 VPWR VGND sg13g2_fill_1
XFILLER_26_749 VPWR VGND sg13g2_fill_2
XFILLER_41_719 VPWR VGND sg13g2_decap_8
XFILLER_40_229 VPWR VGND sg13g2_decap_8
XFILLER_22_933 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_325 VPWR VGND sg13g2_fill_1
XFILLER_0_314 VPWR VGND sg13g2_decap_8
XFILLER_0_358 VPWR VGND sg13g2_decap_8
XFILLER_0_369 VPWR VGND sg13g2_fill_1
XFILLER_17_30 VPWR VGND sg13g2_decap_8
XFILLER_16_248 VPWR VGND sg13g2_decap_8
XFILLER_9_926 VPWR VGND sg13g2_decap_8
XFILLER_13_955 VPWR VGND sg13g2_decap_8
XFILLER_32_1010 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_decap_8
XFILLER_4_631 VPWR VGND sg13g2_decap_4
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_39_307 VPWR VGND sg13g2_decap_8
XFILLER_0_892 VPWR VGND sg13g2_decap_8
Xhold3 sdr_i.mac1.sum_lvl1_ff\[32\] VPWR VGND net203 sg13g2_dlygate4sd3_1
XFILLER_48_863 VPWR VGND sg13g2_decap_8
X_2040_ net456 net797 _0172_ VPWR VGND sg13g2_nor2_1
XFILLER_35_513 VPWR VGND sg13g2_decap_4
XFILLER_23_708 VPWR VGND sg13g2_fill_2
XFILLER_23_719 VPWR VGND sg13g2_fill_1
XFILLER_35_579 VPWR VGND sg13g2_decap_8
X_2942_ net546 VGND VPWR _0133_ sdr_i.DP_4.matrix\[10\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2873_ net301 _0136_ VPWR VGND sg13g2_buf_1
XFILLER_30_251 VPWR VGND sg13g2_decap_8
XFILLER_30_273 VPWR VGND sg13g2_fill_2
X_1824_ _0371_ VPWR _0002_ VGND _1277_ _0368_ sg13g2_o21ai_1
X_1755_ _1322_ net448 _1209_ net453 _1188_ VPWR VGND sg13g2_a22oi_1
Xhold425 ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] VPWR VGND net805 sg13g2_dlygate4sd3_1
Xhold403 _0008_ VPWR VGND net783 sg13g2_dlygate4sd3_1
Xhold436 ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] VPWR VGND net816 sg13g2_dlygate4sd3_1
Xhold414 ppwm_i.u_ppwm.pwm_value\[2\] VPWR VGND net794 sg13g2_dlygate4sd3_1
Xhold447 ppwm_i.u_ppwm.pc\[2\] VPWR VGND net827 sg13g2_dlygate4sd3_1
X_1686_ VPWR _1257_ ppwm_i.u_ppwm.global_counter\[12\] VGND sg13g2_inv_1
Xhold458 ppwm_i.u_ppwm.pwm_value\[4\] VPWR VGND net838 sg13g2_dlygate4sd3_1
X_2307_ _0728_ VPWR _0729_ VGND _1265_ _1295_ sg13g2_o21ai_1
XFILLER_39_841 VPWR VGND sg13g2_decap_8
X_2238_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] net505 net399 _0662_ VPWR VGND sg13g2_mux2_1
X_2169_ _0595_ _1226_ ppwm_i.u_ppwm.global_counter\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_41_505 VPWR VGND sg13g2_decap_8
XFILLER_14_708 VPWR VGND sg13g2_fill_2
XFILLER_26_557 VPWR VGND sg13g2_decap_8
XFILLER_26_579 VPWR VGND sg13g2_decap_8
XFILLER_10_958 VPWR VGND sg13g2_decap_8
XFILLER_5_428 VPWR VGND sg13g2_fill_1
XFILLER_1_601 VPWR VGND sg13g2_decap_8
XFILLER_0_144 VPWR VGND sg13g2_decap_4
XFILLER_49_649 VPWR VGND sg13g2_decap_8
XFILLER_0_177 VPWR VGND sg13g2_decap_4
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_44_321 VPWR VGND sg13g2_decap_4
XFILLER_17_535 VPWR VGND sg13g2_decap_8
XFILLER_45_877 VPWR VGND sg13g2_decap_8
XFILLER_32_505 VPWR VGND sg13g2_fill_2
XFILLER_44_72 VPWR VGND sg13g2_fill_2
XFILLER_25_590 VPWR VGND sg13g2_decap_8
XFILLER_8_211 VPWR VGND sg13g2_fill_1
XFILLER_9_712 VPWR VGND sg13g2_decap_4
XFILLER_13_785 VPWR VGND sg13g2_decap_8
XFILLER_9_778 VPWR VGND sg13g2_fill_1
XFILLER_8_277 VPWR VGND sg13g2_fill_1
XFILLER_5_951 VPWR VGND sg13g2_decap_8
X_1540_ VPWR _1111_ net773 VGND sg13g2_inv_1
X_3210_ net542 VGND VPWR net266 sdr_i.mac2.sum_lvl1_ff\[16\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3141_ net84 VGND VPWR net332 ppwm_i.u_ppwm.u_mem.bit_count\[5\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_39_104 VPWR VGND sg13g2_decap_4
X_3072_ net149 VGND VPWR _0263_ ppwm_i.u_ppwm.u_mem.memory\[48\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_2
XFILLER_36_800 VPWR VGND sg13g2_decap_8
X_2023_ _0167_ net328 _0473_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_1016 VPWR VGND sg13g2_decap_8
XFILLER_36_877 VPWR VGND sg13g2_decap_8
XFILLER_23_538 VPWR VGND sg13g2_fill_2
XFILLER_35_387 VPWR VGND sg13g2_fill_2
X_2925_ net538 VGND VPWR _0116_ sdr_i.DP_3.matrix\[18\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_31_560 VPWR VGND sg13g2_decap_4
X_2856_ net236 _0119_ VPWR VGND sg13g2_buf_1
X_1807_ _0356_ net449 ppwm_i.u_ppwm.u_mem.memory\[58\] net451 ppwm_i.u_ppwm.u_mem.memory\[79\]
+ VPWR VGND sg13g2_a22oi_1
Xhold200 ppwm_i.u_ppwm.u_pwm.cmp_value\[7\] VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold211 _0275_ VPWR VGND net591 sg13g2_dlygate4sd3_1
X_2787_ _1075_ net748 _1073_ VPWR VGND sg13g2_xnor2_1
Xhold233 _0321_ VPWR VGND net613 sg13g2_dlygate4sd3_1
X_1738_ _1305_ net446 _1170_ net454 _1156_ VPWR VGND sg13g2_a22oi_1
Xhold222 _0417_ VPWR VGND net602 sg13g2_dlygate4sd3_1
Xhold244 _0234_ VPWR VGND net624 sg13g2_dlygate4sd3_1
Xhold277 ppwm_i.u_ppwm.u_mem.memory\[52\] VPWR VGND net657 sg13g2_dlygate4sd3_1
Xhold255 ppwm_i.u_ppwm.u_mem.memory\[96\] VPWR VGND net635 sg13g2_dlygate4sd3_1
Xhold266 ppwm_i.u_ppwm.u_mem.memory\[16\] VPWR VGND net646 sg13g2_dlygate4sd3_1
X_1669_ VPWR _1240_ ppwm_i.u_ppwm.u_pwm.counter\[1\] VGND sg13g2_inv_1
Xhold288 _0285_ VPWR VGND net668 sg13g2_dlygate4sd3_1
Xhold299 _0297_ VPWR VGND net679 sg13g2_dlygate4sd3_1
XFILLER_26_365 VPWR VGND sg13g2_fill_1
XFILLER_27_877 VPWR VGND sg13g2_decap_8
XFILLER_38_192 VPWR VGND sg13g2_decap_8
XFILLER_42_825 VPWR VGND sg13g2_decap_8
X_3086__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_49_457 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_decap_4
XFILLER_39_83 VPWR VGND sg13g2_decap_8
XFILLER_49_468 VPWR VGND sg13g2_fill_1
XFILLER_45_685 VPWR VGND sg13g2_decap_8
XFILLER_33_825 VPWR VGND sg13g2_decap_8
XFILLER_9_531 VPWR VGND sg13g2_decap_4
X_2710_ net412 VPWR _1034_ VGND net469 net706 sg13g2_o21ai_1
XFILLER_9_575 VPWR VGND sg13g2_decap_8
X_2641_ VGND VPWR net483 _1163_ _0260_ _0999_ sg13g2_a21oi_1
X_2572_ net433 VPWR _0965_ VGND net498 net647 sg13g2_o21ai_1
X_3124_ net187 VGND VPWR _0315_ ppwm_i.u_ppwm.u_mem.memory\[100\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
X_3055_ net40 VGND VPWR net346 ppwm_i.u_ppwm.u_mem.memory\[31\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_24_803 VPWR VGND sg13g2_fill_1
X_2006_ _0465_ net557 _0158_ VPWR VGND sg13g2_xor2_1
XFILLER_36_641 VPWR VGND sg13g2_fill_1
XFILLER_36_652 VPWR VGND sg13g2_fill_2
XFILLER_24_847 VPWR VGND sg13g2_decap_8
XFILLER_23_324 VPWR VGND sg13g2_decap_8
XFILLER_23_357 VPWR VGND sg13g2_fill_2
X_2908_ net527 VGND VPWR _0099_ sdr_i.DP_2.matrix\[19\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_32_891 VPWR VGND sg13g2_decap_8
X_2839_ net312 _0102_ VPWR VGND sg13g2_buf_1
XFILLER_4_8 VPWR VGND sg13g2_decap_8
Xfanout532 net534 net532 VPWR VGND sg13g2_buf_8
Xfanout521 net524 net521 VPWR VGND sg13g2_buf_8
Xfanout510 net513 net510 VPWR VGND sg13g2_buf_8
Xfanout543 net547 net543 VPWR VGND sg13g2_buf_2
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_46_416 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_38_clk clknet_3_4__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_42_600 VPWR VGND sg13g2_decap_8
XFILLER_42_677 VPWR VGND sg13g2_decap_8
XFILLER_30_839 VPWR VGND sg13g2_decap_8
XFILLER_41_176 VPWR VGND sg13g2_fill_1
XFILLER_23_880 VPWR VGND sg13g2_decap_8
XFILLER_10_541 VPWR VGND sg13g2_decap_8
XFILLER_22_390 VPWR VGND sg13g2_fill_1
XFILLER_41_62 VPWR VGND sg13g2_decap_8
XFILLER_6_523 VPWR VGND sg13g2_fill_1
XFILLER_6_567 VPWR VGND sg13g2_fill_2
XFILLER_29_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_1_283 VPWR VGND sg13g2_fill_1
XFILLER_49_254 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_4
XFILLER_38_917 VPWR VGND sg13g2_decap_8
XFILLER_37_427 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_46_983 VPWR VGND sg13g2_decap_8
XFILLER_33_600 VPWR VGND sg13g2_fill_2
XFILLER_9_350 VPWR VGND sg13g2_decap_8
X_2624_ net425 VPWR _0991_ VGND net482 net606 sg13g2_o21ai_1
X_2555_ VGND VPWR net489 _1206_ _0217_ _0956_ sg13g2_a21oi_1
X_2486_ _0896_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] net393 VPWR VGND sg13g2_xnor2_1
XFILLER_29_906 VPWR VGND sg13g2_decap_8
X_3107_ net160 VGND VPWR _0298_ ppwm_i.u_ppwm.u_mem.memory\[83\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_3038_ net73 VGND VPWR net589 ppwm_i.u_ppwm.u_mem.memory\[14\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_11_305 VPWR VGND sg13g2_decap_4
XFILLER_23_154 VPWR VGND sg13g2_fill_1
XFILLER_11_54 VPWR VGND sg13g2_decap_8
Xfanout373 _0683_ net373 VPWR VGND sg13g2_buf_8
Xfanout384 net385 net384 VPWR VGND sg13g2_buf_8
XFILLER_46_213 VPWR VGND sg13g2_fill_1
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
Xfanout395 _1325_ net395 VPWR VGND sg13g2_buf_8
XFILLER_15_600 VPWR VGND sg13g2_decap_8
XFILLER_15_611 VPWR VGND sg13g2_fill_1
XFILLER_34_419 VPWR VGND sg13g2_decap_8
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_42_463 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_fill_2
XFILLER_7_843 VPWR VGND sg13g2_decap_8
XFILLER_10_393 VPWR VGND sg13g2_decap_8
XFILLER_6_364 VPWR VGND sg13g2_decap_4
X_2340_ VGND VPWR _0755_ _0758_ _0760_ _0759_ sg13g2_a21oi_1
XFILLER_2_592 VPWR VGND sg13g2_decap_8
X_2271_ _0693_ VPWR _0694_ VGND _1229_ net401 sg13g2_o21ai_1
XFILLER_46_780 VPWR VGND sg13g2_decap_8
XFILLER_19_972 VPWR VGND sg13g2_decap_8
XFILLER_37_279 VPWR VGND sg13g2_decap_8
XFILLER_33_430 VPWR VGND sg13g2_decap_4
XFILLER_34_931 VPWR VGND sg13g2_decap_8
XFILLER_33_474 VPWR VGND sg13g2_decap_8
XFILLER_21_658 VPWR VGND sg13g2_decap_8
X_3004__140 VPWR VGND net140 sg13g2_tiehi
X_1986_ net822 ppwm_i.u_ppwm.global_counter\[0\] net326 _0456_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_2607_ VGND VPWR net492 _1180_ _0243_ _0982_ sg13g2_a21oi_1
X_2538_ VGND VPWR _1221_ net381 _0944_ _0672_ sg13g2_a21oi_1
XFILLER_0_529 VPWR VGND sg13g2_fill_1
X_2469_ _0879_ _0880_ net378 _0881_ VPWR VGND sg13g2_nand3_1
XFILLER_24_430 VPWR VGND sg13g2_decap_4
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_25_964 VPWR VGND sg13g2_decap_8
XFILLER_40_934 VPWR VGND sg13g2_decap_8
XFILLER_24_474 VPWR VGND sg13g2_decap_8
XFILLER_22_97 VPWR VGND sg13g2_fill_2
XFILLER_4_846 VPWR VGND sg13g2_decap_8
XFILLER_26_1018 VPWR VGND sg13g2_decap_8
XFILLER_19_224 VPWR VGND sg13g2_decap_4
XFILLER_35_728 VPWR VGND sg13g2_fill_1
XFILLER_16_920 VPWR VGND sg13g2_decap_8
XFILLER_34_227 VPWR VGND sg13g2_decap_8
XFILLER_43_761 VPWR VGND sg13g2_decap_8
XFILLER_31_912 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_16_997 VPWR VGND sg13g2_decap_8
X_1840_ net14 net548 _0382_ _0383_ VPWR VGND sg13g2_and3_2
XFILLER_30_477 VPWR VGND sg13g2_decap_8
XFILLER_31_989 VPWR VGND sg13g2_decap_8
XFILLER_8_99 VPWR VGND sg13g2_decap_8
X_1771_ _1331_ net509 _1337_ _1338_ VPWR VGND sg13g2_a21o_2
XFILLER_7_684 VPWR VGND sg13g2_fill_1
X_2323_ _0744_ _0743_ VPWR VGND sg13g2_inv_2
X_2254_ _0678_ _1229_ _1311_ VPWR VGND sg13g2_nand2_1
X_2185_ VPWR VGND _1217_ _0610_ ppwm_i.u_ppwm.global_counter\[2\] _1216_ _0611_ ppwm_i.u_ppwm.global_counter\[3\]
+ sg13g2_a221oi_1
XFILLER_38_566 VPWR VGND sg13g2_decap_8
XFILLER_41_709 VPWR VGND sg13g2_decap_4
XFILLER_22_912 VPWR VGND sg13g2_decap_8
XFILLER_40_219 VPWR VGND sg13g2_decap_4
XFILLER_21_400 VPWR VGND sg13g2_fill_2
XFILLER_33_271 VPWR VGND sg13g2_decap_4
XFILLER_22_989 VPWR VGND sg13g2_decap_8
X_1969_ _0446_ net304 net226 VPWR VGND sg13g2_nand2_1
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_337 VPWR VGND sg13g2_decap_8
XFILLER_1_849 VPWR VGND sg13g2_decap_8
XFILLER_29_544 VPWR VGND sg13g2_fill_2
XFILLER_29_588 VPWR VGND sg13g2_decap_8
XFILLER_16_227 VPWR VGND sg13g2_decap_8
XFILLER_32_709 VPWR VGND sg13g2_fill_1
XFILLER_13_934 VPWR VGND sg13g2_decap_8
XFILLER_9_905 VPWR VGND sg13g2_decap_8
XFILLER_33_52 VPWR VGND sg13g2_fill_1
XFILLER_33_74 VPWR VGND sg13g2_fill_1
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_0_871 VPWR VGND sg13g2_decap_8
Xhold4 sdr_i.mac2.sum_lvl1_ff\[33\] VPWR VGND net204 sg13g2_dlygate4sd3_1
XFILLER_48_842 VPWR VGND sg13g2_decap_8
XFILLER_47_396 VPWR VGND sg13g2_decap_4
XFILLER_35_525 VPWR VGND sg13g2_fill_1
XFILLER_35_558 VPWR VGND sg13g2_fill_1
X_2941_ net546 VGND VPWR _0132_ sdr_i.DP_4.matrix\[9\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2872_ net234 _0135_ VPWR VGND sg13g2_buf_1
XFILLER_31_786 VPWR VGND sg13g2_decap_8
X_1823_ _0369_ VPWR _0371_ VGND net759 net317 sg13g2_o21ai_1
XFILLER_8_993 VPWR VGND sg13g2_decap_8
X_1754_ VPWR VGND _1174_ _1320_ net444 _1160_ _1321_ net453 sg13g2_a221oi_1
Xhold426 ppwm_i.u_ppwm.global_counter\[4\] VPWR VGND net806 sg13g2_dlygate4sd3_1
Xhold415 _0170_ VPWR VGND net795 sg13g2_dlygate4sd3_1
Xhold404 ppwm_i.u_ppwm.u_pwm.counter\[2\] VPWR VGND net784 sg13g2_dlygate4sd3_1
Xhold437 ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] VPWR VGND net817 sg13g2_dlygate4sd3_1
Xhold459 ppwm_i.u_ppwm.u_pwm.counter\[8\] VPWR VGND net839 sg13g2_dlygate4sd3_1
Xhold448 ppwm_i.u_ppwm.pwm_value\[5\] VPWR VGND net828 sg13g2_dlygate4sd3_1
X_3424_ net549 net11 VPWR VGND sg13g2_buf_1
X_1685_ _1256_ net776 VPWR VGND sg13g2_inv_2
XFILLER_39_820 VPWR VGND sg13g2_decap_8
X_2306_ _0728_ ppwm_i.u_ppwm.global_counter\[12\] net401 VPWR VGND sg13g2_nand2_1
X_2237_ VGND VPWR ppwm_i.u_ppwm.pwm_value\[4\] net399 _0661_ _0660_ sg13g2_a21oi_1
XFILLER_39_897 VPWR VGND sg13g2_decap_8
X_2168_ VPWR VGND _0592_ _0593_ _0588_ net506 _0594_ _1264_ sg13g2_a221oi_1
X_2099_ net768 VPWR _0528_ VGND _0518_ _0527_ sg13g2_o21ai_1
XFILLER_10_937 VPWR VGND sg13g2_decap_8
XFILLER_22_764 VPWR VGND sg13g2_decap_8
XFILLER_6_919 VPWR VGND sg13g2_decap_8
XFILLER_21_274 VPWR VGND sg13g2_fill_2
XFILLER_0_123 VPWR VGND sg13g2_decap_8
XFILLER_1_657 VPWR VGND sg13g2_fill_1
XFILLER_49_628 VPWR VGND sg13g2_decap_8
XFILLER_45_856 VPWR VGND sg13g2_decap_8
X_3128__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_28_96 VPWR VGND sg13g2_decap_8
XFILLER_44_355 VPWR VGND sg13g2_decap_8
XFILLER_32_528 VPWR VGND sg13g2_fill_1
XFILLER_13_731 VPWR VGND sg13g2_decap_4
XFILLER_13_753 VPWR VGND sg13g2_decap_4
XFILLER_40_550 VPWR VGND sg13g2_decap_8
XFILLER_8_201 VPWR VGND sg13g2_fill_1
XFILLER_9_724 VPWR VGND sg13g2_decap_4
XFILLER_9_735 VPWR VGND sg13g2_decap_4
XFILLER_40_594 VPWR VGND sg13g2_decap_8
XFILLER_8_234 VPWR VGND sg13g2_fill_2
XFILLER_12_296 VPWR VGND sg13g2_decap_4
XFILLER_5_930 VPWR VGND sg13g2_decap_8
XFILLER_5_34 VPWR VGND sg13g2_decap_8
XFILLER_5_78 VPWR VGND sg13g2_decap_4
XFILLER_4_495 VPWR VGND sg13g2_decap_8
XFILLER_4_484 VPWR VGND sg13g2_fill_1
X_3140_ net147 VGND VPWR _0331_ ppwm_i.u_ppwm.u_mem.bit_count\[4\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_3071_ net154 VGND VPWR net571 ppwm_i.u_ppwm.u_mem.memory\[47\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2022_ _0473_ _0474_ _0166_ VPWR VGND sg13g2_and2_1
XFILLER_35_300 VPWR VGND sg13g2_decap_8
XFILLER_47_193 VPWR VGND sg13g2_fill_1
XFILLER_36_856 VPWR VGND sg13g2_decap_8
XFILLER_35_377 VPWR VGND sg13g2_fill_1
X_2924_ net546 VGND VPWR _0115_ sdr_i.DP_3.matrix\[10\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2855_ net278 _0118_ VPWR VGND sg13g2_buf_1
X_1806_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[65\] net443 _0355_ net511 sg13g2_a21oi_1
Xhold201 _0175_ VPWR VGND net581 sg13g2_dlygate4sd3_1
X_2786_ _1067_ _1073_ net662 _0330_ VPWR VGND sg13g2_nor3_1
Xhold212 ppwm_i.u_ppwm.u_mem.memory\[46\] VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold234 ppwm_i.u_ppwm.u_mem.memory\[90\] VPWR VGND net614 sg13g2_dlygate4sd3_1
X_1737_ _1304_ _1163_ net441 VPWR VGND sg13g2_nand2_1
Xhold223 _0006_ VPWR VGND net603 sg13g2_dlygate4sd3_1
X_1668_ VPWR _1239_ net520 VGND sg13g2_inv_1
Xhold278 _0267_ VPWR VGND net658 sg13g2_dlygate4sd3_1
Xhold256 ppwm_i.u_ppwm.u_mem.memory\[29\] VPWR VGND net636 sg13g2_dlygate4sd3_1
Xhold245 ppwm_i.u_ppwm.u_mem.memory\[102\] VPWR VGND net625 sg13g2_dlygate4sd3_1
Xhold267 ppwm_i.u_ppwm.u_mem.memory\[11\] VPWR VGND net647 sg13g2_dlygate4sd3_1
Xhold289 ppwm_i.u_ppwm.u_mem.memory\[54\] VPWR VGND net669 sg13g2_dlygate4sd3_1
X_1599_ VPWR _1170_ net698 VGND sg13g2_inv_1
XFILLER_46_609 VPWR VGND sg13g2_fill_2
XFILLER_22_1010 VPWR VGND sg13g2_decap_8
X_2986__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_42_804 VPWR VGND sg13g2_decap_8
XFILLER_26_344 VPWR VGND sg13g2_decap_8
XFILLER_27_856 VPWR VGND sg13g2_decap_8
XFILLER_14_539 VPWR VGND sg13g2_decap_4
XFILLER_26_377 VPWR VGND sg13g2_decap_4
XFILLER_41_325 VPWR VGND sg13g2_decap_4
XFILLER_26_399 VPWR VGND sg13g2_fill_1
XFILLER_41_369 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_fill_1
XFILLER_14_98 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_97 VPWR VGND sg13g2_decap_8
XFILLER_49_414 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_39_62 VPWR VGND sg13g2_fill_1
XFILLER_18_801 VPWR VGND sg13g2_decap_8
XFILLER_29_171 VPWR VGND sg13g2_decap_8
XFILLER_45_642 VPWR VGND sg13g2_fill_2
XFILLER_18_856 VPWR VGND sg13g2_decap_8
XFILLER_33_804 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_8
XFILLER_32_325 VPWR VGND sg13g2_fill_1
XFILLER_41_892 VPWR VGND sg13g2_decap_8
XFILLER_13_583 VPWR VGND sg13g2_fill_2
X_2640_ net426 VPWR _0999_ VGND net483 ppwm_i.u_ppwm.u_mem.memory\[45\] sg13g2_o21ai_1
X_2571_ VGND VPWR net498 _1198_ _0225_ _0964_ sg13g2_a21oi_1
XFILLER_5_771 VPWR VGND sg13g2_decap_8
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_281 VPWR VGND sg13g2_decap_8
X_3123_ net33 VGND VPWR net363 ppwm_i.u_ppwm.u_mem.memory\[99\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_28_609 VPWR VGND sg13g2_decap_4
X_3054_ net42 VGND VPWR net361 ppwm_i.u_ppwm.u_mem.memory\[30\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_36_620 VPWR VGND sg13g2_fill_1
X_2005_ net557 _0465_ _0466_ VPWR VGND sg13g2_and2_1
XFILLER_35_163 VPWR VGND sg13g2_fill_1
XFILLER_35_185 VPWR VGND sg13g2_decap_8
XFILLER_32_870 VPWR VGND sg13g2_decap_8
X_2907_ net525 VGND VPWR _0098_ sdr_i.DP_2.matrix\[18\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2838_ net226 _0101_ VPWR VGND sg13g2_buf_1
X_2769_ VGND VPWR net472 _1099_ _0324_ _1063_ sg13g2_a21oi_1
Xfanout533 net534 net533 VPWR VGND sg13g2_buf_8
Xfanout511 net513 net511 VPWR VGND sg13g2_buf_2
Xfanout522 net524 net522 VPWR VGND sg13g2_buf_8
Xfanout500 net501 net500 VPWR VGND sg13g2_buf_8
X_3014__120 VPWR VGND net120 sg13g2_tiehi
Xfanout544 net546 net544 VPWR VGND sg13g2_buf_8
XFILLER_18_119 VPWR VGND sg13g2_decap_8
XFILLER_26_130 VPWR VGND sg13g2_decap_8
XFILLER_27_631 VPWR VGND sg13g2_decap_8
XFILLER_42_612 VPWR VGND sg13g2_decap_8
XFILLER_42_623 VPWR VGND sg13g2_fill_1
XFILLER_42_667 VPWR VGND sg13g2_fill_1
XFILLER_30_818 VPWR VGND sg13g2_decap_8
XFILLER_41_30 VPWR VGND sg13g2_decap_8
XFILLER_6_557 VPWR VGND sg13g2_fill_1
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_49_233 VPWR VGND sg13g2_decap_8
XFILLER_2_13 VPWR VGND sg13g2_decap_8
XFILLER_37_406 VPWR VGND sg13g2_decap_8
XFILLER_46_962 VPWR VGND sg13g2_decap_8
XFILLER_17_130 VPWR VGND sg13g2_fill_2
XFILLER_18_664 VPWR VGND sg13g2_decap_8
XFILLER_33_656 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_9_340 VPWR VGND sg13g2_decap_4
XFILLER_13_380 VPWR VGND sg13g2_decap_8
XFILLER_9_373 VPWR VGND sg13g2_decap_8
X_2623_ VGND VPWR net487 _1172_ _0251_ _0990_ sg13g2_a21oi_1
X_2554_ net431 VPWR _0956_ VGND net489 net337 sg13g2_o21ai_1
X_2485_ _1215_ net393 _0895_ VPWR VGND sg13g2_nor2_1
X_3106_ net168 VGND VPWR net679 ppwm_i.u_ppwm.u_mem.memory\[82\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_3037_ net75 VGND VPWR _0228_ ppwm_i.u_ppwm.u_mem.memory\[13\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
XFILLER_37_984 VPWR VGND sg13g2_decap_8
XFILLER_36_483 VPWR VGND sg13g2_fill_1
XFILLER_20_884 VPWR VGND sg13g2_decap_8
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
Xfanout374 _0860_ net374 VPWR VGND sg13g2_buf_8
XFILLER_19_439 VPWR VGND sg13g2_fill_1
Xfanout396 _1310_ net396 VPWR VGND sg13g2_buf_8
Xfanout385 _0349_ net385 VPWR VGND sg13g2_buf_8
XFILLER_46_225 VPWR VGND sg13g2_decap_8
XFILLER_27_472 VPWR VGND sg13g2_decap_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_42_431 VPWR VGND sg13g2_fill_1
XFILLER_27_483 VPWR VGND sg13g2_fill_1
XFILLER_36_85 VPWR VGND sg13g2_decap_4
XFILLER_42_453 VPWR VGND sg13g2_fill_1
XFILLER_42_442 VPWR VGND sg13g2_fill_2
XFILLER_14_155 VPWR VGND sg13g2_decap_8
XFILLER_14_177 VPWR VGND sg13g2_decap_8
XFILLER_7_822 VPWR VGND sg13g2_decap_8
XFILLER_7_811 VPWR VGND sg13g2_fill_2
XFILLER_11_895 VPWR VGND sg13g2_decap_8
XFILLER_10_372 VPWR VGND sg13g2_decap_8
XFILLER_6_332 VPWR VGND sg13g2_fill_1
XFILLER_7_899 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_fill_2
X_2270_ _0693_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] net401 VPWR VGND sg13g2_nand2_1
XFILLER_38_737 VPWR VGND sg13g2_decap_8
XFILLER_19_951 VPWR VGND sg13g2_decap_8
XFILLER_37_236 VPWR VGND sg13g2_fill_1
XFILLER_18_461 VPWR VGND sg13g2_fill_1
XFILLER_34_910 VPWR VGND sg13g2_decap_8
XFILLER_21_604 VPWR VGND sg13g2_decap_4
XFILLER_34_987 VPWR VGND sg13g2_decap_8
XFILLER_21_626 VPWR VGND sg13g2_fill_2
XFILLER_21_637 VPWR VGND sg13g2_decap_8
X_1985_ ppwm_i.u_ppwm.global_counter\[0\] net326 _0148_ VPWR VGND sg13g2_xor2_1
X_2606_ net429 VPWR _0982_ VGND net491 net596 sg13g2_o21ai_1
X_2537_ _0942_ VPWR _0943_ VGND _0939_ _0941_ sg13g2_o21ai_1
X_2468_ VGND VPWR _0880_ _0878_ _0875_ sg13g2_or2_1
X_2399_ VPWR _0816_ _0815_ VGND sg13g2_inv_1
XFILLER_28_225 VPWR VGND sg13g2_decap_8
XFILLER_43_239 VPWR VGND sg13g2_decap_8
XFILLER_25_943 VPWR VGND sg13g2_decap_8
XFILLER_37_781 VPWR VGND sg13g2_decap_8
XFILLER_40_913 VPWR VGND sg13g2_decap_8
XFILLER_4_825 VPWR VGND sg13g2_decap_8
XFILLER_47_556 VPWR VGND sg13g2_fill_2
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_16_976 VPWR VGND sg13g2_decap_8
XFILLER_30_445 VPWR VGND sg13g2_fill_2
XFILLER_31_968 VPWR VGND sg13g2_decap_8
X_1770_ VPWR VGND _1336_ net509 _1335_ _1333_ _1337_ _1334_ sg13g2_a221oi_1
X_3035__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_6_140 VPWR VGND sg13g2_fill_1
XFILLER_6_173 VPWR VGND sg13g2_fill_1
X_2322_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] ppwm_i.u_ppwm.pwm_value\[7\] net400 _0743_
+ VPWR VGND sg13g2_mux2_1
X_2253_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0675_ net375 _0670_ _0677_
+ net376 sg13g2_a221oi_1
X_2184_ VPWR VGND _0608_ _0609_ _0607_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] _0610_
+ _1265_ sg13g2_a221oi_1
XFILLER_25_217 VPWR VGND sg13g2_decap_4
XFILLER_25_239 VPWR VGND sg13g2_decap_8
XFILLER_33_250 VPWR VGND sg13g2_decap_8
XFILLER_34_784 VPWR VGND sg13g2_decap_8
XFILLER_22_968 VPWR VGND sg13g2_decap_8
X_1968_ _0445_ _0444_ _0041_ VPWR VGND sg13g2_xor2_1
X_1899_ net293 net294 _0062_ VPWR VGND sg13g2_and2_1
XFILLER_1_828 VPWR VGND sg13g2_decap_8
XFILLER_44_515 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_decap_4
XFILLER_13_913 VPWR VGND sg13g2_decap_8
XFILLER_24_250 VPWR VGND sg13g2_fill_2
XFILLER_25_773 VPWR VGND sg13g2_decap_8
XFILLER_31_209 VPWR VGND sg13g2_fill_2
XFILLER_12_423 VPWR VGND sg13g2_decap_8
XFILLER_40_787 VPWR VGND sg13g2_decap_8
XFILLER_8_449 VPWR VGND sg13g2_decap_8
X_2996__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_3_165 VPWR VGND sg13g2_fill_1
XFILLER_0_850 VPWR VGND sg13g2_decap_8
XFILLER_48_821 VPWR VGND sg13g2_decap_8
XFILLER_47_331 VPWR VGND sg13g2_decap_4
Xhold5 sdr_i.mac1.sum_lvl2_ff\[9\] VPWR VGND net205 sg13g2_dlygate4sd3_1
XFILLER_47_342 VPWR VGND sg13g2_fill_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
X_2940_ net545 VGND VPWR _0131_ sdr_i.DP_4.matrix\[1\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_15_261 VPWR VGND sg13g2_fill_1
XFILLER_16_773 VPWR VGND sg13g2_fill_1
XFILLER_22_209 VPWR VGND sg13g2_decap_8
X_2871_ net294 _0134_ VPWR VGND sg13g2_buf_1
XFILLER_31_743 VPWR VGND sg13g2_decap_4
X_1822_ _0370_ VPWR _0000_ VGND _1278_ _0368_ sg13g2_o21ai_1
XFILLER_30_275 VPWR VGND sg13g2_fill_1
XFILLER_8_972 VPWR VGND sg13g2_decap_8
X_1753_ ppwm_i.u_ppwm.u_mem.memory\[28\] net514 net517 _1320_ VPWR VGND sg13g2_nor3_1
Xhold427 ppwm_i.u_ppwm.global_counter\[8\] VPWR VGND net807 sg13g2_dlygate4sd3_1
Xhold405 ppwm_i.u_ppwm.u_pwm.counter\[4\] VPWR VGND net785 sg13g2_dlygate4sd3_1
Xhold416 ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] VPWR VGND net796 sg13g2_dlygate4sd3_1
X_1684_ VPWR _1255_ net572 VGND sg13g2_inv_1
X_3423_ net548 net10 VPWR VGND sg13g2_buf_1
Xhold449 _0200_ VPWR VGND net829 sg13g2_dlygate4sd3_1
Xhold438 ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] VPWR VGND net818 sg13g2_dlygate4sd3_1
XFILLER_31_0 VPWR VGND sg13g2_decap_8
X_2305_ net393 _0674_ _0727_ VPWR VGND sg13g2_nor2_1
X_2236_ _1215_ net399 _0660_ VPWR VGND sg13g2_nor2_1
XFILLER_39_876 VPWR VGND sg13g2_decap_8
XFILLER_26_537 VPWR VGND sg13g2_decap_8
X_2167_ _1227_ ppwm_i.u_ppwm.global_counter\[2\] _0593_ VPWR VGND sg13g2_nor2_1
X_2098_ _0524_ _0522_ _0527_ VPWR VGND sg13g2_xor2_1
XFILLER_26_548 VPWR VGND sg13g2_fill_1
XFILLER_10_916 VPWR VGND sg13g2_decap_8
XFILLER_16_1018 VPWR VGND sg13g2_decap_8
XFILLER_22_798 VPWR VGND sg13g2_decap_4
XFILLER_5_419 VPWR VGND sg13g2_decap_8
XFILLER_28_75 VPWR VGND sg13g2_decap_8
XFILLER_29_331 VPWR VGND sg13g2_fill_2
XFILLER_45_835 VPWR VGND sg13g2_decap_8
X_3089__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_17_515 VPWR VGND sg13g2_fill_2
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_8_246 VPWR VGND sg13g2_decap_8
XFILLER_12_264 VPWR VGND sg13g2_decap_8
XFILLER_5_986 VPWR VGND sg13g2_decap_8
X_3070_ net158 VGND VPWR _0261_ ppwm_i.u_ppwm.u_mem.memory\[46\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_39_139 VPWR VGND sg13g2_fill_2
X_2021_ _0472_ net798 net804 _0474_ VPWR VGND sg13g2_a21o_1
XFILLER_48_640 VPWR VGND sg13g2_fill_2
XFILLER_36_835 VPWR VGND sg13g2_decap_8
XFILLER_35_389 VPWR VGND sg13g2_fill_1
X_2923_ net546 VGND VPWR _0114_ sdr_i.DP_3.matrix\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2854_ net245 _0117_ VPWR VGND sg13g2_buf_1
X_1805_ _0354_ ppwm_i.u_ppwm.u_mem.memory\[72\] net439 VPWR VGND sg13g2_nand2_1
X_2785_ net661 _1072_ _1074_ VPWR VGND sg13g2_nor2_1
X_1736_ _1303_ _1177_ net448 VPWR VGND sg13g2_nand2_1
Xhold202 ppwm_i.u_ppwm.u_mem.memory\[111\] VPWR VGND net582 sg13g2_dlygate4sd3_1
Xhold213 _0260_ VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold235 _0304_ VPWR VGND net615 sg13g2_dlygate4sd3_1
Xhold224 ppwm_i.u_ppwm.u_mem.memory\[110\] VPWR VGND net604 sg13g2_dlygate4sd3_1
XFILLER_49_19 VPWR VGND sg13g2_decap_8
X_1667_ VPWR _1238_ ppwm_i.u_ppwm.u_pwm.counter\[6\] VGND sg13g2_inv_1
Xhold257 ppwm_i.u_ppwm.u_mem.memory\[69\] VPWR VGND net637 sg13g2_dlygate4sd3_1
Xhold246 _0316_ VPWR VGND net626 sg13g2_dlygate4sd3_1
Xhold268 _0225_ VPWR VGND net648 sg13g2_dlygate4sd3_1
X_1598_ VPWR _1169_ net699 VGND sg13g2_inv_1
Xhold279 ppwm_i.u_ppwm.u_mem.memory\[66\] VPWR VGND net659 sg13g2_dlygate4sd3_1
X_2219_ _0641_ VPWR _0645_ VGND _0642_ _0644_ sg13g2_o21ai_1
XFILLER_45_109 VPWR VGND sg13g2_decap_4
XFILLER_39_673 VPWR VGND sg13g2_decap_8
XFILLER_27_835 VPWR VGND sg13g2_decap_8
X_3199_ net542 VGND VPWR _0067_ sdr_i.mac2.products_ff\[86\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_26_323 VPWR VGND sg13g2_decap_4
XFILLER_41_337 VPWR VGND sg13g2_fill_1
XFILLER_6_717 VPWR VGND sg13g2_fill_2
XFILLER_10_768 VPWR VGND sg13g2_fill_1
XFILLER_10_757 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_30_76 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_1_422 VPWR VGND sg13g2_fill_1
XFILLER_1_477 VPWR VGND sg13g2_decap_4
XFILLER_45_621 VPWR VGND sg13g2_decap_4
XFILLER_29_194 VPWR VGND sg13g2_decap_8
XFILLER_41_871 VPWR VGND sg13g2_decap_8
XFILLER_13_562 VPWR VGND sg13g2_decap_8
XFILLER_5_750 VPWR VGND sg13g2_decap_8
X_2570_ net431 VPWR _0964_ VGND net497 net642 sg13g2_o21ai_1
XFILLER_5_794 VPWR VGND sg13g2_fill_1
X_3122_ net41 VGND VPWR net556 ppwm_i.u_ppwm.u_mem.memory\[98\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_49_993 VPWR VGND sg13g2_decap_8
X_3053_ net44 VGND VPWR net577 ppwm_i.u_ppwm.u_mem.memory\[29\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2004_ _0157_ net335 _0463_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_827 VPWR VGND sg13g2_decap_8
XFILLER_36_665 VPWR VGND sg13g2_fill_2
XFILLER_23_359 VPWR VGND sg13g2_fill_1
X_2906_ net521 VGND VPWR _0097_ sdr_i.DP_2.matrix\[10\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2837_ net275 _0100_ VPWR VGND sg13g2_buf_1
X_2768_ net415 VPWR _1063_ VGND net472 ppwm_i.u_ppwm.u_mem.memory\[109\] sg13g2_o21ai_1
X_1719_ _1286_ net439 _1136_ net443 _1143_ VPWR VGND sg13g2_a22oi_1
X_2699_ VGND VPWR net465 _1134_ _0289_ _1028_ sg13g2_a21oi_1
Xfanout523 net524 net523 VPWR VGND sg13g2_buf_8
Xfanout512 net513 net512 VPWR VGND sg13g2_buf_8
Xfanout501 net690 net501 VPWR VGND sg13g2_buf_8
Xfanout545 net546 net545 VPWR VGND sg13g2_buf_2
Xfanout534 net547 net534 VPWR VGND sg13g2_buf_8
XFILLER_27_621 VPWR VGND sg13g2_fill_2
XFILLER_14_315 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_41_145 VPWR VGND sg13g2_fill_2
XFILLER_22_381 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_6_503 VPWR VGND sg13g2_decap_8
XFILLER_10_576 VPWR VGND sg13g2_decap_8
XFILLER_6_569 VPWR VGND sg13g2_fill_1
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_49_212 VPWR VGND sg13g2_decap_8
XFILLER_1_274 VPWR VGND sg13g2_decap_8
XFILLER_49_289 VPWR VGND sg13g2_decap_8
XFILLER_46_941 VPWR VGND sg13g2_decap_8
XFILLER_18_621 VPWR VGND sg13g2_decap_8
XFILLER_18_643 VPWR VGND sg13g2_decap_8
XFILLER_18_698 VPWR VGND sg13g2_fill_2
XFILLER_21_819 VPWR VGND sg13g2_decap_8
XFILLER_14_893 VPWR VGND sg13g2_decap_8
XFILLER_20_307 VPWR VGND sg13g2_fill_2
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_2622_ net430 VPWR _0990_ VGND net487 net584 sg13g2_o21ai_1
X_2553_ VGND VPWR net490 _1207_ _0216_ _0955_ sg13g2_a21oi_1
X_2484_ VPWR VGND _0894_ net458 _0891_ _1216_ _0208_ net370 sg13g2_a221oi_1
X_3105_ net176 VGND VPWR net701 ppwm_i.u_ppwm.u_mem.memory\[81\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_28_407 VPWR VGND sg13g2_decap_8
XFILLER_49_790 VPWR VGND sg13g2_decap_8
X_3036_ net77 VGND VPWR net610 ppwm_i.u_ppwm.u_mem.memory\[12\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_37_963 VPWR VGND sg13g2_decap_8
XFILLER_12_819 VPWR VGND sg13g2_decap_8
XFILLER_23_189 VPWR VGND sg13g2_decap_4
XFILLER_11_89 VPWR VGND sg13g2_fill_2
XFILLER_47_705 VPWR VGND sg13g2_decap_8
Xfanout375 _0676_ net375 VPWR VGND sg13g2_buf_8
XFILLER_47_716 VPWR VGND sg13g2_fill_1
XFILLER_19_407 VPWR VGND sg13g2_fill_1
Xfanout397 _1310_ net397 VPWR VGND sg13g2_buf_8
Xfanout386 net388 net386 VPWR VGND sg13g2_buf_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_36_64 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
XFILLER_14_112 VPWR VGND sg13g2_decap_4
XFILLER_36_97 VPWR VGND sg13g2_fill_1
XFILLER_14_145 VPWR VGND sg13g2_decap_4
XFILLER_15_646 VPWR VGND sg13g2_fill_1
XFILLER_15_657 VPWR VGND sg13g2_fill_1
X_3047__55 VPWR VGND net55 sg13g2_tiehi
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_7_801 VPWR VGND sg13g2_fill_1
XFILLER_10_340 VPWR VGND sg13g2_decap_4
XFILLER_6_311 VPWR VGND sg13g2_decap_8
XFILLER_7_878 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_fill_2
XFILLER_42_1014 VPWR VGND sg13g2_decap_8
XFILLER_38_716 VPWR VGND sg13g2_decap_8
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_18_440 VPWR VGND sg13g2_fill_2
XFILLER_33_421 VPWR VGND sg13g2_decap_4
XFILLER_34_966 VPWR VGND sg13g2_decap_8
X_1984_ _0455_ _0454_ _0051_ VPWR VGND sg13g2_xor2_1
X_2605_ VGND VPWR net493 _1181_ _0242_ _0981_ sg13g2_a21oi_1
X_2536_ VGND VPWR _0939_ _0941_ _0942_ _0685_ sg13g2_a21oi_1
X_2467_ _0879_ _0875_ _0878_ VPWR VGND sg13g2_nand2_1
X_2398_ _0815_ net503 net391 VPWR VGND sg13g2_xnor2_1
XFILLER_29_738 VPWR VGND sg13g2_decap_4
XFILLER_25_922 VPWR VGND sg13g2_decap_8
X_3019_ net111 VGND VPWR _0210_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_11_104 VPWR VGND sg13g2_decap_8
XFILLER_25_999 VPWR VGND sg13g2_decap_8
XFILLER_40_969 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_decap_4
XFILLER_22_55 VPWR VGND sg13g2_decap_8
XFILLER_22_99 VPWR VGND sg13g2_fill_1
XFILLER_3_336 VPWR VGND sg13g2_fill_1
XFILLER_3_314 VPWR VGND sg13g2_decap_4
XFILLER_47_568 VPWR VGND sg13g2_decap_4
XFILLER_28_782 VPWR VGND sg13g2_decap_8
XFILLER_16_955 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_decap_8
XFILLER_42_295 VPWR VGND sg13g2_decap_8
XFILLER_30_424 VPWR VGND sg13g2_decap_8
XFILLER_31_947 VPWR VGND sg13g2_decap_8
XFILLER_11_671 VPWR VGND sg13g2_decap_8
X_2321_ VPWR VGND net390 _0741_ _0695_ net386 _0742_ _0655_ sg13g2_a221oi_1
X_2252_ _0551_ net380 _0676_ VPWR VGND sg13g2_and2_1
XFILLER_2_380 VPWR VGND sg13g2_decap_8
X_2183_ _1218_ ppwm_i.u_ppwm.global_counter\[1\] _0609_ VPWR VGND sg13g2_nor2_1
XFILLER_19_760 VPWR VGND sg13g2_decap_8
XFILLER_21_402 VPWR VGND sg13g2_fill_1
XFILLER_21_435 VPWR VGND sg13g2_decap_8
XFILLER_22_947 VPWR VGND sg13g2_decap_8
XFILLER_21_468 VPWR VGND sg13g2_decap_8
X_1967_ _0445_ net281 net240 VPWR VGND sg13g2_nand2_1
X_1898_ net290 net296 _0060_ VPWR VGND sg13g2_and2_1
XFILLER_1_807 VPWR VGND sg13g2_decap_8
X_2519_ VGND VPWR _0916_ _0919_ _0926_ _0915_ sg13g2_a21oi_1
XFILLER_25_1020 VPWR VGND sg13g2_decap_8
XFILLER_44_527 VPWR VGND sg13g2_decap_4
XFILLER_17_44 VPWR VGND sg13g2_decap_8
XFILLER_13_969 VPWR VGND sg13g2_decap_8
XFILLER_8_406 VPWR VGND sg13g2_decap_8
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_33_98 VPWR VGND sg13g2_decap_4
XFILLER_48_800 VPWR VGND sg13g2_decap_8
Xhold6 sdr_i.mac1.sum_lvl1_ff\[33\] VPWR VGND net206 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_decap_8
XFILLER_35_538 VPWR VGND sg13g2_fill_2
XFILLER_35_549 VPWR VGND sg13g2_fill_2
X_2870_ net222 _0133_ VPWR VGND sg13g2_buf_1
XFILLER_43_593 VPWR VGND sg13g2_decap_4
XFILLER_15_273 VPWR VGND sg13g2_decap_8
XFILLER_15_295 VPWR VGND sg13g2_decap_4
X_1821_ VGND VPWR _1249_ net759 _0370_ net457 sg13g2_a21oi_1
XFILLER_8_951 VPWR VGND sg13g2_decap_8
X_1752_ VGND VPWR _1167_ net440 _1319_ net461 sg13g2_a21oi_1
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_1683_ _1254_ net780 VPWR VGND sg13g2_inv_2
Xhold406 ppwm_i.u_ppwm.u_pwm.counter\[3\] VPWR VGND net786 sg13g2_dlygate4sd3_1
Xhold417 _0486_ VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold439 ppwm_i.u_ppwm.u_pwm.counter\[7\] VPWR VGND net819 sg13g2_dlygate4sd3_1
Xhold428 ppwm_i.u_ppwm.u_pwm.counter\[6\] VPWR VGND net808 sg13g2_dlygate4sd3_1
X_3422_ net548 net9 VPWR VGND sg13g2_buf_1
X_2304_ VPWR VGND _0659_ _0721_ _0725_ net379 _0726_ _0668_ sg13g2_a221oi_1
X_2235_ net396 net395 net392 _0659_ VGND VPWR _0651_ sg13g2_nor4_2
XFILLER_38_310 VPWR VGND sg13g2_decap_8
XFILLER_39_855 VPWR VGND sg13g2_decap_8
X_2166_ _0591_ VPWR _0592_ VGND _0589_ _0590_ sg13g2_o21ai_1
XFILLER_0_1011 VPWR VGND sg13g2_decap_8
XFILLER_38_365 VPWR VGND sg13g2_decap_8
X_2097_ _0518_ VPWR _0526_ VGND net451 net449 sg13g2_o21ai_1
X_2999_ net150 VGND VPWR _0190_ ppwm_i.u_ppwm.pc\[1\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_21_276 VPWR VGND sg13g2_fill_1
XFILLER_1_615 VPWR VGND sg13g2_decap_4
XFILLER_1_648 VPWR VGND sg13g2_decap_8
XFILLER_45_814 VPWR VGND sg13g2_decap_8
XFILLER_29_398 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_fill_1
XFILLER_12_221 VPWR VGND sg13g2_decap_8
X_3024__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_40_585 VPWR VGND sg13g2_fill_1
XFILLER_8_236 VPWR VGND sg13g2_fill_1
XFILLER_13_799 VPWR VGND sg13g2_decap_4
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_4_475 VPWR VGND sg13g2_decap_8
X_2020_ net798 _0472_ net804 _0473_ VPWR VGND sg13g2_nand3_1
XFILLER_47_140 VPWR VGND sg13g2_fill_1
XFILLER_47_151 VPWR VGND sg13g2_fill_1
XFILLER_36_814 VPWR VGND sg13g2_decap_8
X_2922_ net545 VGND VPWR _0113_ sdr_i.DP_3.matrix\[1\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2853_ net293 _0116_ VPWR VGND sg13g2_buf_1
XFILLER_31_585 VPWR VGND sg13g2_decap_8
XFILLER_31_596 VPWR VGND sg13g2_fill_1
X_1804_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[86\] net460 net449 ppwm_i.u_ppwm.u_mem.memory\[107\]
+ _0353_ net452 sg13g2_a221oi_1
X_2784_ net661 _1072_ _1073_ VPWR VGND sg13g2_and2_1
X_1735_ _1302_ _1300_ _1301_ _1299_ _1297_ VPWR VGND sg13g2_a22oi_1
Xhold214 ppwm_i.u_ppwm.u_mem.memory\[103\] VPWR VGND net594 sg13g2_dlygate4sd3_1
Xhold225 _0324_ VPWR VGND net605 sg13g2_dlygate4sd3_1
Xhold203 _0325_ VPWR VGND net583 sg13g2_dlygate4sd3_1
X_1666_ VPWR _1237_ net819 VGND sg13g2_inv_1
Xhold258 ppwm_i.u_ppwm.u_mem.memory\[49\] VPWR VGND net638 sg13g2_dlygate4sd3_1
Xhold236 ppwm_i.u_ppwm.u_mem.memory\[108\] VPWR VGND net616 sg13g2_dlygate4sd3_1
Xhold247 ppwm_i.u_ppwm.u_mem.memory\[109\] VPWR VGND net627 sg13g2_dlygate4sd3_1
Xhold269 ppwm_i.u_ppwm.u_mem.memory\[101\] VPWR VGND net649 sg13g2_dlygate4sd3_1
X_1597_ VPWR _1168_ net702 VGND sg13g2_inv_1
X_2218_ _0638_ _0643_ _0644_ VPWR VGND sg13g2_and2_1
XFILLER_26_313 VPWR VGND sg13g2_fill_1
X_3198_ net543 VGND VPWR _0066_ sdr_i.mac2.products_ff\[85\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2149_ _0575_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _1256_ VPWR VGND sg13g2_nand2_1
XFILLER_42_839 VPWR VGND sg13g2_decap_8
XFILLER_22_563 VPWR VGND sg13g2_fill_2
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_39_97 VPWR VGND sg13g2_decap_8
XFILLER_17_302 VPWR VGND sg13g2_decap_8
XFILLER_17_324 VPWR VGND sg13g2_decap_8
XFILLER_18_869 VPWR VGND sg13g2_decap_8
XFILLER_45_666 VPWR VGND sg13g2_fill_2
XFILLER_33_839 VPWR VGND sg13g2_decap_8
XFILLER_41_850 VPWR VGND sg13g2_decap_8
XFILLER_13_552 VPWR VGND sg13g2_fill_2
XFILLER_13_585 VPWR VGND sg13g2_fill_1
XFILLER_9_589 VPWR VGND sg13g2_decap_8
X_3121_ net49 VGND VPWR _0312_ ppwm_i.u_ppwm.u_mem.memory\[97\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_49_972 VPWR VGND sg13g2_decap_8
X_3052_ net46 VGND VPWR _0243_ ppwm_i.u_ppwm.u_mem.memory\[28\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_2003_ _1259_ _0463_ _0465_ VPWR VGND sg13g2_nor2_2
X_2905_ net521 VGND VPWR _0096_ sdr_i.DP_2.matrix\[9\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_31_360 VPWR VGND sg13g2_decap_4
X_2836_ net241 _0099_ VPWR VGND sg13g2_buf_1
X_2767_ VGND VPWR net469 _1100_ _0323_ _1062_ sg13g2_a21oi_1
X_2698_ net412 VPWR _1028_ VGND net465 ppwm_i.u_ppwm.u_mem.memory\[74\] sg13g2_o21ai_1
X_1718_ VPWR VGND _1108_ _1281_ net439 _1101_ _1285_ net451 sg13g2_a221oi_1
X_1649_ ppwm_i.u_ppwm.pwm_value\[9\] _1220_ VPWR VGND sg13g2_inv_4
XFILLER_6_90 VPWR VGND sg13g2_decap_8
X_3138__68 VPWR VGND net68 sg13g2_tiehi
Xfanout502 net836 net502 VPWR VGND sg13g2_buf_8
Xfanout524 net547 net524 VPWR VGND sg13g2_buf_8
Xfanout513 net827 net513 VPWR VGND sg13g2_buf_8
Xfanout535 net537 net535 VPWR VGND sg13g2_buf_8
Xfanout546 net547 net546 VPWR VGND sg13g2_buf_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_27_655 VPWR VGND sg13g2_fill_2
XFILLER_27_677 VPWR VGND sg13g2_decap_4
XFILLER_23_894 VPWR VGND sg13g2_decap_8
XFILLER_10_555 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_29_1018 VPWR VGND sg13g2_decap_8
XFILLER_2_37 VPWR VGND sg13g2_decap_8
XFILLER_49_268 VPWR VGND sg13g2_decap_8
XFILLER_46_920 VPWR VGND sg13g2_decap_8
XFILLER_46_997 VPWR VGND sg13g2_decap_8
XFILLER_33_614 VPWR VGND sg13g2_decap_8
XFILLER_13_360 VPWR VGND sg13g2_fill_2
XFILLER_9_320 VPWR VGND sg13g2_fill_1
X_2621_ VGND VPWR net491 _1173_ _0250_ _0989_ sg13g2_a21oi_1
X_2552_ net430 VPWR _0955_ VGND net490 ppwm_i.u_ppwm.u_mem.memory\[1\] sg13g2_o21ai_1
X_2483_ _0894_ _0748_ net374 _0893_ VPWR VGND sg13g2_and3_1
X_3104_ net183 VGND VPWR _0295_ ppwm_i.u_ppwm.u_mem.memory\[80\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_3035_ net79 VGND VPWR _0226_ ppwm_i.u_ppwm.u_mem.memory\[11\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_37_942 VPWR VGND sg13g2_decap_8
XFILLER_24_625 VPWR VGND sg13g2_decap_4
XFILLER_36_496 VPWR VGND sg13g2_decap_4
XFILLER_23_135 VPWR VGND sg13g2_decap_8
XFILLER_24_647 VPWR VGND sg13g2_fill_2
XFILLER_32_691 VPWR VGND sg13g2_decap_8
X_2819_ net304 _0082_ VPWR VGND sg13g2_buf_1
XFILLER_11_68 VPWR VGND sg13g2_decap_8
XFILLER_2_8 VPWR VGND sg13g2_fill_1
Xfanout376 _0673_ net376 VPWR VGND sg13g2_buf_8
Xfanout398 net400 net398 VPWR VGND sg13g2_buf_8
Xfanout387 net388 net387 VPWR VGND sg13g2_buf_2
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_15_625 VPWR VGND sg13g2_decap_8
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_30_617 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_22_190 VPWR VGND sg13g2_fill_1
XFILLER_7_857 VPWR VGND sg13g2_decap_8
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_46_794 VPWR VGND sg13g2_decap_8
XFILLER_33_411 VPWR VGND sg13g2_fill_2
XFILLER_34_945 VPWR VGND sg13g2_decap_8
XFILLER_33_488 VPWR VGND sg13g2_fill_2
X_1983_ _0455_ net303 net225 VPWR VGND sg13g2_nand2_1
XFILLER_9_150 VPWR VGND sg13g2_fill_1
XFILLER_9_183 VPWR VGND sg13g2_decap_8
X_2604_ net429 VPWR _0981_ VGND net493 net550 sg13g2_o21ai_1
X_2535_ _0941_ _1211_ _0335_ VPWR VGND sg13g2_xnor2_1
X_2466_ _0876_ _0877_ _0878_ VPWR VGND sg13g2_and2_1
X_2397_ VGND VPWR _0796_ _0800_ _0814_ _0795_ sg13g2_a21oi_1
XFILLER_29_717 VPWR VGND sg13g2_decap_8
XFILLER_25_901 VPWR VGND sg13g2_decap_8
X_3018_ net113 VGND VPWR _0209_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] clknet_3_6__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_25_978 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_24_466 VPWR VGND sg13g2_decap_4
XFILLER_40_948 VPWR VGND sg13g2_decap_8
XFILLER_22_34 VPWR VGND sg13g2_decap_8
XFILLER_47_514 VPWR VGND sg13g2_decap_8
X_3122__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_47_558 VPWR VGND sg13g2_fill_1
XFILLER_47_86 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_16_934 VPWR VGND sg13g2_decap_8
XFILLER_43_731 VPWR VGND sg13g2_decap_8
XFILLER_42_230 VPWR VGND sg13g2_fill_1
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_42_263 VPWR VGND sg13g2_decap_4
XFILLER_15_455 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_fill_2
XFILLER_31_926 VPWR VGND sg13g2_decap_8
XFILLER_42_274 VPWR VGND sg13g2_decap_8
XFILLER_11_694 VPWR VGND sg13g2_fill_1
XFILLER_3_882 VPWR VGND sg13g2_decap_8
X_2320_ _0740_ VPWR _0741_ VGND _0351_ _0656_ sg13g2_o21ai_1
X_2251_ _1311_ _0674_ _0675_ VPWR VGND sg13g2_nor2_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ _1219_ ppwm_i.u_ppwm.global_counter\[0\] _0608_ VPWR VGND sg13g2_nor2_1
XFILLER_18_282 VPWR VGND sg13g2_fill_1
XFILLER_22_926 VPWR VGND sg13g2_decap_8
X_1966_ _0444_ net273 net241 VPWR VGND sg13g2_nand2_1
X_1897_ _0033_ _0410_ _0411_ VPWR VGND sg13g2_xnor2_1
X_3034__81 VPWR VGND net81 sg13g2_tiehi
X_2518_ VGND VPWR _1213_ net370 _0211_ _0925_ sg13g2_a21oi_1
XFILLER_0_307 VPWR VGND sg13g2_decap_8
X_2449_ _0863_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] net397 VPWR VGND sg13g2_nand2_1
XFILLER_25_742 VPWR VGND sg13g2_decap_8
XFILLER_25_753 VPWR VGND sg13g2_fill_1
XFILLER_13_948 VPWR VGND sg13g2_decap_8
XFILLER_9_919 VPWR VGND sg13g2_decap_8
XFILLER_12_458 VPWR VGND sg13g2_decap_8
XFILLER_32_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_635 VPWR VGND sg13g2_fill_2
XFILLER_4_624 VPWR VGND sg13g2_decap_8
XFILLER_0_885 VPWR VGND sg13g2_decap_8
Xhold7 sdr_i.mac1.products_ff\[137\] VPWR VGND net207 sg13g2_dlygate4sd3_1
XFILLER_48_856 VPWR VGND sg13g2_decap_8
XFILLER_35_517 VPWR VGND sg13g2_fill_1
XFILLER_16_731 VPWR VGND sg13g2_decap_8
XFILLER_16_786 VPWR VGND sg13g2_fill_2
XFILLER_31_712 VPWR VGND sg13g2_decap_8
XFILLER_30_200 VPWR VGND sg13g2_fill_1
X_1820_ _1249_ net457 _0369_ VPWR VGND sg13g2_nor2_1
XFILLER_30_244 VPWR VGND sg13g2_decap_8
XFILLER_31_756 VPWR VGND sg13g2_decap_8
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_30_266 VPWR VGND sg13g2_decap_8
X_1751_ VPWR VGND _1317_ _1231_ _1316_ _1314_ _1318_ _1315_ sg13g2_a221oi_1
X_3001__146 VPWR VGND net146 sg13g2_tiehi
Xhold418 ppwm_i.u_ppwm.global_counter\[17\] VPWR VGND net798 sg13g2_dlygate4sd3_1
X_1682_ VPWR _1253_ net798 VGND sg13g2_inv_1
Xhold407 ppwm_i.u_ppwm.global_counter\[11\] VPWR VGND net787 sg13g2_dlygate4sd3_1
XFILLER_48_1010 VPWR VGND sg13g2_decap_8
Xhold429 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] VPWR VGND net809 sg13g2_dlygate4sd3_1
X_3421_ net549 net8 VPWR VGND sg13g2_buf_1
X_3112__119 VPWR VGND net119 sg13g2_tiehi
X_2303_ VGND VPWR net387 _0723_ _0725_ _0724_ sg13g2_a21oi_1
XFILLER_39_834 VPWR VGND sg13g2_decap_8
X_2234_ VGND VPWR net384 _0655_ _0658_ _0657_ sg13g2_a21oi_1
XFILLER_17_0 VPWR VGND sg13g2_decap_8
X_2165_ _0591_ ppwm_i.u_ppwm.pwm_value\[1\] ppwm_i.u_ppwm.global_counter\[1\] VPWR
+ VGND sg13g2_nand2b_1
X_2096_ _0525_ _1232_ net515 VPWR VGND sg13g2_nand2_1
XFILLER_21_233 VPWR VGND sg13g2_fill_2
X_2998_ net152 VGND VPWR _0189_ ppwm_i.u_ppwm.pc\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_21_266 VPWR VGND sg13g2_decap_4
X_1949_ _0028_ _0434_ net744 VPWR VGND sg13g2_xnor2_1
XFILLER_48_108 VPWR VGND sg13g2_fill_2
XFILLER_0_159 VPWR VGND sg13g2_fill_2
XFILLER_0_137 VPWR VGND sg13g2_decap_8
XFILLER_44_314 VPWR VGND sg13g2_decap_8
XFILLER_44_369 VPWR VGND sg13g2_fill_1
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_44_65 VPWR VGND sg13g2_decap_8
XFILLER_25_583 VPWR VGND sg13g2_decap_8
XFILLER_9_705 VPWR VGND sg13g2_decap_8
XFILLER_9_716 VPWR VGND sg13g2_fill_1
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_4_465 VPWR VGND sg13g2_decap_8
XFILLER_0_682 VPWR VGND sg13g2_decap_8
XFILLER_39_108 VPWR VGND sg13g2_fill_2
XFILLER_48_686 VPWR VGND sg13g2_fill_2
XFILLER_39_1009 VPWR VGND sg13g2_decap_8
XFILLER_35_358 VPWR VGND sg13g2_decap_4
X_2921_ net544 VGND VPWR _0112_ sdr_i.DP_3.matrix\[0\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_16_583 VPWR VGND sg13g2_decap_4
XFILLER_31_531 VPWR VGND sg13g2_decap_8
XFILLER_31_542 VPWR VGND sg13g2_fill_2
XFILLER_31_553 VPWR VGND sg13g2_decap_8
X_2852_ net219 _0115_ VPWR VGND sg13g2_buf_1
X_1803_ _0352_ net439 ppwm_i.u_ppwm.u_mem.memory\[100\] net443 ppwm_i.u_ppwm.u_mem.memory\[93\]
+ VPWR VGND sg13g2_a22oi_1
X_2783_ _1067_ net717 _1072_ _0329_ VPWR VGND sg13g2_nor3_1
X_1734_ VPWR VGND _1135_ net510 net438 _1149_ _1301_ net447 sg13g2_a221oi_1
Xhold204 ppwm_i.u_ppwm.u_mem.memory\[36\] VPWR VGND net584 sg13g2_dlygate4sd3_1
Xhold226 ppwm_i.u_ppwm.u_mem.memory\[37\] VPWR VGND net606 sg13g2_dlygate4sd3_1
Xhold215 _0317_ VPWR VGND net595 sg13g2_dlygate4sd3_1
X_1665_ VPWR _1236_ ppwm_i.u_ppwm.u_pwm.counter\[8\] VGND sg13g2_inv_1
Xhold259 ppwm_i.u_ppwm.u_mem.memory\[50\] VPWR VGND net639 sg13g2_dlygate4sd3_1
Xhold237 ppwm_i.u_ppwm.u_mem.memory\[23\] VPWR VGND net617 sg13g2_dlygate4sd3_1
Xhold248 ppwm_i.u_ppwm.u_mem.memory\[6\] VPWR VGND net628 sg13g2_dlygate4sd3_1
X_1596_ VPWR _1167_ net682 VGND sg13g2_inv_1
XFILLER_39_620 VPWR VGND sg13g2_decap_4
X_2217_ VGND VPWR _1210_ ppwm_i.u_ppwm.pwm_value\[9\] _0643_ net381 sg13g2_a21oi_1
XFILLER_22_1024 VPWR VGND sg13g2_decap_4
X_3197_ net543 VGND VPWR _0047_ sdr_i.mac2.products_ff\[69\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2148_ VPWR VGND _0572_ _0573_ _0571_ _1217_ _0574_ ppwm_i.u_ppwm.global_counter\[12\]
+ sg13g2_a221oi_1
XFILLER_38_174 VPWR VGND sg13g2_fill_2
XFILLER_38_185 VPWR VGND sg13g2_decap_8
X_2079_ net766 _0511_ _0512_ VPWR VGND sg13g2_nor2_1
XFILLER_42_818 VPWR VGND sg13g2_decap_8
XFILLER_26_358 VPWR VGND sg13g2_decap_8
XFILLER_35_892 VPWR VGND sg13g2_decap_8
XFILLER_22_542 VPWR VGND sg13g2_decap_8
XFILLER_6_719 VPWR VGND sg13g2_fill_1
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_49_428 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_39_76 VPWR VGND sg13g2_decap_8
XFILLER_18_815 VPWR VGND sg13g2_decap_8
XFILLER_44_111 VPWR VGND sg13g2_decap_8
XFILLER_29_185 VPWR VGND sg13g2_decap_4
XFILLER_33_818 VPWR VGND sg13g2_decap_8
XFILLER_26_892 VPWR VGND sg13g2_decap_8
XFILLER_9_524 VPWR VGND sg13g2_decap_8
XFILLER_40_394 VPWR VGND sg13g2_decap_8
XFILLER_40_383 VPWR VGND sg13g2_decap_8
XFILLER_4_240 VPWR VGND sg13g2_decap_4
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_295 VPWR VGND sg13g2_decap_8
X_3120_ net56 VGND VPWR _0311_ ppwm_i.u_ppwm.u_mem.memory\[96\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_49_951 VPWR VGND sg13g2_decap_8
X_3051_ net48 VGND VPWR _0242_ ppwm_i.u_ppwm.u_mem.memory\[27\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
X_2002_ _0463_ _0464_ _0156_ VPWR VGND sg13g2_and2_1
XFILLER_36_634 VPWR VGND sg13g2_decap_8
XFILLER_23_317 VPWR VGND sg13g2_decap_8
X_2904_ net523 VGND VPWR _0095_ sdr_i.DP_2.matrix\[1\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_32_884 VPWR VGND sg13g2_decap_8
X_2835_ net281 _0098_ VPWR VGND sg13g2_buf_1
XFILLER_31_383 VPWR VGND sg13g2_decap_4
X_2766_ net419 VPWR _1062_ VGND net474 net616 sg13g2_o21ai_1
X_2697_ VGND VPWR net466 _1135_ _0288_ _1027_ sg13g2_a21oi_1
X_1717_ VGND VPWR _1115_ net443 _1284_ net460 sg13g2_a21oi_1
X_1648_ _1219_ net812 VPWR VGND sg13g2_inv_2
Xfanout503 net833 net503 VPWR VGND sg13g2_buf_8
Xfanout514 net516 net514 VPWR VGND sg13g2_buf_8
X_1579_ VPWR _1150_ net728 VGND sg13g2_inv_1
Xfanout547 rst_n_sdr net547 VPWR VGND sg13g2_buf_8
Xfanout525 net527 net525 VPWR VGND sg13g2_buf_8
Xfanout536 net537 net536 VPWR VGND sg13g2_buf_8
XFILLER_39_450 VPWR VGND sg13g2_decap_8
X_3059__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_26_144 VPWR VGND sg13g2_fill_1
XFILLER_23_840 VPWR VGND sg13g2_decap_4
XFILLER_23_873 VPWR VGND sg13g2_decap_8
XFILLER_10_534 VPWR VGND sg13g2_decap_8
XFILLER_2_700 VPWR VGND sg13g2_fill_2
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_49_247 VPWR VGND sg13g2_decap_8
XFILLER_46_976 VPWR VGND sg13g2_decap_8
XFILLER_32_103 VPWR VGND sg13g2_decap_8
XFILLER_14_851 VPWR VGND sg13g2_fill_1
XFILLER_13_394 VPWR VGND sg13g2_decap_8
X_2620_ net428 VPWR _0989_ VGND net491 ppwm_i.u_ppwm.u_mem.memory\[35\] sg13g2_o21ai_1
X_2551_ VGND VPWR net495 _1208_ _0215_ _0954_ sg13g2_a21oi_1
X_2482_ _0892_ VPWR _0893_ VGND net383 _0750_ sg13g2_o21ai_1
X_3103_ net191 VGND VPWR _0294_ ppwm_i.u_ppwm.u_mem.memory\[79\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_3034_ net81 VGND VPWR net648 ppwm_i.u_ppwm.u_mem.memory\[10\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_37_921 VPWR VGND sg13g2_decap_8
XFILLER_37_998 VPWR VGND sg13g2_decap_8
XFILLER_23_147 VPWR VGND sg13g2_decap_8
XFILLER_32_670 VPWR VGND sg13g2_decap_8
XFILLER_20_898 VPWR VGND sg13g2_decap_8
X_2818_ net240 _0081_ VPWR VGND sg13g2_buf_1
X_2749_ VGND VPWR net478 _1109_ _0314_ _1053_ sg13g2_a21oi_1
XFILLER_3_508 VPWR VGND sg13g2_fill_2
Xfanout399 net400 net399 VPWR VGND sg13g2_buf_8
Xfanout377 _0684_ net377 VPWR VGND sg13g2_buf_8
Xfanout388 net389 net388 VPWR VGND sg13g2_buf_1
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_27_431 VPWR VGND sg13g2_decap_8
XFILLER_27_442 VPWR VGND sg13g2_fill_2
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_10_386 VPWR VGND sg13g2_decap_8
XFILLER_7_836 VPWR VGND sg13g2_decap_8
XFILLER_6_357 VPWR VGND sg13g2_decap_8
XFILLER_2_552 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_46_773 VPWR VGND sg13g2_decap_8
XFILLER_34_924 VPWR VGND sg13g2_decap_8
X_1982_ _0454_ net310 net264 VPWR VGND sg13g2_nand2_1
X_2603_ VGND VPWR net493 _1182_ _0241_ _0980_ sg13g2_a21oi_1
X_2534_ _0940_ net841 net390 VPWR VGND sg13g2_nand2_1
XFILLER_6_891 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_fill_2
XFILLER_5_390 VPWR VGND sg13g2_fill_1
X_2465_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] VPWR _0877_ VGND net407 net405 sg13g2_o21ai_1
X_2396_ _0812_ _0813_ _0201_ VPWR VGND sg13g2_nor2_1
X_3011__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_28_239 VPWR VGND sg13g2_fill_1
X_3017_ net115 VGND VPWR _0208_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
XFILLER_36_261 VPWR VGND sg13g2_decap_8
XFILLER_37_795 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_25_957 VPWR VGND sg13g2_decap_8
XFILLER_40_927 VPWR VGND sg13g2_decap_8
XFILLER_4_839 VPWR VGND sg13g2_decap_8
XFILLER_19_217 VPWR VGND sg13g2_fill_2
XFILLER_16_913 VPWR VGND sg13g2_decap_8
XFILLER_15_412 VPWR VGND sg13g2_fill_2
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_42_242 VPWR VGND sg13g2_decap_8
XFILLER_31_905 VPWR VGND sg13g2_decap_8
XFILLER_6_187 VPWR VGND sg13g2_fill_1
XFILLER_40_7 VPWR VGND sg13g2_fill_2
XFILLER_3_861 VPWR VGND sg13g2_decap_8
X_2250_ _0674_ _0651_ _0672_ VPWR VGND sg13g2_nand2_1
X_2181_ _0607_ _1218_ ppwm_i.u_ppwm.global_counter\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_38_526 VPWR VGND sg13g2_decap_8
XFILLER_19_751 VPWR VGND sg13g2_decap_4
XFILLER_38_559 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_34_721 VPWR VGND sg13g2_decap_8
XFILLER_22_905 VPWR VGND sg13g2_decap_8
XFILLER_15_990 VPWR VGND sg13g2_decap_8
XFILLER_33_264 VPWR VGND sg13g2_decap_8
XFILLER_34_798 VPWR VGND sg13g2_decap_8
X_1965_ net553 VPWR _0029_ VGND _0412_ _0414_ sg13g2_o21ai_1
XFILLER_30_993 VPWR VGND sg13g2_decap_8
X_1896_ sdr_i.mac2.products_ff\[1\] sdr_i.mac2.products_ff\[18\] _0411_ VPWR VGND
+ sg13g2_xor2_1
X_2517_ net436 VPWR _0925_ VGND _0921_ _0924_ sg13g2_o21ai_1
X_2448_ VPWR VGND _1309_ _1219_ _1306_ net508 _0862_ _1302_ sg13g2_a221oi_1
X_2379_ net390 VPWR _0797_ VGND ppwm_i.u_ppwm.pwm_value\[5\] net505 sg13g2_o21ai_1
XFILLER_29_537 VPWR VGND sg13g2_decap_8
XFILLER_25_721 VPWR VGND sg13g2_decap_8
XFILLER_13_927 VPWR VGND sg13g2_decap_8
XFILLER_24_286 VPWR VGND sg13g2_fill_2
XFILLER_25_787 VPWR VGND sg13g2_fill_2
XFILLER_12_448 VPWR VGND sg13g2_decap_4
XFILLER_21_982 VPWR VGND sg13g2_decap_8
XFILLER_20_492 VPWR VGND sg13g2_decap_8
XFILLER_4_614 VPWR VGND sg13g2_decap_4
XFILLER_4_647 VPWR VGND sg13g2_decap_4
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_864 VPWR VGND sg13g2_decap_8
XFILLER_48_835 VPWR VGND sg13g2_decap_8
Xhold8 sdr_i.mac2.sum_lvl2_ff\[8\] VPWR VGND net208 sg13g2_dlygate4sd3_1
XFILLER_47_389 VPWR VGND sg13g2_decap_8
XFILLER_28_570 VPWR VGND sg13g2_decap_8
XFILLER_43_562 VPWR VGND sg13g2_decap_8
XFILLER_43_540 VPWR VGND sg13g2_fill_2
XFILLER_31_779 VPWR VGND sg13g2_decap_8
X_1750_ VPWR VGND _1153_ net510 net447 _1132_ _1317_ net450 sg13g2_a221oi_1
XFILLER_12_982 VPWR VGND sg13g2_decap_8
X_1681_ VPWR _1252_ ppwm_i.u_ppwm.global_counter\[18\] VGND sg13g2_inv_1
XFILLER_8_986 VPWR VGND sg13g2_decap_8
XFILLER_7_485 VPWR VGND sg13g2_fill_1
Xhold408 ppwm_i.u_ppwm.pc\[0\] VPWR VGND net788 sg13g2_dlygate4sd3_1
Xhold419 _0165_ VPWR VGND net799 sg13g2_dlygate4sd3_1
X_3420_ net549 net7 VPWR VGND sg13g2_buf_1
X_2302_ net387 _0697_ _0724_ VPWR VGND sg13g2_nor2_1
XFILLER_39_813 VPWR VGND sg13g2_decap_8
X_2233_ net384 _0656_ _0657_ VPWR VGND sg13g2_nor2_1
X_2164_ _0590_ ppwm_i.u_ppwm.pwm_value\[0\] ppwm_i.u_ppwm.global_counter\[0\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_19_570 VPWR VGND sg13g2_decap_8
XFILLER_19_592 VPWR VGND sg13g2_decap_8
X_2095_ net397 net515 _0524_ VPWR VGND sg13g2_xor2_1
XFILLER_0_82 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_decap_4
XFILLER_21_212 VPWR VGND sg13g2_decap_8
XFILLER_22_757 VPWR VGND sg13g2_decap_8
X_2997_ net153 VGND VPWR net567 ppwm_i.u_ppwm.period_start clknet_leaf_20_clk sg13g2_dfrbpq_2
X_1948_ net743 sdr_i.mac1.sum_lvl2_ff\[5\] _0435_ VPWR VGND sg13g2_xor2_1
XFILLER_30_790 VPWR VGND sg13g2_decap_8
X_1879_ net299 net277 _0046_ VPWR VGND sg13g2_and2_1
XFILLER_0_116 VPWR VGND sg13g2_decap_8
XFILLER_28_89 VPWR VGND sg13g2_decap_8
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_44_348 VPWR VGND sg13g2_decap_8
XFILLER_25_540 VPWR VGND sg13g2_decap_8
XFILLER_25_551 VPWR VGND sg13g2_fill_1
XFILLER_13_724 VPWR VGND sg13g2_decap_8
XFILLER_13_735 VPWR VGND sg13g2_fill_1
XFILLER_40_543 VPWR VGND sg13g2_decap_8
X_3063__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_13_757 VPWR VGND sg13g2_fill_1
XFILLER_8_227 VPWR VGND sg13g2_decap_8
XFILLER_8_216 VPWR VGND sg13g2_decap_8
XFILLER_9_728 VPWR VGND sg13g2_fill_2
XFILLER_21_790 VPWR VGND sg13g2_fill_1
XFILLER_5_923 VPWR VGND sg13g2_decap_8
XFILLER_5_27 VPWR VGND sg13g2_fill_2
XFILLER_4_433 VPWR VGND sg13g2_decap_4
XFILLER_10_8 VPWR VGND sg13g2_fill_1
XFILLER_36_849 VPWR VGND sg13g2_decap_8
XFILLER_44_893 VPWR VGND sg13g2_decap_8
XFILLER_16_562 VPWR VGND sg13g2_decap_8
X_2920_ net521 VGND VPWR _0111_ sdr_i.DP_2.matrix\[73\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_43_392 VPWR VGND sg13g2_decap_8
X_2851_ net290 _0114_ VPWR VGND sg13g2_buf_1
X_2782_ net716 _1070_ _1072_ VPWR VGND sg13g2_and2_1
X_1802_ _0351_ net392 net385 VPWR VGND sg13g2_nand2_2
X_1733_ _1300_ net442 _1142_ net450 _1128_ VPWR VGND sg13g2_a22oi_1
Xhold205 _0250_ VPWR VGND net585 sg13g2_dlygate4sd3_1
Xhold216 ppwm_i.u_ppwm.u_mem.memory\[28\] VPWR VGND net596 sg13g2_dlygate4sd3_1
Xhold227 ppwm_i.u_ppwm.u_mem.memory\[75\] VPWR VGND net607 sg13g2_dlygate4sd3_1
Xhold238 _0237_ VPWR VGND net618 sg13g2_dlygate4sd3_1
Xhold249 _0220_ VPWR VGND net629 sg13g2_dlygate4sd3_1
X_1664_ VPWR _1235_ net715 VGND sg13g2_inv_1
X_1595_ VPWR _1166_ ppwm_i.u_ppwm.u_mem.memory\[43\] VGND sg13g2_inv_1
X_2216_ VGND VPWR net399 _0568_ _0642_ _0551_ sg13g2_a21oi_1
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
X_3196_ net542 VGND VPWR _0046_ sdr_i.mac2.products_ff\[68\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_39_698 VPWR VGND sg13g2_decap_8
XFILLER_27_849 VPWR VGND sg13g2_decap_8
X_2147_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _1256_ _0573_ VPWR VGND sg13g2_nor2_1
X_2078_ net455 _0510_ _0511_ _0185_ VPWR VGND sg13g2_nor3_1
XFILLER_35_871 VPWR VGND sg13g2_decap_8
XFILLER_10_705 VPWR VGND sg13g2_fill_1
XFILLER_30_46 VPWR VGND sg13g2_fill_2
XFILLER_49_407 VPWR VGND sg13g2_decap_8
XFILLER_39_44 VPWR VGND sg13g2_decap_4
XFILLER_44_101 VPWR VGND sg13g2_fill_2
XFILLER_29_164 VPWR VGND sg13g2_decap_8
XFILLER_26_871 VPWR VGND sg13g2_decap_8
XFILLER_13_521 VPWR VGND sg13g2_fill_1
XFILLER_41_885 VPWR VGND sg13g2_decap_8
XFILLER_13_576 VPWR VGND sg13g2_decap_8
XFILLER_5_764 VPWR VGND sg13g2_decap_8
XFILLER_4_252 VPWR VGND sg13g2_fill_2
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_930 VPWR VGND sg13g2_decap_8
XFILLER_0_480 VPWR VGND sg13g2_decap_8
XFILLER_0_491 VPWR VGND sg13g2_fill_1
X_3050_ net50 VGND VPWR net551 ppwm_i.u_ppwm.u_mem.memory\[26\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_48_462 VPWR VGND sg13g2_fill_2
X_2001_ _0462_ net654 net807 _0464_ VPWR VGND sg13g2_a21o_1
XFILLER_35_101 VPWR VGND sg13g2_fill_2
XFILLER_35_112 VPWR VGND sg13g2_decap_4
XFILLER_17_882 VPWR VGND sg13g2_decap_8
XFILLER_16_392 VPWR VGND sg13g2_fill_2
X_2903_ net523 VGND VPWR _0094_ sdr_i.DP_2.matrix\[0\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_32_863 VPWR VGND sg13g2_decap_8
X_2834_ net237 _0097_ VPWR VGND sg13g2_buf_1
X_3077__129 VPWR VGND net129 sg13g2_tiehi
X_2765_ VGND VPWR net479 _1101_ _0322_ _1061_ sg13g2_a21oi_1
X_2696_ net416 VPWR _1027_ VGND net473 ppwm_i.u_ppwm.u_mem.memory\[73\] sg13g2_o21ai_1
X_1716_ net517 net514 _1283_ VPWR VGND sg13g2_nor2b_2
X_1647_ _1218_ net826 VPWR VGND sg13g2_inv_2
Xfanout504 net830 net504 VPWR VGND sg13g2_buf_8
Xfanout515 net825 net515 VPWR VGND sg13g2_buf_8
X_1578_ VPWR _1149_ net619 VGND sg13g2_inv_1
Xfanout548 net1 net548 VPWR VGND sg13g2_buf_2
Xfanout526 net527 net526 VPWR VGND sg13g2_buf_8
Xfanout537 net541 net537 VPWR VGND sg13g2_buf_8
X_3179_ net524 VGND VPWR net203 sdr_i.mac1.sum_lvl2_ff\[8\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_15_808 VPWR VGND sg13g2_fill_2
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_14_329 VPWR VGND sg13g2_fill_2
XFILLER_25_79 VPWR VGND sg13g2_decap_4
XFILLER_35_690 VPWR VGND sg13g2_fill_1
XFILLER_22_395 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_244 VPWR VGND sg13g2_fill_2
XFILLER_49_226 VPWR VGND sg13g2_decap_8
XFILLER_46_955 VPWR VGND sg13g2_decap_8
XFILLER_18_657 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_fill_1
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_33_649 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
XFILLER_9_344 VPWR VGND sg13g2_fill_1
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
XFILLER_5_550 VPWR VGND sg13g2_fill_1
X_2550_ net429 VPWR _0954_ VGND net495 ppwm_i.u_ppwm.u_mem.memory\[0\] sg13g2_o21ai_1
X_2481_ VGND VPWR _1226_ net383 _0892_ _0672_ sg13g2_a21oi_1
X_3102_ net31 VGND VPWR net365 ppwm_i.u_ppwm.u_mem.memory\[78\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_37_900 VPWR VGND sg13g2_decap_8
X_3033_ net83 VGND VPWR _0224_ ppwm_i.u_ppwm.u_mem.memory\[9\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
XFILLER_37_977 VPWR VGND sg13g2_decap_8
XFILLER_20_822 VPWR VGND sg13g2_fill_1
XFILLER_20_877 VPWR VGND sg13g2_decap_8
X_2817_ net273 _0080_ VPWR VGND sg13g2_buf_1
X_2748_ net418 VPWR _1053_ VGND net478 ppwm_i.u_ppwm.u_mem.memory\[99\] sg13g2_o21ai_1
X_2679_ VGND VPWR net477 _1144_ _0279_ _1018_ sg13g2_a21oi_1
Xfanout389 _0348_ net389 VPWR VGND sg13g2_buf_2
Xfanout378 _0684_ net378 VPWR VGND sg13g2_buf_8
XFILLER_46_218 VPWR VGND sg13g2_decap_8
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_36_78 VPWR VGND sg13g2_decap_8
XFILLER_11_800 VPWR VGND sg13g2_decap_8
XFILLER_23_660 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_fill_2
XFILLER_23_671 VPWR VGND sg13g2_fill_1
XFILLER_6_325 VPWR VGND sg13g2_decap_8
XFILLER_11_888 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_410 VPWR VGND sg13g2_fill_1
XFILLER_46_730 VPWR VGND sg13g2_fill_1
XFILLER_19_944 VPWR VGND sg13g2_decap_8
XFILLER_34_903 VPWR VGND sg13g2_decap_8
XFILLER_45_284 VPWR VGND sg13g2_decap_4
XFILLER_21_619 VPWR VGND sg13g2_decap_8
X_2982__182 VPWR VGND net182 sg13g2_tiehi
X_1981_ _0453_ _0452_ _0049_ VPWR VGND sg13g2_xor2_1
XFILLER_14_660 VPWR VGND sg13g2_fill_2
XFILLER_14_693 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_40_clk clknet_3_4__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_2602_ net432 VPWR _0980_ VGND net500 ppwm_i.u_ppwm.u_mem.memory\[26\] sg13g2_o21ai_1
X_2533_ VGND VPWR _0900_ _0936_ _0939_ _0938_ sg13g2_a21oi_1
XFILLER_6_870 VPWR VGND sg13g2_decap_8
X_2464_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] net407 net405 _0876_ VPWR VGND sg13g2_or3_1
X_2395_ net423 VPWR _0813_ VGND _0802_ _0811_ sg13g2_o21ai_1
XFILLER_3_1022 VPWR VGND sg13g2_decap_8
X_3131__76 VPWR VGND net76 sg13g2_tiehi
X_3016_ net116 VGND VPWR _0207_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
XFILLER_37_774 VPWR VGND sg13g2_decap_8
XFILLER_25_936 VPWR VGND sg13g2_decap_8
XFILLER_40_906 VPWR VGND sg13g2_decap_8
XFILLER_24_446 VPWR VGND sg13g2_fill_1
XFILLER_20_630 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_31_clk clknet_3_5__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
XFILLER_4_818 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_fill_2
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_16_969 VPWR VGND sg13g2_decap_8
XFILLER_24_980 VPWR VGND sg13g2_decap_8
XFILLER_30_438 VPWR VGND sg13g2_decap_8
XFILLER_11_630 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_22_clk clknet_3_6__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_6_111 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_decap_8
XFILLER_3_840 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_fill_2
X_2180_ _1212_ ppwm_i.u_ppwm.global_counter\[7\] _0606_ VPWR VGND sg13g2_nor2_1
XFILLER_2_394 VPWR VGND sg13g2_decap_4
XFILLER_19_774 VPWR VGND sg13g2_decap_4
XFILLER_34_700 VPWR VGND sg13g2_decap_8
XFILLER_46_593 VPWR VGND sg13g2_decap_8
XFILLER_33_243 VPWR VGND sg13g2_decap_8
X_1964_ _0443_ _0442_ _0061_ VPWR VGND sg13g2_xor2_1
XFILLER_21_449 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_13_clk clknet_3_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
XFILLER_30_972 VPWR VGND sg13g2_decap_8
X_1895_ net254 sdr_i.mac2.products_ff\[17\] _0032_ VPWR VGND sg13g2_xor2_1
X_2516_ _0807_ net374 _0805_ _0924_ VPWR VGND _0923_ sg13g2_nand4_1
X_2447_ _0861_ net374 VPWR VGND sg13g2_inv_2
X_2378_ _0796_ net504 net391 VPWR VGND sg13g2_xnor2_1
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_17_25 VPWR VGND sg13g2_fill_1
XFILLER_17_58 VPWR VGND sg13g2_decap_4
XFILLER_13_906 VPWR VGND sg13g2_decap_8
XFILLER_25_766 VPWR VGND sg13g2_decap_8
XFILLER_33_13 VPWR VGND sg13g2_fill_1
XFILLER_21_961 VPWR VGND sg13g2_decap_8
XFILLER_3_114 VPWR VGND sg13g2_decap_8
XFILLER_0_843 VPWR VGND sg13g2_decap_8
XFILLER_48_814 VPWR VGND sg13g2_decap_8
Xhold9 sdr_i.mac2.sum_lvl2_ff\[9\] VPWR VGND net209 sg13g2_dlygate4sd3_1
XFILLER_47_335 VPWR VGND sg13g2_fill_2
XFILLER_15_221 VPWR VGND sg13g2_decap_4
XFILLER_16_766 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_fill_1
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_30_279 VPWR VGND sg13g2_fill_2
XFILLER_8_965 VPWR VGND sg13g2_decap_8
X_1680_ VPWR _1251_ ppwm_i.u_ppwm.global_counter\[19\] VGND sg13g2_inv_1
Xhold409 ppwm_i.u_ppwm.global_counter\[3\] VPWR VGND net789 sg13g2_dlygate4sd3_1
X_2301_ VPWR _0723_ _0722_ VGND sg13g2_inv_1
XFILLER_3_681 VPWR VGND sg13g2_fill_2
XFILLER_3_670 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2232_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] ppwm_i.u_ppwm.pwm_value\[2\] net398 _0656_
+ VPWR VGND sg13g2_mux2_1
XFILLER_39_869 VPWR VGND sg13g2_decap_8
X_2163_ ppwm_i.u_ppwm.pwm_value\[1\] ppwm_i.u_ppwm.global_counter\[1\] _0589_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_38_346 VPWR VGND sg13g2_fill_2
XFILLER_38_379 VPWR VGND sg13g2_decap_4
XFILLER_0_61 VPWR VGND sg13g2_decap_8
X_3101__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_0_1025 VPWR VGND sg13g2_decap_4
X_2094_ net515 net396 _0523_ VPWR VGND sg13g2_and2_1
XFILLER_34_552 VPWR VGND sg13g2_decap_8
XFILLER_10_909 VPWR VGND sg13g2_decap_8
XFILLER_22_747 VPWR VGND sg13g2_decap_4
X_2996_ net155 VGND VPWR _0187_ ppwm_i.u_ppwm.u_pwm.counter\[9\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
X_1947_ net305 sdr_i.mac1.sum_lvl2_ff\[4\] _0027_ VPWR VGND sg13g2_xor2_1
X_1878_ net282 net283 _0044_ VPWR VGND sg13g2_and2_1
XFILLER_45_828 VPWR VGND sg13g2_decap_8
XFILLER_17_508 VPWR VGND sg13g2_decap_8
XFILLER_28_68 VPWR VGND sg13g2_decap_8
XFILLER_29_357 VPWR VGND sg13g2_decap_4
XFILLER_13_703 VPWR VGND sg13g2_fill_1
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_40_577 VPWR VGND sg13g2_fill_2
X_3104__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_20_290 VPWR VGND sg13g2_decap_4
XFILLER_4_412 VPWR VGND sg13g2_decap_8
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_0_662 VPWR VGND sg13g2_fill_2
XFILLER_47_121 VPWR VGND sg13g2_decap_8
XFILLER_36_828 VPWR VGND sg13g2_decap_8
XFILLER_18_90 VPWR VGND sg13g2_decap_8
XFILLER_44_872 VPWR VGND sg13g2_decap_8
X_2850_ net223 _0113_ VPWR VGND sg13g2_buf_1
XFILLER_43_382 VPWR VGND sg13g2_fill_1
XFILLER_31_544 VPWR VGND sg13g2_fill_1
XFILLER_15_1011 VPWR VGND sg13g2_decap_8
X_1801_ net390 net387 _0350_ VPWR VGND sg13g2_nor2_2
XFILLER_8_740 VPWR VGND sg13g2_decap_8
X_2781_ net716 _1070_ _1071_ VPWR VGND sg13g2_nor2_1
X_1732_ VPWR VGND _1107_ _1298_ net438 _1100_ _1299_ net450 sg13g2_a221oi_1
X_1663_ VPWR _1234_ net752 VGND sg13g2_inv_1
Xhold217 ppwm_i.u_ppwm.u_mem.memory\[95\] VPWR VGND net597 sg13g2_dlygate4sd3_1
Xhold206 ppwm_i.u_ppwm.u_mem.memory\[25\] VPWR VGND net586 sg13g2_dlygate4sd3_1
Xhold239 ppwm_i.u_ppwm.u_mem.memory\[60\] VPWR VGND net619 sg13g2_dlygate4sd3_1
Xhold228 _0289_ VPWR VGND net608 sg13g2_dlygate4sd3_1
X_1594_ VPWR _1165_ net356 VGND sg13g2_inv_1
X_2215_ _0641_ net402 _0640_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_644 VPWR VGND sg13g2_fill_2
X_3195_ net540 VGND VPWR _0065_ sdr_i.mac2.products_ff\[52\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_39_666 VPWR VGND sg13g2_decap_8
XFILLER_27_828 VPWR VGND sg13g2_decap_8
XFILLER_26_338 VPWR VGND sg13g2_fill_2
X_2146_ _0572_ _1258_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _1257_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2077_ net819 net808 net520 _0504_ _0511_ VPWR VGND sg13g2_and4_1
XFILLER_35_850 VPWR VGND sg13g2_decap_8
XFILLER_22_500 VPWR VGND sg13g2_decap_8
X_2979_ net188 VGND VPWR net795 ppwm_i.u_ppwm.u_pwm.cmp_value\[2\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_2_949 VPWR VGND sg13g2_decap_8
XFILLER_29_132 VPWR VGND sg13g2_decap_4
XFILLER_45_625 VPWR VGND sg13g2_fill_1
XFILLER_45_614 VPWR VGND sg13g2_decap_8
XFILLER_45_647 VPWR VGND sg13g2_decap_4
XFILLER_17_338 VPWR VGND sg13g2_fill_2
XFILLER_26_850 VPWR VGND sg13g2_decap_8
XFILLER_13_500 VPWR VGND sg13g2_fill_1
XFILLER_38_1022 VPWR VGND sg13g2_decap_8
XFILLER_41_864 VPWR VGND sg13g2_decap_8
XFILLER_40_341 VPWR VGND sg13g2_decap_4
XFILLER_40_330 VPWR VGND sg13g2_decap_8
XFILLER_5_743 VPWR VGND sg13g2_decap_8
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_49_986 VPWR VGND sg13g2_decap_8
X_2000_ net654 _0462_ net807 _0463_ VPWR VGND sg13g2_nand3_1
X_2902_ net521 VGND VPWR _0093_ sdr_i.DP_1.matrix\[73\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_32_842 VPWR VGND sg13g2_decap_8
XFILLER_31_330 VPWR VGND sg13g2_decap_4
X_2833_ net274 _0096_ VPWR VGND sg13g2_buf_1
X_2764_ net420 VPWR _1061_ VGND net479 net612 sg13g2_o21ai_1
X_1715_ net514 net517 _1282_ VPWR VGND sg13g2_nor2b_2
X_2695_ VGND VPWR net479 _1136_ _0287_ _1026_ sg13g2_a21oi_1
XFILLER_6_60 VPWR VGND sg13g2_decap_8
X_1646_ _1217_ net811 VPWR VGND sg13g2_inv_2
X_1577_ VPWR _1148_ net590 VGND sg13g2_inv_1
Xfanout505 net838 net505 VPWR VGND sg13g2_buf_8
Xfanout538 net540 net538 VPWR VGND sg13g2_buf_8
Xfanout516 ppwm_i.u_ppwm.pc\[1\] net516 VPWR VGND sg13g2_buf_2
Xfanout527 net547 net527 VPWR VGND sg13g2_buf_8
Xfanout549 net1 net549 VPWR VGND sg13g2_buf_1
XFILLER_39_485 VPWR VGND sg13g2_decap_4
X_3178_ net531 VGND VPWR net747 sdr_i.mac1.sum_lvl2_ff\[5\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2129_ net507 ppwm_i.u_ppwm.global_counter\[11\] _0555_ VPWR VGND sg13g2_nor2b_1
XFILLER_14_308 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_4
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_41_138 VPWR VGND sg13g2_decap_8
X_3021__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_10_514 VPWR VGND sg13g2_fill_1
XFILLER_22_374 VPWR VGND sg13g2_decap_8
XFILLER_10_569 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_fill_1
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_49_205 VPWR VGND sg13g2_decap_8
XFILLER_46_934 VPWR VGND sg13g2_decap_8
XFILLER_18_636 VPWR VGND sg13g2_decap_8
XFILLER_33_628 VPWR VGND sg13g2_decap_4
XFILLER_41_650 VPWR VGND sg13g2_decap_4
XFILLER_9_301 VPWR VGND sg13g2_fill_2
XFILLER_14_886 VPWR VGND sg13g2_decap_8
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
X_2480_ _0889_ _0890_ net378 _0891_ VPWR VGND sg13g2_nand3_1
XFILLER_49_5 VPWR VGND sg13g2_decap_8
X_3101_ net35 VGND VPWR net653 ppwm_i.u_ppwm.u_mem.memory\[77\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_49_783 VPWR VGND sg13g2_decap_8
X_3032_ net85 VGND VPWR net562 ppwm_i.u_ppwm.u_mem.memory\[8\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_36_411 VPWR VGND sg13g2_fill_1
XFILLER_37_956 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_4
XFILLER_36_455 VPWR VGND sg13g2_decap_8
XFILLER_17_691 VPWR VGND sg13g2_decap_8
X_2816_ net220 _0079_ VPWR VGND sg13g2_buf_1
XFILLER_20_845 VPWR VGND sg13g2_decap_4
X_2747_ VGND VPWR net476 _1110_ _0313_ _1052_ sg13g2_a21oi_1
X_2678_ net417 VPWR _1018_ VGND net477 ppwm_i.u_ppwm.u_mem.memory\[64\] sg13g2_o21ai_1
X_1629_ VPWR _1200_ net561 VGND sg13g2_inv_1
X_3170__195 VPWR VGND net195 sg13g2_tiehi
Xfanout379 _0653_ net379 VPWR VGND sg13g2_buf_8
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_36_57 VPWR VGND sg13g2_decap_8
XFILLER_14_105 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_fill_2
XFILLER_15_639 VPWR VGND sg13g2_decap_8
XFILLER_14_149 VPWR VGND sg13g2_fill_2
XFILLER_11_823 VPWR VGND sg13g2_fill_1
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_10_344 VPWR VGND sg13g2_fill_1
XFILLER_10_311 VPWR VGND sg13g2_fill_2
XFILLER_42_1007 VPWR VGND sg13g2_decap_8
XFILLER_19_923 VPWR VGND sg13g2_decap_8
XFILLER_45_263 VPWR VGND sg13g2_fill_2
XFILLER_18_499 VPWR VGND sg13g2_fill_2
XFILLER_34_959 VPWR VGND sg13g2_decap_8
X_1980_ _0453_ net311 net244 VPWR VGND sg13g2_nand2_1
XFILLER_14_650 VPWR VGND sg13g2_fill_1
XFILLER_33_447 VPWR VGND sg13g2_decap_4
XFILLER_14_672 VPWR VGND sg13g2_decap_8
XFILLER_41_480 VPWR VGND sg13g2_fill_1
XFILLER_9_197 VPWR VGND sg13g2_decap_4
X_2601_ VGND VPWR net497 _1183_ _0240_ _0979_ sg13g2_a21oi_1
X_2532_ _0938_ _0917_ _0937_ VPWR VGND sg13g2_nand2_1
XFILLER_47_2 VPWR VGND sg13g2_fill_1
X_2463_ _0867_ _0862_ _0868_ _0875_ VPWR VGND sg13g2_a21o_2
X_2394_ net504 net371 _0812_ VPWR VGND sg13g2_nor2_1
XFILLER_3_83 VPWR VGND sg13g2_decap_4
XFILLER_3_1001 VPWR VGND sg13g2_decap_8
X_3015_ net118 VGND VPWR _0206_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_25_915 VPWR VGND sg13g2_decap_8
XFILLER_36_274 VPWR VGND sg13g2_decap_4
XFILLER_20_664 VPWR VGND sg13g2_fill_1
XFILLER_22_48 VPWR VGND sg13g2_decap_8
XFILLER_3_318 VPWR VGND sg13g2_fill_2
XFILLER_47_528 VPWR VGND sg13g2_decap_4
XFILLER_19_219 VPWR VGND sg13g2_fill_1
XFILLER_28_720 VPWR VGND sg13g2_decap_8
XFILLER_28_753 VPWR VGND sg13g2_decap_4
XFILLER_28_775 VPWR VGND sg13g2_decap_8
XFILLER_15_414 VPWR VGND sg13g2_fill_1
XFILLER_16_948 VPWR VGND sg13g2_decap_8
XFILLER_43_789 VPWR VGND sg13g2_decap_8
XFILLER_42_288 VPWR VGND sg13g2_decap_8
XFILLER_11_642 VPWR VGND sg13g2_decap_8
XFILLER_11_664 VPWR VGND sg13g2_decap_8
XFILLER_10_163 VPWR VGND sg13g2_fill_1
XFILLER_3_896 VPWR VGND sg13g2_decap_8
XFILLER_2_362 VPWR VGND sg13g2_fill_2
XFILLER_19_720 VPWR VGND sg13g2_decap_8
XFILLER_19_731 VPWR VGND sg13g2_fill_2
XFILLER_46_550 VPWR VGND sg13g2_decap_8
XFILLER_21_428 VPWR VGND sg13g2_decap_8
X_1963_ _0443_ net296 net219 VPWR VGND sg13g2_nand2_1
XFILLER_30_951 VPWR VGND sg13g2_decap_8
X_1894_ _0410_ net757 net254 VPWR VGND sg13g2_nand2_1
X_2515_ _0922_ VPWR _0923_ VGND net381 _0809_ sg13g2_o21ai_1
X_2446_ _0860_ net768 _0681_ _0859_ VPWR VGND sg13g2_and3_2
XFILLER_25_1013 VPWR VGND sg13g2_decap_8
X_2377_ _1223_ net391 _0795_ VPWR VGND sg13g2_nor2_1
XFILLER_17_37 VPWR VGND sg13g2_decap_8
XFILLER_37_561 VPWR VGND sg13g2_fill_2
XFILLER_21_940 VPWR VGND sg13g2_decap_8
XFILLER_24_288 VPWR VGND sg13g2_fill_1
XFILLER_32_1017 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_137 VPWR VGND sg13g2_fill_1
XFILLER_0_822 VPWR VGND sg13g2_decap_8
XFILLER_0_899 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_decap_8
XFILLER_15_266 VPWR VGND sg13g2_decap_8
XFILLER_31_726 VPWR VGND sg13g2_fill_1
XFILLER_43_597 VPWR VGND sg13g2_fill_1
XFILLER_12_940 VPWR VGND sg13g2_decap_8
XFILLER_15_299 VPWR VGND sg13g2_fill_2
XFILLER_30_258 VPWR VGND sg13g2_decap_4
XFILLER_8_944 VPWR VGND sg13g2_decap_8
XFILLER_23_91 VPWR VGND sg13g2_decap_4
X_3031__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_48_1024 VPWR VGND sg13g2_decap_4
X_2300_ net502 ppwm_i.u_ppwm.pwm_value\[6\] net399 _0722_ VPWR VGND sg13g2_mux2_1
X_2231_ VGND VPWR _0654_ _0655_ net400 net507 sg13g2_a21oi_2
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_848 VPWR VGND sg13g2_decap_8
X_2162_ _0588_ _1227_ ppwm_i.u_ppwm.global_counter\[2\] VPWR VGND sg13g2_nand2_1
X_2093_ net518 net401 _0522_ VPWR VGND sg13g2_and2_1
XFILLER_0_1004 VPWR VGND sg13g2_decap_8
XFILLER_34_542 VPWR VGND sg13g2_decap_4
X_2995_ net157 VGND VPWR _0186_ ppwm_i.u_ppwm.u_pwm.counter\[8\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
X_1946_ _0434_ sdr_i.mac1.sum_lvl2_ff\[4\] net305 VPWR VGND sg13g2_nand2_1
X_1877_ net304 net275 _0042_ VPWR VGND sg13g2_and2_1
XFILLER_1_608 VPWR VGND sg13g2_decap_8
XFILLER_1_619 VPWR VGND sg13g2_fill_2
X_2429_ _0844_ _1220_ net391 VPWR VGND sg13g2_xnor2_1
XFILLER_45_807 VPWR VGND sg13g2_decap_8
XFILLER_29_347 VPWR VGND sg13g2_fill_1
XFILLER_25_564 VPWR VGND sg13g2_fill_2
XFILLER_40_512 VPWR VGND sg13g2_decap_8
XFILLER_25_597 VPWR VGND sg13g2_fill_2
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_5_29 VPWR VGND sg13g2_fill_1
X_3070__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_645 VPWR VGND sg13g2_fill_1
XFILLER_47_100 VPWR VGND sg13g2_decap_8
XFILLER_0_696 VPWR VGND sg13g2_decap_8
XFILLER_36_807 VPWR VGND sg13g2_decap_8
XFILLER_29_892 VPWR VGND sg13g2_decap_8
XFILLER_44_851 VPWR VGND sg13g2_decap_8
XFILLER_43_361 VPWR VGND sg13g2_fill_1
XFILLER_43_350 VPWR VGND sg13g2_decap_8
XFILLER_43_372 VPWR VGND sg13g2_fill_1
X_1800_ VGND VPWR _0349_ _0347_ _0341_ sg13g2_or2_1
X_2780_ _1067_ net340 _1070_ _0328_ VPWR VGND sg13g2_nor3_1
X_1731_ ppwm_i.u_ppwm.u_mem.memory\[88\] net515 net518 _1298_ VPWR VGND sg13g2_nor3_1
XFILLER_8_796 VPWR VGND sg13g2_decap_4
X_1662_ VPWR _1233_ net512 VGND sg13g2_inv_1
Xhold207 _0239_ VPWR VGND net587 sg13g2_dlygate4sd3_1
X_2979__188 VPWR VGND net188 sg13g2_tiehi
Xhold218 _0309_ VPWR VGND net598 sg13g2_dlygate4sd3_1
Xhold229 ppwm_i.u_ppwm.u_mem.memory\[13\] VPWR VGND net609 sg13g2_dlygate4sd3_1
X_1593_ VPWR _1164_ net611 VGND sg13g2_inv_1
XFILLER_39_601 VPWR VGND sg13g2_decap_4
X_2214_ VPWR VGND _0584_ _0551_ _0583_ _1210_ _0640_ ppwm_i.u_ppwm.global_counter\[19\]
+ sg13g2_a221oi_1
X_3194_ net540 VGND VPWR _0064_ sdr_i.mac2.products_ff\[51\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_38_100 VPWR VGND sg13g2_decap_8
X_2145_ _0570_ VPWR _0571_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _1258_ sg13g2_o21ai_1
X_2076_ _1237_ _0509_ _0510_ VPWR VGND sg13g2_and2_1
XFILLER_38_199 VPWR VGND sg13g2_decap_8
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_34_372 VPWR VGND sg13g2_decap_4
XFILLER_22_556 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_fill_2
X_2978_ net190 VGND VPWR net579 ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_1929_ _0018_ _0424_ _0425_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_48 VPWR VGND sg13g2_fill_1
XFILLER_2_928 VPWR VGND sg13g2_decap_8
XFILLER_29_111 VPWR VGND sg13g2_fill_1
XFILLER_17_317 VPWR VGND sg13g2_decap_8
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_41_843 VPWR VGND sg13g2_decap_8
XFILLER_25_372 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_fill_2
XFILLER_5_700 VPWR VGND sg13g2_decap_8
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_decap_8
XFILLER_48_431 VPWR VGND sg13g2_fill_2
Xhold90 sdr_i.DP_3.matrix\[9\] VPWR VGND net290 sg13g2_dlygate4sd3_1
XFILLER_35_103 VPWR VGND sg13g2_fill_1
XFILLER_35_136 VPWR VGND sg13g2_fill_2
XFILLER_36_659 VPWR VGND sg13g2_fill_2
XFILLER_44_692 VPWR VGND sg13g2_decap_8
X_2901_ net521 VGND VPWR _0092_ sdr_i.DP_1.matrix\[72\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_32_821 VPWR VGND sg13g2_decap_8
XFILLER_31_353 VPWR VGND sg13g2_decap_8
X_2832_ net252 _0095_ VPWR VGND sg13g2_buf_1
XFILLER_32_898 VPWR VGND sg13g2_decap_8
X_2763_ VGND VPWR net480 _1102_ _0321_ _1060_ sg13g2_a21oi_1
X_1714_ ppwm_i.u_ppwm.u_mem.memory\[87\] net515 net518 _1281_ VPWR VGND sg13g2_nor3_1
X_2694_ net417 VPWR _1026_ VGND net477 net559 sg13g2_o21ai_1
XFILLER_6_83 VPWR VGND sg13g2_decap_8
X_1645_ _1216_ net816 VPWR VGND sg13g2_inv_2
X_2992__163 VPWR VGND net163 sg13g2_tiehi
X_1576_ VPWR _1147_ net660 VGND sg13g2_inv_1
Xfanout506 net770 net506 VPWR VGND sg13g2_buf_8
Xfanout539 net540 net539 VPWR VGND sg13g2_buf_8
Xfanout528 net530 net528 VPWR VGND sg13g2_buf_8
Xfanout517 net519 net517 VPWR VGND sg13g2_buf_8
XFILLER_6_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_464 VPWR VGND sg13g2_fill_2
X_3177_ net531 VGND VPWR net268 sdr_i.mac1.sum_lvl2_ff\[4\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_2128_ _0554_ net507 ppwm_i.u_ppwm.global_counter\[11\] VPWR VGND sg13g2_nand2b_1
XFILLER_42_629 VPWR VGND sg13g2_fill_1
XFILLER_42_607 VPWR VGND sg13g2_fill_1
X_2059_ _0499_ net715 net707 net769 VPWR VGND sg13g2_and3_1
XFILLER_23_887 VPWR VGND sg13g2_decap_8
XFILLER_10_548 VPWR VGND sg13g2_decap_8
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_1_246 VPWR VGND sg13g2_fill_1
XFILLER_46_913 VPWR VGND sg13g2_decap_8
XFILLER_45_401 VPWR VGND sg13g2_decap_4
XFILLER_26_670 VPWR VGND sg13g2_decap_8
XFILLER_41_695 VPWR VGND sg13g2_decap_8
XFILLER_40_150 VPWR VGND sg13g2_decap_8
XFILLER_9_313 VPWR VGND sg13g2_decap_8
XFILLER_13_353 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_9_357 VPWR VGND sg13g2_fill_2
XFILLER_5_530 VPWR VGND sg13g2_decap_4
X_3100_ net39 VGND VPWR _0291_ ppwm_i.u_ppwm.u_mem.memory\[76\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_49_762 VPWR VGND sg13g2_decap_8
X_3031_ net87 VGND VPWR net693 ppwm_i.u_ppwm.u_mem.memory\[7\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_37_935 VPWR VGND sg13g2_decap_8
XFILLER_48_283 VPWR VGND sg13g2_fill_1
XFILLER_48_272 VPWR VGND sg13g2_decap_8
XFILLER_36_423 VPWR VGND sg13g2_decap_4
X_3056__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_17_670 VPWR VGND sg13g2_decap_8
XFILLER_23_128 VPWR VGND sg13g2_decap_8
XFILLER_24_629 VPWR VGND sg13g2_fill_1
X_3124__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_32_684 VPWR VGND sg13g2_decap_8
X_2815_ net285 _0078_ VPWR VGND sg13g2_buf_1
XFILLER_9_891 VPWR VGND sg13g2_decap_8
X_2746_ net416 VPWR _1052_ VGND net476 ppwm_i.u_ppwm.u_mem.memory\[98\] sg13g2_o21ai_1
X_2677_ VGND VPWR net473 _1145_ _0278_ _1017_ sg13g2_a21oi_1
X_1628_ VPWR _1199_ net642 VGND sg13g2_inv_1
X_1559_ VPWR _1130_ net364 VGND sg13g2_inv_1
XFILLER_46_209 VPWR VGND sg13g2_decap_4
X_3229_ net525 VGND VPWR net260 sdr_i.mac2.total_sum\[0\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_15_607 VPWR VGND sg13g2_decap_4
XFILLER_23_640 VPWR VGND sg13g2_fill_2
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_10_367 VPWR VGND sg13g2_fill_1
XFILLER_2_500 VPWR VGND sg13g2_decap_4
Xhold390 ppwm_i.u_ppwm.pwm_value\[3\] VPWR VGND net770 sg13g2_dlygate4sd3_1
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_46_787 VPWR VGND sg13g2_decap_8
XFILLER_45_242 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_33_404 VPWR VGND sg13g2_decap_8
XFILLER_34_938 VPWR VGND sg13g2_decap_8
XFILLER_42_993 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_fill_1
XFILLER_9_176 VPWR VGND sg13g2_decap_8
X_2600_ net433 VPWR _0979_ VGND net497 net586 sg13g2_o21ai_1
X_2531_ net390 VPWR _0937_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] net502 sg13g2_o21ai_1
X_2462_ VPWR VGND _0701_ net458 _0874_ _1218_ _0206_ net370 sg13g2_a221oi_1
X_2393_ _0805_ _0807_ _0683_ _0811_ VPWR VGND _0810_ sg13g2_nand4_1
XFILLER_3_62 VPWR VGND sg13g2_decap_8
XFILLER_49_581 VPWR VGND sg13g2_decap_8
X_3014_ net120 VGND VPWR _0205_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_2
XFILLER_24_459 VPWR VGND sg13g2_decap_8
XFILLER_33_993 VPWR VGND sg13g2_decap_8
XFILLER_32_481 VPWR VGND sg13g2_decap_8
XFILLER_22_27 VPWR VGND sg13g2_decap_8
X_2729_ VGND VPWR net464 _1119_ _0304_ _1043_ sg13g2_a21oi_1
XFILLER_47_507 VPWR VGND sg13g2_decap_8
XFILLER_47_79 VPWR VGND sg13g2_decap_8
XFILLER_28_732 VPWR VGND sg13g2_decap_8
XFILLER_27_253 VPWR VGND sg13g2_fill_1
XFILLER_43_724 VPWR VGND sg13g2_decap_8
X_3066__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_16_927 VPWR VGND sg13g2_decap_8
XFILLER_43_768 VPWR VGND sg13g2_decap_8
XFILLER_42_223 VPWR VGND sg13g2_decap_8
XFILLER_31_919 VPWR VGND sg13g2_decap_8
XFILLER_42_256 VPWR VGND sg13g2_decap_8
X_3107__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_30_418 VPWR VGND sg13g2_fill_2
XFILLER_23_492 VPWR VGND sg13g2_decap_4
X_3028__93 VPWR VGND net93 sg13g2_tiehi
X_3043__63 VPWR VGND net63 sg13g2_tiehi
X_3073__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_3_875 VPWR VGND sg13g2_decap_8
XFILLER_18_275 VPWR VGND sg13g2_decap_8
XFILLER_22_919 VPWR VGND sg13g2_decap_8
X_1962_ _0442_ net290 net222 VPWR VGND sg13g2_nand2_1
XFILLER_42_790 VPWR VGND sg13g2_decap_8
XFILLER_30_930 VPWR VGND sg13g2_decap_8
X_1893_ _0037_ _0408_ net755 VPWR VGND sg13g2_xnor2_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2514_ VGND VPWR _1223_ net381 _0922_ _0672_ sg13g2_a21oi_1
X_2445_ VGND VPWR _0859_ _0680_ net380 sg13g2_or2_1
X_2376_ _0794_ _0793_ _0200_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_540 VPWR VGND sg13g2_decap_8
XFILLER_25_735 VPWR VGND sg13g2_decap_8
XFILLER_24_212 VPWR VGND sg13g2_decap_4
XFILLER_37_595 VPWR VGND sg13g2_fill_2
XFILLER_40_705 VPWR VGND sg13g2_decap_4
XFILLER_33_790 VPWR VGND sg13g2_decap_8
XFILLER_21_996 VPWR VGND sg13g2_decap_8
XFILLER_0_801 VPWR VGND sg13g2_decap_8
XFILLER_0_878 VPWR VGND sg13g2_decap_8
XFILLER_48_849 VPWR VGND sg13g2_decap_8
XFILLER_47_326 VPWR VGND sg13g2_fill_1
XFILLER_28_584 VPWR VGND sg13g2_fill_2
XFILLER_31_705 VPWR VGND sg13g2_decap_8
XFILLER_30_237 VPWR VGND sg13g2_decap_8
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_48_1003 VPWR VGND sg13g2_decap_8
XFILLER_2_171 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_fill_2
X_2230_ _1218_ net398 _0654_ VPWR VGND sg13g2_nor2_1
XFILLER_39_827 VPWR VGND sg13g2_decap_8
X_2161_ _0587_ ppwm_i.u_ppwm.global_counter\[8\] _1221_ ppwm_i.u_ppwm.global_counter\[9\]
+ _1220_ VPWR VGND sg13g2_a22oi_1
X_2092_ VGND VPWR net518 _0520_ _0189_ _0521_ sg13g2_a21oi_1
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_0_96 VPWR VGND sg13g2_decap_8
XFILLER_22_716 VPWR VGND sg13g2_fill_2
X_2994_ net159 VGND VPWR _0185_ ppwm_i.u_ppwm.u_pwm.counter\[7\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
XFILLER_21_226 VPWR VGND sg13g2_decap_8
X_1945_ _0026_ _0432_ _0433_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_248 VPWR VGND sg13g2_fill_2
XFILLER_21_259 VPWR VGND sg13g2_decap_8
X_1876_ net273 net281 _0040_ VPWR VGND sg13g2_and2_1
X_2428_ _0843_ _0842_ _0203_ VPWR VGND sg13g2_nor2b_1
X_2359_ _0778_ ppwm_i.u_ppwm.pwm_value\[5\] net391 VPWR VGND sg13g2_xnor2_1
XFILLER_38_882 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_25_576 VPWR VGND sg13g2_decap_8
XFILLER_40_579 VPWR VGND sg13g2_fill_1
XFILLER_40_557 VPWR VGND sg13g2_decap_8
XFILLER_5_937 VPWR VGND sg13g2_decap_8
XFILLER_0_675 VPWR VGND sg13g2_decap_8
XFILLER_29_871 VPWR VGND sg13g2_decap_8
XFILLER_35_307 VPWR VGND sg13g2_fill_1
XFILLER_44_830 VPWR VGND sg13g2_decap_8
X_3095__58 VPWR VGND net58 sg13g2_tiehi
XFILLER_16_576 VPWR VGND sg13g2_decap_8
XFILLER_16_587 VPWR VGND sg13g2_fill_2
XFILLER_31_524 VPWR VGND sg13g2_decap_8
XFILLER_8_720 VPWR VGND sg13g2_fill_1
XFILLER_12_771 VPWR VGND sg13g2_fill_1
XFILLER_11_281 VPWR VGND sg13g2_fill_1
XFILLER_11_292 VPWR VGND sg13g2_fill_2
XFILLER_12_793 VPWR VGND sg13g2_decap_8
X_1730_ VGND VPWR _1114_ net442 _1297_ net460 sg13g2_a21oi_1
X_1661_ _1232_ net768 VPWR VGND sg13g2_inv_2
Xhold208 ppwm_i.u_ppwm.u_mem.memory\[15\] VPWR VGND net588 sg13g2_dlygate4sd3_1
XFILLER_7_296 VPWR VGND sg13g2_fill_1
Xhold219 ppwm_i.u_ppwm.u_mem.memory\[24\] VPWR VGND net599 sg13g2_dlygate4sd3_1
X_1592_ VPWR _1163_ net592 VGND sg13g2_inv_1
XFILLER_3_480 VPWR VGND sg13g2_fill_1
X_3193_ net539 VGND VPWR _0063_ sdr_i.mac2.products_ff\[35\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_39_613 VPWR VGND sg13g2_decap_8
X_2213_ _0639_ net397 net385 VPWR VGND sg13g2_nand2_2
XFILLER_39_646 VPWR VGND sg13g2_fill_1
XFILLER_22_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
X_2144_ ppwm_i.u_ppwm.global_counter\[10\] ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0570_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_38_145 VPWR VGND sg13g2_fill_2
X_2075_ _0184_ net422 _0508_ _0509_ VPWR VGND sg13g2_and3_1
XFILLER_34_351 VPWR VGND sg13g2_fill_2
XFILLER_35_885 VPWR VGND sg13g2_decap_8
XFILLER_22_535 VPWR VGND sg13g2_decap_8
X_2977_ net192 VGND VPWR net323 ppwm_i.u_ppwm.u_pwm.cmp_value\[0\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_1928_ sdr_i.mac1.products_ff\[35\] sdr_i.mac1.products_ff\[52\] _0425_ VPWR VGND
+ sg13g2_xor2_1
X_1859_ _0395_ _0394_ _0065_ VPWR VGND sg13g2_xor2_1
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_39_58 VPWR VGND sg13g2_decap_4
XFILLER_18_808 VPWR VGND sg13g2_decap_8
XFILLER_45_605 VPWR VGND sg13g2_decap_4
XFILLER_29_178 VPWR VGND sg13g2_decap_8
XFILLER_41_822 VPWR VGND sg13g2_decap_8
XFILLER_26_885 VPWR VGND sg13g2_decap_8
XFILLER_9_517 VPWR VGND sg13g2_decap_8
XFILLER_41_899 VPWR VGND sg13g2_decap_8
XFILLER_40_376 VPWR VGND sg13g2_decap_8
XFILLER_4_233 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_4
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_4_288 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_944 VPWR VGND sg13g2_decap_8
Xhold80 sdr_i.DP_4.matrix\[0\] VPWR VGND net280 sg13g2_dlygate4sd3_1
Xhold91 sdr_i.mac2.sum_lvl1_ff\[0\] VPWR VGND net291 sg13g2_dlygate4sd3_1
XFILLER_36_627 VPWR VGND sg13g2_decap_8
XFILLER_32_800 VPWR VGND sg13g2_decap_8
X_2900_ net528 VGND VPWR _0091_ sdr_i.DP_1.matrix\[64\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_17_896 VPWR VGND sg13g2_decap_8
XFILLER_32_877 VPWR VGND sg13g2_decap_8
X_3007__134 VPWR VGND net134 sg13g2_tiehi
X_2831_ net287 _0094_ VPWR VGND sg13g2_buf_1
XFILLER_31_387 VPWR VGND sg13g2_fill_2
X_2762_ net417 VPWR _1060_ VGND net480 ppwm_i.u_ppwm.u_mem.memory\[106\] sg13g2_o21ai_1
XFILLER_31_398 VPWR VGND sg13g2_decap_4
X_1713_ net514 net517 _1280_ VPWR VGND sg13g2_nor2_1
X_2693_ VGND VPWR net485 _1137_ _0286_ _1025_ sg13g2_a21oi_1
X_1644_ net818 _1215_ VPWR VGND sg13g2_inv_4
X_1575_ VPWR _1146_ net650 VGND sg13g2_inv_1
Xfanout529 net530 net529 VPWR VGND sg13g2_buf_8
Xfanout518 net788 net518 VPWR VGND sg13g2_buf_8
Xfanout507 net831 net507 VPWR VGND sg13g2_buf_8
X_3176_ net533 VGND VPWR net738 sdr_i.mac1.sum_lvl2_ff\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_27_638 VPWR VGND sg13g2_fill_2
X_2127_ ppwm_i.u_ppwm.pwm_value\[3\] _1256_ _0553_ VPWR VGND sg13g2_nor2_1
XFILLER_42_619 VPWR VGND sg13g2_decap_4
X_2058_ VGND VPWR ppwm_i.u_ppwm.mem_write_done ppwm_i.u_ppwm.u_pwm.counter\[0\] _0498_
+ net707 sg13g2_a21oi_1
XFILLER_23_833 VPWR VGND sg13g2_fill_2
XFILLER_35_671 VPWR VGND sg13g2_fill_2
XFILLER_23_844 VPWR VGND sg13g2_fill_2
XFILLER_41_37 VPWR VGND sg13g2_fill_1
XFILLER_1_203 VPWR VGND sg13g2_fill_2
XFILLER_46_969 VPWR VGND sg13g2_decap_8
XFILLER_17_159 VPWR VGND sg13g2_fill_2
XFILLER_14_833 VPWR VGND sg13g2_fill_1
XFILLER_13_387 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_decap_8
XFILLER_49_741 VPWR VGND sg13g2_decap_8
XFILLER_48_251 VPWR VGND sg13g2_decap_8
X_3030_ net89 VGND VPWR _0221_ ppwm_i.u_ppwm.u_mem.memory\[6\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
XFILLER_37_914 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_43_clk clknet_3_1__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
XFILLER_32_630 VPWR VGND sg13g2_fill_2
X_2814_ net229 _0077_ VPWR VGND sg13g2_buf_1
XFILLER_31_173 VPWR VGND sg13g2_fill_2
XFILLER_31_195 VPWR VGND sg13g2_decap_8
XFILLER_9_870 VPWR VGND sg13g2_decap_8
X_2745_ VGND VPWR net468 _1111_ _0312_ _1051_ sg13g2_a21oi_1
X_2676_ net416 VPWR _1017_ VGND net473 net650 sg13g2_o21ai_1
X_1627_ VPWR _1198_ net647 VGND sg13g2_inv_1
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
X_1558_ VPWR _1129_ net706 VGND sg13g2_inv_1
X_3228_ net526 VGND VPWR net209 sdr_i.mac2.sum_lvl3_ff\[3\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_925 VPWR VGND sg13g2_decap_8
XFILLER_39_262 VPWR VGND sg13g2_decap_8
X_3159_ net530 VGND VPWR _0053_ sdr_i.mac1.products_ff\[120\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_27_424 VPWR VGND sg13g2_decap_8
XFILLER_27_479 VPWR VGND sg13g2_decap_4
XFILLER_42_449 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_34_clk clknet_3_5__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_23_696 VPWR VGND sg13g2_decap_8
XFILLER_7_829 VPWR VGND sg13g2_decap_8
XFILLER_6_306 VPWR VGND sg13g2_fill_1
XFILLER_22_195 VPWR VGND sg13g2_decap_8
XFILLER_10_379 VPWR VGND sg13g2_decap_8
XFILLER_2_545 VPWR VGND sg13g2_decap_8
Xhold380 _0000_ VPWR VGND net760 sg13g2_dlygate4sd3_1
XFILLER_2_578 VPWR VGND sg13g2_decap_8
Xhold391 _0483_ VPWR VGND net771 sg13g2_dlygate4sd3_1
XFILLER_19_958 VPWR VGND sg13g2_decap_8
XFILLER_46_766 VPWR VGND sg13g2_decap_8
XFILLER_34_917 VPWR VGND sg13g2_decap_8
XFILLER_45_265 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_25_clk clknet_3_7__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_26_70 VPWR VGND sg13g2_decap_4
XFILLER_42_972 VPWR VGND sg13g2_decap_8
XFILLER_13_140 VPWR VGND sg13g2_decap_4
XFILLER_41_471 VPWR VGND sg13g2_decap_8
X_2530_ _0896_ _0908_ _0916_ _0927_ _0936_ VPWR VGND sg13g2_and4_1
XFILLER_6_884 VPWR VGND sg13g2_decap_8
X_2461_ _0707_ net370 _0871_ _0873_ _0874_ VPWR VGND sg13g2_nor4_1
X_2392_ _0810_ _0809_ net376 net375 net502 VPWR VGND sg13g2_a22oi_1
XFILLER_3_30 VPWR VGND sg13g2_decap_8
XFILLER_49_560 VPWR VGND sg13g2_decap_8
XFILLER_3_96 VPWR VGND sg13g2_fill_1
X_3013_ net122 VGND VPWR _0204_ ppwm_i.u_ppwm.pwm_value\[9\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_37_744 VPWR VGND sg13g2_fill_2
XFILLER_36_254 VPWR VGND sg13g2_decap_8
XFILLER_37_788 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_3_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_20_600 VPWR VGND sg13g2_fill_2
XFILLER_33_972 VPWR VGND sg13g2_decap_8
X_2728_ net413 VPWR _1043_ VGND net464 ppwm_i.u_ppwm.u_mem.memory\[89\] sg13g2_o21ai_1
X_2659_ VGND VPWR net481 _1154_ _0269_ _1008_ sg13g2_a21oi_1
XFILLER_16_906 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_fill_1
XFILLER_42_202 VPWR VGND sg13g2_decap_8
XFILLER_43_747 VPWR VGND sg13g2_fill_1
XFILLER_42_235 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_24_994 VPWR VGND sg13g2_decap_8
XFILLER_7_604 VPWR VGND sg13g2_fill_1
XFILLER_6_125 VPWR VGND sg13g2_decap_4
XFILLER_3_854 VPWR VGND sg13g2_decap_8
XFILLER_38_508 VPWR VGND sg13g2_fill_2
XFILLER_18_243 VPWR VGND sg13g2_decap_8
XFILLER_19_744 VPWR VGND sg13g2_decap_8
XFILLER_19_788 VPWR VGND sg13g2_fill_2
XFILLER_34_714 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_fill_1
X_3080__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_33_257 VPWR VGND sg13g2_decap_8
XFILLER_15_983 VPWR VGND sg13g2_decap_8
X_1961_ _0012_ _0440_ net723 VPWR VGND sg13g2_xnor2_1
X_1892_ net754 sdr_i.mac2.products_ff\[86\] _0409_ VPWR VGND sg13g2_xor2_1
XFILLER_30_986 VPWR VGND sg13g2_decap_8
X_2513_ VGND VPWR _0916_ _0919_ _0921_ _0920_ sg13g2_a21oi_1
Xclkbuf_leaf_5_clk clknet_3_0__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2444_ VGND VPWR _1229_ net383 _0858_ _0857_ sg13g2_a21oi_1
X_2375_ net422 VPWR _0794_ VGND net828 net371 sg13g2_o21ai_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
X_2989__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_24_202 VPWR VGND sg13g2_fill_1
XFILLER_24_246 VPWR VGND sg13g2_decap_4
XFILLER_24_279 VPWR VGND sg13g2_fill_2
XFILLER_21_975 VPWR VGND sg13g2_decap_8
XFILLER_4_607 VPWR VGND sg13g2_decap_8
XFILLER_4_618 VPWR VGND sg13g2_fill_2
XFILLER_0_857 VPWR VGND sg13g2_decap_8
XFILLER_48_828 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_20 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_28_563 VPWR VGND sg13g2_decap_8
XFILLER_43_533 VPWR VGND sg13g2_decap_8
XFILLER_43_555 VPWR VGND sg13g2_decap_8
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_7_445 VPWR VGND sg13g2_fill_1
XFILLER_7_478 VPWR VGND sg13g2_decap_8
XFILLER_2_150 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_39_806 VPWR VGND sg13g2_decap_8
X_2160_ _0586_ ppwm_i.u_ppwm.pwm_value\[9\] _1259_ VPWR VGND sg13g2_nand2_1
X_2091_ net427 VPWR _0521_ VGND net518 _0520_ sg13g2_o21ai_1
XFILLER_19_541 VPWR VGND sg13g2_fill_2
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_fill_2
XFILLER_19_563 VPWR VGND sg13g2_decap_8
XFILLER_0_75 VPWR VGND sg13g2_decap_8
XFILLER_19_585 VPWR VGND sg13g2_decap_8
XFILLER_34_522 VPWR VGND sg13g2_decap_4
XFILLER_22_706 VPWR VGND sg13g2_fill_2
XFILLER_34_577 VPWR VGND sg13g2_fill_2
X_2993_ net161 VGND VPWR _0184_ ppwm_i.u_ppwm.u_pwm.counter\[6\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
XFILLER_34_599 VPWR VGND sg13g2_decap_8
X_1944_ sdr_i.mac1.sum_lvl1_ff\[17\] sdr_i.mac1.sum_lvl1_ff\[25\] _0433_ VPWR VGND
+ sg13g2_xor2_1
XFILLER_30_783 VPWR VGND sg13g2_decap_8
X_1875_ net2 net1 rst_n_sdr VPWR VGND sg13g2_and2_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_2427_ net424 VPWR _0843_ VGND net814 net372 sg13g2_o21ai_1
X_2358_ VGND VPWR _0755_ _0758_ _0777_ _0754_ sg13g2_a21oi_1
XFILLER_29_338 VPWR VGND sg13g2_fill_1
X_2289_ net424 VPWR _0712_ VGND net507 net371 sg13g2_o21ai_1
XFILLER_38_861 VPWR VGND sg13g2_decap_8
XFILLER_25_533 VPWR VGND sg13g2_decap_8
XFILLER_13_717 VPWR VGND sg13g2_decap_8
XFILLER_25_566 VPWR VGND sg13g2_fill_1
XFILLER_40_536 VPWR VGND sg13g2_decap_8
XFILLER_12_205 VPWR VGND sg13g2_fill_2
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_21_794 VPWR VGND sg13g2_decap_8
XFILLER_5_916 VPWR VGND sg13g2_decap_8
XFILLER_4_437 VPWR VGND sg13g2_fill_1
XFILLER_4_426 VPWR VGND sg13g2_decap_8
XFILLER_29_850 VPWR VGND sg13g2_decap_8
XFILLER_28_393 VPWR VGND sg13g2_decap_8
XFILLER_16_555 VPWR VGND sg13g2_decap_8
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_31_503 VPWR VGND sg13g2_decap_4
XFILLER_12_750 VPWR VGND sg13g2_decap_4
XFILLER_15_1025 VPWR VGND sg13g2_decap_4
XFILLER_8_754 VPWR VGND sg13g2_fill_1
XFILLER_8_776 VPWR VGND sg13g2_fill_2
X_1660_ net508 _1231_ VPWR VGND sg13g2_inv_4
X_1591_ _1162_ net703 VPWR VGND sg13g2_inv_2
Xhold209 _0229_ VPWR VGND net589 sg13g2_dlygate4sd3_1
XFILLER_4_993 VPWR VGND sg13g2_decap_8
X_2212_ _0637_ VPWR _0638_ VGND _0634_ _0636_ sg13g2_o21ai_1
X_3192_ net540 VGND VPWR _0062_ sdr_i.mac2.products_ff\[34\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2143_ _0569_ _1211_ ppwm_i.u_ppwm.global_counter\[18\] VPWR VGND sg13g2_nand2_1
X_2074_ net520 _0504_ net808 _0509_ VPWR VGND sg13g2_nand3_1
XFILLER_19_371 VPWR VGND sg13g2_fill_2
XFILLER_19_393 VPWR VGND sg13g2_decap_8
XFILLER_34_330 VPWR VGND sg13g2_decap_8
XFILLER_35_864 VPWR VGND sg13g2_decap_8
XFILLER_22_514 VPWR VGND sg13g2_decap_4
X_2976_ net423 VGND VPWR net329 ppwm_i.u_ppwm.global_counter\[19\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
X_1927_ net313 sdr_i.mac1.products_ff\[51\] _0017_ VPWR VGND sg13g2_xor2_1
X_1858_ _0395_ net278 net228 VPWR VGND sg13g2_nand2_1
XFILLER_30_39 VPWR VGND sg13g2_decap_8
X_1789_ VPWR VGND _1113_ net460 net442 _1120_ _0338_ net447 sg13g2_a221oi_1
XFILLER_39_37 VPWR VGND sg13g2_decap_8
XFILLER_39_48 VPWR VGND sg13g2_fill_1
XFILLER_41_801 VPWR VGND sg13g2_decap_8
XFILLER_25_352 VPWR VGND sg13g2_decap_8
XFILLER_26_864 VPWR VGND sg13g2_decap_8
XFILLER_13_514 VPWR VGND sg13g2_decap_8
XFILLER_41_878 VPWR VGND sg13g2_decap_8
XFILLER_13_569 VPWR VGND sg13g2_decap_8
XFILLER_5_757 VPWR VGND sg13g2_decap_8
X_2978__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_49_923 VPWR VGND sg13g2_decap_8
XFILLER_0_473 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_48_433 VPWR VGND sg13g2_fill_1
Xhold92 _0013_ VPWR VGND net292 sg13g2_dlygate4sd3_1
Xhold81 sdr_i.DP_2.matrix\[18\] VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold70 _0011_ VPWR VGND net270 sg13g2_dlygate4sd3_1
XFILLER_35_138 VPWR VGND sg13g2_fill_1
XFILLER_17_875 VPWR VGND sg13g2_decap_8
X_2830_ net232 _0093_ VPWR VGND sg13g2_buf_1
XFILLER_31_311 VPWR VGND sg13g2_decap_4
XFILLER_32_856 VPWR VGND sg13g2_decap_8
X_2761_ VGND VPWR net479 _1103_ _0320_ _1059_ sg13g2_a21oi_1
XFILLER_8_551 VPWR VGND sg13g2_decap_8
X_2692_ net426 VPWR _1025_ VGND net485 ppwm_i.u_ppwm.u_mem.memory\[71\] sg13g2_o21ai_1
X_1712_ _1279_ net768 net419 VPWR VGND sg13g2_nand2_1
XFILLER_6_52 VPWR VGND sg13g2_decap_4
X_1643_ _1214_ net821 VPWR VGND sg13g2_inv_2
X_1574_ VPWR _1145_ ppwm_i.u_ppwm.u_mem.memory\[64\] VGND sg13g2_inv_1
Xfanout519 ppwm_i.u_ppwm.pc\[0\] net519 VPWR VGND sg13g2_buf_2
Xfanout508 net509 net508 VPWR VGND sg13g2_buf_8
X_3175_ net533 VGND VPWR net216 sdr_i.mac1.sum_lvl2_ff\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2126_ _0552_ ppwm_i.u_ppwm.global_counter\[18\] _1221_ ppwm_i.u_ppwm.global_counter\[19\]
+ _1220_ VPWR VGND sg13g2_a22oi_1
X_2057_ net455 _0497_ _0178_ VPWR VGND sg13g2_nor2_1
XFILLER_22_322 VPWR VGND sg13g2_decap_4
XFILLER_22_388 VPWR VGND sg13g2_fill_2
X_2959_ net422 VGND VPWR net711 ppwm_i.u_ppwm.global_counter\[2\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
XFILLER_41_49 VPWR VGND sg13g2_decap_4
XFILLER_49_219 VPWR VGND sg13g2_decap_8
XFILLER_46_948 VPWR VGND sg13g2_decap_8
X_3069__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_18_628 VPWR VGND sg13g2_decap_4
XFILLER_45_458 VPWR VGND sg13g2_fill_1
XFILLER_14_812 VPWR VGND sg13g2_fill_2
XFILLER_25_182 VPWR VGND sg13g2_decap_8
XFILLER_9_359 VPWR VGND sg13g2_fill_1
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
X_3076__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_60 VPWR VGND sg13g2_fill_1
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_1_793 VPWR VGND sg13g2_decap_8
XFILLER_49_797 VPWR VGND sg13g2_decap_8
XFILLER_31_141 VPWR VGND sg13g2_decap_4
X_2813_ net276 _0076_ VPWR VGND sg13g2_buf_1
X_2744_ net412 VPWR _1051_ VGND net468 net680 sg13g2_o21ai_1
X_2675_ VGND VPWR net466 _1146_ _0277_ _1016_ sg13g2_a21oi_1
X_1626_ VPWR _1197_ net686 VGND sg13g2_inv_1
X_1557_ VPWR _1128_ net700 VGND sg13g2_inv_1
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
X_3227_ net532 VGND VPWR net208 sdr_i.mac2.sum_lvl3_ff\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_904 VPWR VGND sg13g2_decap_8
X_3158_ net530 VGND VPWR _0052_ sdr_i.mac1.products_ff\[119\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_36_27 VPWR VGND sg13g2_fill_2
X_2109_ _0536_ VPWR _0537_ VGND _0518_ _0535_ sg13g2_o21ai_1
XFILLER_43_929 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_fill_2
X_3089_ net82 VGND VPWR _0280_ ppwm_i.u_ppwm.u_mem.memory\[65\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_3055__40 VPWR VGND net40 sg13g2_tiehi
XFILLER_23_653 VPWR VGND sg13g2_decap_8
XFILLER_10_358 VPWR VGND sg13g2_decap_4
XFILLER_6_318 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_decap_4
Xhold381 sdr_i.mac1.products_ff\[103\] VPWR VGND net761 sg13g2_dlygate4sd3_1
Xhold370 _0320_ VPWR VGND net750 sg13g2_dlygate4sd3_1
Xhold392 _0171_ VPWR VGND net772 sg13g2_dlygate4sd3_1
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_18_436 VPWR VGND sg13g2_decap_4
XFILLER_42_951 VPWR VGND sg13g2_decap_8
XFILLER_14_686 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_10_881 VPWR VGND sg13g2_decap_8
XFILLER_6_863 VPWR VGND sg13g2_decap_8
X_2460_ VGND VPWR _1228_ net383 _0873_ _0872_ sg13g2_a21oi_1
XFILLER_5_395 VPWR VGND sg13g2_fill_1
X_2391_ _0808_ VPWR _0809_ VGND _1261_ net402 sg13g2_o21ai_1
X_3116__88 VPWR VGND net88 sg13g2_tiehi
X_3012_ net124 VGND VPWR net815 ppwm_i.u_ppwm.pwm_value\[8\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_3_1015 VPWR VGND sg13g2_decap_8
XFILLER_37_712 VPWR VGND sg13g2_decap_8
XFILLER_18_981 VPWR VGND sg13g2_decap_8
XFILLER_25_929 VPWR VGND sg13g2_decap_8
XFILLER_17_480 VPWR VGND sg13g2_decap_8
XFILLER_33_951 VPWR VGND sg13g2_decap_8
X_2727_ VGND VPWR net468 _1120_ _0303_ _1042_ sg13g2_a21oi_1
X_2658_ net425 VPWR _1008_ VGND net481 net669 sg13g2_o21ai_1
X_1609_ VPWR _1180_ net636 VGND sg13g2_inv_1
X_2589_ VGND VPWR net499 _1189_ _0234_ _0973_ sg13g2_a21oi_1
XFILLER_27_200 VPWR VGND sg13g2_fill_2
XFILLER_28_789 VPWR VGND sg13g2_decap_4
XFILLER_27_288 VPWR VGND sg13g2_fill_1
XFILLER_24_973 VPWR VGND sg13g2_decap_8
XFILLER_11_601 VPWR VGND sg13g2_fill_2
XFILLER_6_104 VPWR VGND sg13g2_decap_8
XFILLER_11_678 VPWR VGND sg13g2_fill_1
XFILLER_6_159 VPWR VGND sg13g2_decap_8
XFILLER_12_84 VPWR VGND sg13g2_fill_1
XFILLER_3_833 VPWR VGND sg13g2_decap_8
XFILLER_2_387 VPWR VGND sg13g2_fill_2
XFILLER_2_398 VPWR VGND sg13g2_fill_2
XFILLER_18_222 VPWR VGND sg13g2_decap_8
XFILLER_19_767 VPWR VGND sg13g2_decap_8
XFILLER_46_564 VPWR VGND sg13g2_decap_4
XFILLER_19_778 VPWR VGND sg13g2_fill_2
XFILLER_33_236 VPWR VGND sg13g2_decap_8
XFILLER_34_737 VPWR VGND sg13g2_fill_2
XFILLER_15_962 VPWR VGND sg13g2_decap_8
XFILLER_18_1023 VPWR VGND sg13g2_decap_4
X_1960_ net722 sdr_i.mac2.sum_lvl1_ff\[25\] _0441_ VPWR VGND sg13g2_xor2_1
XFILLER_30_965 VPWR VGND sg13g2_decap_8
X_1891_ net265 sdr_i.mac2.products_ff\[85\] _0036_ VPWR VGND sg13g2_xor2_1
X_2512_ net378 VPWR _0920_ VGND _0916_ _0919_ sg13g2_o21ai_1
XFILLER_6_682 VPWR VGND sg13g2_fill_2
X_2443_ net383 _0670_ _0857_ VPWR VGND sg13g2_nor2_1
X_2374_ _0781_ _0789_ net371 _0793_ VPWR VGND _0792_ sg13g2_nand4_1
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_597 VPWR VGND sg13g2_fill_1
XFILLER_20_442 VPWR VGND sg13g2_fill_2
XFILLER_21_954 VPWR VGND sg13g2_decap_8
X_3137__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_0_836 VPWR VGND sg13g2_decap_8
XFILLER_48_807 VPWR VGND sg13g2_decap_8
XFILLER_47_306 VPWR VGND sg13g2_decap_4
XFILLER_43_501 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_21 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_15_214 VPWR VGND sg13g2_decap_8
XFILLER_11_431 VPWR VGND sg13g2_fill_2
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_7_402 VPWR VGND sg13g2_decap_8
XFILLER_11_475 VPWR VGND sg13g2_fill_1
XFILLER_8_958 VPWR VGND sg13g2_decap_8
XFILLER_38_317 VPWR VGND sg13g2_fill_2
XFILLER_47_840 VPWR VGND sg13g2_decap_8
X_2090_ _1232_ _0519_ _0520_ VPWR VGND sg13g2_nor2_1
XFILLER_0_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_372 VPWR VGND sg13g2_fill_1
XFILLER_22_718 VPWR VGND sg13g2_fill_1
X_2992_ net163 VGND VPWR _0183_ ppwm_i.u_ppwm.u_pwm.counter\[5\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_1
X_1943_ net267 sdr_i.mac1.sum_lvl1_ff\[24\] _0025_ VPWR VGND sg13g2_xor2_1
X_1874_ _0405_ _0404_ _0075_ VPWR VGND sg13g2_xor2_1
XFILLER_6_490 VPWR VGND sg13g2_fill_2
X_3017__115 VPWR VGND net115 sg13g2_tiehi
X_2426_ _0835_ _0838_ net372 _0842_ VPWR VGND _0841_ sg13g2_nand4_1
XFILLER_9_1010 VPWR VGND sg13g2_decap_8
X_2357_ _0775_ _0776_ _0199_ VPWR VGND sg13g2_nor2_1
X_2288_ _0701_ _0706_ net371 _0711_ VPWR VGND _0710_ sg13g2_nand4_1
XFILLER_38_840 VPWR VGND sg13g2_decap_8
XFILLER_25_512 VPWR VGND sg13g2_decap_8
XFILLER_25_556 VPWR VGND sg13g2_decap_4
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_20_250 VPWR VGND sg13g2_decap_8
XFILLER_20_283 VPWR VGND sg13g2_decap_8
XFILLER_4_405 VPWR VGND sg13g2_decap_8
XFILLER_20_294 VPWR VGND sg13g2_fill_2
XFILLER_0_611 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_47_114 VPWR VGND sg13g2_fill_2
XFILLER_16_501 VPWR VGND sg13g2_fill_2
XFILLER_28_372 VPWR VGND sg13g2_decap_8
XFILLER_44_865 VPWR VGND sg13g2_decap_8
XFILLER_43_320 VPWR VGND sg13g2_fill_1
XFILLER_15_1004 VPWR VGND sg13g2_decap_8
XFILLER_31_548 VPWR VGND sg13g2_fill_1
XFILLER_12_762 VPWR VGND sg13g2_decap_8
XFILLER_11_294 VPWR VGND sg13g2_fill_1
X_1590_ VPWR _1161_ net570 VGND sg13g2_inv_1
XFILLER_4_972 VPWR VGND sg13g2_decap_8
X_3191_ net546 VGND VPWR _0061_ sdr_i.mac2.products_ff\[18\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2211_ _0637_ _1221_ ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] _1220_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\]
+ VPWR VGND sg13g2_a22oi_1
X_2142_ _0568_ _0552_ _0567_ _1251_ ppwm_i.u_ppwm.pwm_value\[9\] VPWR VGND sg13g2_a22oi_1
X_2073_ _0504_ net520 net808 _0508_ VPWR VGND sg13g2_a21o_1
XFILLER_38_147 VPWR VGND sg13g2_fill_1
XFILLER_35_843 VPWR VGND sg13g2_decap_8
XFILLER_34_353 VPWR VGND sg13g2_fill_1
X_2975_ net436 VGND VPWR _0166_ ppwm_i.u_ppwm.global_counter\[18\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
X_1926_ _0424_ net778 net313 VPWR VGND sg13g2_nand2_1
X_1857_ _0394_ net301 net236 VPWR VGND sg13g2_nand2_1
X_1788_ _0337_ net438 _1106_ net452 _1099_ VPWR VGND sg13g2_a22oi_1
X_2409_ net423 VPWR _0826_ VGND net503 net372 sg13g2_o21ai_1
XFILLER_29_136 VPWR VGND sg13g2_fill_1
XFILLER_17_309 VPWR VGND sg13g2_decap_4
XFILLER_26_843 VPWR VGND sg13g2_decap_8
XFILLER_38_1015 VPWR VGND sg13g2_decap_8
XFILLER_41_857 VPWR VGND sg13g2_decap_8
XFILLER_13_548 VPWR VGND sg13g2_decap_4
XFILLER_25_386 VPWR VGND sg13g2_fill_2
XFILLER_5_736 VPWR VGND sg13g2_decap_8
XFILLER_49_902 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_0_496 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_fill_1
XFILLER_49_979 VPWR VGND sg13g2_decap_8
Xhold60 _0007_ VPWR VGND net260 sg13g2_dlygate4sd3_1
Xhold82 sdr_i.DP_3.matrix\[54\] VPWR VGND net282 sg13g2_dlygate4sd3_1
XFILLER_36_618 VPWR VGND sg13g2_fill_2
Xhold71 sdr_i.DP_3.matrix\[63\] VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold93 sdr_i.DP_3.matrix\[18\] VPWR VGND net293 sg13g2_dlygate4sd3_1
XFILLER_16_342 VPWR VGND sg13g2_decap_8
XFILLER_45_81 VPWR VGND sg13g2_decap_8
XFILLER_31_334 VPWR VGND sg13g2_fill_1
XFILLER_32_835 VPWR VGND sg13g2_decap_8
X_3091__74 VPWR VGND net74 sg13g2_tiehi
X_2760_ net416 VPWR _1059_ VGND net475 net749 sg13g2_o21ai_1
X_2691_ VGND VPWR net473 _1138_ _0285_ _1024_ sg13g2_a21oi_1
X_1711_ net510 net450 net508 _1278_ VPWR VGND sg13g2_nand3_1
X_1642_ VPWR _1213_ net502 VGND sg13g2_inv_1
XFILLER_6_97 VPWR VGND sg13g2_decap_8
X_1573_ VPWR _1144_ net347 VGND sg13g2_inv_1
Xfanout509 net835 net509 VPWR VGND sg13g2_buf_8
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
X_3174_ net522 VGND VPWR net207 sdr_i.mac1.sum_lvl1_ff\[33\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_27_607 VPWR VGND sg13g2_fill_2
X_2125_ _0551_ _1311_ net388 VPWR VGND sg13g2_nand2_2
XFILLER_25_18 VPWR VGND sg13g2_decap_8
X_2056_ _0497_ net715 net769 VPWR VGND sg13g2_xnor2_1
XFILLER_22_301 VPWR VGND sg13g2_decap_4
XFILLER_25_29 VPWR VGND sg13g2_fill_2
XFILLER_10_507 VPWR VGND sg13g2_decap_8
XFILLER_22_367 VPWR VGND sg13g2_decap_8
X_2958_ net421 VGND VPWR net824 ppwm_i.u_ppwm.global_counter\[1\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
X_1909_ sdr_i.mac1.sum_lvl3_ff\[1\] net552 _0415_ VPWR VGND sg13g2_xor2_1
X_2889_ net527 VGND VPWR _0080_ sdr_i.DP_1.matrix\[18\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_46_927 VPWR VGND sg13g2_decap_8
XFILLER_26_684 VPWR VGND sg13g2_fill_1
XFILLER_41_643 VPWR VGND sg13g2_decap_8
XFILLER_41_665 VPWR VGND sg13g2_decap_8
XFILLER_14_879 VPWR VGND sg13g2_decap_8
XFILLER_40_164 VPWR VGND sg13g2_fill_1
XFILLER_15_95 VPWR VGND sg13g2_fill_2
Xoutput4 net4 uio_oe[0] VPWR VGND sg13g2_buf_1
XFILLER_1_772 VPWR VGND sg13g2_decap_8
XFILLER_0_271 VPWR VGND sg13g2_decap_8
XFILLER_49_776 VPWR VGND sg13g2_decap_8
XFILLER_0_293 VPWR VGND sg13g2_decap_8
XFILLER_37_949 VPWR VGND sg13g2_decap_8
XFILLER_45_982 VPWR VGND sg13g2_decap_8
XFILLER_44_470 VPWR VGND sg13g2_fill_2
XFILLER_17_684 VPWR VGND sg13g2_decap_8
XFILLER_31_120 VPWR VGND sg13g2_decap_8
XFILLER_32_654 VPWR VGND sg13g2_decap_4
XFILLER_20_849 VPWR VGND sg13g2_fill_1
X_2812_ VGND VPWR net712 _1095_ _0334_ _1096_ sg13g2_a21oi_1
XFILLER_32_698 VPWR VGND sg13g2_decap_8
X_2743_ VGND VPWR net464 _1112_ _0311_ _1050_ sg13g2_a21oi_1
X_2674_ net412 VPWR _1016_ VGND net466 net660 sg13g2_o21ai_1
X_1625_ VPWR _1196_ net609 VGND sg13g2_inv_1
X_1556_ VPWR _1127_ ppwm_i.u_ppwm.u_mem.memory\[82\] VGND sg13g2_inv_1
X_3119__64 VPWR VGND net64 sg13g2_tiehi
X_3226_ net537 VGND VPWR net765 sdr_i.mac2.sum_lvl3_ff\[1\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3157_ net528 VGND VPWR _0051_ sdr_i.mac1.products_ff\[103\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_27_404 VPWR VGND sg13g2_decap_4
XFILLER_43_908 VPWR VGND sg13g2_decap_8
X_2108_ VGND VPWR _0518_ _0533_ _0536_ _1232_ sg13g2_a21oi_1
X_3088_ net86 VGND VPWR net348 ppwm_i.u_ppwm.u_mem.memory\[64\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_36_982 VPWR VGND sg13g2_decap_8
X_2039_ _0485_ VPWR _0486_ VGND net505 net409 sg13g2_o21ai_1
XFILLER_35_481 VPWR VGND sg13g2_decap_4
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
XFILLER_10_304 VPWR VGND sg13g2_decap_8
XFILLER_22_153 VPWR VGND sg13g2_decap_4
XFILLER_22_175 VPWR VGND sg13g2_fill_2
XFILLER_22_186 VPWR VGND sg13g2_decap_4
Xhold371 ppwm_i.u_ppwm.u_mem.bit_count\[0\] VPWR VGND net751 sg13g2_dlygate4sd3_1
Xhold360 _0039_ VPWR VGND net740 sg13g2_dlygate4sd3_1
Xhold382 _0429_ VPWR VGND net762 sg13g2_dlygate4sd3_1
Xhold393 ppwm_i.u_ppwm.u_mem.memory\[98\] VPWR VGND net773 sg13g2_dlygate4sd3_1
XFILLER_19_916 VPWR VGND sg13g2_decap_8
XFILLER_18_459 VPWR VGND sg13g2_fill_2
XFILLER_45_256 VPWR VGND sg13g2_decap_8
XFILLER_27_982 VPWR VGND sg13g2_decap_8
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_26_492 VPWR VGND sg13g2_fill_1
XFILLER_13_120 VPWR VGND sg13g2_fill_2
XFILLER_14_643 VPWR VGND sg13g2_decap_8
XFILLER_41_495 VPWR VGND sg13g2_decap_4
XFILLER_9_146 VPWR VGND sg13g2_decap_4
XFILLER_6_842 VPWR VGND sg13g2_decap_8
X_2390_ _0808_ ppwm_i.u_ppwm.global_counter\[16\] net403 VPWR VGND sg13g2_nand2_1
XFILLER_1_580 VPWR VGND sg13g2_decap_8
XFILLER_3_87 VPWR VGND sg13g2_fill_1
XFILLER_3_76 VPWR VGND sg13g2_decap_8
X_3011_ net126 VGND VPWR net834 ppwm_i.u_ppwm.pwm_value\[7\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_25_908 VPWR VGND sg13g2_decap_8
XFILLER_18_960 VPWR VGND sg13g2_decap_8
XFILLER_36_278 VPWR VGND sg13g2_fill_1
XFILLER_33_930 VPWR VGND sg13g2_decap_8
XFILLER_20_602 VPWR VGND sg13g2_fill_1
XFILLER_9_691 VPWR VGND sg13g2_decap_8
X_2726_ net414 VPWR _1042_ VGND net469 net354 sg13g2_o21ai_1
X_2657_ VGND VPWR net481 _1155_ _0268_ _1007_ sg13g2_a21oi_1
X_1608_ VPWR _1179_ net576 VGND sg13g2_inv_1
X_2588_ net432 VPWR _0973_ VGND net499 ppwm_i.u_ppwm.u_mem.memory\[19\] sg13g2_o21ai_1
X_1539_ VPWR _1110_ net555 VGND sg13g2_inv_1
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
X_3209_ net544 VGND VPWR net730 sdr_i.mac2.sum_lvl1_ff\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_28_746 VPWR VGND sg13g2_decap_8
XFILLER_28_757 VPWR VGND sg13g2_fill_1
X_3130__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_24_952 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_4
XFILLER_11_657 VPWR VGND sg13g2_decap_8
XFILLER_6_138 VPWR VGND sg13g2_fill_2
XFILLER_3_812 VPWR VGND sg13g2_decap_8
XFILLER_3_889 VPWR VGND sg13g2_decap_8
Xhold190 ppwm_i.u_ppwm.u_mem.memory\[48\] VPWR VGND net570 sg13g2_dlygate4sd3_1
XFILLER_19_713 VPWR VGND sg13g2_decap_8
XFILLER_15_941 VPWR VGND sg13g2_decap_8
XFILLER_18_1002 VPWR VGND sg13g2_decap_8
XFILLER_30_944 VPWR VGND sg13g2_decap_8
X_1890_ _0408_ sdr_i.mac2.products_ff\[85\] net265 VPWR VGND sg13g2_nand2_1
X_2511_ _0917_ VPWR _0919_ VGND _0899_ _0918_ sg13g2_o21ai_1
XFILLER_6_661 VPWR VGND sg13g2_decap_8
X_2442_ VGND VPWR _0847_ _0855_ _0204_ _0856_ sg13g2_a21oi_1
X_2373_ _0792_ _0791_ net376 net375 ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_25_1006 VPWR VGND sg13g2_decap_8
XFILLER_38_2 VPWR VGND sg13g2_fill_1
XFILLER_37_554 VPWR VGND sg13g2_decap_8
XFILLER_25_749 VPWR VGND sg13g2_decap_4
XFILLER_21_933 VPWR VGND sg13g2_decap_8
XFILLER_32_292 VPWR VGND sg13g2_decap_4
X_3025__99 VPWR VGND net99 sg13g2_tiehi
X_2709_ VGND VPWR net477 _1129_ _0294_ _1033_ sg13g2_a21oi_1
X_3040__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_0_815 VPWR VGND sg13g2_decap_8
XFILLER_28_521 VPWR VGND sg13g2_decap_8
XFILLER_16_738 VPWR VGND sg13g2_fill_1
Xtiny_wrapper_22 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_31_719 VPWR VGND sg13g2_decap_8
XFILLER_12_933 VPWR VGND sg13g2_decap_8
XFILLER_23_281 VPWR VGND sg13g2_decap_8
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_7_425 VPWR VGND sg13g2_decap_8
XFILLER_23_84 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_fill_2
XFILLER_48_1017 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_141 VPWR VGND sg13g2_fill_1
X_3098__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_19_543 VPWR VGND sg13g2_fill_1
X_2988__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_34_546 VPWR VGND sg13g2_fill_2
X_2991_ net165 VGND VPWR _0182_ ppwm_i.u_ppwm.u_pwm.counter\[4\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
XFILLER_34_579 VPWR VGND sg13g2_fill_1
X_1942_ _0432_ net746 net267 VPWR VGND sg13g2_nand2_1
XFILLER_30_741 VPWR VGND sg13g2_fill_1
XFILLER_9_97 VPWR VGND sg13g2_fill_2
X_1873_ _0405_ net276 net252 VPWR VGND sg13g2_nand2_1
XFILLER_31_1010 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_4
X_2425_ _0841_ _0840_ _0673_ _0676_ ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] VPWR VGND
+ sg13g2_a22oi_1
X_2356_ net421 VPWR _0776_ VGND net505 net371 sg13g2_o21ai_1
X_2287_ VPWR VGND net376 _0707_ _0709_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _0710_
+ net375 sg13g2_a221oi_1
XFILLER_37_362 VPWR VGND sg13g2_fill_2
XFILLER_38_896 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_fill_1
XFILLER_40_505 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_fill_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_689 VPWR VGND sg13g2_decap_8
XFILLER_18_40 VPWR VGND sg13g2_fill_1
XFILLER_29_885 VPWR VGND sg13g2_decap_8
XFILLER_44_844 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_24_590 VPWR VGND sg13g2_fill_2
X_3079__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_11_251 VPWR VGND sg13g2_fill_1
XFILLER_8_778 VPWR VGND sg13g2_fill_1
XFILLER_7_277 VPWR VGND sg13g2_fill_1
XFILLER_4_951 VPWR VGND sg13g2_decap_8
X_2210_ _0635_ VPWR _0636_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] _1221_ sg13g2_o21ai_1
XFILLER_3_494 VPWR VGND sg13g2_decap_8
X_3190_ net546 VGND VPWR _0060_ sdr_i.mac2.products_ff\[17\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2141_ _0566_ VPWR _0567_ VGND _0563_ _0565_ sg13g2_o21ai_1
X_2072_ VGND VPWR net520 _0504_ _0183_ _0507_ sg13g2_a21oi_1
XFILLER_47_660 VPWR VGND sg13g2_decap_8
XFILLER_19_373 VPWR VGND sg13g2_fill_1
XFILLER_35_822 VPWR VGND sg13g2_decap_8
XFILLER_34_365 VPWR VGND sg13g2_decap_8
XFILLER_34_376 VPWR VGND sg13g2_fill_1
XFILLER_35_899 VPWR VGND sg13g2_decap_8
X_2974_ net436 VGND VPWR net799 ppwm_i.u_ppwm.global_counter\[17\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_22_549 VPWR VGND sg13g2_decap_8
X_1925_ _0014_ _0422_ _0423_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_582 VPWR VGND sg13g2_decap_8
X_1856_ _0393_ _0392_ _0063_ VPWR VGND sg13g2_xor2_1
XFILLER_30_593 VPWR VGND sg13g2_fill_2
X_1787_ VGND VPWR _0336_ net406 net407 sg13g2_or2_1
XFILLER_39_28 VPWR VGND sg13g2_fill_1
X_2408_ VGND VPWR _0817_ _0818_ _0825_ _0824_ sg13g2_a21oi_1
X_2339_ net377 VPWR _0759_ VGND _0755_ _0758_ sg13g2_o21ai_1
XFILLER_44_118 VPWR VGND sg13g2_fill_1
XFILLER_26_811 VPWR VGND sg13g2_decap_8
XFILLER_38_671 VPWR VGND sg13g2_fill_2
XFILLER_26_899 VPWR VGND sg13g2_decap_8
XFILLER_41_836 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_0_453 VPWR VGND sg13g2_fill_2
XFILLER_49_958 VPWR VGND sg13g2_decap_8
Xhold50 sdr_i.DP_3.matrix\[64\] VPWR VGND net250 sg13g2_dlygate4sd3_1
Xhold61 sdr_i.mac1.sum_lvl3_ff\[0\] VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold72 sdr_i.DP_1.matrix\[72\] VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold83 sdr_i.DP_4.matrix\[54\] VPWR VGND net283 sg13g2_dlygate4sd3_1
Xhold94 sdr_i.DP_4.matrix\[18\] VPWR VGND net294 sg13g2_dlygate4sd3_1
XFILLER_29_671 VPWR VGND sg13g2_decap_8
XFILLER_35_129 VPWR VGND sg13g2_decap_8
XFILLER_44_641 VPWR VGND sg13g2_decap_4
XFILLER_45_60 VPWR VGND sg13g2_decap_8
XFILLER_44_685 VPWR VGND sg13g2_decap_8
XFILLER_16_376 VPWR VGND sg13g2_fill_2
XFILLER_32_814 VPWR VGND sg13g2_decap_8
XFILLER_31_324 VPWR VGND sg13g2_fill_1
XFILLER_31_346 VPWR VGND sg13g2_decap_8
X_2690_ net416 VPWR _1024_ VGND net473 net667 sg13g2_o21ai_1
X_1710_ _1277_ net508 net510 net450 VPWR VGND sg13g2_and3_1
X_1641_ _1212_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] VPWR VGND sg13g2_inv_2
X_1572_ VPWR _1143_ net659 VGND sg13g2_inv_1
XFILLER_4_781 VPWR VGND sg13g2_fill_2
XFILLER_6_1003 VPWR VGND sg13g2_decap_8
X_3173_ net522 VGND VPWR net201 sdr_i.mac1.sum_lvl1_ff\[32\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_39_457 VPWR VGND sg13g2_decap_8
X_2124_ net349 VPWR _0550_ VGND net394 _0548_ sg13g2_o21ai_1
X_2055_ net455 _0496_ _0177_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_46_clk clknet_3_1__leaf_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
X_2957_ net421 VGND VPWR net327 ppwm_i.u_ppwm.global_counter\[0\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
XFILLER_31_891 VPWR VGND sg13g2_decap_8
X_2888_ net521 VGND VPWR _0079_ sdr_i.DP_1.matrix\[10\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1908_ net552 sdr_i.mac1.sum_lvl3_ff\[1\] _0414_ VPWR VGND sg13g2_nor2_1
XFILLER_30_390 VPWR VGND sg13g2_decap_8
X_1839_ _0378_ _0376_ _0381_ _0383_ VPWR VGND sg13g2_a21o_1
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_46_906 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_4
XFILLER_45_405 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_37_clk clknet_3_4__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_38_490 VPWR VGND sg13g2_fill_2
XFILLER_14_814 VPWR VGND sg13g2_fill_1
XFILLER_26_663 VPWR VGND sg13g2_decap_8
XFILLER_41_622 VPWR VGND sg13g2_decap_8
XFILLER_25_162 VPWR VGND sg13g2_decap_8
XFILLER_9_306 VPWR VGND sg13g2_decap_8
XFILLER_13_346 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_41_688 VPWR VGND sg13g2_decap_8
XFILLER_22_891 VPWR VGND sg13g2_decap_8
XFILLER_31_51 VPWR VGND sg13g2_fill_1
XFILLER_5_534 VPWR VGND sg13g2_fill_1
XFILLER_31_95 VPWR VGND sg13g2_decap_8
Xoutput5 net5 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_49_755 VPWR VGND sg13g2_decap_8
XFILLER_48_265 VPWR VGND sg13g2_decap_8
XFILLER_36_416 VPWR VGND sg13g2_decap_8
XFILLER_36_427 VPWR VGND sg13g2_fill_2
XFILLER_37_928 VPWR VGND sg13g2_decap_8
X_3083__106 VPWR VGND net106 sg13g2_tiehi
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_decap_8
XFILLER_44_493 VPWR VGND sg13g2_decap_4
XFILLER_16_195 VPWR VGND sg13g2_decap_4
X_2811_ net414 VPWR _1096_ VGND net712 _1095_ sg13g2_o21ai_1
XFILLER_32_677 VPWR VGND sg13g2_decap_8
XFILLER_12_390 VPWR VGND sg13g2_fill_1
X_2742_ net414 VPWR _1050_ VGND net464 net635 sg13g2_o21ai_1
XFILLER_9_884 VPWR VGND sg13g2_decap_8
XFILLER_8_383 VPWR VGND sg13g2_fill_2
X_2673_ VGND VPWR net462 _1147_ _0276_ _1015_ sg13g2_a21oi_1
X_1624_ VPWR _1195_ net666 VGND sg13g2_inv_1
X_1555_ VPWR _1126_ net678 VGND sg13g2_inv_1
X_3225_ net536 VGND VPWR net298 sdr_i.mac2.sum_lvl3_ff\[0\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3156_ net528 VGND VPWR _0050_ sdr_i.mac1.products_ff\[102\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_28_939 VPWR VGND sg13g2_decap_8
XFILLER_39_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_19_clk clknet_3_6__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_3087_ net90 VGND VPWR net651 ppwm_i.u_ppwm.u_mem.memory\[63\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_2107_ _0532_ _0530_ _0535_ VPWR VGND sg13g2_xor2_1
XFILLER_27_438 VPWR VGND sg13g2_decap_4
XFILLER_36_29 VPWR VGND sg13g2_fill_1
XFILLER_42_408 VPWR VGND sg13g2_fill_1
X_2038_ _0485_ _1244_ net410 VPWR VGND sg13g2_nand2_1
XFILLER_36_961 VPWR VGND sg13g2_decap_8
XFILLER_23_622 VPWR VGND sg13g2_decap_8
Xhold350 _0035_ VPWR VGND net730 sg13g2_dlygate4sd3_1
Xhold361 sdr_i.mac1.products_ff\[68\] VPWR VGND net741 sg13g2_dlygate4sd3_1
Xhold372 ppwm_i.u_ppwm.u_pwm.counter\[9\] VPWR VGND net752 sg13g2_dlygate4sd3_1
Xhold383 _0022_ VPWR VGND net763 sg13g2_dlygate4sd3_1
XFILLER_2_559 VPWR VGND sg13g2_fill_2
Xhold394 sdr_i.mac1.sum_lvl3_ff\[2\] VPWR VGND net774 sg13g2_dlygate4sd3_1
XFILLER_18_416 VPWR VGND sg13g2_decap_4
XFILLER_45_213 VPWR VGND sg13g2_fill_2
XFILLER_27_961 VPWR VGND sg13g2_decap_8
XFILLER_26_460 VPWR VGND sg13g2_fill_2
XFILLER_42_986 VPWR VGND sg13g2_decap_8
XFILLER_41_452 VPWR VGND sg13g2_fill_1
XFILLER_42_50 VPWR VGND sg13g2_decap_8
XFILLER_9_169 VPWR VGND sg13g2_decap_8
XFILLER_5_331 VPWR VGND sg13g2_fill_1
XFILLER_6_898 VPWR VGND sg13g2_decap_8
XFILLER_5_386 VPWR VGND sg13g2_decap_4
XFILLER_3_55 VPWR VGND sg13g2_decap_8
XFILLER_49_574 VPWR VGND sg13g2_fill_2
X_3010_ net128 VGND VPWR _0201_ ppwm_i.u_ppwm.pwm_value\[6\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_36_202 VPWR VGND sg13g2_fill_1
XFILLER_36_268 VPWR VGND sg13g2_fill_2
X_3037__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_32_474 VPWR VGND sg13g2_decap_8
XFILLER_33_986 VPWR VGND sg13g2_decap_8
XFILLER_9_670 VPWR VGND sg13g2_fill_2
X_2725_ VGND VPWR net474 _1121_ _0302_ _1041_ sg13g2_a21oi_1
X_2656_ net425 VPWR _1007_ VGND net482 net726 sg13g2_o21ai_1
Xclkbuf_leaf_8_clk clknet_3_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_1607_ VPWR _1178_ net360 VGND sg13g2_inv_1
X_2587_ VGND VPWR net498 _1190_ _0233_ _0972_ sg13g2_a21oi_1
X_1538_ VPWR _1109_ net362 VGND sg13g2_inv_1
X_3208_ net540 VGND VPWR net214 sdr_i.mac2.sum_lvl1_ff\[8\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3139_ net37 VGND VPWR net663 ppwm_i.u_ppwm.u_mem.bit_count\[3\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_27_202 VPWR VGND sg13g2_fill_1
XFILLER_42_216 VPWR VGND sg13g2_decap_8
XFILLER_24_931 VPWR VGND sg13g2_decap_8
XFILLER_42_249 VPWR VGND sg13g2_decap_8
XFILLER_11_603 VPWR VGND sg13g2_fill_1
XFILLER_7_629 VPWR VGND sg13g2_decap_8
Xhold180 _0286_ VPWR VGND net560 sg13g2_dlygate4sd3_1
XFILLER_3_868 VPWR VGND sg13g2_decap_8
Xhold191 _0262_ VPWR VGND net571 sg13g2_dlygate4sd3_1
XFILLER_46_588 VPWR VGND sg13g2_fill_1
XFILLER_15_920 VPWR VGND sg13g2_decap_8
XFILLER_42_783 VPWR VGND sg13g2_decap_8
XFILLER_15_997 VPWR VGND sg13g2_decap_8
XFILLER_30_923 VPWR VGND sg13g2_decap_8
X_2510_ _0918_ _0896_ _0908_ VPWR VGND sg13g2_nand2_1
X_2441_ net423 VPWR _0856_ VGND net793 net372 sg13g2_o21ai_1
X_2372_ _0790_ VPWR _0791_ VGND _1262_ net402 sg13g2_o21ai_1
XFILLER_49_393 VPWR VGND sg13g2_decap_8
XFILLER_37_533 VPWR VGND sg13g2_decap_8
XFILLER_25_728 VPWR VGND sg13g2_decap_8
XFILLER_37_588 VPWR VGND sg13g2_decap_8
XFILLER_40_709 VPWR VGND sg13g2_fill_1
XFILLER_21_912 VPWR VGND sg13g2_decap_8
XFILLER_33_783 VPWR VGND sg13g2_decap_8
XFILLER_32_271 VPWR VGND sg13g2_decap_8
XFILLER_21_989 VPWR VGND sg13g2_decap_8
XFILLER_20_499 VPWR VGND sg13g2_fill_2
X_2708_ net418 VPWR _1033_ VGND net477 net364 sg13g2_o21ai_1
X_2639_ VGND VPWR net481 _1164_ _0259_ _0998_ sg13g2_a21oi_1
XFILLER_47_319 VPWR VGND sg13g2_decap_8
Xtiny_wrapper_23 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_28_577 VPWR VGND sg13g2_decap_8
XFILLER_43_569 VPWR VGND sg13g2_fill_1
XFILLER_12_912 VPWR VGND sg13g2_decap_8
XFILLER_11_411 VPWR VGND sg13g2_fill_1
XFILLER_11_433 VPWR VGND sg13g2_fill_1
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_7_437 VPWR VGND sg13g2_fill_2
XFILLER_11_499 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_fill_2
XFILLER_2_164 VPWR VGND sg13g2_decap_8
XFILLER_38_319 VPWR VGND sg13g2_fill_1
Xfanout490 net500 net490 VPWR VGND sg13g2_buf_2
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_19_577 VPWR VGND sg13g2_decap_4
XFILLER_19_599 VPWR VGND sg13g2_decap_8
XFILLER_0_89 VPWR VGND sg13g2_decap_8
XFILLER_15_750 VPWR VGND sg13g2_decap_8
XFILLER_21_219 VPWR VGND sg13g2_decap_8
X_2990_ net167 VGND VPWR _0181_ ppwm_i.u_ppwm.u_pwm.counter\[3\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_2
XFILLER_42_580 VPWR VGND sg13g2_fill_2
XFILLER_9_43 VPWR VGND sg13g2_decap_4
X_1941_ _0024_ _0430_ net737 VPWR VGND sg13g2_xnor2_1
X_1872_ _0404_ net287 net229 VPWR VGND sg13g2_nand2_1
XFILLER_30_797 VPWR VGND sg13g2_decap_8
X_2424_ _0839_ VPWR _0840_ VGND _1260_ net402 sg13g2_o21ai_1
X_2355_ _0760_ _0770_ _0774_ _0775_ VPWR VGND sg13g2_nor3_1
X_2286_ _0708_ VPWR _0709_ VGND _1258_ net398 sg13g2_o21ai_1
XFILLER_38_875 VPWR VGND sg13g2_decap_8
XFILLER_25_547 VPWR VGND sg13g2_decap_4
X_3143__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_21_775 VPWR VGND sg13g2_fill_1
XFILLER_0_668 VPWR VGND sg13g2_decap_8
X_3111__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_47_116 VPWR VGND sg13g2_fill_1
XFILLER_47_149 VPWR VGND sg13g2_fill_2
XFILLER_47_138 VPWR VGND sg13g2_fill_2
XFILLER_29_864 VPWR VGND sg13g2_decap_8
XFILLER_44_823 VPWR VGND sg13g2_decap_8
XFILLER_43_300 VPWR VGND sg13g2_fill_2
XFILLER_43_311 VPWR VGND sg13g2_decap_8
XFILLER_16_569 VPWR VGND sg13g2_decap_8
XFILLER_31_517 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_8_713 VPWR VGND sg13g2_decap_8
XFILLER_4_930 VPWR VGND sg13g2_decap_8
X_2140_ _0566_ _1253_ net503 _1252_ ppwm_i.u_ppwm.pwm_value\[8\] VPWR VGND sg13g2_a22oi_1
X_2071_ net422 VPWR _0507_ VGND net520 _0504_ sg13g2_o21ai_1
XFILLER_35_801 VPWR VGND sg13g2_decap_8
XFILLER_46_193 VPWR VGND sg13g2_decap_8
XFILLER_46_171 VPWR VGND sg13g2_decap_8
X_3094__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_34_344 VPWR VGND sg13g2_decap_8
XFILLER_35_878 VPWR VGND sg13g2_decap_8
X_2973_ net436 VGND VPWR net781 ppwm_i.u_ppwm.global_counter\[16\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
X_1924_ sdr_i.mac2.sum_lvl1_ff\[1\] sdr_i.mac2.sum_lvl1_ff\[9\] _0423_ VPWR VGND sg13g2_xor2_1
XFILLER_30_561 VPWR VGND sg13g2_decap_8
X_1855_ _0393_ net293 net234 VPWR VGND sg13g2_nand2_1
X_1786_ net407 net406 _0335_ VPWR VGND sg13g2_nor2_2
X_2407_ _0821_ _0823_ _0683_ _0824_ VPWR VGND sg13g2_nand3_1
XFILLER_29_116 VPWR VGND sg13g2_decap_8
X_2338_ _0756_ _0713_ _0757_ _0758_ VPWR VGND sg13g2_a21o_2
X_2269_ _0692_ net396 _0652_ VPWR VGND sg13g2_nand2_2
XFILLER_37_193 VPWR VGND sg13g2_decap_4
XFILLER_41_815 VPWR VGND sg13g2_decap_8
XFILLER_25_366 VPWR VGND sg13g2_fill_2
XFILLER_26_878 VPWR VGND sg13g2_decap_8
XFILLER_25_388 VPWR VGND sg13g2_fill_1
XFILLER_40_369 VPWR VGND sg13g2_decap_8
X_3221__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_4_226 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_fill_2
XFILLER_20_64 VPWR VGND sg13g2_fill_1
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_0_432 VPWR VGND sg13g2_decap_8
XFILLER_49_937 VPWR VGND sg13g2_decap_8
XFILLER_0_487 VPWR VGND sg13g2_decap_4
Xhold40 sdr_i.DP_1.matrix\[19\] VPWR VGND net240 sg13g2_dlygate4sd3_1
Xhold62 _0030_ VPWR VGND net262 sg13g2_dlygate4sd3_1
XFILLER_21_1010 VPWR VGND sg13g2_decap_8
Xhold73 sdr_i.DP_1.matrix\[18\] VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold51 sdr_i.DP_4.matrix\[37\] VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold95 sdr_i.DP_1.matrix\[36\] VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold84 sdr_i.DP_2.matrix\[72\] VPWR VGND net284 sg13g2_dlygate4sd3_1
XFILLER_28_193 VPWR VGND sg13g2_decap_4
XFILLER_44_664 VPWR VGND sg13g2_decap_4
XFILLER_43_152 VPWR VGND sg13g2_decap_8
XFILLER_17_889 VPWR VGND sg13g2_decap_8
XFILLER_12_572 VPWR VGND sg13g2_decap_8
XFILLER_40_892 VPWR VGND sg13g2_decap_8
XFILLER_12_583 VPWR VGND sg13g2_fill_2
X_1640_ _1211_ net809 VPWR VGND sg13g2_inv_2
XFILLER_8_598 VPWR VGND sg13g2_fill_2
X_1571_ VPWR _1142_ net671 VGND sg13g2_inv_1
XFILLER_3_281 VPWR VGND sg13g2_decap_8
XFILLER_39_414 VPWR VGND sg13g2_decap_8
XFILLER_39_403 VPWR VGND sg13g2_fill_2
X_3172_ net197 VGND VPWR net325 ppwm_i.u_ppwm.u_mem.state_q\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_2123_ net394 _0548_ _0549_ VPWR VGND sg13g2_nor2_1
XFILLER_47_491 VPWR VGND sg13g2_fill_2
X_2054_ _0495_ VPWR _0496_ VGND net793 net411 sg13g2_o21ai_1
XFILLER_35_620 VPWR VGND sg13g2_decap_4
XFILLER_35_653 VPWR VGND sg13g2_decap_4
XFILLER_35_686 VPWR VGND sg13g2_decap_4
XFILLER_22_336 VPWR VGND sg13g2_decap_4
X_2956_ net533 VGND VPWR _0147_ sdr_i.DP_4.matrix\[73\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_31_870 VPWR VGND sg13g2_decap_8
X_2887_ net521 VGND VPWR _0078_ sdr_i.DP_1.matrix\[9\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1907_ _0413_ net552 sdr_i.mac1.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
X_1838_ _0378_ _0381_ _0376_ _0382_ VPWR VGND sg13g2_nand3_1
X_1769_ VPWR VGND _1166_ net461 net440 _1173_ _1336_ net444 sg13g2_a221oi_1
XFILLER_39_981 VPWR VGND sg13g2_decap_8
XFILLER_26_631 VPWR VGND sg13g2_decap_4
XFILLER_25_141 VPWR VGND sg13g2_decap_8
XFILLER_14_826 VPWR VGND sg13g2_decap_8
XFILLER_40_122 VPWR VGND sg13g2_decap_8
XFILLER_25_196 VPWR VGND sg13g2_decap_8
XFILLER_22_870 VPWR VGND sg13g2_decap_8
XFILLER_5_546 VPWR VGND sg13g2_decap_4
XFILLER_31_74 VPWR VGND sg13g2_decap_8
Xoutput6 net6 uio_oe[2] VPWR VGND sg13g2_buf_1
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_49_734 VPWR VGND sg13g2_decap_8
XFILLER_0_251 VPWR VGND sg13g2_decap_8
XFILLER_48_244 VPWR VGND sg13g2_decap_8
XFILLER_37_907 VPWR VGND sg13g2_decap_8
XFILLER_45_940 VPWR VGND sg13g2_decap_8
XFILLER_44_472 VPWR VGND sg13g2_fill_1
XFILLER_32_623 VPWR VGND sg13g2_decap_8
X_2810_ _1095_ _1093_ net840 net725 _1234_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_818 VPWR VGND sg13g2_decap_4
XFILLER_9_863 VPWR VGND sg13g2_decap_8
XFILLER_13_892 VPWR VGND sg13g2_decap_8
X_2741_ VGND VPWR net468 _1113_ _0310_ _1049_ sg13g2_a21oi_1
XFILLER_31_188 VPWR VGND sg13g2_decap_8
X_2672_ net413 VPWR _1015_ VGND net462 net590 sg13g2_o21ai_1
X_1623_ VPWR _1194_ net588 VGND sg13g2_inv_1
X_1554_ VPWR _1125_ net681 VGND sg13g2_inv_1
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_3224_ net536 VGND VPWR net204 sdr_i.mac2.sum_lvl2_ff\[9\] clknet_leaf_10_clk sg13g2_dfrbpq_1
.ends

