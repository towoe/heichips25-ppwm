magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755323502
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 27819 37568 27861 37577
rect 27819 37528 27820 37568
rect 27860 37528 27861 37568
rect 27819 37519 27861 37528
rect 27619 37400 27677 37401
rect 27619 37360 27628 37400
rect 27668 37360 27677 37400
rect 27619 37359 27677 37360
rect 30979 37400 31037 37401
rect 30979 37360 30988 37400
rect 31028 37360 31037 37400
rect 30979 37359 31037 37360
rect 31755 37400 31797 37409
rect 31755 37360 31756 37400
rect 31796 37360 31797 37400
rect 31755 37351 31797 37360
rect 32419 37400 32477 37401
rect 32419 37360 32428 37400
rect 32468 37360 32477 37400
rect 32419 37359 32477 37360
rect 27531 37232 27573 37241
rect 27531 37192 27532 37232
rect 27572 37192 27573 37232
rect 27531 37183 27573 37192
rect 30891 37232 30933 37241
rect 30891 37192 30892 37232
rect 30932 37192 30933 37232
rect 30891 37183 30933 37192
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 31651 36896 31709 36897
rect 31651 36856 31660 36896
rect 31700 36856 31709 36896
rect 31651 36855 31709 36856
rect 33291 36812 33333 36821
rect 33291 36772 33292 36812
rect 33332 36772 33333 36812
rect 33291 36763 33333 36772
rect 12547 36728 12605 36729
rect 12547 36688 12556 36728
rect 12596 36688 12605 36728
rect 12547 36687 12605 36688
rect 12651 36728 12693 36737
rect 12651 36688 12652 36728
rect 12692 36688 12693 36728
rect 12651 36679 12693 36688
rect 12843 36728 12885 36737
rect 12843 36688 12844 36728
rect 12884 36688 12885 36728
rect 12843 36679 12885 36688
rect 13699 36728 13757 36729
rect 13699 36688 13708 36728
rect 13748 36688 13757 36728
rect 13699 36687 13757 36688
rect 16099 36728 16157 36729
rect 16099 36688 16108 36728
rect 16148 36688 16157 36728
rect 16099 36687 16157 36688
rect 25603 36728 25661 36729
rect 25603 36688 25612 36728
rect 25652 36688 25661 36728
rect 25603 36687 25661 36688
rect 25707 36728 25749 36737
rect 25707 36688 25708 36728
rect 25748 36688 25749 36728
rect 25707 36679 25749 36688
rect 25899 36728 25941 36737
rect 25899 36688 25900 36728
rect 25940 36688 25941 36728
rect 25899 36679 25941 36688
rect 26091 36728 26133 36737
rect 26091 36688 26092 36728
rect 26132 36688 26133 36728
rect 26091 36679 26133 36688
rect 26187 36728 26229 36737
rect 26187 36688 26188 36728
rect 26228 36688 26229 36728
rect 26187 36679 26229 36688
rect 26283 36728 26325 36737
rect 26283 36688 26284 36728
rect 26324 36688 26325 36728
rect 26283 36679 26325 36688
rect 26379 36728 26421 36737
rect 26379 36688 26380 36728
rect 26420 36688 26421 36728
rect 26379 36679 26421 36688
rect 27715 36728 27773 36729
rect 27715 36688 27724 36728
rect 27764 36688 27773 36728
rect 27715 36687 27773 36688
rect 28003 36728 28061 36729
rect 28003 36688 28012 36728
rect 28052 36688 28061 36728
rect 28003 36687 28061 36688
rect 28683 36728 28725 36737
rect 28683 36688 28684 36728
rect 28724 36688 28725 36728
rect 28683 36679 28725 36688
rect 28963 36728 29021 36729
rect 28963 36688 28972 36728
rect 29012 36688 29021 36728
rect 28963 36687 29021 36688
rect 30499 36728 30557 36729
rect 30499 36688 30508 36728
rect 30548 36688 30557 36728
rect 30499 36687 30557 36688
rect 30787 36728 30845 36729
rect 30787 36688 30796 36728
rect 30836 36688 30845 36728
rect 30787 36687 30845 36688
rect 32323 36728 32381 36729
rect 32323 36688 32332 36728
rect 32372 36688 32381 36728
rect 32323 36687 32381 36688
rect 32611 36728 32669 36729
rect 32611 36688 32620 36728
rect 32660 36688 32669 36728
rect 32611 36687 32669 36688
rect 36067 36728 36125 36729
rect 36067 36688 36076 36728
rect 36116 36688 36125 36728
rect 36067 36687 36125 36688
rect 40003 36728 40061 36729
rect 40003 36688 40012 36728
rect 40052 36688 40061 36728
rect 40003 36687 40061 36688
rect 41059 36728 41117 36729
rect 41059 36688 41068 36728
rect 41108 36688 41117 36728
rect 41059 36687 41117 36688
rect 9963 36560 10005 36569
rect 9963 36520 9964 36560
rect 10004 36520 10005 36560
rect 9963 36511 10005 36520
rect 12843 36560 12885 36569
rect 12843 36520 12844 36560
rect 12884 36520 12885 36560
rect 12843 36511 12885 36520
rect 13899 36560 13941 36569
rect 13899 36520 13900 36560
rect 13940 36520 13941 36560
rect 13899 36511 13941 36520
rect 16299 36560 16341 36569
rect 16299 36520 16300 36560
rect 16340 36520 16341 36560
rect 16299 36511 16341 36520
rect 24939 36560 24981 36569
rect 24939 36520 24940 36560
rect 24980 36520 24981 36560
rect 24939 36511 24981 36520
rect 25899 36560 25941 36569
rect 25899 36520 25900 36560
rect 25940 36520 25941 36560
rect 25899 36511 25941 36520
rect 29643 36560 29685 36569
rect 29643 36520 29644 36560
rect 29684 36520 29685 36560
rect 29643 36511 29685 36520
rect 33483 36560 33525 36569
rect 33483 36520 33484 36560
rect 33524 36520 33525 36560
rect 33483 36511 33525 36520
rect 36459 36560 36501 36569
rect 36459 36520 36460 36560
rect 36500 36520 36501 36560
rect 36459 36511 36501 36520
rect 39147 36560 39189 36569
rect 39147 36520 39148 36560
rect 39188 36520 39189 36560
rect 39147 36511 39189 36520
rect 13027 36476 13085 36477
rect 13027 36436 13036 36476
rect 13076 36436 13085 36476
rect 13027 36435 13085 36436
rect 15427 36476 15485 36477
rect 15427 36436 15436 36476
rect 15476 36436 15485 36476
rect 15427 36435 15485 36436
rect 27043 36476 27101 36477
rect 27043 36436 27052 36476
rect 27092 36436 27101 36476
rect 27043 36435 27101 36436
rect 29067 36476 29109 36485
rect 29067 36436 29068 36476
rect 29108 36436 29109 36476
rect 29067 36427 29109 36436
rect 29827 36476 29885 36477
rect 29827 36436 29836 36476
rect 29876 36436 29885 36476
rect 29827 36435 29885 36436
rect 31459 36476 31517 36477
rect 31459 36436 31468 36476
rect 31508 36436 31517 36476
rect 31459 36435 31517 36436
rect 35395 36476 35453 36477
rect 35395 36436 35404 36476
rect 35444 36436 35453 36476
rect 35395 36435 35453 36436
rect 39331 36476 39389 36477
rect 39331 36436 39340 36476
rect 39380 36436 39389 36476
rect 39331 36435 39389 36436
rect 40387 36476 40445 36477
rect 40387 36436 40396 36476
rect 40436 36436 40445 36476
rect 40387 36435 40445 36436
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 12555 36140 12597 36149
rect 12555 36100 12556 36140
rect 12596 36100 12597 36140
rect 12555 36091 12597 36100
rect 29443 36140 29501 36141
rect 29443 36100 29452 36140
rect 29492 36100 29501 36140
rect 29443 36099 29501 36100
rect 32035 36140 32093 36141
rect 32035 36100 32044 36140
rect 32084 36100 32093 36140
rect 32035 36099 32093 36100
rect 32235 36140 32277 36149
rect 32235 36100 32236 36140
rect 32276 36100 32277 36140
rect 32235 36091 32277 36100
rect 35595 36140 35637 36149
rect 35595 36100 35596 36140
rect 35636 36100 35637 36140
rect 35595 36091 35637 36100
rect 19755 36056 19797 36065
rect 19755 36016 19756 36056
rect 19796 36016 19797 36056
rect 19755 36007 19797 36016
rect 23883 36056 23925 36065
rect 23883 36016 23884 36056
rect 23924 36016 23925 36056
rect 23883 36007 23925 36016
rect 9859 35888 9917 35889
rect 9859 35848 9868 35888
rect 9908 35848 9917 35888
rect 9859 35847 9917 35848
rect 10723 35888 10781 35889
rect 10723 35848 10732 35888
rect 10772 35848 10781 35888
rect 10723 35847 10781 35848
rect 12451 35888 12509 35889
rect 12451 35848 12460 35888
rect 12500 35848 12509 35888
rect 12451 35847 12509 35848
rect 12747 35888 12789 35897
rect 12747 35848 12748 35888
rect 12788 35848 12789 35888
rect 12747 35839 12789 35848
rect 13123 35888 13181 35889
rect 13123 35848 13132 35888
rect 13172 35848 13181 35888
rect 13123 35847 13181 35848
rect 13987 35888 14045 35889
rect 13987 35848 13996 35888
rect 14036 35848 14045 35888
rect 13987 35847 14045 35848
rect 15339 35888 15381 35897
rect 15339 35848 15340 35888
rect 15380 35848 15381 35888
rect 15339 35839 15381 35848
rect 15715 35888 15773 35889
rect 15715 35848 15724 35888
rect 15764 35848 15773 35888
rect 15715 35847 15773 35848
rect 16579 35888 16637 35889
rect 16579 35848 16588 35888
rect 16628 35848 16637 35888
rect 16579 35847 16637 35848
rect 19555 35888 19613 35889
rect 19555 35848 19564 35888
rect 19604 35848 19613 35888
rect 19555 35847 19613 35848
rect 21763 35888 21821 35889
rect 21763 35848 21772 35888
rect 21812 35848 21821 35888
rect 21763 35847 21821 35848
rect 24459 35888 24501 35897
rect 24459 35848 24460 35888
rect 24500 35848 24501 35888
rect 24459 35839 24501 35848
rect 24835 35888 24893 35889
rect 24835 35848 24844 35888
rect 24884 35848 24893 35888
rect 24835 35847 24893 35848
rect 25699 35888 25757 35889
rect 25699 35848 25708 35888
rect 25748 35848 25757 35888
rect 25699 35847 25757 35848
rect 27427 35888 27485 35889
rect 27427 35848 27436 35888
rect 27476 35848 27485 35888
rect 27427 35847 27485 35848
rect 28291 35888 28349 35889
rect 28291 35848 28300 35888
rect 28340 35848 28349 35888
rect 28291 35847 28349 35848
rect 29643 35888 29685 35897
rect 29643 35848 29644 35888
rect 29684 35848 29685 35888
rect 29643 35839 29685 35848
rect 30019 35888 30077 35889
rect 30019 35848 30028 35888
rect 30068 35848 30077 35888
rect 30019 35847 30077 35848
rect 30883 35888 30941 35889
rect 30883 35848 30892 35888
rect 30932 35848 30941 35888
rect 30883 35847 30941 35848
rect 32235 35888 32277 35897
rect 32235 35848 32236 35888
rect 32276 35848 32277 35888
rect 32235 35839 32277 35848
rect 32427 35888 32469 35897
rect 32427 35848 32428 35888
rect 32468 35848 32469 35888
rect 32427 35839 32469 35848
rect 32515 35888 32573 35889
rect 32515 35848 32524 35888
rect 32564 35848 32573 35888
rect 32515 35847 32573 35848
rect 32715 35888 32757 35897
rect 32715 35848 32716 35888
rect 32756 35848 32757 35888
rect 32715 35839 32757 35848
rect 33091 35888 33149 35889
rect 33091 35848 33100 35888
rect 33140 35848 33149 35888
rect 33091 35847 33149 35848
rect 33955 35888 34013 35889
rect 33955 35848 33964 35888
rect 34004 35848 34013 35888
rect 33955 35847 34013 35848
rect 35203 35888 35261 35889
rect 35203 35848 35212 35888
rect 35252 35848 35261 35888
rect 35203 35847 35261 35848
rect 36739 35888 36797 35889
rect 36739 35848 36748 35888
rect 36788 35848 36797 35888
rect 36739 35847 36797 35848
rect 37603 35888 37661 35889
rect 37603 35848 37612 35888
rect 37652 35848 37661 35888
rect 37603 35847 37661 35848
rect 37995 35888 38037 35897
rect 37995 35848 37996 35888
rect 38036 35848 38037 35888
rect 37995 35839 38037 35848
rect 38187 35888 38229 35897
rect 38187 35848 38188 35888
rect 38228 35848 38229 35888
rect 38187 35839 38229 35848
rect 38851 35888 38909 35889
rect 38851 35848 38860 35888
rect 38900 35848 38909 35888
rect 38851 35847 38909 35848
rect 39051 35888 39093 35897
rect 39051 35848 39052 35888
rect 39092 35848 39093 35888
rect 39051 35839 39093 35848
rect 39427 35888 39485 35889
rect 39427 35848 39436 35888
rect 39476 35848 39485 35888
rect 39427 35847 39485 35848
rect 40291 35888 40349 35889
rect 40291 35848 40300 35888
rect 40340 35848 40349 35888
rect 40291 35847 40349 35848
rect 9483 35804 9525 35813
rect 9483 35764 9484 35804
rect 9524 35764 9525 35804
rect 9483 35755 9525 35764
rect 27051 35804 27093 35813
rect 27051 35764 27052 35804
rect 27092 35764 27093 35804
rect 27051 35755 27093 35764
rect 11875 35720 11933 35721
rect 11875 35680 11884 35720
rect 11924 35680 11933 35720
rect 11875 35679 11933 35680
rect 15139 35720 15197 35721
rect 15139 35680 15148 35720
rect 15188 35680 15197 35720
rect 15139 35679 15197 35680
rect 17731 35720 17789 35721
rect 17731 35680 17740 35720
rect 17780 35680 17789 35720
rect 17731 35679 17789 35680
rect 18883 35720 18941 35721
rect 18883 35680 18892 35720
rect 18932 35680 18941 35720
rect 18883 35679 18941 35680
rect 21091 35720 21149 35721
rect 21091 35680 21100 35720
rect 21140 35680 21149 35720
rect 21091 35679 21149 35680
rect 26851 35720 26909 35721
rect 26851 35680 26860 35720
rect 26900 35680 26909 35720
rect 26851 35679 26909 35680
rect 32035 35720 32093 35721
rect 32035 35680 32044 35720
rect 32084 35680 32093 35720
rect 32035 35679 32093 35680
rect 41443 35720 41501 35721
rect 41443 35680 41452 35720
rect 41492 35680 41501 35720
rect 41443 35679 41501 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 8995 35384 9053 35385
rect 8995 35344 9004 35384
rect 9044 35344 9053 35384
rect 8995 35343 9053 35344
rect 12259 35384 12317 35385
rect 12259 35344 12268 35384
rect 12308 35344 12317 35384
rect 12259 35343 12317 35344
rect 27235 35384 27293 35385
rect 27235 35344 27244 35384
rect 27284 35344 27293 35384
rect 27235 35343 27293 35344
rect 37611 35384 37653 35393
rect 37611 35344 37612 35384
rect 37652 35344 37653 35384
rect 37611 35335 37653 35344
rect 38467 35384 38525 35385
rect 38467 35344 38476 35384
rect 38516 35344 38525 35384
rect 38467 35343 38525 35344
rect 5931 35300 5973 35309
rect 5931 35260 5932 35300
rect 5972 35260 5973 35300
rect 5931 35251 5973 35260
rect 13995 35300 14037 35309
rect 13995 35260 13996 35300
rect 14036 35260 14037 35300
rect 13995 35251 14037 35260
rect 18795 35300 18837 35309
rect 18795 35260 18796 35300
rect 18836 35260 18837 35300
rect 18795 35251 18837 35260
rect 23403 35300 23445 35309
rect 23403 35260 23404 35300
rect 23444 35260 23445 35300
rect 23403 35251 23445 35260
rect 26379 35300 26421 35309
rect 26379 35260 26380 35300
rect 26420 35260 26421 35300
rect 26379 35251 26421 35260
rect 29739 35300 29781 35309
rect 29739 35260 29740 35300
rect 29780 35260 29781 35300
rect 29739 35251 29781 35260
rect 31371 35300 31413 35309
rect 31371 35260 31372 35300
rect 31412 35260 31413 35300
rect 31371 35251 31413 35260
rect 33195 35300 33237 35309
rect 33195 35260 33196 35300
rect 33236 35260 33237 35300
rect 33195 35251 33237 35260
rect 34635 35300 34677 35309
rect 34635 35260 34636 35300
rect 34676 35260 34677 35300
rect 34635 35251 34677 35260
rect 36075 35300 36117 35309
rect 36075 35260 36076 35300
rect 36116 35260 36117 35300
rect 36075 35251 36117 35260
rect 39051 35300 39093 35309
rect 39051 35260 39052 35300
rect 39092 35260 39093 35300
rect 39051 35251 39093 35260
rect 39435 35300 39477 35309
rect 39435 35260 39436 35300
rect 39476 35260 39477 35300
rect 39435 35251 39477 35260
rect 5347 35216 5405 35217
rect 5347 35176 5356 35216
rect 5396 35176 5405 35216
rect 5347 35175 5405 35176
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5643 35216 5685 35225
rect 5643 35176 5644 35216
rect 5684 35176 5685 35216
rect 5643 35167 5685 35176
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 6027 35216 6069 35225
rect 6027 35176 6028 35216
rect 6068 35176 6069 35216
rect 6027 35167 6069 35176
rect 6115 35216 6173 35217
rect 6115 35176 6124 35216
rect 6164 35176 6173 35216
rect 6115 35175 6173 35176
rect 6979 35216 7037 35217
rect 6979 35176 6988 35216
rect 7028 35176 7037 35216
rect 6979 35175 7037 35176
rect 8323 35216 8381 35217
rect 8323 35176 8332 35216
rect 8372 35176 8381 35216
rect 8323 35175 8381 35176
rect 8803 35216 8861 35217
rect 8803 35176 8812 35216
rect 8852 35176 8861 35216
rect 8803 35175 8861 35176
rect 8907 35216 8949 35225
rect 8907 35176 8908 35216
rect 8948 35176 8949 35216
rect 8907 35167 8949 35176
rect 9099 35216 9141 35225
rect 9099 35176 9100 35216
rect 9140 35176 9141 35216
rect 9099 35167 9141 35176
rect 9291 35216 9333 35225
rect 9291 35176 9292 35216
rect 9332 35176 9333 35216
rect 9291 35167 9333 35176
rect 9667 35216 9725 35217
rect 9667 35176 9676 35216
rect 9716 35176 9725 35216
rect 9667 35175 9725 35176
rect 10531 35216 10589 35217
rect 10531 35176 10540 35216
rect 10580 35176 10589 35216
rect 10531 35175 10589 35176
rect 12931 35216 12989 35217
rect 12931 35176 12940 35216
rect 12980 35176 12989 35216
rect 12931 35175 12989 35176
rect 13795 35216 13853 35217
rect 13795 35176 13804 35216
rect 13844 35176 13853 35216
rect 13795 35175 13853 35176
rect 14083 35216 14141 35217
rect 14083 35176 14092 35216
rect 14132 35176 14141 35216
rect 14083 35175 14141 35176
rect 14283 35216 14325 35225
rect 14283 35176 14284 35216
rect 14324 35176 14325 35216
rect 14283 35167 14325 35176
rect 14379 35216 14421 35225
rect 14379 35176 14380 35216
rect 14420 35176 14421 35216
rect 14379 35167 14421 35176
rect 14475 35216 14517 35225
rect 14475 35176 14476 35216
rect 14516 35176 14517 35216
rect 14475 35167 14517 35176
rect 14571 35216 14613 35225
rect 14571 35176 14572 35216
rect 14612 35176 14613 35216
rect 14571 35167 14613 35176
rect 15427 35216 15485 35217
rect 15427 35176 15436 35216
rect 15476 35176 15485 35216
rect 15427 35175 15485 35176
rect 16291 35216 16349 35217
rect 16291 35176 16300 35216
rect 16340 35176 16349 35216
rect 16291 35175 16349 35176
rect 16491 35216 16533 35225
rect 16491 35176 16492 35216
rect 16532 35176 16533 35216
rect 16491 35167 16533 35176
rect 16683 35216 16725 35225
rect 16683 35176 16684 35216
rect 16724 35176 16725 35216
rect 16683 35167 16725 35176
rect 16771 35216 16829 35217
rect 16771 35176 16780 35216
rect 16820 35176 16829 35216
rect 16771 35175 16829 35176
rect 16971 35216 17013 35225
rect 16971 35176 16972 35216
rect 17012 35176 17013 35216
rect 16971 35167 17013 35176
rect 17067 35216 17109 35225
rect 17067 35176 17068 35216
rect 17108 35176 17109 35216
rect 17067 35167 17109 35176
rect 17163 35216 17205 35225
rect 17163 35176 17164 35216
rect 17204 35176 17205 35216
rect 17163 35167 17205 35176
rect 17259 35216 17301 35225
rect 17259 35176 17260 35216
rect 17300 35176 17301 35216
rect 17259 35167 17301 35176
rect 18307 35216 18365 35217
rect 18307 35176 18316 35216
rect 18356 35176 18365 35216
rect 18307 35175 18365 35176
rect 19171 35216 19229 35217
rect 19171 35176 19180 35216
rect 19220 35176 19229 35216
rect 19171 35175 19229 35176
rect 20035 35216 20093 35217
rect 20035 35176 20044 35216
rect 20084 35176 20093 35216
rect 20035 35175 20093 35176
rect 22243 35216 22301 35217
rect 22243 35176 22252 35216
rect 22292 35176 22301 35216
rect 22243 35175 22301 35176
rect 23779 35216 23837 35217
rect 23779 35176 23788 35216
rect 23828 35176 23837 35216
rect 23779 35175 23837 35176
rect 24643 35216 24701 35217
rect 24643 35176 24652 35216
rect 24692 35176 24701 35216
rect 24643 35175 24701 35176
rect 25987 35216 26045 35217
rect 25987 35176 25996 35216
rect 26036 35176 26045 35216
rect 25987 35175 26045 35176
rect 26091 35216 26133 35225
rect 26091 35176 26092 35216
rect 26132 35176 26133 35216
rect 26091 35167 26133 35176
rect 26283 35216 26325 35225
rect 26283 35176 26284 35216
rect 26324 35176 26325 35216
rect 26283 35167 26325 35176
rect 26475 35216 26517 35225
rect 26475 35176 26476 35216
rect 26516 35176 26517 35216
rect 26475 35167 26517 35176
rect 26563 35216 26621 35217
rect 26563 35176 26572 35216
rect 26612 35176 26621 35216
rect 26563 35175 26621 35176
rect 26755 35216 26813 35217
rect 26755 35176 26764 35216
rect 26804 35176 26813 35216
rect 26755 35175 26813 35176
rect 26859 35216 26901 35225
rect 26859 35176 26860 35216
rect 26900 35176 26901 35216
rect 26859 35167 26901 35176
rect 27051 35216 27093 35225
rect 27051 35176 27052 35216
rect 27092 35176 27093 35216
rect 27051 35167 27093 35176
rect 27907 35216 27965 35217
rect 27907 35176 27916 35216
rect 27956 35176 27965 35216
rect 27907 35175 27965 35176
rect 29539 35216 29597 35217
rect 29539 35176 29548 35216
rect 29588 35176 29597 35216
rect 29539 35175 29597 35176
rect 29643 35216 29685 35225
rect 29643 35176 29644 35216
rect 29684 35176 29685 35216
rect 29643 35167 29685 35176
rect 29835 35216 29877 35225
rect 29835 35176 29836 35216
rect 29876 35176 29877 35216
rect 29835 35167 29877 35176
rect 30411 35216 30453 35225
rect 30411 35176 30412 35216
rect 30452 35176 30453 35216
rect 30411 35167 30453 35176
rect 30507 35216 30549 35225
rect 30507 35176 30508 35216
rect 30548 35176 30549 35216
rect 30507 35167 30549 35176
rect 30603 35216 30645 35225
rect 30603 35176 30604 35216
rect 30644 35176 30645 35216
rect 30603 35167 30645 35176
rect 30699 35216 30741 35225
rect 30699 35176 30700 35216
rect 30740 35176 30741 35216
rect 30699 35167 30741 35176
rect 30979 35216 31037 35217
rect 30979 35176 30988 35216
rect 31028 35176 31037 35216
rect 30979 35175 31037 35176
rect 31275 35216 31317 35225
rect 31275 35176 31276 35216
rect 31316 35176 31317 35216
rect 31275 35167 31317 35176
rect 31939 35216 31997 35217
rect 31939 35176 31948 35216
rect 31988 35176 31997 35216
rect 31939 35175 31997 35176
rect 32899 35216 32957 35217
rect 32899 35176 32908 35216
rect 32948 35176 32957 35216
rect 32899 35175 32957 35176
rect 33091 35216 33149 35217
rect 33091 35176 33100 35216
rect 33140 35176 33149 35216
rect 33091 35175 33149 35176
rect 34251 35216 34293 35225
rect 34251 35176 34252 35216
rect 34292 35176 34293 35216
rect 34251 35167 34293 35176
rect 34723 35216 34781 35217
rect 34723 35176 34732 35216
rect 34772 35176 34781 35216
rect 34723 35175 34781 35176
rect 35299 35216 35357 35217
rect 35299 35176 35308 35216
rect 35348 35176 35357 35216
rect 35299 35175 35357 35176
rect 35403 35216 35445 35225
rect 35403 35176 35404 35216
rect 35444 35176 35445 35216
rect 35403 35167 35445 35176
rect 35595 35216 35637 35225
rect 35595 35176 35596 35216
rect 35636 35176 35637 35216
rect 35595 35167 35637 35176
rect 35787 35216 35829 35225
rect 35787 35176 35788 35216
rect 35828 35176 35829 35216
rect 35787 35167 35829 35176
rect 35883 35216 35925 35225
rect 35883 35176 35884 35216
rect 35924 35176 35925 35216
rect 35883 35167 35925 35176
rect 35979 35216 36021 35225
rect 35979 35176 35980 35216
rect 36020 35176 36021 35216
rect 35979 35167 36021 35176
rect 36931 35216 36989 35217
rect 36931 35176 36940 35216
rect 36980 35176 36989 35216
rect 36931 35175 36989 35176
rect 38083 35216 38141 35217
rect 38083 35176 38092 35216
rect 38132 35176 38141 35216
rect 38083 35175 38141 35176
rect 38379 35216 38421 35225
rect 38379 35176 38380 35216
rect 38420 35176 38421 35216
rect 38379 35167 38421 35176
rect 38571 35216 38613 35225
rect 38571 35176 38572 35216
rect 38612 35176 38613 35216
rect 38571 35167 38613 35176
rect 38659 35216 38717 35217
rect 38659 35176 38668 35216
rect 38708 35176 38717 35216
rect 38659 35175 38717 35176
rect 39139 35216 39197 35217
rect 39139 35176 39148 35216
rect 39188 35176 39197 35216
rect 39139 35175 39197 35176
rect 39339 35216 39381 35225
rect 39339 35176 39340 35216
rect 39380 35176 39381 35216
rect 39339 35167 39381 35176
rect 39531 35216 39573 35225
rect 39531 35176 39532 35216
rect 39572 35176 39573 35216
rect 39531 35167 39573 35176
rect 39619 35216 39677 35217
rect 39619 35176 39628 35216
rect 39668 35176 39677 35216
rect 39619 35175 39677 35176
rect 40107 35216 40149 35225
rect 40107 35176 40108 35216
rect 40148 35176 40149 35216
rect 40107 35167 40149 35176
rect 40291 35216 40349 35217
rect 40291 35176 40300 35216
rect 40340 35176 40349 35216
rect 40291 35175 40349 35176
rect 40875 35216 40917 35225
rect 40875 35176 40876 35216
rect 40916 35176 40917 35216
rect 40875 35167 40917 35176
rect 41251 35216 41309 35217
rect 41251 35176 41260 35216
rect 41300 35176 41309 35216
rect 41251 35175 41309 35176
rect 42115 35216 42173 35217
rect 42115 35176 42124 35216
rect 42164 35176 42173 35216
rect 42115 35175 42173 35176
rect 44419 35216 44477 35217
rect 44419 35176 44428 35216
rect 44468 35176 44477 35216
rect 44419 35175 44477 35176
rect 11691 35132 11733 35141
rect 11691 35092 11692 35132
rect 11732 35092 11733 35132
rect 11691 35083 11733 35092
rect 25803 35132 25845 35141
rect 25803 35092 25804 35132
rect 25844 35092 25845 35132
rect 25803 35083 25845 35092
rect 28483 35132 28541 35133
rect 28483 35092 28492 35132
rect 28532 35092 28541 35132
rect 28483 35091 28541 35092
rect 37227 35132 37269 35141
rect 37227 35092 37228 35132
rect 37268 35092 37269 35132
rect 37227 35083 37269 35092
rect 4491 35048 4533 35057
rect 4491 35008 4492 35048
rect 4532 35008 4533 35048
rect 4491 34999 4533 35008
rect 7179 35048 7221 35057
rect 7179 35008 7180 35048
rect 7220 35008 7221 35048
rect 7179 34999 7221 35008
rect 12075 35048 12117 35057
rect 12075 35008 12076 35048
rect 12116 35008 12117 35048
rect 12075 34999 12117 35008
rect 17451 35048 17493 35057
rect 17451 35008 17452 35048
rect 17492 35008 17493 35048
rect 17451 34999 17493 35008
rect 22443 35048 22485 35057
rect 22443 35008 22444 35048
rect 22484 35008 22485 35048
rect 22443 34999 22485 35008
rect 27051 35048 27093 35057
rect 27051 35008 27052 35048
rect 27092 35008 27093 35048
rect 27051 34999 27093 35008
rect 28299 35048 28341 35057
rect 28299 35008 28300 35048
rect 28340 35008 28341 35048
rect 28299 34999 28341 35008
rect 28875 35048 28917 35057
rect 28875 35008 28876 35048
rect 28916 35008 28917 35048
rect 28875 34999 28917 35008
rect 29259 35048 29301 35057
rect 29259 35008 29260 35048
rect 29300 35008 29301 35048
rect 29259 34999 29301 35008
rect 30219 35048 30261 35057
rect 30219 35008 30220 35048
rect 30260 35008 30261 35048
rect 30219 34999 30261 35008
rect 35115 35048 35157 35057
rect 35115 35008 35116 35048
rect 35156 35008 35157 35048
rect 35115 34999 35157 35008
rect 40683 35048 40725 35057
rect 40683 35008 40684 35048
rect 40724 35008 40725 35048
rect 40683 34999 40725 35008
rect 5643 34964 5685 34973
rect 5643 34924 5644 34964
rect 5684 34924 5685 34964
rect 5643 34915 5685 34924
rect 6307 34964 6365 34965
rect 6307 34924 6316 34964
rect 6356 34924 6365 34964
rect 6307 34923 6365 34924
rect 7651 34964 7709 34965
rect 7651 34924 7660 34964
rect 7700 34924 7709 34964
rect 7651 34923 7709 34924
rect 12259 34964 12317 34965
rect 12259 34924 12268 34964
rect 12308 34924 12317 34964
rect 12259 34923 12317 34924
rect 13123 34964 13181 34965
rect 13123 34924 13132 34964
rect 13172 34924 13181 34964
rect 13123 34923 13181 34924
rect 14755 34964 14813 34965
rect 14755 34924 14764 34964
rect 14804 34924 14813 34964
rect 14755 34923 14813 34924
rect 15619 34964 15677 34965
rect 15619 34924 15628 34964
rect 15668 34924 15677 34964
rect 15619 34923 15677 34924
rect 16491 34964 16533 34973
rect 16491 34924 16492 34964
rect 16532 34924 16533 34964
rect 16491 34915 16533 34924
rect 18411 34964 18453 34973
rect 18411 34924 18412 34964
rect 18452 34924 18453 34964
rect 18411 34915 18453 34924
rect 21187 34964 21245 34965
rect 21187 34924 21196 34964
rect 21236 34924 21245 34964
rect 21187 34923 21245 34924
rect 21571 34964 21629 34965
rect 21571 34924 21580 34964
rect 21620 34924 21629 34964
rect 21571 34923 21629 34924
rect 31651 34964 31709 34965
rect 31651 34924 31660 34964
rect 31700 34924 31709 34964
rect 31651 34923 31709 34924
rect 32235 34964 32277 34973
rect 32235 34924 32236 34964
rect 32276 34924 32277 34964
rect 32235 34915 32277 34924
rect 33867 34964 33909 34973
rect 33867 34924 33868 34964
rect 33908 34924 33909 34964
rect 33867 34915 33909 34924
rect 35595 34964 35637 34973
rect 35595 34924 35596 34964
rect 35636 34924 35637 34964
rect 35595 34915 35637 34924
rect 36259 34964 36317 34965
rect 36259 34924 36268 34964
rect 36308 34924 36317 34964
rect 36259 34923 36317 34924
rect 40203 34964 40245 34973
rect 40203 34924 40204 34964
rect 40244 34924 40245 34964
rect 40203 34915 40245 34924
rect 43275 34964 43317 34973
rect 43275 34924 43276 34964
rect 43316 34924 43317 34964
rect 43275 34915 43317 34924
rect 43747 34964 43805 34965
rect 43747 34924 43756 34964
rect 43796 34924 43805 34964
rect 43747 34923 43805 34924
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 6019 34628 6077 34629
rect 6019 34588 6028 34628
rect 6068 34588 6077 34628
rect 6019 34587 6077 34588
rect 9387 34628 9429 34637
rect 9387 34588 9388 34628
rect 9428 34588 9429 34628
rect 9387 34579 9429 34588
rect 10923 34628 10965 34637
rect 10923 34588 10924 34628
rect 10964 34588 10965 34628
rect 10923 34579 10965 34588
rect 18307 34628 18365 34629
rect 18307 34588 18316 34628
rect 18356 34588 18365 34628
rect 18307 34587 18365 34588
rect 24075 34628 24117 34637
rect 24075 34588 24076 34628
rect 24116 34588 24117 34628
rect 24075 34579 24117 34588
rect 32523 34628 32565 34637
rect 32523 34588 32524 34628
rect 32564 34588 32565 34628
rect 32523 34579 32565 34588
rect 41443 34628 41501 34629
rect 41443 34588 41452 34628
rect 41492 34588 41501 34628
rect 41443 34587 41501 34588
rect 2571 34544 2613 34553
rect 2571 34504 2572 34544
rect 2612 34504 2613 34544
rect 2571 34495 2613 34504
rect 10443 34544 10485 34553
rect 10443 34504 10444 34544
rect 10484 34504 10485 34544
rect 10443 34495 10485 34504
rect 14179 34544 14237 34545
rect 14179 34504 14188 34544
rect 14228 34504 14237 34544
rect 14179 34503 14237 34504
rect 28579 34544 28637 34545
rect 28579 34504 28588 34544
rect 28628 34504 28637 34544
rect 28579 34503 28637 34504
rect 42603 34544 42645 34553
rect 42603 34504 42604 34544
rect 42644 34504 42645 34544
rect 42603 34495 42645 34504
rect 43659 34544 43701 34553
rect 43659 34504 43660 34544
rect 43700 34504 43701 34544
rect 43659 34495 43701 34504
rect 18123 34460 18165 34469
rect 18123 34420 18124 34460
rect 18164 34420 18165 34460
rect 18123 34411 18165 34420
rect 42123 34460 42165 34469
rect 42123 34420 42124 34460
rect 42164 34420 42165 34460
rect 19363 34418 19421 34419
rect 3627 34376 3669 34385
rect 3627 34336 3628 34376
rect 3668 34336 3669 34376
rect 3627 34327 3669 34336
rect 4003 34376 4061 34377
rect 4003 34336 4012 34376
rect 4052 34336 4061 34376
rect 4003 34335 4061 34336
rect 4867 34376 4925 34377
rect 4867 34336 4876 34376
rect 4916 34336 4925 34376
rect 4867 34335 4925 34336
rect 6219 34376 6261 34385
rect 6219 34336 6220 34376
rect 6260 34336 6261 34376
rect 6219 34327 6261 34336
rect 6595 34376 6653 34377
rect 6595 34336 6604 34376
rect 6644 34336 6653 34376
rect 6595 34335 6653 34336
rect 7459 34376 7517 34377
rect 7459 34336 7468 34376
rect 7508 34336 7517 34376
rect 7459 34335 7517 34336
rect 8803 34376 8861 34377
rect 8803 34336 8812 34376
rect 8852 34336 8861 34376
rect 8803 34335 8861 34336
rect 8907 34376 8949 34385
rect 8907 34336 8908 34376
rect 8948 34336 8949 34376
rect 8907 34327 8949 34336
rect 9091 34376 9149 34377
rect 9091 34336 9100 34376
rect 9140 34336 9149 34376
rect 9091 34335 9149 34336
rect 9195 34376 9237 34385
rect 9195 34336 9196 34376
rect 9236 34336 9237 34376
rect 9195 34327 9237 34336
rect 9387 34376 9429 34385
rect 9387 34336 9388 34376
rect 9428 34336 9429 34376
rect 9387 34327 9429 34336
rect 9571 34376 9629 34377
rect 9571 34336 9580 34376
rect 9620 34336 9629 34376
rect 9571 34335 9629 34336
rect 10251 34376 10293 34385
rect 10251 34336 10252 34376
rect 10292 34336 10293 34376
rect 10251 34327 10293 34336
rect 10819 34376 10877 34377
rect 10819 34336 10828 34376
rect 10868 34336 10877 34376
rect 10819 34335 10877 34336
rect 11203 34376 11261 34377
rect 11203 34336 11212 34376
rect 11252 34336 11261 34376
rect 11203 34335 11261 34336
rect 11499 34376 11541 34385
rect 11499 34336 11500 34376
rect 11540 34336 11541 34376
rect 11499 34327 11541 34336
rect 11595 34376 11637 34385
rect 11595 34336 11596 34376
rect 11636 34336 11637 34376
rect 11595 34327 11637 34336
rect 11691 34376 11733 34385
rect 11691 34336 11692 34376
rect 11732 34336 11733 34376
rect 11691 34327 11733 34336
rect 11883 34376 11925 34385
rect 11883 34336 11884 34376
rect 11924 34336 11925 34376
rect 11883 34327 11925 34336
rect 11979 34376 12021 34385
rect 11979 34336 11980 34376
rect 12020 34336 12021 34376
rect 11979 34327 12021 34336
rect 12075 34376 12117 34385
rect 12075 34336 12076 34376
rect 12116 34336 12117 34376
rect 12075 34327 12117 34336
rect 12171 34376 12213 34385
rect 12171 34336 12172 34376
rect 12212 34336 12213 34376
rect 12171 34327 12213 34336
rect 12363 34376 12405 34385
rect 12363 34336 12364 34376
rect 12404 34336 12405 34376
rect 12363 34327 12405 34336
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 12555 34376 12597 34385
rect 12555 34336 12556 34376
rect 12596 34336 12597 34376
rect 12555 34327 12597 34336
rect 12939 34376 12981 34385
rect 12939 34336 12940 34376
rect 12980 34336 12981 34376
rect 12939 34327 12981 34336
rect 13035 34376 13077 34385
rect 13035 34336 13036 34376
rect 13076 34336 13077 34376
rect 13035 34327 13077 34336
rect 13131 34376 13173 34385
rect 13131 34336 13132 34376
rect 13172 34336 13173 34376
rect 13131 34327 13173 34336
rect 13227 34376 13269 34385
rect 13227 34336 13228 34376
rect 13268 34336 13269 34376
rect 13227 34327 13269 34336
rect 13507 34376 13565 34377
rect 13507 34336 13516 34376
rect 13556 34336 13565 34376
rect 13507 34335 13565 34336
rect 13803 34376 13845 34385
rect 13803 34336 13804 34376
rect 13844 34336 13845 34376
rect 13803 34327 13845 34336
rect 14371 34376 14429 34377
rect 14371 34336 14380 34376
rect 14420 34336 14429 34376
rect 14371 34335 14429 34336
rect 14475 34376 14517 34385
rect 14475 34336 14476 34376
rect 14516 34336 14517 34376
rect 14475 34327 14517 34336
rect 14659 34376 14717 34377
rect 14659 34336 14668 34376
rect 14708 34336 14717 34376
rect 14659 34335 14717 34336
rect 14763 34376 14805 34385
rect 14763 34336 14764 34376
rect 14804 34336 14805 34376
rect 14763 34327 14805 34336
rect 14955 34376 14997 34385
rect 14955 34336 14956 34376
rect 14996 34336 14997 34376
rect 14955 34327 14997 34336
rect 15147 34376 15189 34385
rect 15147 34336 15148 34376
rect 15188 34336 15189 34376
rect 15147 34327 15189 34336
rect 15339 34376 15381 34385
rect 15339 34336 15340 34376
rect 15380 34336 15381 34376
rect 15339 34327 15381 34336
rect 15427 34376 15485 34377
rect 15427 34336 15436 34376
rect 15476 34336 15485 34376
rect 15427 34335 15485 34336
rect 16099 34376 16157 34377
rect 16099 34336 16108 34376
rect 16148 34336 16157 34376
rect 16099 34335 16157 34336
rect 16963 34376 17021 34377
rect 16963 34336 16972 34376
rect 17012 34336 17021 34376
rect 19275 34376 19317 34385
rect 19363 34378 19372 34418
rect 19412 34378 19421 34418
rect 42123 34411 42165 34420
rect 19363 34377 19421 34378
rect 16963 34335 17021 34336
rect 18979 34351 19037 34352
rect 18979 34311 18988 34351
rect 19028 34311 19037 34351
rect 19275 34336 19276 34376
rect 19316 34336 19317 34376
rect 19275 34327 19317 34336
rect 19467 34376 19509 34385
rect 19467 34336 19468 34376
rect 19508 34336 19509 34376
rect 19467 34327 19509 34336
rect 21387 34376 21429 34385
rect 21387 34336 21388 34376
rect 21428 34336 21429 34376
rect 21387 34327 21429 34336
rect 21763 34376 21821 34377
rect 21763 34336 21772 34376
rect 21812 34336 21821 34376
rect 21763 34335 21821 34336
rect 22627 34376 22685 34377
rect 22627 34336 22636 34376
rect 22676 34336 22685 34376
rect 22627 34335 22685 34336
rect 24163 34376 24221 34377
rect 24163 34336 24172 34376
rect 24212 34336 24221 34376
rect 24163 34335 24221 34336
rect 24363 34376 24405 34385
rect 24363 34336 24364 34376
rect 24404 34336 24405 34376
rect 24363 34327 24405 34336
rect 25027 34376 25085 34377
rect 25027 34336 25036 34376
rect 25076 34336 25085 34376
rect 25027 34335 25085 34336
rect 25419 34376 25461 34385
rect 25419 34336 25420 34376
rect 25460 34336 25461 34376
rect 25419 34327 25461 34336
rect 25515 34376 25557 34385
rect 25515 34336 25516 34376
rect 25556 34336 25557 34376
rect 25515 34327 25557 34336
rect 25611 34376 25653 34385
rect 25611 34336 25612 34376
rect 25652 34336 25653 34376
rect 25611 34327 25653 34336
rect 25707 34376 25749 34385
rect 25707 34336 25708 34376
rect 25748 34336 25749 34376
rect 25707 34327 25749 34336
rect 25891 34376 25949 34377
rect 25891 34336 25900 34376
rect 25940 34336 25949 34376
rect 25891 34335 25949 34336
rect 26851 34376 26909 34377
rect 26851 34336 26860 34376
rect 26900 34336 26909 34376
rect 26851 34335 26909 34336
rect 27339 34376 27381 34385
rect 27339 34336 27340 34376
rect 27380 34336 27381 34376
rect 27339 34327 27381 34336
rect 27435 34376 27477 34385
rect 27435 34336 27436 34376
rect 27476 34336 27477 34376
rect 27435 34327 27477 34336
rect 27531 34376 27573 34385
rect 27531 34336 27532 34376
rect 27572 34336 27573 34376
rect 27531 34327 27573 34336
rect 27627 34376 27669 34385
rect 27627 34336 27628 34376
rect 27668 34336 27669 34376
rect 27627 34327 27669 34336
rect 27907 34376 27965 34377
rect 27907 34336 27916 34376
rect 27956 34336 27965 34376
rect 27907 34335 27965 34336
rect 28203 34376 28245 34385
rect 28203 34336 28204 34376
rect 28244 34336 28245 34376
rect 28203 34327 28245 34336
rect 28299 34376 28341 34385
rect 28299 34336 28300 34376
rect 28340 34336 28341 34376
rect 28299 34327 28341 34336
rect 28771 34376 28829 34377
rect 28771 34336 28780 34376
rect 28820 34336 28829 34376
rect 28771 34335 28829 34336
rect 29835 34376 29877 34385
rect 29835 34336 29836 34376
rect 29876 34336 29877 34376
rect 29835 34327 29877 34336
rect 29931 34376 29973 34385
rect 29931 34336 29932 34376
rect 29972 34336 29973 34376
rect 29931 34327 29973 34336
rect 30027 34376 30069 34385
rect 30027 34336 30028 34376
rect 30068 34336 30069 34376
rect 30027 34327 30069 34336
rect 30123 34376 30165 34385
rect 30123 34336 30124 34376
rect 30164 34336 30165 34376
rect 30123 34327 30165 34336
rect 31267 34376 31325 34377
rect 31267 34336 31276 34376
rect 31316 34336 31325 34376
rect 31267 34335 31325 34336
rect 31651 34376 31709 34377
rect 31651 34336 31660 34376
rect 31700 34336 31709 34376
rect 31651 34335 31709 34336
rect 31755 34376 31797 34385
rect 31755 34336 31756 34376
rect 31796 34336 31797 34376
rect 31755 34327 31797 34336
rect 31947 34376 31989 34385
rect 31947 34336 31948 34376
rect 31988 34336 31989 34376
rect 31947 34327 31989 34336
rect 32227 34376 32285 34377
rect 32227 34336 32236 34376
rect 32276 34336 32285 34376
rect 32227 34335 32285 34336
rect 33187 34376 33245 34377
rect 33187 34336 33196 34376
rect 33236 34336 33245 34376
rect 33187 34335 33245 34336
rect 33387 34376 33429 34385
rect 33387 34336 33388 34376
rect 33428 34336 33429 34376
rect 33387 34327 33429 34336
rect 33763 34376 33821 34377
rect 33763 34336 33772 34376
rect 33812 34336 33821 34376
rect 33763 34335 33821 34336
rect 34627 34376 34685 34377
rect 34627 34336 34636 34376
rect 34676 34336 34685 34376
rect 34627 34335 34685 34336
rect 35979 34376 36021 34385
rect 35979 34336 35980 34376
rect 36020 34336 36021 34376
rect 35979 34327 36021 34336
rect 36355 34376 36413 34377
rect 36355 34336 36364 34376
rect 36404 34336 36413 34376
rect 36355 34335 36413 34336
rect 37219 34376 37277 34377
rect 37219 34336 37228 34376
rect 37268 34336 37277 34376
rect 37219 34335 37277 34336
rect 38859 34376 38901 34385
rect 38859 34336 38860 34376
rect 38900 34336 38901 34376
rect 38859 34327 38901 34336
rect 38955 34376 38997 34385
rect 38955 34336 38956 34376
rect 38996 34336 38997 34376
rect 38955 34327 38997 34336
rect 39051 34376 39093 34385
rect 39051 34336 39052 34376
rect 39092 34336 39093 34376
rect 39051 34327 39093 34336
rect 39147 34376 39189 34385
rect 39147 34336 39148 34376
rect 39188 34336 39189 34376
rect 39147 34327 39189 34336
rect 39339 34376 39381 34385
rect 39339 34336 39340 34376
rect 39380 34336 39381 34376
rect 39339 34327 39381 34336
rect 39435 34376 39477 34385
rect 39435 34336 39436 34376
rect 39476 34336 39477 34376
rect 39435 34327 39477 34336
rect 39531 34376 39573 34385
rect 39531 34336 39532 34376
rect 39572 34336 39573 34376
rect 39531 34327 39573 34336
rect 39627 34376 39669 34385
rect 39627 34336 39628 34376
rect 39668 34336 39669 34376
rect 39627 34327 39669 34336
rect 39819 34376 39861 34385
rect 39819 34336 39820 34376
rect 39860 34336 39861 34376
rect 39819 34327 39861 34336
rect 40011 34376 40053 34385
rect 40011 34336 40012 34376
rect 40052 34336 40053 34376
rect 40011 34327 40053 34336
rect 40099 34376 40157 34377
rect 40099 34336 40108 34376
rect 40148 34336 40157 34376
rect 40099 34335 40157 34336
rect 40395 34376 40437 34385
rect 40395 34336 40396 34376
rect 40436 34336 40437 34376
rect 40395 34327 40437 34336
rect 40491 34376 40533 34385
rect 40491 34336 40492 34376
rect 40532 34336 40533 34376
rect 40491 34327 40533 34336
rect 40587 34376 40629 34385
rect 40587 34336 40588 34376
rect 40628 34336 40629 34376
rect 40587 34327 40629 34336
rect 40771 34376 40829 34377
rect 40771 34336 40780 34376
rect 40820 34336 40829 34376
rect 40771 34335 40829 34336
rect 41643 34376 41685 34385
rect 41643 34336 41644 34376
rect 41684 34336 41685 34376
rect 41643 34327 41685 34336
rect 41835 34376 41877 34385
rect 41835 34336 41836 34376
rect 41876 34336 41877 34376
rect 41835 34327 41877 34336
rect 41923 34376 41981 34377
rect 41923 34336 41932 34376
rect 41972 34336 41981 34376
rect 41923 34335 41981 34336
rect 42211 34376 42269 34377
rect 42211 34336 42220 34376
rect 42260 34336 42269 34376
rect 42211 34335 42269 34336
rect 42795 34376 42837 34385
rect 42795 34336 42796 34376
rect 42836 34336 42837 34376
rect 42795 34327 42837 34336
rect 42891 34376 42933 34385
rect 42891 34336 42892 34376
rect 42932 34336 42933 34376
rect 42891 34327 42933 34336
rect 42987 34376 43029 34385
rect 42987 34336 42988 34376
rect 43028 34336 43029 34376
rect 42987 34327 43029 34336
rect 44515 34376 44573 34377
rect 44515 34336 44524 34376
rect 44564 34336 44573 34376
rect 44515 34335 44573 34336
rect 18979 34310 19037 34311
rect 13899 34292 13941 34301
rect 13899 34252 13900 34292
rect 13940 34252 13941 34292
rect 13899 34243 13941 34252
rect 14859 34292 14901 34301
rect 14859 34252 14860 34292
rect 14900 34252 14901 34292
rect 14859 34243 14901 34252
rect 15723 34292 15765 34301
rect 15723 34252 15724 34292
rect 15764 34252 15765 34292
rect 15723 34243 15765 34252
rect 39915 34292 39957 34301
rect 39915 34252 39916 34292
rect 39956 34252 39957 34292
rect 39915 34243 39957 34252
rect 8611 34208 8669 34209
rect 8611 34168 8620 34208
rect 8660 34168 8669 34208
rect 8611 34167 8669 34168
rect 11115 34208 11157 34217
rect 11115 34168 11116 34208
rect 11156 34168 11157 34208
rect 11115 34159 11157 34168
rect 11395 34208 11453 34209
rect 11395 34168 11404 34208
rect 11444 34168 11453 34208
rect 11395 34167 11453 34168
rect 12643 34208 12701 34209
rect 12643 34168 12652 34208
rect 12692 34168 12701 34208
rect 12643 34167 12701 34168
rect 15235 34208 15293 34209
rect 15235 34168 15244 34208
rect 15284 34168 15293 34208
rect 15235 34167 15293 34168
rect 19171 34208 19229 34209
rect 19171 34168 19180 34208
rect 19220 34168 19229 34208
rect 19171 34167 19229 34168
rect 23779 34208 23837 34209
rect 23779 34168 23788 34208
rect 23828 34168 23837 34208
rect 23779 34167 23837 34168
rect 29443 34208 29501 34209
rect 29443 34168 29452 34208
rect 29492 34168 29501 34208
rect 29443 34167 29501 34168
rect 30795 34208 30837 34217
rect 30795 34168 30796 34208
rect 30836 34168 30837 34208
rect 30795 34159 30837 34168
rect 31843 34208 31901 34209
rect 31843 34168 31852 34208
rect 31892 34168 31901 34208
rect 31843 34167 31901 34168
rect 35779 34208 35837 34209
rect 35779 34168 35788 34208
rect 35828 34168 35837 34208
rect 35779 34167 35837 34168
rect 38371 34208 38429 34209
rect 38371 34168 38380 34208
rect 38420 34168 38429 34208
rect 38371 34167 38429 34168
rect 40291 34208 40349 34209
rect 40291 34168 40300 34208
rect 40340 34168 40349 34208
rect 40291 34167 40349 34168
rect 41731 34208 41789 34209
rect 41731 34168 41740 34208
rect 41780 34168 41789 34208
rect 41731 34167 41789 34168
rect 43075 34208 43133 34209
rect 43075 34168 43084 34208
rect 43124 34168 43133 34208
rect 43075 34167 43133 34168
rect 43843 34208 43901 34209
rect 43843 34168 43852 34208
rect 43892 34168 43901 34208
rect 43843 34167 43901 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 4587 33872 4629 33881
rect 4587 33832 4588 33872
rect 4628 33832 4629 33872
rect 4587 33823 4629 33832
rect 6307 33872 6365 33873
rect 6307 33832 6316 33872
rect 6356 33832 6365 33872
rect 6307 33831 6365 33832
rect 9483 33872 9525 33881
rect 9483 33832 9484 33872
rect 9524 33832 9525 33872
rect 9483 33823 9525 33832
rect 11779 33872 11837 33873
rect 11779 33832 11788 33872
rect 11828 33832 11837 33872
rect 11779 33831 11837 33832
rect 18787 33872 18845 33873
rect 18787 33832 18796 33872
rect 18836 33832 18845 33872
rect 18787 33831 18845 33832
rect 21763 33872 21821 33873
rect 21763 33832 21772 33872
rect 21812 33832 21821 33872
rect 21763 33831 21821 33832
rect 33859 33872 33917 33873
rect 33859 33832 33868 33872
rect 33908 33832 33917 33872
rect 33859 33831 33917 33832
rect 36355 33872 36413 33873
rect 36355 33832 36364 33872
rect 36404 33832 36413 33872
rect 36355 33831 36413 33832
rect 45955 33872 46013 33873
rect 45955 33832 45964 33872
rect 46004 33832 46013 33872
rect 45955 33831 46013 33832
rect 4875 33788 4917 33797
rect 4875 33748 4876 33788
rect 4916 33748 4917 33788
rect 4875 33739 4917 33748
rect 6979 33788 7037 33789
rect 6979 33748 6988 33788
rect 7028 33748 7037 33788
rect 6979 33747 7037 33748
rect 9003 33788 9045 33797
rect 9003 33748 9004 33788
rect 9044 33748 9045 33788
rect 9003 33739 9045 33748
rect 17643 33788 17685 33797
rect 17643 33748 17644 33788
rect 17684 33748 17685 33788
rect 17643 33739 17685 33748
rect 25995 33788 26037 33797
rect 25995 33748 25996 33788
rect 26036 33748 26037 33788
rect 25995 33739 26037 33748
rect 30411 33788 30453 33797
rect 30411 33748 30412 33788
rect 30452 33748 30453 33788
rect 30411 33739 30453 33748
rect 32419 33788 32477 33789
rect 32419 33748 32428 33788
rect 32468 33748 32477 33788
rect 32419 33747 32477 33748
rect 42115 33788 42173 33789
rect 42115 33748 42124 33788
rect 42164 33748 42173 33788
rect 42115 33747 42173 33748
rect 1995 33704 2037 33713
rect 1995 33664 1996 33704
rect 2036 33664 2037 33704
rect 1995 33655 2037 33664
rect 2371 33704 2429 33705
rect 2371 33664 2380 33704
rect 2420 33664 2429 33704
rect 2371 33663 2429 33664
rect 3235 33704 3293 33705
rect 3235 33664 3244 33704
rect 3284 33664 3293 33704
rect 3235 33663 3293 33664
rect 4675 33704 4733 33705
rect 4675 33664 4684 33704
rect 4724 33664 4733 33704
rect 4675 33663 4733 33664
rect 4971 33704 5013 33713
rect 4971 33664 4972 33704
rect 5012 33664 5013 33704
rect 4971 33655 5013 33664
rect 5067 33704 5109 33713
rect 5067 33664 5068 33704
rect 5108 33664 5109 33704
rect 5067 33655 5109 33664
rect 5163 33704 5205 33713
rect 5163 33664 5164 33704
rect 5204 33664 5205 33704
rect 5163 33655 5205 33664
rect 5355 33704 5397 33713
rect 5355 33664 5356 33704
rect 5396 33664 5397 33704
rect 5355 33655 5397 33664
rect 6019 33704 6077 33705
rect 6019 33664 6028 33704
rect 6068 33664 6077 33704
rect 6019 33663 6077 33664
rect 6411 33704 6453 33713
rect 6411 33664 6412 33704
rect 6452 33664 6453 33704
rect 6411 33655 6453 33664
rect 6507 33704 6549 33713
rect 6507 33664 6508 33704
rect 6548 33664 6549 33704
rect 6507 33655 6549 33664
rect 6603 33704 6645 33713
rect 6603 33664 6604 33704
rect 6644 33664 6645 33704
rect 6603 33655 6645 33664
rect 7843 33704 7901 33705
rect 7843 33664 7852 33704
rect 7892 33664 7901 33704
rect 7843 33663 7901 33664
rect 8611 33704 8669 33705
rect 8611 33664 8620 33704
rect 8660 33664 8669 33704
rect 8611 33663 8669 33664
rect 8907 33704 8949 33713
rect 8907 33664 8908 33704
rect 8948 33664 8949 33704
rect 8907 33655 8949 33664
rect 10435 33704 10493 33705
rect 10435 33664 10444 33704
rect 10484 33664 10493 33704
rect 10435 33663 10493 33664
rect 10627 33704 10685 33705
rect 10627 33664 10636 33704
rect 10676 33664 10685 33704
rect 10627 33663 10685 33664
rect 11587 33704 11645 33705
rect 11587 33664 11596 33704
rect 11636 33664 11645 33704
rect 11587 33663 11645 33664
rect 12931 33704 12989 33705
rect 12931 33664 12940 33704
rect 12980 33664 12989 33704
rect 12931 33663 12989 33664
rect 13795 33704 13853 33705
rect 13795 33664 13804 33704
rect 13844 33664 13853 33704
rect 13795 33663 13853 33664
rect 14187 33704 14229 33713
rect 14187 33664 14188 33704
rect 14228 33664 14229 33704
rect 14187 33655 14229 33664
rect 14379 33704 14421 33713
rect 14379 33664 14380 33704
rect 14420 33664 14421 33704
rect 14379 33655 14421 33664
rect 15043 33704 15101 33705
rect 15043 33664 15052 33704
rect 15092 33664 15101 33704
rect 15043 33663 15101 33664
rect 15907 33704 15965 33705
rect 15907 33664 15916 33704
rect 15956 33664 15965 33704
rect 15907 33663 15965 33664
rect 17739 33704 17781 33713
rect 17739 33664 17740 33704
rect 17780 33664 17781 33704
rect 17739 33655 17781 33664
rect 18019 33704 18077 33705
rect 18019 33664 18028 33704
rect 18068 33664 18077 33704
rect 18019 33663 18077 33664
rect 18595 33704 18653 33705
rect 18595 33664 18604 33704
rect 18644 33664 18653 33704
rect 18595 33663 18653 33664
rect 18699 33704 18741 33713
rect 18699 33664 18700 33704
rect 18740 33664 18741 33704
rect 18699 33655 18741 33664
rect 18891 33704 18933 33713
rect 18891 33664 18892 33704
rect 18932 33664 18933 33704
rect 18891 33655 18933 33664
rect 19275 33704 19317 33713
rect 19275 33664 19276 33704
rect 19316 33664 19317 33704
rect 19275 33655 19317 33664
rect 20323 33704 20381 33705
rect 20323 33664 20332 33704
rect 20372 33664 20381 33704
rect 20323 33663 20381 33664
rect 20899 33704 20957 33705
rect 20899 33664 20908 33704
rect 20948 33664 20957 33704
rect 20899 33663 20957 33664
rect 21099 33704 21141 33713
rect 21099 33664 21100 33704
rect 21140 33664 21141 33704
rect 21099 33655 21141 33664
rect 21195 33704 21237 33713
rect 21195 33664 21196 33704
rect 21236 33664 21237 33704
rect 21195 33655 21237 33664
rect 21291 33704 21333 33713
rect 21291 33664 21292 33704
rect 21332 33664 21333 33704
rect 21291 33655 21333 33664
rect 21387 33704 21429 33713
rect 21387 33664 21388 33704
rect 21428 33664 21429 33704
rect 21387 33655 21429 33664
rect 21571 33704 21629 33705
rect 21571 33664 21580 33704
rect 21620 33664 21629 33704
rect 21571 33663 21629 33664
rect 21675 33704 21717 33713
rect 21675 33664 21676 33704
rect 21716 33664 21717 33704
rect 21675 33655 21717 33664
rect 21867 33704 21909 33713
rect 21867 33664 21868 33704
rect 21908 33664 21909 33704
rect 21867 33655 21909 33664
rect 24163 33704 24221 33705
rect 24163 33664 24172 33704
rect 24212 33664 24221 33704
rect 24163 33663 24221 33664
rect 25603 33704 25661 33705
rect 25603 33664 25612 33704
rect 25652 33664 25661 33704
rect 25603 33663 25661 33664
rect 25899 33704 25941 33713
rect 25899 33664 25900 33704
rect 25940 33664 25941 33704
rect 25899 33655 25941 33664
rect 26755 33704 26813 33705
rect 26755 33664 26764 33704
rect 26804 33664 26813 33704
rect 26755 33663 26813 33664
rect 27627 33704 27669 33713
rect 27627 33664 27628 33704
rect 27668 33664 27669 33704
rect 27627 33655 27669 33664
rect 29155 33704 29213 33705
rect 29155 33664 29164 33704
rect 29204 33664 29213 33704
rect 29155 33663 29213 33664
rect 30019 33704 30077 33705
rect 30019 33664 30028 33704
rect 30068 33664 30077 33704
rect 30019 33663 30077 33664
rect 30595 33704 30653 33705
rect 30595 33664 30604 33704
rect 30644 33664 30653 33704
rect 30595 33663 30653 33664
rect 32131 33704 32189 33705
rect 32131 33664 32140 33704
rect 32180 33664 32189 33704
rect 32131 33663 32189 33664
rect 33195 33704 33237 33713
rect 33195 33664 33196 33704
rect 33236 33664 33237 33704
rect 33195 33655 33237 33664
rect 33667 33704 33725 33705
rect 33667 33664 33676 33704
rect 33716 33664 33725 33704
rect 33667 33663 33725 33664
rect 33771 33704 33813 33713
rect 33771 33664 33772 33704
rect 33812 33664 33813 33704
rect 33771 33655 33813 33664
rect 33963 33704 34005 33713
rect 33963 33664 33964 33704
rect 34004 33664 34005 33704
rect 33963 33655 34005 33664
rect 34155 33704 34197 33713
rect 34155 33664 34156 33704
rect 34196 33664 34197 33704
rect 34155 33655 34197 33664
rect 34251 33704 34293 33713
rect 34251 33664 34252 33704
rect 34292 33664 34293 33704
rect 34251 33655 34293 33664
rect 34347 33704 34389 33713
rect 34347 33664 34348 33704
rect 34388 33664 34389 33704
rect 34347 33655 34389 33664
rect 34443 33704 34485 33713
rect 34443 33664 34444 33704
rect 34484 33664 34485 33704
rect 34443 33655 34485 33664
rect 36459 33704 36501 33713
rect 36459 33664 36460 33704
rect 36500 33664 36501 33704
rect 36459 33655 36501 33664
rect 36555 33704 36597 33713
rect 36555 33664 36556 33704
rect 36596 33664 36597 33704
rect 36555 33655 36597 33664
rect 36651 33704 36693 33713
rect 36651 33664 36652 33704
rect 36692 33664 36693 33704
rect 36651 33655 36693 33664
rect 36835 33704 36893 33705
rect 36835 33664 36844 33704
rect 36884 33664 36893 33704
rect 36835 33663 36893 33664
rect 37987 33704 38045 33705
rect 37987 33664 37996 33704
rect 38036 33664 38045 33704
rect 37987 33663 38045 33664
rect 38091 33704 38133 33713
rect 38091 33664 38092 33704
rect 38132 33664 38133 33704
rect 38091 33655 38133 33664
rect 38283 33704 38325 33713
rect 38283 33664 38284 33704
rect 38324 33664 38325 33704
rect 38283 33655 38325 33664
rect 38475 33704 38517 33713
rect 38475 33664 38476 33704
rect 38516 33664 38517 33704
rect 38475 33655 38517 33664
rect 38563 33704 38621 33705
rect 38563 33664 38572 33704
rect 38612 33664 38621 33704
rect 38563 33663 38621 33664
rect 38763 33704 38805 33713
rect 38763 33664 38764 33704
rect 38804 33664 38805 33704
rect 38763 33655 38805 33664
rect 38859 33704 38901 33713
rect 38859 33664 38860 33704
rect 38900 33664 38901 33704
rect 38859 33655 38901 33664
rect 38955 33704 38997 33713
rect 38955 33664 38956 33704
rect 38996 33664 38997 33704
rect 38955 33655 38997 33664
rect 39051 33704 39093 33713
rect 39051 33664 39052 33704
rect 39092 33664 39093 33704
rect 39051 33655 39093 33664
rect 39235 33704 39293 33705
rect 39235 33664 39244 33704
rect 39284 33664 39293 33704
rect 39235 33663 39293 33664
rect 40107 33704 40149 33713
rect 40107 33664 40108 33704
rect 40148 33664 40149 33704
rect 40107 33655 40149 33664
rect 40771 33704 40829 33705
rect 40771 33664 40780 33704
rect 40820 33664 40829 33704
rect 40771 33663 40829 33664
rect 41155 33704 41213 33705
rect 41155 33664 41164 33704
rect 41204 33664 41213 33704
rect 41155 33663 41213 33664
rect 42891 33704 42933 33713
rect 42891 33664 42892 33704
rect 42932 33664 42933 33704
rect 42891 33655 42933 33664
rect 43363 33704 43421 33705
rect 43363 33664 43372 33704
rect 43412 33664 43421 33704
rect 43363 33663 43421 33664
rect 43563 33704 43605 33713
rect 43563 33664 43564 33704
rect 43604 33664 43605 33704
rect 43563 33655 43605 33664
rect 43939 33704 43997 33705
rect 43939 33664 43948 33704
rect 43988 33664 43997 33704
rect 43939 33663 43997 33664
rect 44803 33704 44861 33705
rect 44803 33664 44812 33704
rect 44852 33664 44861 33704
rect 44803 33663 44861 33664
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 9667 33620 9725 33621
rect 9667 33580 9676 33620
rect 9716 33580 9725 33620
rect 9667 33579 9725 33580
rect 20043 33620 20085 33629
rect 20043 33580 20044 33620
rect 20084 33580 20085 33620
rect 20043 33571 20085 33580
rect 20811 33620 20853 33629
rect 20811 33580 20812 33620
rect 20852 33580 20853 33620
rect 20811 33571 20853 33580
rect 25027 33620 25085 33621
rect 25027 33580 25036 33620
rect 25076 33580 25085 33620
rect 25027 33579 25085 33580
rect 28011 33620 28053 33629
rect 28011 33580 28012 33620
rect 28052 33580 28053 33620
rect 28011 33571 28053 33580
rect 37515 33620 37557 33629
rect 37515 33580 37516 33620
rect 37556 33580 37557 33620
rect 37515 33571 37557 33580
rect 24363 33536 24405 33545
rect 24363 33496 24364 33536
rect 24404 33496 24405 33536
rect 24363 33487 24405 33496
rect 27435 33536 27477 33545
rect 27435 33496 27436 33536
rect 27476 33496 27477 33536
rect 27435 33487 27477 33496
rect 34635 33536 34677 33545
rect 34635 33496 34636 33536
rect 34676 33496 34677 33536
rect 34635 33487 34677 33496
rect 39907 33536 39965 33537
rect 39907 33496 39916 33536
rect 39956 33496 39965 33536
rect 39907 33495 39965 33496
rect 9283 33452 9341 33453
rect 9283 33412 9292 33452
rect 9332 33412 9341 33452
rect 9283 33411 9341 33412
rect 10915 33452 10973 33453
rect 10915 33412 10924 33452
rect 10964 33412 10973 33452
rect 10915 33411 10973 33412
rect 11779 33452 11837 33453
rect 11779 33412 11788 33452
rect 11828 33412 11837 33452
rect 11779 33411 11837 33412
rect 15235 33452 15293 33453
rect 15235 33412 15244 33452
rect 15284 33412 15293 33452
rect 15235 33411 15293 33412
rect 17347 33452 17405 33453
rect 17347 33412 17356 33452
rect 17396 33412 17405 33452
rect 17347 33411 17405 33412
rect 19467 33452 19509 33461
rect 19467 33412 19468 33452
rect 19508 33412 19509 33452
rect 19467 33403 19509 33412
rect 20427 33452 20469 33461
rect 20427 33412 20428 33452
rect 20468 33412 20469 33452
rect 20427 33403 20469 33412
rect 23491 33452 23549 33453
rect 23491 33412 23500 33452
rect 23540 33412 23549 33452
rect 23491 33411 23549 33412
rect 26275 33452 26333 33453
rect 26275 33412 26284 33452
rect 26324 33412 26333 33452
rect 26275 33411 26333 33412
rect 31267 33452 31325 33453
rect 31267 33412 31276 33452
rect 31316 33412 31325 33452
rect 31267 33411 31325 33412
rect 31459 33452 31517 33453
rect 31459 33412 31468 33452
rect 31508 33412 31517 33452
rect 31459 33411 31517 33412
rect 38283 33452 38325 33461
rect 38283 33412 38284 33452
rect 38324 33412 38325 33452
rect 38283 33403 38325 33412
rect 41827 33452 41885 33453
rect 41827 33412 41836 33452
rect 41876 33412 41885 33452
rect 41827 33411 41885 33412
rect 43275 33452 43317 33461
rect 43275 33412 43276 33452
rect 43316 33412 43317 33452
rect 43275 33403 43317 33412
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 4491 33116 4533 33125
rect 4491 33076 4492 33116
rect 4532 33076 4533 33116
rect 4491 33067 4533 33076
rect 12939 33116 12981 33125
rect 12939 33076 12940 33116
rect 12980 33076 12981 33116
rect 12939 33067 12981 33076
rect 13803 33116 13845 33125
rect 13803 33076 13804 33116
rect 13844 33076 13845 33116
rect 13803 33067 13845 33076
rect 20331 33116 20373 33125
rect 20331 33076 20332 33116
rect 20372 33076 20373 33116
rect 20331 33067 20373 33076
rect 30219 33116 30261 33125
rect 30219 33076 30220 33116
rect 30260 33076 30261 33116
rect 30219 33067 30261 33076
rect 44131 33116 44189 33117
rect 44131 33076 44140 33116
rect 44180 33076 44189 33116
rect 44131 33075 44189 33076
rect 1707 33032 1749 33041
rect 1707 32992 1708 33032
rect 1748 32992 1749 33032
rect 1707 32983 1749 32992
rect 2379 33032 2421 33041
rect 2379 32992 2380 33032
rect 2420 32992 2421 33032
rect 2379 32983 2421 32992
rect 5163 33032 5205 33041
rect 5163 32992 5164 33032
rect 5204 32992 5205 33032
rect 5163 32983 5205 32992
rect 7083 33032 7125 33041
rect 7083 32992 7084 33032
rect 7124 32992 7125 33032
rect 7083 32983 7125 32992
rect 21387 33032 21429 33041
rect 21387 32992 21388 33032
rect 21428 32992 21429 33032
rect 21387 32983 21429 32992
rect 28675 33032 28733 33033
rect 28675 32992 28684 33032
rect 28724 32992 28733 33032
rect 28675 32991 28733 32992
rect 34635 33032 34677 33041
rect 34635 32992 34636 33032
rect 34676 32992 34677 33032
rect 34635 32983 34677 32992
rect 36931 33032 36989 33033
rect 36931 32992 36940 33032
rect 36980 32992 36989 33032
rect 36931 32991 36989 32992
rect 41067 33032 41109 33041
rect 41067 32992 41068 33032
rect 41108 32992 41109 33032
rect 41067 32983 41109 32992
rect 44811 33032 44853 33041
rect 44811 32992 44812 33032
rect 44852 32992 44853 33032
rect 44811 32983 44853 32992
rect 47883 33032 47925 33041
rect 47883 32992 47884 33032
rect 47924 32992 47925 33032
rect 47883 32983 47925 32992
rect 3051 32948 3093 32957
rect 3051 32908 3052 32948
rect 3092 32908 3093 32948
rect 3051 32899 3093 32908
rect 11979 32948 12021 32957
rect 11979 32908 11980 32948
rect 12020 32908 12021 32948
rect 11979 32899 12021 32908
rect 17259 32948 17301 32957
rect 17259 32908 17260 32948
rect 17300 32908 17301 32948
rect 17259 32899 17301 32908
rect 18603 32948 18645 32957
rect 18603 32908 18604 32948
rect 18644 32908 18645 32948
rect 18603 32899 18645 32908
rect 18699 32948 18741 32957
rect 18699 32908 18700 32948
rect 18740 32908 18741 32948
rect 18699 32899 18741 32908
rect 25707 32948 25749 32957
rect 25707 32908 25708 32948
rect 25748 32908 25749 32948
rect 25707 32899 25749 32908
rect 40299 32948 40341 32957
rect 40299 32908 40300 32948
rect 40340 32908 40341 32948
rect 40299 32899 40341 32908
rect 17643 32873 17685 32882
rect 2083 32864 2141 32865
rect 2083 32824 2092 32864
rect 2132 32824 2141 32864
rect 2083 32823 2141 32824
rect 2187 32864 2229 32873
rect 2187 32824 2188 32864
rect 2228 32824 2229 32864
rect 2187 32815 2229 32824
rect 2379 32864 2421 32873
rect 2379 32824 2380 32864
rect 2420 32824 2421 32864
rect 2379 32815 2421 32824
rect 2571 32864 2613 32873
rect 2571 32824 2572 32864
rect 2612 32824 2613 32864
rect 2571 32815 2613 32824
rect 2667 32864 2709 32873
rect 2667 32824 2668 32864
rect 2708 32824 2709 32864
rect 2667 32815 2709 32824
rect 2763 32864 2805 32873
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 2859 32864 2901 32873
rect 2859 32824 2860 32864
rect 2900 32824 2901 32864
rect 2859 32815 2901 32824
rect 3715 32864 3773 32865
rect 3715 32824 3724 32864
rect 3764 32824 3773 32864
rect 3715 32823 3773 32824
rect 4011 32864 4053 32873
rect 4011 32824 4012 32864
rect 4052 32824 4053 32864
rect 4011 32815 4053 32824
rect 4107 32864 4149 32873
rect 4107 32824 4108 32864
rect 4148 32824 4149 32864
rect 4107 32815 4149 32824
rect 4203 32864 4245 32873
rect 4203 32824 4204 32864
rect 4244 32824 4245 32864
rect 4203 32815 4245 32824
rect 4299 32864 4341 32873
rect 4299 32824 4300 32864
rect 4340 32824 4341 32864
rect 4299 32815 4341 32824
rect 4491 32864 4533 32873
rect 4491 32824 4492 32864
rect 4532 32824 4533 32864
rect 4491 32815 4533 32824
rect 4683 32864 4725 32873
rect 4683 32824 4684 32864
rect 4724 32824 4725 32864
rect 4683 32815 4725 32824
rect 4771 32864 4829 32865
rect 4771 32824 4780 32864
rect 4820 32824 4829 32864
rect 4771 32823 4829 32824
rect 6019 32864 6077 32865
rect 6019 32824 6028 32864
rect 6068 32824 6077 32864
rect 6019 32823 6077 32824
rect 6411 32864 6453 32873
rect 6411 32824 6412 32864
rect 6452 32824 6453 32864
rect 6411 32815 6453 32824
rect 6507 32864 6549 32873
rect 6507 32824 6508 32864
rect 6548 32824 6549 32864
rect 6507 32815 6549 32824
rect 6603 32864 6645 32873
rect 6603 32824 6604 32864
rect 6644 32824 6645 32864
rect 6603 32815 6645 32824
rect 6787 32864 6845 32865
rect 6787 32824 6796 32864
rect 6836 32824 6845 32864
rect 6787 32823 6845 32824
rect 6891 32864 6933 32873
rect 6891 32824 6892 32864
rect 6932 32824 6933 32864
rect 6891 32815 6933 32824
rect 7083 32864 7125 32873
rect 7083 32824 7084 32864
rect 7124 32824 7125 32864
rect 7083 32815 7125 32824
rect 7267 32864 7325 32865
rect 7267 32824 7276 32864
rect 7316 32824 7325 32864
rect 7267 32823 7325 32824
rect 8131 32864 8189 32865
rect 8131 32824 8140 32864
rect 8180 32824 8189 32864
rect 8131 32823 8189 32824
rect 8995 32864 9053 32865
rect 8995 32824 9004 32864
rect 9044 32824 9053 32864
rect 8995 32823 9053 32824
rect 9955 32864 10013 32865
rect 9955 32824 9964 32864
rect 10004 32824 10013 32864
rect 9955 32823 10013 32824
rect 10243 32864 10301 32865
rect 10243 32824 10252 32864
rect 10292 32824 10301 32864
rect 10243 32823 10301 32824
rect 10435 32864 10493 32865
rect 10435 32824 10444 32864
rect 10484 32824 10493 32864
rect 10435 32823 10493 32824
rect 11107 32864 11165 32865
rect 11107 32824 11116 32864
rect 11156 32824 11165 32864
rect 11107 32823 11165 32824
rect 13219 32864 13277 32865
rect 13219 32824 13228 32864
rect 13268 32824 13277 32864
rect 13219 32823 13277 32824
rect 13507 32864 13565 32865
rect 13507 32824 13516 32864
rect 13556 32824 13565 32864
rect 13507 32823 13565 32824
rect 13611 32864 13653 32873
rect 13611 32824 13612 32864
rect 13652 32824 13653 32864
rect 13611 32815 13653 32824
rect 13803 32864 13845 32873
rect 13803 32824 13804 32864
rect 13844 32824 13845 32864
rect 13803 32815 13845 32824
rect 14659 32864 14717 32865
rect 14659 32824 14668 32864
rect 14708 32824 14717 32864
rect 14659 32823 14717 32824
rect 14859 32864 14901 32873
rect 14859 32824 14860 32864
rect 14900 32824 14901 32864
rect 14859 32815 14901 32824
rect 15235 32864 15293 32865
rect 15235 32824 15244 32864
rect 15284 32824 15293 32864
rect 15235 32823 15293 32824
rect 16099 32864 16157 32865
rect 16099 32824 16108 32864
rect 16148 32824 16157 32864
rect 17643 32833 17644 32873
rect 17684 32833 17685 32873
rect 17643 32824 17685 32833
rect 18115 32864 18173 32865
rect 18115 32824 18124 32864
rect 18164 32824 18173 32864
rect 16099 32823 16157 32824
rect 18115 32823 18173 32824
rect 19083 32864 19125 32873
rect 19083 32824 19084 32864
rect 19124 32824 19125 32864
rect 19083 32815 19125 32824
rect 19179 32864 19221 32873
rect 19179 32824 19180 32864
rect 19220 32824 19221 32864
rect 19179 32815 19221 32824
rect 19467 32864 19509 32873
rect 19467 32824 19468 32864
rect 19508 32824 19509 32864
rect 19467 32815 19509 32824
rect 19659 32864 19701 32873
rect 19659 32824 19660 32864
rect 19700 32824 19701 32864
rect 19659 32815 19701 32824
rect 19747 32864 19805 32865
rect 19747 32824 19756 32864
rect 19796 32824 19805 32864
rect 19747 32823 19805 32824
rect 20035 32864 20093 32865
rect 20035 32824 20044 32864
rect 20084 32824 20093 32864
rect 20035 32823 20093 32824
rect 23307 32864 23349 32873
rect 23307 32824 23308 32864
rect 23348 32824 23349 32864
rect 23307 32815 23349 32824
rect 23683 32864 23741 32865
rect 23683 32824 23692 32864
rect 23732 32824 23741 32864
rect 23683 32823 23741 32824
rect 24547 32864 24605 32865
rect 24547 32824 24556 32864
rect 24596 32824 24605 32864
rect 24547 32823 24605 32824
rect 25995 32864 26037 32873
rect 25995 32824 25996 32864
rect 26036 32824 26037 32864
rect 25995 32815 26037 32824
rect 26091 32864 26133 32873
rect 26091 32824 26092 32864
rect 26132 32824 26133 32864
rect 26091 32815 26133 32824
rect 26187 32864 26229 32873
rect 26187 32824 26188 32864
rect 26228 32824 26229 32864
rect 26187 32815 26229 32824
rect 26371 32864 26429 32865
rect 26371 32824 26380 32864
rect 26420 32824 26429 32864
rect 26371 32823 26429 32824
rect 27051 32864 27093 32873
rect 27051 32824 27052 32864
rect 27092 32824 27093 32864
rect 27051 32815 27093 32824
rect 27235 32864 27293 32865
rect 27235 32824 27244 32864
rect 27284 32824 27293 32864
rect 27235 32823 27293 32824
rect 27531 32864 27573 32873
rect 27531 32824 27532 32864
rect 27572 32824 27573 32864
rect 27531 32815 27573 32824
rect 27627 32864 27669 32873
rect 27627 32824 27628 32864
rect 27668 32824 27669 32864
rect 27627 32815 27669 32824
rect 27723 32864 27765 32873
rect 27723 32824 27724 32864
rect 27764 32824 27765 32864
rect 27723 32815 27765 32824
rect 28003 32864 28061 32865
rect 28003 32824 28012 32864
rect 28052 32824 28061 32864
rect 28003 32823 28061 32824
rect 29059 32864 29117 32865
rect 29059 32824 29068 32864
rect 29108 32824 29117 32864
rect 29059 32823 29117 32824
rect 29163 32864 29205 32873
rect 29163 32824 29164 32864
rect 29204 32824 29205 32864
rect 29163 32815 29205 32824
rect 29355 32864 29397 32873
rect 29355 32824 29356 32864
rect 29396 32824 29397 32864
rect 29355 32815 29397 32824
rect 30499 32864 30557 32865
rect 30499 32824 30508 32864
rect 30548 32824 30557 32864
rect 30499 32823 30557 32824
rect 30883 32864 30941 32865
rect 30883 32824 30892 32864
rect 30932 32824 30941 32864
rect 30883 32823 30941 32824
rect 31083 32864 31125 32873
rect 31083 32824 31084 32864
rect 31124 32824 31125 32864
rect 31083 32815 31125 32824
rect 31459 32864 31517 32865
rect 31459 32824 31468 32864
rect 31508 32824 31517 32864
rect 31459 32823 31517 32824
rect 32323 32864 32381 32865
rect 32323 32824 32332 32864
rect 32372 32824 32381 32864
rect 32323 32823 32381 32824
rect 34435 32864 34493 32865
rect 34435 32824 34444 32864
rect 34484 32824 34493 32864
rect 34435 32823 34493 32824
rect 36067 32864 36125 32865
rect 36067 32824 36076 32864
rect 36116 32824 36125 32864
rect 36067 32823 36125 32824
rect 37323 32864 37365 32873
rect 37323 32824 37324 32864
rect 37364 32824 37365 32864
rect 37323 32815 37365 32824
rect 37603 32864 37661 32865
rect 37603 32824 37612 32864
rect 37652 32824 37661 32864
rect 37603 32823 37661 32824
rect 37899 32864 37941 32873
rect 37899 32824 37900 32864
rect 37940 32824 37941 32864
rect 37899 32815 37941 32824
rect 38275 32864 38333 32865
rect 38275 32824 38284 32864
rect 38324 32824 38333 32864
rect 38275 32823 38333 32824
rect 39139 32864 39197 32865
rect 39139 32824 39148 32864
rect 39188 32824 39197 32864
rect 39139 32823 39197 32824
rect 40483 32864 40541 32865
rect 40483 32824 40492 32864
rect 40532 32824 40541 32864
rect 40483 32823 40541 32824
rect 40683 32864 40725 32873
rect 40683 32824 40684 32864
rect 40724 32824 40725 32864
rect 40683 32815 40725 32824
rect 41259 32864 41301 32873
rect 41259 32824 41260 32864
rect 41300 32824 41301 32864
rect 41259 32815 41301 32824
rect 41355 32864 41397 32873
rect 41355 32824 41356 32864
rect 41396 32824 41397 32864
rect 41355 32815 41397 32824
rect 41451 32864 41493 32873
rect 41451 32824 41452 32864
rect 41492 32824 41493 32864
rect 41451 32815 41493 32824
rect 41547 32864 41589 32873
rect 41547 32824 41548 32864
rect 41588 32824 41589 32864
rect 41547 32815 41589 32824
rect 41739 32864 41781 32873
rect 41739 32824 41740 32864
rect 41780 32824 41781 32864
rect 41739 32815 41781 32824
rect 42115 32864 42173 32865
rect 42115 32824 42124 32864
rect 42164 32824 42173 32864
rect 42115 32823 42173 32824
rect 42979 32864 43037 32865
rect 42979 32824 42988 32864
rect 43028 32824 43037 32864
rect 42979 32823 43037 32824
rect 45667 32864 45725 32865
rect 45667 32824 45676 32864
rect 45716 32824 45725 32864
rect 45667 32823 45725 32824
rect 47683 32864 47741 32865
rect 47683 32824 47692 32864
rect 47732 32824 47741 32864
rect 47683 32823 47741 32824
rect 5355 32780 5397 32789
rect 5355 32740 5356 32780
rect 5396 32740 5397 32780
rect 5355 32731 5397 32740
rect 8811 32780 8853 32789
rect 8811 32740 8812 32780
rect 8852 32740 8853 32780
rect 8811 32731 8853 32740
rect 17451 32780 17493 32789
rect 17451 32740 17452 32780
rect 17492 32740 17493 32780
rect 17451 32731 17493 32740
rect 20899 32780 20957 32781
rect 20899 32740 20908 32780
rect 20948 32740 20957 32780
rect 20899 32739 20957 32740
rect 37227 32780 37269 32789
rect 37227 32740 37228 32780
rect 37268 32740 37269 32780
rect 37227 32731 37269 32740
rect 40587 32780 40629 32789
rect 40587 32740 40588 32780
rect 40628 32740 40629 32780
rect 40587 32731 40629 32740
rect 6307 32696 6365 32697
rect 6307 32656 6316 32696
rect 6356 32656 6365 32696
rect 6307 32655 6365 32656
rect 7939 32696 7997 32697
rect 7939 32656 7948 32696
rect 7988 32656 7997 32696
rect 7939 32655 7997 32656
rect 13987 32696 14045 32697
rect 13987 32656 13996 32696
rect 14036 32656 14045 32696
rect 13987 32655 14045 32656
rect 19555 32696 19613 32697
rect 19555 32656 19564 32696
rect 19604 32656 19613 32696
rect 19555 32655 19613 32656
rect 25891 32696 25949 32697
rect 25891 32656 25900 32696
rect 25940 32656 25949 32696
rect 25891 32655 25949 32656
rect 27339 32696 27381 32705
rect 27339 32656 27340 32696
rect 27380 32656 27381 32696
rect 27339 32647 27381 32656
rect 27811 32696 27869 32697
rect 27811 32656 27820 32696
rect 27860 32656 27869 32696
rect 27811 32655 27869 32656
rect 29251 32696 29309 32697
rect 29251 32656 29260 32696
rect 29300 32656 29309 32696
rect 29251 32655 29309 32656
rect 30795 32696 30837 32705
rect 30795 32656 30796 32696
rect 30836 32656 30837 32696
rect 30795 32647 30837 32656
rect 33475 32696 33533 32697
rect 33475 32656 33484 32696
rect 33524 32656 33533 32696
rect 33475 32655 33533 32656
rect 33763 32696 33821 32697
rect 33763 32656 33772 32696
rect 33812 32656 33821 32696
rect 33763 32655 33821 32656
rect 36739 32696 36797 32697
rect 36739 32656 36748 32696
rect 36788 32656 36797 32696
rect 36739 32655 36797 32656
rect 44995 32696 45053 32697
rect 44995 32656 45004 32696
rect 45044 32656 45053 32696
rect 44995 32655 45053 32656
rect 47011 32696 47069 32697
rect 47011 32656 47020 32696
rect 47060 32656 47069 32696
rect 47011 32655 47069 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 4099 32360 4157 32361
rect 4099 32320 4108 32360
rect 4148 32320 4157 32360
rect 4099 32319 4157 32320
rect 7363 32360 7421 32361
rect 7363 32320 7372 32360
rect 7412 32320 7421 32360
rect 7363 32319 7421 32320
rect 7563 32360 7605 32369
rect 7563 32320 7564 32360
rect 7604 32320 7605 32360
rect 7563 32311 7605 32320
rect 7939 32360 7997 32361
rect 7939 32320 7948 32360
rect 7988 32320 7997 32360
rect 7939 32319 7997 32320
rect 14275 32360 14333 32361
rect 14275 32320 14284 32360
rect 14324 32320 14333 32360
rect 14275 32319 14333 32320
rect 14955 32360 14997 32369
rect 14955 32320 14956 32360
rect 14996 32320 14997 32360
rect 14955 32311 14997 32320
rect 15139 32360 15197 32361
rect 15139 32320 15148 32360
rect 15188 32320 15197 32360
rect 15139 32319 15197 32320
rect 18211 32360 18269 32361
rect 18211 32320 18220 32360
rect 18260 32320 18269 32360
rect 18211 32319 18269 32320
rect 19075 32360 19133 32361
rect 19075 32320 19084 32360
rect 19124 32320 19133 32360
rect 19075 32319 19133 32320
rect 20131 32360 20189 32361
rect 20131 32320 20140 32360
rect 20180 32320 20189 32360
rect 20131 32319 20189 32320
rect 23587 32360 23645 32361
rect 23587 32320 23596 32360
rect 23636 32320 23645 32360
rect 23587 32319 23645 32320
rect 27235 32360 27293 32361
rect 27235 32320 27244 32360
rect 27284 32320 27293 32360
rect 27235 32319 27293 32320
rect 28491 32360 28533 32369
rect 28491 32320 28492 32360
rect 28532 32320 28533 32360
rect 28491 32311 28533 32320
rect 31843 32360 31901 32361
rect 31843 32320 31852 32360
rect 31892 32320 31901 32360
rect 31843 32319 31901 32320
rect 36067 32360 36125 32361
rect 36067 32320 36076 32360
rect 36116 32320 36125 32360
rect 36067 32319 36125 32320
rect 37707 32360 37749 32369
rect 37707 32320 37708 32360
rect 37748 32320 37749 32360
rect 37707 32311 37749 32320
rect 40203 32360 40245 32369
rect 40203 32320 40204 32360
rect 40244 32320 40245 32360
rect 40203 32311 40245 32320
rect 42115 32360 42173 32361
rect 42115 32320 42124 32360
rect 42164 32320 42173 32360
rect 42115 32319 42173 32320
rect 43947 32360 43989 32369
rect 43947 32320 43948 32360
rect 43988 32320 43989 32360
rect 43947 32311 43989 32320
rect 47107 32360 47165 32361
rect 47107 32320 47116 32360
rect 47156 32320 47165 32360
rect 47107 32319 47165 32320
rect 1323 32276 1365 32285
rect 1323 32236 1324 32276
rect 1364 32236 1365 32276
rect 1323 32227 1365 32236
rect 4971 32276 5013 32285
rect 4971 32236 4972 32276
rect 5012 32236 5013 32276
rect 4971 32227 5013 32236
rect 8427 32276 8469 32285
rect 8427 32236 8428 32276
rect 8468 32236 8469 32276
rect 8427 32227 8469 32236
rect 22539 32276 22581 32285
rect 22539 32236 22540 32276
rect 22580 32236 22581 32276
rect 22539 32227 22581 32236
rect 33675 32276 33717 32285
rect 33675 32236 33676 32276
rect 33716 32236 33717 32276
rect 33675 32227 33717 32236
rect 44715 32276 44757 32285
rect 44715 32236 44716 32276
rect 44756 32236 44757 32276
rect 44715 32227 44757 32236
rect 4771 32217 4829 32218
rect 1699 32192 1757 32193
rect 1699 32152 1708 32192
rect 1748 32152 1757 32192
rect 1699 32151 1757 32152
rect 2563 32192 2621 32193
rect 2563 32152 2572 32192
rect 2612 32152 2621 32192
rect 4771 32177 4780 32217
rect 4820 32177 4829 32217
rect 4771 32176 4829 32177
rect 5347 32192 5405 32193
rect 2563 32151 2621 32152
rect 5347 32152 5356 32192
rect 5396 32152 5405 32192
rect 5347 32151 5405 32152
rect 6211 32192 6269 32193
rect 6211 32152 6220 32192
rect 6260 32152 6269 32192
rect 6211 32151 6269 32152
rect 7651 32192 7709 32193
rect 7651 32152 7660 32192
rect 7700 32152 7709 32192
rect 7651 32151 7709 32152
rect 8043 32192 8085 32201
rect 8043 32152 8044 32192
rect 8084 32152 8085 32192
rect 8043 32143 8085 32152
rect 8139 32192 8181 32201
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8235 32192 8277 32201
rect 8235 32152 8236 32192
rect 8276 32152 8277 32192
rect 8235 32143 8277 32152
rect 8803 32192 8861 32193
rect 8803 32152 8812 32192
rect 8852 32152 8861 32192
rect 8803 32151 8861 32152
rect 9667 32192 9725 32193
rect 9667 32152 9676 32192
rect 9716 32152 9725 32192
rect 9667 32151 9725 32152
rect 11011 32192 11069 32193
rect 11011 32152 11020 32192
rect 11060 32152 11069 32192
rect 11011 32151 11069 32152
rect 11883 32192 11925 32201
rect 11883 32152 11884 32192
rect 11924 32152 11925 32192
rect 11883 32143 11925 32152
rect 12259 32192 12317 32193
rect 12259 32152 12268 32192
rect 12308 32152 12317 32192
rect 12259 32151 12317 32152
rect 13123 32192 13181 32193
rect 13123 32152 13132 32192
rect 13172 32152 13181 32192
rect 13123 32151 13181 32152
rect 14851 32192 14909 32193
rect 14851 32152 14860 32192
rect 14900 32152 14909 32192
rect 14851 32151 14909 32152
rect 15339 32192 15381 32201
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15235 32150 15293 32151
rect 3723 32108 3765 32117
rect 3723 32068 3724 32108
rect 3764 32068 3765 32108
rect 3723 32059 3765 32068
rect 10827 32108 10869 32117
rect 15235 32110 15244 32150
rect 15284 32110 15293 32150
rect 15339 32143 15381 32152
rect 15435 32192 15477 32201
rect 15435 32152 15436 32192
rect 15476 32152 15477 32192
rect 15435 32143 15477 32152
rect 15627 32192 15669 32201
rect 15627 32152 15628 32192
rect 15668 32152 15669 32192
rect 15627 32143 15669 32152
rect 15723 32192 15765 32201
rect 15723 32152 15724 32192
rect 15764 32152 15765 32192
rect 15723 32143 15765 32152
rect 15819 32192 15861 32201
rect 15819 32152 15820 32192
rect 15860 32152 15861 32192
rect 15819 32143 15861 32152
rect 15915 32192 15957 32201
rect 15915 32152 15916 32192
rect 15956 32152 15957 32192
rect 15915 32143 15957 32152
rect 16107 32192 16149 32201
rect 16107 32152 16108 32192
rect 16148 32152 16149 32192
rect 16107 32143 16149 32152
rect 16771 32192 16829 32193
rect 16771 32152 16780 32192
rect 16820 32152 16829 32192
rect 16771 32151 16829 32152
rect 17635 32192 17693 32193
rect 17635 32152 17644 32192
rect 17684 32152 17693 32192
rect 17635 32151 17693 32152
rect 17931 32192 17973 32201
rect 17931 32152 17932 32192
rect 17972 32152 17973 32192
rect 17931 32143 17973 32152
rect 18027 32192 18069 32201
rect 18027 32152 18028 32192
rect 18068 32152 18069 32192
rect 18027 32143 18069 32152
rect 18123 32192 18165 32201
rect 18123 32152 18124 32192
rect 18164 32152 18165 32192
rect 18123 32143 18165 32152
rect 18403 32192 18461 32193
rect 18403 32152 18412 32192
rect 18452 32152 18461 32192
rect 18403 32151 18461 32152
rect 19267 32192 19325 32193
rect 19267 32152 19276 32192
rect 19316 32152 19325 32192
rect 19267 32151 19325 32152
rect 19947 32192 19989 32201
rect 19947 32152 19948 32192
rect 19988 32152 19989 32192
rect 19947 32143 19989 32152
rect 21283 32192 21341 32193
rect 21283 32152 21292 32192
rect 21332 32152 21341 32192
rect 21283 32151 21341 32152
rect 22147 32192 22205 32193
rect 22147 32152 22156 32192
rect 22196 32152 22205 32192
rect 22147 32151 22205 32152
rect 23499 32192 23541 32201
rect 23499 32152 23500 32192
rect 23540 32152 23541 32192
rect 23499 32143 23541 32152
rect 23691 32192 23733 32201
rect 23691 32152 23692 32192
rect 23732 32152 23733 32192
rect 23691 32143 23733 32152
rect 23779 32192 23837 32193
rect 23779 32152 23788 32192
rect 23828 32152 23837 32192
rect 23779 32151 23837 32152
rect 24843 32192 24885 32201
rect 24843 32152 24844 32192
rect 24884 32152 24885 32192
rect 24843 32143 24885 32152
rect 25219 32192 25277 32193
rect 25219 32152 25228 32192
rect 25268 32152 25277 32192
rect 25219 32151 25277 32152
rect 26083 32192 26141 32193
rect 26083 32152 26092 32192
rect 26132 32152 26141 32192
rect 26083 32151 26141 32152
rect 27523 32192 27581 32193
rect 27523 32152 27532 32192
rect 27572 32152 27581 32192
rect 27523 32151 27581 32152
rect 27819 32192 27861 32201
rect 27819 32152 27820 32192
rect 27860 32152 27861 32192
rect 27819 32143 27861 32152
rect 27915 32192 27957 32201
rect 27915 32152 27916 32192
rect 27956 32152 27957 32192
rect 27915 32143 27957 32152
rect 28387 32192 28445 32193
rect 28387 32152 28396 32192
rect 28436 32152 28445 32192
rect 28387 32151 28445 32152
rect 29347 32192 29405 32193
rect 29347 32152 29356 32192
rect 29396 32152 29405 32192
rect 29347 32151 29405 32152
rect 30499 32192 30557 32193
rect 30499 32152 30508 32192
rect 30548 32152 30557 32192
rect 30499 32151 30557 32152
rect 30883 32192 30941 32193
rect 30883 32152 30892 32192
rect 30932 32152 30941 32192
rect 30883 32151 30941 32152
rect 31179 32192 31221 32201
rect 31179 32152 31180 32192
rect 31220 32152 31221 32192
rect 31179 32143 31221 32152
rect 31275 32192 31317 32201
rect 31275 32152 31276 32192
rect 31316 32152 31317 32192
rect 31275 32143 31317 32152
rect 31947 32192 31989 32201
rect 31947 32152 31948 32192
rect 31988 32152 31989 32192
rect 31947 32143 31989 32152
rect 32043 32192 32085 32201
rect 32043 32152 32044 32192
rect 32084 32152 32085 32192
rect 32043 32143 32085 32152
rect 32139 32192 32181 32201
rect 32139 32152 32140 32192
rect 32180 32152 32181 32192
rect 32139 32143 32181 32152
rect 32331 32192 32373 32201
rect 32331 32152 32332 32192
rect 32372 32152 32373 32192
rect 32331 32143 32373 32152
rect 32427 32192 32469 32201
rect 32427 32152 32428 32192
rect 32468 32152 32469 32192
rect 32427 32143 32469 32152
rect 32523 32192 32565 32201
rect 32523 32152 32524 32192
rect 32564 32152 32565 32192
rect 32523 32143 32565 32152
rect 32619 32192 32661 32201
rect 32619 32152 32620 32192
rect 32660 32152 32661 32192
rect 32619 32143 32661 32152
rect 33475 32192 33533 32193
rect 33475 32152 33484 32192
rect 33524 32152 33533 32192
rect 33475 32151 33533 32152
rect 34051 32192 34109 32193
rect 34051 32152 34060 32192
rect 34100 32152 34109 32192
rect 34051 32151 34109 32152
rect 34915 32192 34973 32193
rect 34915 32152 34924 32192
rect 34964 32152 34973 32192
rect 34915 32151 34973 32152
rect 36643 32192 36701 32193
rect 36643 32152 36652 32192
rect 36692 32152 36701 32192
rect 36643 32151 36701 32152
rect 37603 32192 37661 32193
rect 37603 32152 37612 32192
rect 37652 32152 37661 32192
rect 37603 32151 37661 32152
rect 37987 32192 38045 32193
rect 37987 32152 37996 32192
rect 38036 32152 38045 32192
rect 37987 32151 38045 32152
rect 38179 32192 38237 32193
rect 38179 32152 38188 32192
rect 38228 32152 38237 32192
rect 38179 32151 38237 32152
rect 39235 32192 39293 32193
rect 39235 32152 39244 32192
rect 39284 32152 39293 32192
rect 39235 32151 39293 32152
rect 40099 32192 40157 32193
rect 40099 32152 40108 32192
rect 40148 32152 40157 32192
rect 40099 32151 40157 32152
rect 40483 32192 40541 32193
rect 40483 32152 40492 32192
rect 40532 32152 40541 32192
rect 40483 32151 40541 32152
rect 41443 32192 41501 32193
rect 41443 32152 41452 32192
rect 41492 32152 41501 32192
rect 41443 32151 41501 32152
rect 41923 32192 41981 32193
rect 41923 32152 41932 32192
rect 41972 32152 41981 32192
rect 41923 32151 41981 32152
rect 42027 32192 42069 32201
rect 42027 32152 42028 32192
rect 42068 32152 42069 32192
rect 42027 32143 42069 32152
rect 42219 32192 42261 32201
rect 42219 32152 42220 32192
rect 42260 32152 42261 32192
rect 42219 32143 42261 32152
rect 42403 32192 42461 32193
rect 42403 32152 42412 32192
rect 42452 32152 42461 32192
rect 42403 32151 42461 32152
rect 42507 32192 42549 32201
rect 42507 32152 42508 32192
rect 42548 32152 42549 32192
rect 42507 32143 42549 32152
rect 42699 32192 42741 32201
rect 42699 32152 42700 32192
rect 42740 32152 42741 32192
rect 42699 32143 42741 32152
rect 42891 32192 42933 32201
rect 42891 32152 42892 32192
rect 42932 32152 42933 32192
rect 42891 32143 42933 32152
rect 42987 32192 43029 32201
rect 42987 32152 42988 32192
rect 43028 32152 43029 32192
rect 42987 32143 43029 32152
rect 43083 32192 43125 32201
rect 43083 32152 43084 32192
rect 43124 32152 43125 32192
rect 43083 32143 43125 32152
rect 43179 32192 43221 32201
rect 43179 32152 43180 32192
rect 43220 32152 43221 32192
rect 43179 32143 43221 32152
rect 43459 32192 43517 32193
rect 43459 32152 43468 32192
rect 43508 32152 43517 32192
rect 43459 32151 43517 32152
rect 45091 32192 45149 32193
rect 45091 32152 45100 32192
rect 45140 32152 45149 32192
rect 45091 32151 45149 32152
rect 45955 32192 46013 32193
rect 45955 32152 45964 32192
rect 46004 32152 46013 32192
rect 45955 32151 46013 32152
rect 48067 32192 48125 32193
rect 48067 32152 48076 32192
rect 48116 32152 48125 32192
rect 48067 32151 48125 32152
rect 48267 32192 48309 32201
rect 48267 32152 48268 32192
rect 48308 32152 48309 32192
rect 48267 32143 48309 32152
rect 48363 32192 48405 32201
rect 48363 32152 48364 32192
rect 48404 32152 48405 32192
rect 48363 32143 48405 32152
rect 48459 32192 48501 32201
rect 48459 32152 48460 32192
rect 48500 32152 48501 32192
rect 48459 32143 48501 32152
rect 48555 32192 48597 32201
rect 48555 32152 48556 32192
rect 48596 32152 48597 32192
rect 48555 32143 48597 32152
rect 49795 32192 49853 32193
rect 49795 32152 49804 32192
rect 49844 32152 49853 32192
rect 49795 32151 49853 32152
rect 15235 32109 15293 32110
rect 10827 32068 10828 32108
rect 10868 32068 10869 32108
rect 10827 32059 10869 32068
rect 14667 32024 14709 32033
rect 14667 31984 14668 32024
rect 14708 31984 14709 32024
rect 14667 31975 14709 31984
rect 38379 32024 38421 32033
rect 38379 31984 38380 32024
rect 38420 31984 38421 32024
rect 38379 31975 38421 31984
rect 39051 32024 39093 32033
rect 39051 31984 39052 32024
rect 39092 31984 39093 32024
rect 39051 31975 39093 31984
rect 4099 31940 4157 31941
rect 4099 31900 4108 31940
rect 4148 31900 4157 31940
rect 4099 31899 4157 31900
rect 7363 31940 7421 31941
rect 7363 31900 7372 31940
rect 7412 31900 7421 31940
rect 7363 31899 7421 31900
rect 11683 31940 11741 31941
rect 11683 31900 11692 31940
rect 11732 31900 11741 31940
rect 11683 31899 11741 31900
rect 16963 31940 17021 31941
rect 16963 31900 16972 31940
rect 17012 31900 17021 31940
rect 16963 31899 17021 31900
rect 28195 31940 28253 31941
rect 28195 31900 28204 31940
rect 28244 31900 28253 31940
rect 28195 31899 28253 31900
rect 28675 31940 28733 31941
rect 28675 31900 28684 31940
rect 28724 31900 28733 31940
rect 28675 31899 28733 31900
rect 30027 31940 30069 31949
rect 30027 31900 30028 31940
rect 30068 31900 30069 31940
rect 30027 31891 30069 31900
rect 31555 31940 31613 31941
rect 31555 31900 31564 31940
rect 31604 31900 31613 31940
rect 31555 31899 31613 31900
rect 32803 31940 32861 31941
rect 32803 31900 32812 31940
rect 32852 31900 32861 31940
rect 32803 31899 32861 31900
rect 36555 31940 36597 31949
rect 36555 31900 36556 31940
rect 36596 31900 36597 31940
rect 36555 31891 36597 31900
rect 39907 31940 39965 31941
rect 39907 31900 39916 31940
rect 39956 31900 39965 31940
rect 39907 31899 39965 31900
rect 42699 31940 42741 31949
rect 42699 31900 42700 31940
rect 42740 31900 42741 31940
rect 42699 31891 42741 31900
rect 47107 31940 47165 31941
rect 47107 31900 47116 31940
rect 47156 31900 47165 31940
rect 47107 31899 47165 31900
rect 47395 31940 47453 31941
rect 47395 31900 47404 31940
rect 47444 31900 47453 31940
rect 47395 31899 47453 31900
rect 49123 31940 49181 31941
rect 49123 31900 49132 31940
rect 49172 31900 49181 31940
rect 49123 31899 49181 31900
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 11499 31604 11541 31613
rect 11499 31564 11500 31604
rect 11540 31564 11541 31604
rect 11499 31555 11541 31564
rect 12267 31604 12309 31613
rect 12267 31564 12268 31604
rect 12308 31564 12309 31604
rect 12267 31555 12309 31564
rect 42027 31604 42069 31613
rect 42027 31564 42028 31604
rect 42068 31564 42069 31604
rect 42027 31555 42069 31564
rect 49699 31604 49757 31605
rect 49699 31564 49708 31604
rect 49748 31564 49757 31604
rect 49699 31563 49757 31564
rect 1899 31520 1941 31529
rect 1899 31480 1900 31520
rect 1940 31480 1941 31520
rect 1899 31471 1941 31480
rect 3435 31520 3477 31529
rect 3435 31480 3436 31520
rect 3476 31480 3477 31520
rect 3435 31471 3477 31480
rect 5547 31520 5589 31529
rect 5547 31480 5548 31520
rect 5588 31480 5589 31520
rect 5547 31471 5589 31480
rect 6699 31520 6741 31529
rect 6699 31480 6700 31520
rect 6740 31480 6741 31520
rect 6699 31471 6741 31480
rect 7371 31520 7413 31529
rect 7371 31480 7372 31520
rect 7412 31480 7413 31520
rect 7371 31471 7413 31480
rect 7659 31520 7701 31529
rect 7659 31480 7660 31520
rect 7700 31480 7701 31520
rect 7659 31471 7701 31480
rect 7851 31520 7893 31529
rect 7851 31480 7852 31520
rect 7892 31480 7893 31520
rect 7851 31471 7893 31480
rect 8331 31520 8373 31529
rect 8331 31480 8332 31520
rect 8372 31480 8373 31520
rect 8331 31471 8373 31480
rect 9963 31520 10005 31529
rect 9963 31480 9964 31520
rect 10004 31480 10005 31520
rect 9963 31471 10005 31480
rect 10443 31520 10485 31529
rect 10443 31480 10444 31520
rect 10484 31480 10485 31520
rect 10443 31471 10485 31480
rect 11691 31520 11733 31529
rect 11691 31480 11692 31520
rect 11732 31480 11733 31520
rect 11691 31471 11733 31480
rect 14083 31520 14141 31521
rect 14083 31480 14092 31520
rect 14132 31480 14141 31520
rect 14083 31479 14141 31480
rect 16779 31520 16821 31529
rect 16779 31480 16780 31520
rect 16820 31480 16821 31520
rect 16779 31471 16821 31480
rect 19363 31520 19421 31521
rect 19363 31480 19372 31520
rect 19412 31480 19421 31520
rect 19363 31479 19421 31480
rect 19755 31520 19797 31529
rect 19755 31480 19756 31520
rect 19796 31480 19797 31520
rect 19755 31471 19797 31480
rect 20811 31520 20853 31529
rect 20811 31480 20812 31520
rect 20852 31480 20853 31520
rect 20811 31471 20853 31480
rect 23019 31520 23061 31529
rect 23019 31480 23020 31520
rect 23060 31480 23061 31520
rect 23019 31471 23061 31480
rect 24075 31520 24117 31529
rect 24075 31480 24076 31520
rect 24116 31480 24117 31520
rect 24075 31471 24117 31480
rect 24555 31520 24597 31529
rect 24555 31480 24556 31520
rect 24596 31480 24597 31520
rect 24555 31471 24597 31480
rect 28779 31520 28821 31529
rect 28779 31480 28780 31520
rect 28820 31480 28821 31520
rect 28779 31471 28821 31480
rect 33099 31520 33141 31529
rect 33099 31480 33100 31520
rect 33140 31480 33141 31520
rect 33099 31471 33141 31480
rect 34539 31520 34581 31529
rect 34539 31480 34540 31520
rect 34580 31480 34581 31520
rect 34539 31471 34581 31480
rect 45099 31520 45141 31529
rect 45099 31480 45100 31520
rect 45140 31480 45141 31520
rect 45099 31471 45141 31480
rect 46443 31520 46485 31529
rect 46443 31480 46444 31520
rect 46484 31480 46485 31520
rect 46443 31471 46485 31480
rect 10819 31436 10877 31437
rect 10819 31396 10828 31436
rect 10868 31396 10877 31436
rect 10819 31395 10877 31396
rect 13323 31436 13365 31445
rect 13323 31396 13324 31436
rect 13364 31396 13365 31436
rect 13323 31387 13365 31396
rect 3523 31352 3581 31353
rect 3523 31312 3532 31352
rect 3572 31312 3581 31352
rect 3523 31311 3581 31312
rect 3811 31352 3869 31353
rect 3811 31312 3820 31352
rect 3860 31312 3869 31352
rect 3811 31311 3869 31312
rect 4011 31352 4053 31361
rect 4011 31312 4012 31352
rect 4052 31312 4053 31352
rect 4011 31303 4053 31312
rect 4107 31352 4149 31361
rect 4107 31312 4108 31352
rect 4148 31312 4149 31352
rect 4107 31303 4149 31312
rect 4203 31352 4245 31361
rect 4203 31312 4204 31352
rect 4244 31312 4245 31352
rect 4203 31303 4245 31312
rect 4299 31352 4341 31361
rect 4299 31312 4300 31352
rect 4340 31312 4341 31352
rect 4299 31303 4341 31312
rect 4491 31352 4533 31361
rect 4491 31312 4492 31352
rect 4532 31312 4533 31352
rect 4491 31303 4533 31312
rect 4683 31352 4725 31361
rect 4683 31312 4684 31352
rect 4724 31312 4725 31352
rect 4683 31303 4725 31312
rect 4771 31352 4829 31353
rect 4771 31312 4780 31352
rect 4820 31312 4829 31352
rect 4771 31311 4829 31312
rect 4963 31352 5021 31353
rect 4963 31312 4972 31352
rect 5012 31312 5021 31352
rect 4963 31311 5021 31312
rect 5067 31352 5109 31361
rect 5067 31312 5068 31352
rect 5108 31312 5109 31352
rect 5067 31303 5109 31312
rect 5251 31352 5309 31353
rect 5251 31312 5260 31352
rect 5300 31312 5309 31352
rect 5251 31311 5309 31312
rect 5355 31352 5397 31361
rect 5355 31312 5356 31352
rect 5396 31312 5397 31352
rect 5355 31303 5397 31312
rect 5547 31352 5589 31361
rect 5547 31312 5548 31352
rect 5588 31312 5589 31352
rect 5547 31303 5589 31312
rect 6123 31352 6165 31361
rect 6123 31312 6124 31352
rect 6164 31312 6165 31352
rect 6123 31303 6165 31312
rect 6979 31352 7037 31353
rect 6979 31312 6988 31352
rect 7028 31312 7037 31352
rect 6979 31311 7037 31312
rect 7555 31352 7613 31353
rect 7555 31312 7564 31352
rect 7604 31312 7613 31352
rect 7555 31311 7613 31312
rect 7939 31352 7997 31353
rect 7939 31312 7948 31352
rect 7988 31312 7997 31352
rect 7939 31311 7997 31312
rect 8515 31352 8573 31353
rect 8515 31312 8524 31352
rect 8564 31312 8573 31352
rect 8515 31311 8573 31312
rect 8619 31352 8661 31361
rect 8619 31312 8620 31352
rect 8660 31312 8661 31352
rect 8619 31303 8661 31312
rect 8811 31352 8853 31361
rect 8811 31312 8812 31352
rect 8852 31312 8853 31352
rect 8811 31303 8853 31312
rect 9667 31352 9725 31353
rect 9667 31312 9676 31352
rect 9716 31312 9725 31352
rect 9667 31311 9725 31312
rect 10051 31352 10109 31353
rect 10051 31312 10060 31352
rect 10100 31312 10109 31352
rect 10051 31311 10109 31312
rect 11883 31352 11925 31361
rect 11883 31312 11884 31352
rect 11924 31312 11925 31352
rect 11883 31303 11925 31312
rect 12267 31352 12309 31361
rect 12267 31312 12268 31352
rect 12308 31312 12309 31352
rect 12267 31303 12309 31312
rect 12459 31352 12501 31361
rect 12459 31312 12460 31352
rect 12500 31312 12501 31352
rect 12459 31303 12501 31312
rect 12547 31352 12605 31353
rect 12547 31312 12556 31352
rect 12596 31312 12605 31352
rect 12547 31311 12605 31312
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 12843 31352 12885 31361
rect 12843 31312 12844 31352
rect 12884 31312 12885 31352
rect 12843 31303 12885 31312
rect 12939 31352 12981 31361
rect 12939 31312 12940 31352
rect 12980 31312 12981 31352
rect 12939 31303 12981 31312
rect 13035 31352 13077 31361
rect 13035 31312 13036 31352
rect 13076 31312 13077 31352
rect 13035 31303 13077 31312
rect 13219 31352 13277 31353
rect 13219 31312 13228 31352
rect 13268 31312 13277 31352
rect 13219 31311 13277 31312
rect 13603 31352 13661 31353
rect 13603 31312 13612 31352
rect 13652 31312 13661 31352
rect 13603 31311 13661 31312
rect 13795 31352 13853 31353
rect 13795 31312 13804 31352
rect 13844 31312 13853 31352
rect 13795 31311 13853 31312
rect 14379 31352 14421 31361
rect 14379 31312 14380 31352
rect 14420 31312 14421 31352
rect 14379 31303 14421 31312
rect 14475 31352 14517 31361
rect 14475 31312 14476 31352
rect 14516 31312 14517 31352
rect 14475 31303 14517 31312
rect 14755 31352 14813 31353
rect 14755 31312 14764 31352
rect 14804 31312 14813 31352
rect 14755 31311 14813 31312
rect 15243 31352 15285 31361
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 15907 31352 15965 31353
rect 15907 31312 15916 31352
rect 15956 31312 15965 31352
rect 15907 31311 15965 31312
rect 16195 31352 16253 31353
rect 16195 31312 16204 31352
rect 16244 31312 16253 31352
rect 16195 31311 16253 31312
rect 16483 31352 16541 31353
rect 16483 31312 16492 31352
rect 16532 31312 16541 31352
rect 16483 31311 16541 31312
rect 16587 31352 16629 31361
rect 16587 31312 16588 31352
rect 16628 31312 16629 31352
rect 16587 31303 16629 31312
rect 16779 31352 16821 31361
rect 16779 31312 16780 31352
rect 16820 31312 16821 31352
rect 16779 31303 16821 31312
rect 16971 31352 17013 31361
rect 16971 31312 16972 31352
rect 17012 31312 17013 31352
rect 16971 31303 17013 31312
rect 17347 31352 17405 31353
rect 17347 31312 17356 31352
rect 17396 31312 17405 31352
rect 17347 31311 17405 31312
rect 18211 31352 18269 31353
rect 18211 31312 18220 31352
rect 18260 31312 18269 31352
rect 18211 31311 18269 31312
rect 20611 31352 20669 31353
rect 20611 31312 20620 31352
rect 20660 31312 20669 31352
rect 20611 31311 20669 31312
rect 20811 31352 20853 31361
rect 20811 31312 20812 31352
rect 20852 31312 20853 31352
rect 20811 31303 20853 31312
rect 21003 31352 21045 31361
rect 21003 31312 21004 31352
rect 21044 31312 21045 31352
rect 21003 31303 21045 31312
rect 21091 31352 21149 31353
rect 21091 31312 21100 31352
rect 21140 31312 21149 31352
rect 21091 31311 21149 31312
rect 21283 31352 21341 31353
rect 21283 31312 21292 31352
rect 21332 31312 21341 31352
rect 21283 31311 21341 31312
rect 24163 31352 24221 31353
rect 24163 31312 24172 31352
rect 24212 31312 24221 31352
rect 24163 31311 24221 31312
rect 25411 31352 25469 31353
rect 25411 31312 25420 31352
rect 25460 31312 25469 31352
rect 25411 31311 25469 31312
rect 25899 31352 25941 31361
rect 25899 31312 25900 31352
rect 25940 31312 25941 31352
rect 25899 31303 25941 31312
rect 26091 31352 26133 31361
rect 26091 31312 26092 31352
rect 26132 31312 26133 31352
rect 26091 31303 26133 31312
rect 26179 31352 26237 31353
rect 26179 31312 26188 31352
rect 26228 31312 26237 31352
rect 26179 31311 26237 31312
rect 26371 31352 26429 31353
rect 26371 31312 26380 31352
rect 26420 31312 26429 31352
rect 26371 31311 26429 31312
rect 27051 31352 27093 31361
rect 27051 31312 27052 31352
rect 27092 31312 27093 31352
rect 27051 31303 27093 31312
rect 27339 31352 27381 31361
rect 27339 31312 27340 31352
rect 27380 31312 27381 31352
rect 27339 31303 27381 31312
rect 27435 31352 27477 31361
rect 27435 31312 27436 31352
rect 27476 31312 27477 31352
rect 27435 31303 27477 31312
rect 27531 31352 27573 31361
rect 27531 31312 27532 31352
rect 27572 31312 27573 31352
rect 27531 31303 27573 31312
rect 27627 31352 27669 31361
rect 27627 31312 27628 31352
rect 27668 31312 27669 31352
rect 27627 31303 27669 31312
rect 27811 31352 27869 31353
rect 27811 31312 27820 31352
rect 27860 31312 27869 31352
rect 27811 31311 27869 31312
rect 27915 31352 27957 31361
rect 27915 31312 27916 31352
rect 27956 31312 27957 31352
rect 27915 31303 27957 31312
rect 28107 31352 28149 31361
rect 28107 31312 28108 31352
rect 28148 31312 28149 31352
rect 28107 31303 28149 31312
rect 28291 31352 28349 31353
rect 28291 31312 28300 31352
rect 28340 31312 28349 31352
rect 28291 31311 28349 31312
rect 28971 31352 29013 31361
rect 28971 31312 28972 31352
rect 29012 31312 29013 31352
rect 28971 31303 29013 31312
rect 29347 31352 29405 31353
rect 29347 31312 29356 31352
rect 29396 31312 29405 31352
rect 29347 31311 29405 31312
rect 30211 31352 30269 31353
rect 30211 31312 30220 31352
rect 30260 31312 30269 31352
rect 30211 31311 30269 31312
rect 31555 31352 31613 31353
rect 31555 31312 31564 31352
rect 31604 31312 31613 31352
rect 31555 31311 31613 31312
rect 32515 31352 32573 31353
rect 32515 31312 32524 31352
rect 32564 31312 32573 31352
rect 32515 31311 32573 31312
rect 33283 31352 33341 31353
rect 33283 31312 33292 31352
rect 33332 31312 33341 31352
rect 33283 31311 33341 31312
rect 33387 31352 33429 31361
rect 33387 31312 33388 31352
rect 33428 31312 33429 31352
rect 33387 31303 33429 31312
rect 33579 31352 33621 31361
rect 33579 31312 33580 31352
rect 33620 31312 33621 31352
rect 33579 31303 33621 31312
rect 33867 31352 33909 31361
rect 33867 31312 33868 31352
rect 33908 31312 33909 31352
rect 33867 31303 33909 31312
rect 33963 31352 34005 31361
rect 33963 31312 33964 31352
rect 34004 31312 34005 31352
rect 33963 31303 34005 31312
rect 34059 31352 34101 31361
rect 34059 31312 34060 31352
rect 34100 31312 34101 31352
rect 34059 31303 34101 31312
rect 34243 31352 34301 31353
rect 34243 31312 34252 31352
rect 34292 31312 34301 31352
rect 34243 31311 34301 31312
rect 34347 31352 34389 31361
rect 34347 31312 34348 31352
rect 34388 31312 34389 31352
rect 34347 31303 34389 31312
rect 34539 31352 34581 31361
rect 34539 31312 34540 31352
rect 34580 31312 34581 31352
rect 34539 31303 34581 31312
rect 35019 31352 35061 31361
rect 35019 31312 35020 31352
rect 35060 31312 35061 31352
rect 35019 31303 35061 31312
rect 35395 31352 35453 31353
rect 35395 31312 35404 31352
rect 35444 31312 35453 31352
rect 35395 31311 35453 31312
rect 36259 31352 36317 31353
rect 36259 31312 36268 31352
rect 36308 31312 36317 31352
rect 36259 31311 36317 31312
rect 38283 31352 38325 31361
rect 38283 31312 38284 31352
rect 38324 31312 38325 31352
rect 38283 31303 38325 31312
rect 39715 31352 39773 31353
rect 39715 31312 39724 31352
rect 39764 31312 39773 31352
rect 39715 31311 39773 31312
rect 40579 31352 40637 31353
rect 40579 31312 40588 31352
rect 40628 31312 40637 31352
rect 40579 31311 40637 31312
rect 41923 31352 41981 31353
rect 41923 31312 41932 31352
rect 41972 31312 41981 31352
rect 41923 31311 41981 31312
rect 42883 31352 42941 31353
rect 42883 31312 42892 31352
rect 42932 31312 42941 31352
rect 42883 31311 42941 31312
rect 43075 31352 43133 31353
rect 43075 31312 43084 31352
rect 43124 31312 43133 31352
rect 43075 31311 43133 31312
rect 44611 31352 44669 31353
rect 44611 31312 44620 31352
rect 44660 31312 44669 31352
rect 44611 31311 44669 31312
rect 44803 31352 44861 31353
rect 44803 31312 44812 31352
rect 44852 31312 44861 31352
rect 44803 31311 44861 31312
rect 44907 31352 44949 31361
rect 44907 31312 44908 31352
rect 44948 31312 44949 31352
rect 44907 31303 44949 31312
rect 45099 31352 45141 31361
rect 45099 31312 45100 31352
rect 45140 31312 45141 31352
rect 45099 31303 45141 31312
rect 45283 31352 45341 31353
rect 45283 31312 45292 31352
rect 45332 31312 45341 31352
rect 45283 31311 45341 31312
rect 45579 31352 45621 31361
rect 45579 31312 45580 31352
rect 45620 31312 45621 31352
rect 45579 31303 45621 31312
rect 45675 31352 45717 31361
rect 45675 31312 45676 31352
rect 45716 31312 45717 31352
rect 45675 31303 45717 31312
rect 45771 31352 45813 31361
rect 45771 31312 45772 31352
rect 45812 31312 45813 31352
rect 45771 31303 45813 31312
rect 45867 31352 45909 31361
rect 45867 31312 45868 31352
rect 45908 31312 45909 31352
rect 45867 31303 45909 31312
rect 46251 31352 46293 31361
rect 46251 31312 46252 31352
rect 46292 31312 46293 31352
rect 46251 31303 46293 31312
rect 47307 31352 47349 31361
rect 47307 31312 47308 31352
rect 47348 31312 47349 31352
rect 47307 31303 47349 31312
rect 47683 31352 47741 31353
rect 47683 31312 47692 31352
rect 47732 31312 47741 31352
rect 47683 31311 47741 31312
rect 48547 31352 48605 31353
rect 48547 31312 48556 31352
rect 48596 31312 48605 31352
rect 48547 31311 48605 31312
rect 8715 31268 8757 31277
rect 8715 31228 8716 31268
rect 8756 31228 8757 31268
rect 8715 31219 8757 31228
rect 13899 31268 13941 31277
rect 13899 31228 13900 31268
rect 13940 31228 13941 31268
rect 13899 31219 13941 31228
rect 25995 31268 26037 31277
rect 25995 31228 25996 31268
rect 26036 31228 26037 31268
rect 25995 31219 26037 31228
rect 28011 31268 28053 31277
rect 28011 31228 28012 31268
rect 28052 31228 28053 31268
rect 28011 31219 28053 31228
rect 28395 31268 28437 31277
rect 28395 31228 28396 31268
rect 28436 31228 28437 31268
rect 28395 31219 28437 31228
rect 33483 31268 33525 31277
rect 33483 31228 33484 31268
rect 33524 31228 33525 31268
rect 33483 31219 33525 31228
rect 39339 31268 39381 31277
rect 39339 31228 39340 31268
rect 39380 31228 39381 31268
rect 39339 31219 39381 31228
rect 45387 31268 45429 31277
rect 45387 31228 45388 31268
rect 45428 31228 45429 31268
rect 45387 31219 45429 31228
rect 3723 31184 3765 31193
rect 3723 31144 3724 31184
rect 3764 31144 3765 31184
rect 3723 31135 3765 31144
rect 4579 31184 4637 31185
rect 4579 31144 4588 31184
rect 4628 31144 4637 31184
rect 4579 31143 4637 31144
rect 8995 31184 9053 31185
rect 8995 31144 9004 31184
rect 9044 31144 9053 31184
rect 8995 31143 9053 31144
rect 13515 31184 13557 31193
rect 13515 31144 13516 31184
rect 13556 31144 13557 31184
rect 13515 31135 13557 31144
rect 16107 31184 16149 31193
rect 16107 31144 16108 31184
rect 16148 31144 16149 31184
rect 16107 31135 16149 31144
rect 19939 31184 19997 31185
rect 19939 31144 19948 31184
rect 19988 31144 19997 31184
rect 19939 31143 19997 31144
rect 21387 31184 21429 31193
rect 21387 31144 21388 31184
rect 21428 31144 21429 31184
rect 21387 31135 21429 31144
rect 24739 31184 24797 31185
rect 24739 31144 24748 31184
rect 24788 31144 24797 31184
rect 24739 31143 24797 31144
rect 31363 31184 31421 31185
rect 31363 31144 31372 31184
rect 31412 31144 31421 31184
rect 31363 31143 31421 31144
rect 32227 31184 32285 31185
rect 32227 31144 32236 31184
rect 32276 31144 32285 31184
rect 32227 31143 32285 31144
rect 32427 31184 32469 31193
rect 32427 31144 32428 31184
rect 32468 31144 32469 31184
rect 32427 31135 32469 31144
rect 33763 31184 33821 31185
rect 33763 31144 33772 31184
rect 33812 31144 33821 31184
rect 33763 31143 33821 31144
rect 37411 31184 37469 31185
rect 37411 31144 37420 31184
rect 37460 31144 37469 31184
rect 37411 31143 37469 31144
rect 38667 31184 38709 31193
rect 38667 31144 38668 31184
rect 38708 31144 38709 31184
rect 38667 31135 38709 31144
rect 41731 31184 41789 31185
rect 41731 31144 41740 31184
rect 41780 31144 41789 31184
rect 41731 31143 41789 31144
rect 42211 31184 42269 31185
rect 42211 31144 42220 31184
rect 42260 31144 42269 31184
rect 42211 31143 42269 31144
rect 43747 31184 43805 31185
rect 43747 31144 43756 31184
rect 43796 31144 43805 31184
rect 43747 31143 43805 31144
rect 43939 31184 43997 31185
rect 43939 31144 43948 31184
rect 43988 31144 43997 31184
rect 43939 31143 43997 31144
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 4003 30848 4061 30849
rect 4003 30808 4012 30848
rect 4052 30808 4061 30848
rect 4003 30807 4061 30808
rect 4867 30848 4925 30849
rect 4867 30808 4876 30848
rect 4916 30808 4925 30848
rect 4867 30807 4925 30808
rect 12931 30848 12989 30849
rect 12931 30808 12940 30848
rect 12980 30808 12989 30848
rect 12931 30807 12989 30808
rect 25027 30848 25085 30849
rect 25027 30808 25036 30848
rect 25076 30808 25085 30848
rect 25027 30807 25085 30808
rect 31075 30848 31133 30849
rect 31075 30808 31084 30848
rect 31124 30808 31133 30848
rect 31075 30807 31133 30808
rect 31275 30848 31317 30857
rect 31275 30808 31276 30848
rect 31316 30808 31317 30848
rect 31275 30799 31317 30808
rect 31563 30848 31605 30857
rect 31563 30808 31564 30848
rect 31604 30808 31605 30848
rect 31563 30799 31605 30808
rect 38659 30848 38717 30849
rect 38659 30808 38668 30848
rect 38708 30808 38717 30848
rect 38659 30807 38717 30808
rect 40971 30848 41013 30857
rect 40971 30808 40972 30848
rect 41012 30808 41013 30848
rect 40971 30799 41013 30808
rect 44611 30848 44669 30849
rect 44611 30808 44620 30848
rect 44660 30808 44669 30848
rect 44611 30807 44669 30808
rect 47203 30848 47261 30849
rect 47203 30808 47212 30848
rect 47252 30808 47261 30848
rect 47203 30807 47261 30808
rect 8619 30764 8661 30773
rect 8619 30724 8620 30764
rect 8660 30724 8661 30764
rect 8619 30715 8661 30724
rect 27723 30764 27765 30773
rect 27723 30724 27724 30764
rect 27764 30724 27765 30764
rect 27723 30715 27765 30724
rect 42219 30764 42261 30773
rect 42219 30724 42220 30764
rect 42260 30724 42261 30764
rect 42219 30715 42261 30724
rect 1323 30680 1365 30689
rect 1323 30640 1324 30680
rect 1364 30640 1365 30680
rect 1323 30631 1365 30640
rect 1699 30680 1757 30681
rect 1699 30640 1708 30680
rect 1748 30640 1757 30680
rect 1699 30639 1757 30640
rect 2563 30680 2621 30681
rect 2563 30640 2572 30680
rect 2612 30640 2621 30680
rect 2563 30639 2621 30640
rect 4675 30680 4733 30681
rect 4675 30640 4684 30680
rect 4724 30640 4733 30680
rect 4675 30639 4733 30640
rect 5539 30680 5597 30681
rect 5539 30640 5548 30680
rect 5588 30640 5597 30680
rect 5539 30639 5597 30640
rect 6595 30680 6653 30681
rect 6595 30640 6604 30680
rect 6644 30640 6653 30680
rect 6595 30639 6653 30640
rect 6891 30680 6933 30689
rect 6891 30640 6892 30680
rect 6932 30640 6933 30680
rect 6891 30631 6933 30640
rect 6987 30680 7029 30689
rect 6987 30640 6988 30680
rect 7028 30640 7029 30680
rect 6987 30631 7029 30640
rect 7371 30680 7413 30689
rect 7371 30640 7372 30680
rect 7412 30640 7413 30680
rect 7371 30631 7413 30640
rect 7939 30680 7997 30681
rect 7939 30640 7948 30680
rect 7988 30640 7997 30680
rect 9667 30680 9725 30681
rect 7939 30639 7997 30640
rect 8427 30666 8469 30675
rect 8427 30626 8428 30666
rect 8468 30626 8469 30666
rect 9667 30640 9676 30680
rect 9716 30640 9725 30680
rect 9667 30639 9725 30640
rect 10923 30680 10965 30689
rect 10923 30640 10924 30680
rect 10964 30640 10965 30680
rect 10923 30631 10965 30640
rect 11019 30680 11061 30689
rect 11019 30640 11020 30680
rect 11060 30640 11061 30680
rect 11019 30631 11061 30640
rect 11115 30680 11157 30689
rect 11115 30640 11116 30680
rect 11156 30640 11157 30680
rect 11115 30631 11157 30640
rect 11211 30680 11253 30689
rect 11211 30640 11212 30680
rect 11252 30640 11253 30680
rect 11211 30631 11253 30640
rect 12067 30680 12125 30681
rect 12067 30640 12076 30680
rect 12116 30640 12125 30680
rect 12067 30639 12125 30640
rect 12259 30680 12317 30681
rect 12259 30640 12268 30680
rect 12308 30640 12317 30680
rect 12259 30639 12317 30640
rect 13123 30680 13181 30681
rect 13123 30640 13132 30680
rect 13172 30640 13181 30680
rect 13123 30639 13181 30640
rect 13323 30680 13365 30689
rect 13323 30640 13324 30680
rect 13364 30640 13365 30680
rect 13323 30631 13365 30640
rect 13507 30680 13565 30681
rect 13507 30640 13516 30680
rect 13556 30640 13565 30680
rect 13507 30639 13565 30640
rect 13611 30680 13653 30689
rect 13611 30640 13612 30680
rect 13652 30640 13653 30680
rect 13611 30631 13653 30640
rect 13803 30680 13845 30689
rect 13803 30640 13804 30680
rect 13844 30640 13845 30680
rect 13803 30631 13845 30640
rect 13987 30680 14045 30681
rect 13987 30640 13996 30680
rect 14036 30640 14045 30680
rect 13987 30639 14045 30640
rect 14947 30680 15005 30681
rect 14947 30640 14956 30680
rect 14996 30640 15005 30680
rect 14947 30639 15005 30640
rect 15907 30680 15965 30681
rect 15907 30640 15916 30680
rect 15956 30640 15965 30680
rect 15907 30639 15965 30640
rect 19651 30680 19709 30681
rect 19651 30640 19660 30680
rect 19700 30640 19709 30680
rect 19651 30639 19709 30640
rect 19947 30680 19989 30689
rect 19947 30640 19948 30680
rect 19988 30640 19989 30680
rect 19947 30631 19989 30640
rect 20323 30680 20381 30681
rect 20323 30640 20332 30680
rect 20372 30640 20381 30680
rect 20323 30639 20381 30640
rect 21187 30680 21245 30681
rect 21187 30640 21196 30680
rect 21236 30640 21245 30680
rect 21187 30639 21245 30640
rect 22635 30680 22677 30689
rect 22635 30640 22636 30680
rect 22676 30640 22677 30680
rect 22635 30631 22677 30640
rect 23011 30680 23069 30681
rect 23011 30640 23020 30680
rect 23060 30640 23069 30680
rect 23011 30639 23069 30640
rect 23875 30680 23933 30681
rect 23875 30640 23884 30680
rect 23924 30640 23933 30680
rect 23875 30639 23933 30640
rect 25515 30680 25557 30689
rect 25515 30640 25516 30680
rect 25556 30640 25557 30680
rect 25515 30631 25557 30640
rect 25611 30680 25653 30689
rect 25611 30640 25612 30680
rect 25652 30640 25653 30680
rect 25611 30631 25653 30640
rect 25707 30680 25749 30689
rect 25707 30640 25708 30680
rect 25748 30640 25749 30680
rect 25707 30631 25749 30640
rect 25803 30680 25845 30689
rect 25803 30640 25804 30680
rect 25844 30640 25845 30680
rect 25803 30631 25845 30640
rect 25987 30680 26045 30681
rect 25987 30640 25996 30680
rect 26036 30640 26045 30680
rect 25987 30639 26045 30640
rect 26947 30680 27005 30681
rect 26947 30640 26956 30680
rect 26996 30640 27005 30680
rect 26947 30639 27005 30640
rect 27331 30680 27389 30681
rect 27331 30640 27340 30680
rect 27380 30640 27389 30680
rect 27331 30639 27389 30640
rect 27627 30680 27669 30689
rect 27627 30640 27628 30680
rect 27668 30640 27669 30680
rect 27627 30631 27669 30640
rect 28395 30680 28437 30689
rect 28395 30640 28396 30680
rect 28436 30640 28437 30680
rect 28395 30631 28437 30640
rect 28491 30680 28533 30689
rect 28491 30640 28492 30680
rect 28532 30640 28533 30680
rect 28491 30631 28533 30640
rect 28587 30680 28629 30689
rect 28587 30640 28588 30680
rect 28628 30640 28629 30680
rect 28587 30631 28629 30640
rect 28683 30680 28725 30689
rect 28683 30640 28684 30680
rect 28724 30640 28725 30680
rect 28683 30631 28725 30640
rect 29731 30680 29789 30681
rect 29731 30640 29740 30680
rect 29780 30640 29789 30680
rect 29731 30639 29789 30640
rect 30595 30680 30653 30681
rect 30595 30640 30604 30680
rect 30644 30640 30653 30680
rect 30595 30639 30653 30640
rect 30795 30680 30837 30689
rect 30795 30640 30796 30680
rect 30836 30640 30837 30680
rect 30795 30631 30837 30640
rect 30891 30680 30933 30689
rect 30891 30640 30892 30680
rect 30932 30640 30933 30680
rect 30891 30631 30933 30640
rect 30987 30680 31029 30689
rect 30987 30640 30988 30680
rect 31028 30640 31029 30680
rect 30987 30631 31029 30640
rect 31363 30680 31421 30681
rect 31363 30640 31372 30680
rect 31412 30640 31421 30680
rect 31363 30639 31421 30640
rect 31651 30680 31709 30681
rect 31651 30640 31660 30680
rect 31700 30640 31709 30680
rect 31651 30639 31709 30640
rect 32419 30680 32477 30681
rect 32419 30640 32428 30680
rect 32468 30640 32477 30680
rect 32419 30639 32477 30640
rect 34243 30680 34301 30681
rect 34243 30640 34252 30680
rect 34292 30640 34301 30680
rect 34243 30639 34301 30640
rect 35107 30680 35165 30681
rect 35107 30640 35116 30680
rect 35156 30640 35165 30680
rect 35107 30639 35165 30640
rect 35307 30680 35349 30689
rect 35307 30640 35308 30680
rect 35348 30640 35349 30680
rect 35307 30631 35349 30640
rect 35403 30680 35445 30689
rect 35403 30640 35404 30680
rect 35444 30640 35445 30680
rect 35403 30631 35445 30640
rect 35499 30680 35541 30689
rect 35499 30640 35500 30680
rect 35540 30640 35541 30680
rect 35499 30631 35541 30640
rect 35595 30680 35637 30689
rect 35595 30640 35596 30680
rect 35636 30640 35637 30680
rect 35595 30631 35637 30640
rect 36643 30680 36701 30681
rect 36643 30640 36652 30680
rect 36692 30640 36701 30680
rect 36643 30639 36701 30640
rect 37027 30680 37085 30681
rect 37027 30640 37036 30680
rect 37076 30640 37085 30680
rect 37027 30639 37085 30640
rect 37227 30680 37269 30689
rect 37227 30640 37228 30680
rect 37268 30640 37269 30680
rect 37227 30631 37269 30640
rect 38083 30680 38141 30681
rect 38083 30640 38092 30680
rect 38132 30640 38141 30680
rect 38083 30639 38141 30640
rect 38187 30680 38229 30689
rect 38187 30640 38188 30680
rect 38228 30640 38229 30680
rect 38187 30631 38229 30640
rect 38379 30680 38421 30689
rect 38379 30640 38380 30680
rect 38420 30640 38421 30680
rect 38379 30631 38421 30640
rect 38571 30680 38613 30689
rect 38571 30640 38572 30680
rect 38612 30640 38613 30680
rect 38571 30631 38613 30640
rect 38763 30680 38805 30689
rect 38763 30640 38764 30680
rect 38804 30640 38805 30680
rect 38763 30631 38805 30640
rect 38851 30680 38909 30681
rect 38851 30640 38860 30680
rect 38900 30640 38909 30680
rect 38851 30639 38909 30640
rect 39051 30680 39093 30689
rect 39051 30640 39052 30680
rect 39092 30640 39093 30680
rect 39051 30631 39093 30640
rect 39147 30680 39189 30689
rect 39147 30640 39148 30680
rect 39188 30640 39189 30680
rect 39147 30631 39189 30640
rect 39243 30680 39285 30689
rect 39243 30640 39244 30680
rect 39284 30640 39285 30680
rect 39243 30631 39285 30640
rect 39339 30680 39381 30689
rect 39339 30640 39340 30680
rect 39380 30640 39381 30680
rect 39339 30631 39381 30640
rect 39523 30680 39581 30681
rect 39523 30640 39532 30680
rect 39572 30640 39581 30680
rect 39523 30639 39581 30640
rect 40483 30680 40541 30681
rect 40483 30640 40492 30680
rect 40532 30640 40541 30680
rect 40483 30639 40541 30640
rect 41643 30680 41685 30689
rect 41643 30640 41644 30680
rect 41684 30640 41685 30680
rect 41643 30631 41685 30640
rect 41739 30680 41781 30689
rect 41739 30640 41740 30680
rect 41780 30640 41781 30680
rect 41739 30631 41781 30640
rect 41835 30680 41877 30689
rect 41835 30640 41836 30680
rect 41876 30640 41877 30680
rect 41835 30631 41877 30640
rect 41931 30680 41973 30689
rect 41931 30640 41932 30680
rect 41972 30640 41973 30680
rect 41931 30631 41973 30640
rect 42595 30680 42653 30681
rect 42595 30640 42604 30680
rect 42644 30640 42653 30680
rect 42595 30639 42653 30640
rect 43459 30680 43517 30681
rect 43459 30640 43468 30680
rect 43508 30640 43517 30680
rect 43459 30639 43517 30640
rect 44811 30680 44853 30689
rect 44811 30640 44812 30680
rect 44852 30640 44853 30680
rect 44811 30631 44853 30640
rect 45003 30680 45045 30689
rect 45003 30640 45004 30680
rect 45044 30640 45045 30680
rect 45003 30631 45045 30640
rect 45091 30680 45149 30681
rect 45091 30640 45100 30680
rect 45140 30640 45149 30680
rect 45091 30639 45149 30640
rect 46531 30680 46589 30681
rect 46531 30640 46540 30680
rect 46580 30640 46589 30680
rect 46531 30639 46589 30640
rect 46819 30680 46877 30681
rect 46819 30640 46828 30680
rect 46868 30640 46877 30680
rect 46819 30639 46877 30640
rect 47011 30680 47069 30681
rect 47011 30640 47020 30680
rect 47060 30640 47069 30680
rect 47011 30639 47069 30640
rect 47115 30680 47157 30689
rect 47115 30640 47116 30680
rect 47156 30640 47157 30680
rect 47115 30631 47157 30640
rect 47307 30680 47349 30689
rect 47307 30640 47308 30680
rect 47348 30640 47349 30680
rect 47307 30631 47349 30640
rect 47691 30680 47733 30689
rect 47691 30640 47692 30680
rect 47732 30640 47733 30680
rect 47691 30631 47733 30640
rect 47787 30680 47829 30689
rect 47787 30640 47788 30680
rect 47828 30640 47829 30680
rect 47787 30631 47829 30640
rect 47883 30680 47925 30689
rect 47883 30640 47884 30680
rect 47924 30640 47925 30680
rect 47883 30631 47925 30640
rect 47979 30680 48021 30689
rect 47979 30640 47980 30680
rect 48020 30640 48021 30680
rect 47979 30631 48021 30640
rect 48267 30680 48309 30689
rect 48267 30640 48268 30680
rect 48308 30640 48309 30680
rect 48267 30631 48309 30640
rect 48459 30680 48501 30689
rect 48459 30640 48460 30680
rect 48500 30640 48501 30680
rect 48459 30631 48501 30640
rect 48547 30680 48605 30681
rect 48547 30640 48556 30680
rect 48596 30640 48605 30680
rect 48547 30639 48605 30640
rect 48931 30680 48989 30681
rect 48931 30640 48940 30680
rect 48980 30640 48989 30680
rect 48931 30639 48989 30640
rect 8427 30617 8469 30626
rect 3723 30596 3765 30605
rect 3723 30556 3724 30596
rect 3764 30556 3765 30596
rect 3723 30547 3765 30556
rect 7467 30596 7509 30605
rect 7467 30556 7468 30596
rect 7508 30556 7509 30596
rect 7467 30547 7509 30556
rect 16291 30596 16349 30597
rect 16291 30556 16300 30596
rect 16340 30556 16349 30596
rect 16291 30555 16349 30556
rect 31939 30596 31997 30597
rect 31939 30556 31948 30596
rect 31988 30556 31997 30596
rect 31939 30555 31997 30556
rect 35979 30596 36021 30605
rect 35979 30556 35980 30596
rect 36020 30556 36021 30596
rect 35979 30547 36021 30556
rect 9867 30512 9909 30521
rect 9867 30472 9868 30512
rect 9908 30472 9909 30512
rect 9867 30463 9909 30472
rect 13803 30512 13845 30521
rect 13803 30472 13804 30512
rect 13844 30472 13845 30512
rect 13803 30463 13845 30472
rect 17451 30512 17493 30521
rect 17451 30472 17452 30512
rect 17492 30472 17493 30512
rect 17451 30463 17493 30472
rect 45291 30512 45333 30521
rect 45291 30472 45292 30512
rect 45332 30472 45333 30512
rect 45291 30463 45333 30472
rect 48267 30512 48309 30521
rect 48267 30472 48268 30512
rect 48308 30472 48309 30512
rect 48267 30463 48309 30472
rect 49995 30512 50037 30521
rect 49995 30472 49996 30512
rect 50036 30472 50037 30512
rect 49995 30463 50037 30472
rect 50187 30512 50229 30521
rect 50187 30472 50188 30512
rect 50228 30472 50229 30512
rect 50187 30463 50229 30472
rect 4003 30428 4061 30429
rect 4003 30388 4012 30428
rect 4052 30388 4061 30428
rect 4003 30387 4061 30388
rect 5923 30428 5981 30429
rect 5923 30388 5932 30428
rect 5972 30388 5981 30428
rect 5923 30387 5981 30388
rect 8995 30428 9053 30429
rect 8995 30388 9004 30428
rect 9044 30388 9053 30428
rect 8995 30387 9053 30388
rect 11395 30428 11453 30429
rect 11395 30388 11404 30428
rect 11444 30388 11453 30428
rect 11395 30387 11453 30388
rect 13227 30428 13269 30437
rect 13227 30388 13228 30428
rect 13268 30388 13269 30428
rect 13227 30379 13269 30388
rect 14659 30428 14717 30429
rect 14659 30388 14668 30428
rect 14708 30388 14717 30428
rect 14659 30387 14717 30388
rect 16107 30428 16149 30437
rect 16107 30388 16108 30428
rect 16148 30388 16149 30428
rect 16107 30379 16149 30388
rect 18987 30428 19029 30437
rect 18987 30388 18988 30428
rect 19028 30388 19029 30428
rect 18987 30379 19029 30388
rect 22347 30428 22389 30437
rect 22347 30388 22348 30428
rect 22388 30388 22389 30428
rect 22347 30379 22389 30388
rect 28003 30428 28061 30429
rect 28003 30388 28012 30428
rect 28052 30388 28061 30428
rect 28003 30387 28061 30388
rect 29059 30428 29117 30429
rect 29059 30388 29068 30428
rect 29108 30388 29117 30428
rect 29059 30387 29117 30388
rect 29923 30428 29981 30429
rect 29923 30388 29932 30428
rect 29972 30388 29981 30428
rect 29923 30387 29981 30388
rect 32715 30428 32757 30437
rect 32715 30388 32716 30428
rect 32756 30388 32757 30428
rect 32715 30379 32757 30388
rect 33571 30428 33629 30429
rect 33571 30388 33580 30428
rect 33620 30388 33629 30428
rect 33571 30387 33629 30388
rect 34435 30428 34493 30429
rect 34435 30388 34444 30428
rect 34484 30388 34493 30428
rect 34435 30387 34493 30388
rect 37131 30428 37173 30437
rect 37131 30388 37132 30428
rect 37172 30388 37173 30428
rect 37131 30379 37173 30388
rect 38379 30428 38421 30437
rect 38379 30388 38380 30428
rect 38420 30388 38421 30428
rect 38379 30379 38421 30388
rect 40195 30428 40253 30429
rect 40195 30388 40204 30428
rect 40244 30388 40253 30428
rect 40195 30387 40253 30388
rect 44811 30428 44853 30437
rect 44811 30388 44812 30428
rect 44852 30388 44853 30428
rect 44811 30379 44853 30388
rect 46443 30428 46485 30437
rect 46443 30388 46444 30428
rect 46484 30388 46485 30428
rect 46443 30379 46485 30388
rect 46731 30428 46773 30437
rect 46731 30388 46732 30428
rect 46772 30388 46773 30428
rect 46731 30379 46773 30388
rect 49603 30428 49661 30429
rect 49603 30388 49612 30428
rect 49652 30388 49661 30428
rect 49603 30387 49661 30388
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 8035 30092 8093 30093
rect 8035 30052 8044 30092
rect 8084 30052 8093 30092
rect 8035 30051 8093 30052
rect 11595 30092 11637 30101
rect 11595 30052 11596 30092
rect 11636 30052 11637 30092
rect 11595 30043 11637 30052
rect 23307 30092 23349 30101
rect 23307 30052 23308 30092
rect 23348 30052 23349 30092
rect 23307 30043 23349 30052
rect 24163 30092 24221 30093
rect 24163 30052 24172 30092
rect 24212 30052 24221 30092
rect 24163 30051 24221 30052
rect 31267 30092 31325 30093
rect 31267 30052 31276 30092
rect 31316 30052 31325 30092
rect 31267 30051 31325 30052
rect 35587 30092 35645 30093
rect 35587 30052 35596 30092
rect 35636 30052 35645 30092
rect 35587 30051 35645 30052
rect 36267 30092 36309 30101
rect 36267 30052 36268 30092
rect 36308 30052 36309 30092
rect 36267 30043 36309 30052
rect 1035 30008 1077 30017
rect 1035 29968 1036 30008
rect 1076 29968 1077 30008
rect 1035 29959 1077 29968
rect 12835 30008 12893 30009
rect 12835 29968 12844 30008
rect 12884 29968 12893 30008
rect 12835 29967 12893 29968
rect 13795 30008 13853 30009
rect 13795 29968 13804 30008
rect 13844 29968 13853 30008
rect 13795 29967 13853 29968
rect 19467 30008 19509 30017
rect 19467 29968 19468 30008
rect 19508 29968 19509 30008
rect 19467 29959 19509 29968
rect 22347 30008 22389 30017
rect 22347 29968 22348 30008
rect 22388 29968 22389 30008
rect 22347 29959 22389 29968
rect 26947 30008 27005 30009
rect 26947 29968 26956 30008
rect 26996 29968 27005 30008
rect 26947 29967 27005 29968
rect 38755 30008 38813 30009
rect 38755 29968 38764 30008
rect 38804 29968 38813 30008
rect 38755 29967 38813 29968
rect 42307 30008 42365 30009
rect 42307 29968 42316 30008
rect 42356 29968 42365 30008
rect 42307 29967 42365 29968
rect 46915 30008 46973 30009
rect 46915 29968 46924 30008
rect 46964 29968 46973 30008
rect 46915 29967 46973 29968
rect 3627 29924 3669 29933
rect 3627 29884 3628 29924
rect 3668 29884 3669 29924
rect 3627 29875 3669 29884
rect 5067 29924 5109 29933
rect 5067 29884 5068 29924
rect 5108 29884 5109 29924
rect 5067 29875 5109 29884
rect 11307 29924 11349 29933
rect 11307 29884 11308 29924
rect 11348 29884 11349 29924
rect 11307 29875 11349 29884
rect 17355 29924 17397 29933
rect 17355 29884 17356 29924
rect 17396 29884 17397 29924
rect 17355 29875 17397 29884
rect 42123 29924 42165 29933
rect 42123 29884 42124 29924
rect 42164 29884 42165 29924
rect 42123 29875 42165 29884
rect 6123 29854 6165 29863
rect 1227 29840 1269 29849
rect 1227 29800 1228 29840
rect 1268 29800 1269 29840
rect 1227 29791 1269 29800
rect 1603 29840 1661 29841
rect 1603 29800 1612 29840
rect 1652 29800 1661 29840
rect 1603 29799 1661 29800
rect 2467 29840 2525 29841
rect 2467 29800 2476 29840
rect 2516 29800 2525 29840
rect 2467 29799 2525 29800
rect 4107 29840 4149 29849
rect 4107 29800 4108 29840
rect 4148 29800 4149 29840
rect 4107 29791 4149 29800
rect 4203 29840 4245 29849
rect 4203 29800 4204 29840
rect 4244 29800 4245 29840
rect 4203 29791 4245 29800
rect 4299 29840 4341 29849
rect 4299 29800 4300 29840
rect 4340 29800 4341 29840
rect 4299 29791 4341 29800
rect 4587 29840 4629 29849
rect 4587 29800 4588 29840
rect 4628 29800 4629 29840
rect 4587 29791 4629 29800
rect 4683 29840 4725 29849
rect 4683 29800 4684 29840
rect 4724 29800 4725 29840
rect 4683 29791 4725 29800
rect 5163 29840 5205 29849
rect 5163 29800 5164 29840
rect 5204 29800 5205 29840
rect 5163 29791 5205 29800
rect 5635 29840 5693 29841
rect 5635 29800 5644 29840
rect 5684 29800 5693 29840
rect 6123 29814 6124 29854
rect 6164 29814 6165 29854
rect 6123 29805 6165 29814
rect 6499 29840 6557 29841
rect 5635 29799 5693 29800
rect 6499 29800 6508 29840
rect 6548 29800 6557 29840
rect 6499 29799 6557 29800
rect 7563 29840 7605 29849
rect 7563 29800 7564 29840
rect 7604 29800 7605 29840
rect 7563 29791 7605 29800
rect 7659 29840 7701 29849
rect 7659 29800 7660 29840
rect 7700 29800 7701 29840
rect 7659 29791 7701 29800
rect 7755 29840 7797 29849
rect 7755 29800 7756 29840
rect 7796 29800 7797 29840
rect 7755 29791 7797 29800
rect 7851 29840 7893 29849
rect 7851 29800 7852 29840
rect 7892 29800 7893 29840
rect 7851 29791 7893 29800
rect 8707 29840 8765 29841
rect 8707 29800 8716 29840
rect 8756 29800 8765 29840
rect 8707 29799 8765 29800
rect 8907 29840 8949 29849
rect 8907 29800 8908 29840
rect 8948 29800 8949 29840
rect 8907 29791 8949 29800
rect 9283 29840 9341 29841
rect 9283 29800 9292 29840
rect 9332 29800 9341 29840
rect 9283 29799 9341 29800
rect 10147 29840 10205 29841
rect 10147 29800 10156 29840
rect 10196 29800 10205 29840
rect 10147 29799 10205 29800
rect 11595 29840 11637 29849
rect 11595 29800 11596 29840
rect 11636 29800 11637 29840
rect 11595 29791 11637 29800
rect 11787 29840 11829 29849
rect 11787 29800 11788 29840
rect 11828 29800 11829 29840
rect 11787 29791 11829 29800
rect 11875 29840 11933 29841
rect 11875 29800 11884 29840
rect 11924 29800 11933 29840
rect 11875 29799 11933 29800
rect 12163 29840 12221 29841
rect 12163 29800 12172 29840
rect 12212 29800 12221 29840
rect 12163 29799 12221 29800
rect 12459 29840 12501 29849
rect 12459 29800 12460 29840
rect 12500 29800 12501 29840
rect 12459 29791 12501 29800
rect 12555 29840 12597 29849
rect 12555 29800 12556 29840
rect 12596 29800 12597 29840
rect 12555 29791 12597 29800
rect 13123 29840 13181 29841
rect 13123 29800 13132 29840
rect 13172 29800 13181 29840
rect 13123 29799 13181 29800
rect 13419 29840 13461 29849
rect 13419 29800 13420 29840
rect 13460 29800 13461 29840
rect 13419 29791 13461 29800
rect 13515 29840 13557 29849
rect 13515 29800 13516 29840
rect 13556 29800 13557 29840
rect 13515 29791 13557 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 14179 29840 14237 29841
rect 14179 29800 14188 29840
rect 14228 29800 14237 29840
rect 14179 29799 14237 29800
rect 14475 29840 14517 29849
rect 14475 29800 14476 29840
rect 14516 29800 14517 29840
rect 14475 29791 14517 29800
rect 14571 29840 14613 29849
rect 14571 29800 14572 29840
rect 14612 29800 14613 29840
rect 14571 29791 14613 29800
rect 14667 29840 14709 29849
rect 14667 29800 14668 29840
rect 14708 29800 14709 29840
rect 14667 29791 14709 29800
rect 14763 29840 14805 29849
rect 14763 29800 14764 29840
rect 14804 29800 14805 29840
rect 14763 29791 14805 29800
rect 14955 29840 14997 29849
rect 14955 29800 14956 29840
rect 14996 29800 14997 29840
rect 14955 29791 14997 29800
rect 15331 29840 15389 29841
rect 15331 29800 15340 29840
rect 15380 29800 15389 29840
rect 15331 29799 15389 29800
rect 16195 29840 16253 29841
rect 16195 29800 16204 29840
rect 16244 29800 16253 29840
rect 16195 29799 16253 29800
rect 18603 29840 18645 29849
rect 18603 29800 18604 29840
rect 18644 29800 18645 29840
rect 18603 29791 18645 29800
rect 18699 29840 18741 29849
rect 18699 29800 18700 29840
rect 18740 29800 18741 29840
rect 18699 29791 18741 29800
rect 18795 29840 18837 29849
rect 18795 29800 18796 29840
rect 18836 29800 18837 29840
rect 18795 29791 18837 29800
rect 18891 29840 18933 29849
rect 18891 29800 18892 29840
rect 18932 29800 18933 29840
rect 18891 29791 18933 29800
rect 19171 29840 19229 29841
rect 19171 29800 19180 29840
rect 19220 29800 19229 29840
rect 19171 29799 19229 29800
rect 20131 29840 20189 29841
rect 20131 29800 20140 29840
rect 20180 29800 20189 29840
rect 20131 29799 20189 29800
rect 20419 29840 20477 29841
rect 20419 29800 20428 29840
rect 20468 29800 20477 29840
rect 20419 29799 20477 29800
rect 21955 29840 22013 29841
rect 21955 29800 21964 29840
rect 22004 29800 22013 29840
rect 21955 29799 22013 29800
rect 23011 29840 23069 29841
rect 23011 29800 23020 29840
rect 23060 29800 23069 29840
rect 23011 29799 23069 29800
rect 25315 29840 25373 29841
rect 25315 29800 25324 29840
rect 25364 29800 25373 29840
rect 25315 29799 25373 29800
rect 26179 29840 26237 29841
rect 26179 29800 26188 29840
rect 26228 29800 26237 29840
rect 26179 29799 26237 29800
rect 27339 29840 27381 29849
rect 27339 29800 27340 29840
rect 27380 29800 27381 29840
rect 27339 29791 27381 29800
rect 27619 29840 27677 29841
rect 27619 29800 27628 29840
rect 27668 29800 27677 29840
rect 27619 29799 27677 29800
rect 28579 29840 28637 29841
rect 28579 29800 28588 29840
rect 28628 29800 28637 29840
rect 28579 29799 28637 29800
rect 28875 29840 28917 29849
rect 28875 29800 28876 29840
rect 28916 29800 28917 29840
rect 28875 29791 28917 29800
rect 29251 29840 29309 29841
rect 29251 29800 29260 29840
rect 29300 29800 29309 29840
rect 29251 29799 29309 29800
rect 30115 29840 30173 29841
rect 30115 29800 30124 29840
rect 30164 29800 30173 29840
rect 30115 29799 30173 29800
rect 31467 29840 31509 29849
rect 31467 29800 31468 29840
rect 31508 29800 31509 29840
rect 31467 29791 31509 29800
rect 31659 29840 31701 29849
rect 31659 29800 31660 29840
rect 31700 29800 31701 29840
rect 31659 29791 31701 29800
rect 31747 29840 31805 29841
rect 31747 29800 31756 29840
rect 31796 29800 31805 29840
rect 31747 29799 31805 29800
rect 31939 29840 31997 29841
rect 31939 29800 31948 29840
rect 31988 29800 31997 29840
rect 31939 29799 31997 29800
rect 32899 29840 32957 29841
rect 32899 29800 32908 29840
rect 32948 29800 32957 29840
rect 32899 29799 32957 29800
rect 33195 29840 33237 29849
rect 33195 29800 33196 29840
rect 33236 29800 33237 29840
rect 33195 29791 33237 29800
rect 33571 29840 33629 29841
rect 33571 29800 33580 29840
rect 33620 29800 33629 29840
rect 33571 29799 33629 29800
rect 34435 29840 34493 29841
rect 34435 29800 34444 29840
rect 34484 29800 34493 29840
rect 34435 29799 34493 29800
rect 35971 29840 36029 29841
rect 35971 29800 35980 29840
rect 36020 29800 36029 29840
rect 35971 29799 36029 29800
rect 36075 29840 36117 29849
rect 36075 29800 36076 29840
rect 36116 29800 36117 29840
rect 36075 29791 36117 29800
rect 36267 29840 36309 29849
rect 36267 29800 36268 29840
rect 36308 29800 36309 29840
rect 36267 29791 36309 29800
rect 37123 29840 37181 29841
rect 37123 29800 37132 29840
rect 37172 29800 37181 29840
rect 37123 29799 37181 29800
rect 37419 29840 37461 29849
rect 37419 29800 37420 29840
rect 37460 29800 37461 29840
rect 37419 29791 37461 29800
rect 37515 29840 37557 29849
rect 37515 29800 37516 29840
rect 37556 29800 37557 29840
rect 37515 29791 37557 29800
rect 37611 29840 37653 29849
rect 37611 29800 37612 29840
rect 37652 29800 37653 29840
rect 37611 29791 37653 29800
rect 38283 29840 38325 29849
rect 38283 29800 38284 29840
rect 38324 29800 38325 29840
rect 38283 29791 38325 29800
rect 38379 29840 38421 29849
rect 38379 29800 38380 29840
rect 38420 29800 38421 29840
rect 38379 29791 38421 29800
rect 38475 29840 38517 29849
rect 38475 29800 38476 29840
rect 38516 29800 38517 29840
rect 38475 29791 38517 29800
rect 38571 29840 38613 29849
rect 38571 29800 38572 29840
rect 38612 29800 38613 29840
rect 38571 29791 38613 29800
rect 39051 29840 39093 29849
rect 39051 29800 39052 29840
rect 39092 29800 39093 29840
rect 39051 29791 39093 29800
rect 39147 29840 39189 29849
rect 39147 29800 39148 29840
rect 39188 29800 39189 29840
rect 39147 29791 39189 29800
rect 39427 29840 39485 29841
rect 39427 29800 39436 29840
rect 39476 29800 39485 29840
rect 39427 29799 39485 29800
rect 39723 29840 39765 29849
rect 39723 29800 39724 29840
rect 39764 29800 39765 29840
rect 39723 29791 39765 29800
rect 40099 29840 40157 29841
rect 40099 29800 40108 29840
rect 40148 29800 40157 29840
rect 40099 29799 40157 29800
rect 40963 29840 41021 29841
rect 40963 29800 40972 29840
rect 41012 29800 41021 29840
rect 40963 29799 41021 29800
rect 42979 29840 43037 29841
rect 42979 29800 42988 29840
rect 43028 29800 43037 29840
rect 42979 29799 43037 29800
rect 43179 29840 43221 29849
rect 43179 29800 43180 29840
rect 43220 29800 43221 29840
rect 43179 29791 43221 29800
rect 43275 29840 43317 29849
rect 43275 29800 43276 29840
rect 43316 29800 43317 29840
rect 43275 29791 43317 29800
rect 43371 29840 43413 29849
rect 43371 29800 43372 29840
rect 43412 29800 43413 29840
rect 43371 29791 43413 29800
rect 43651 29840 43709 29841
rect 43651 29800 43660 29840
rect 43700 29800 43709 29840
rect 43651 29799 43709 29800
rect 44899 29840 44957 29841
rect 44899 29800 44908 29840
rect 44948 29800 44957 29840
rect 44899 29799 44957 29800
rect 45763 29840 45821 29841
rect 45763 29800 45772 29840
rect 45812 29800 45821 29840
rect 45763 29799 45821 29800
rect 47779 29840 47837 29841
rect 47779 29800 47788 29840
rect 47828 29800 47837 29840
rect 47779 29799 47837 29800
rect 48547 29840 48605 29841
rect 48547 29800 48556 29840
rect 48596 29800 48605 29840
rect 48547 29799 48605 29800
rect 49411 29840 49469 29841
rect 49411 29800 49420 29840
rect 49460 29800 49469 29840
rect 49411 29799 49469 29800
rect 14091 29756 14133 29765
rect 14091 29716 14092 29756
rect 14132 29716 14133 29756
rect 14091 29707 14133 29716
rect 26571 29756 26613 29765
rect 26571 29716 26572 29756
rect 26612 29716 26613 29756
rect 26571 29707 26613 29716
rect 27243 29756 27285 29765
rect 27243 29716 27244 29756
rect 27284 29716 27285 29756
rect 27243 29707 27285 29716
rect 27915 29756 27957 29765
rect 27915 29716 27916 29756
rect 27956 29716 27957 29756
rect 27915 29707 27957 29716
rect 44331 29756 44373 29765
rect 44331 29716 44332 29756
rect 44372 29716 44373 29756
rect 44331 29707 44373 29716
rect 44523 29756 44565 29765
rect 44523 29716 44524 29756
rect 44564 29716 44565 29756
rect 44523 29707 44565 29716
rect 48171 29756 48213 29765
rect 48171 29716 48172 29756
rect 48212 29716 48213 29756
rect 48171 29707 48213 29716
rect 4003 29672 4061 29673
rect 4003 29632 4012 29672
rect 4052 29632 4061 29672
rect 4003 29631 4061 29632
rect 6315 29672 6357 29681
rect 6315 29632 6316 29672
rect 6356 29632 6357 29672
rect 6315 29623 6357 29632
rect 7171 29672 7229 29673
rect 7171 29632 7180 29672
rect 7220 29632 7229 29672
rect 7171 29631 7229 29632
rect 21091 29672 21149 29673
rect 21091 29632 21100 29672
rect 21140 29632 21149 29672
rect 21091 29631 21149 29632
rect 21283 29672 21341 29673
rect 21283 29632 21292 29672
rect 21332 29632 21341 29672
rect 21283 29631 21341 29632
rect 23499 29672 23541 29681
rect 23499 29632 23500 29672
rect 23540 29632 23541 29672
rect 23499 29623 23541 29632
rect 31555 29672 31613 29673
rect 31555 29632 31564 29672
rect 31604 29632 31613 29672
rect 31555 29631 31613 29632
rect 36451 29672 36509 29673
rect 36451 29632 36460 29672
rect 36500 29632 36509 29672
rect 36451 29631 36509 29632
rect 37699 29672 37757 29673
rect 37699 29632 37708 29672
rect 37748 29632 37757 29672
rect 37699 29631 37757 29632
rect 43459 29672 43517 29673
rect 43459 29632 43468 29672
rect 43508 29632 43517 29672
rect 43459 29631 43517 29632
rect 47107 29672 47165 29673
rect 47107 29632 47116 29672
rect 47156 29632 47165 29672
rect 47107 29631 47165 29632
rect 50563 29672 50621 29673
rect 50563 29632 50572 29672
rect 50612 29632 50621 29672
rect 50563 29631 50621 29632
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 5539 29336 5597 29337
rect 5539 29296 5548 29336
rect 5588 29296 5597 29336
rect 5539 29295 5597 29296
rect 6019 29336 6077 29337
rect 6019 29296 6028 29336
rect 6068 29296 6077 29336
rect 6019 29295 6077 29296
rect 13315 29336 13373 29337
rect 13315 29296 13324 29336
rect 13364 29296 13373 29336
rect 13315 29295 13373 29296
rect 20515 29336 20573 29337
rect 20515 29296 20524 29336
rect 20564 29296 20573 29336
rect 20515 29295 20573 29296
rect 33195 29336 33237 29345
rect 33195 29296 33196 29336
rect 33236 29296 33237 29336
rect 33195 29287 33237 29296
rect 33571 29336 33629 29337
rect 33571 29296 33580 29336
rect 33620 29296 33629 29336
rect 33571 29295 33629 29296
rect 41259 29336 41301 29345
rect 41259 29296 41260 29336
rect 41300 29296 41301 29336
rect 41259 29287 41301 29296
rect 42507 29336 42549 29345
rect 42507 29296 42508 29336
rect 42548 29296 42549 29336
rect 42507 29287 42549 29296
rect 45099 29336 45141 29345
rect 45099 29296 45100 29336
rect 45140 29296 45141 29336
rect 45099 29287 45141 29296
rect 47595 29336 47637 29345
rect 47595 29296 47596 29336
rect 47636 29296 47637 29336
rect 47595 29287 47637 29296
rect 49219 29336 49277 29337
rect 49219 29296 49228 29336
rect 49268 29296 49277 29336
rect 49219 29295 49277 29296
rect 3243 29252 3285 29261
rect 2763 29210 2805 29219
rect 2763 29170 2764 29210
rect 2804 29170 2805 29210
rect 3243 29212 3244 29252
rect 3284 29212 3285 29252
rect 3243 29203 3285 29212
rect 5259 29252 5301 29261
rect 5259 29212 5260 29252
rect 5300 29212 5301 29252
rect 5259 29203 5301 29212
rect 8427 29252 8469 29261
rect 8427 29212 8428 29252
rect 8468 29212 8469 29252
rect 8427 29203 8469 29212
rect 10923 29252 10965 29261
rect 10923 29212 10924 29252
rect 10964 29212 10965 29252
rect 10923 29203 10965 29212
rect 14379 29252 14421 29261
rect 14379 29212 14380 29252
rect 14420 29212 14421 29252
rect 14379 29203 14421 29212
rect 22923 29252 22965 29261
rect 22923 29212 22924 29252
rect 22964 29212 22965 29252
rect 35979 29252 36021 29261
rect 22923 29203 22965 29212
rect 27915 29210 27957 29219
rect 2763 29161 2805 29170
rect 2955 29168 2997 29177
rect 2955 29128 2956 29168
rect 2996 29128 2997 29168
rect 2955 29119 2997 29128
rect 3043 29168 3101 29169
rect 3043 29128 3052 29168
rect 3092 29128 3101 29168
rect 3043 29127 3101 29128
rect 3339 29168 3381 29177
rect 3339 29128 3340 29168
rect 3380 29128 3381 29168
rect 3339 29119 3381 29128
rect 3435 29168 3477 29177
rect 3435 29128 3436 29168
rect 3476 29128 3477 29168
rect 3435 29119 3477 29128
rect 3531 29168 3573 29177
rect 3531 29128 3532 29168
rect 3572 29128 3573 29168
rect 3531 29119 3573 29128
rect 3715 29168 3773 29169
rect 3715 29128 3724 29168
rect 3764 29128 3773 29168
rect 3715 29127 3773 29128
rect 4675 29168 4733 29169
rect 4675 29128 4684 29168
rect 4724 29128 4733 29168
rect 4675 29127 4733 29128
rect 5059 29168 5117 29169
rect 5059 29128 5068 29168
rect 5108 29128 5117 29168
rect 5059 29127 5117 29128
rect 5163 29168 5205 29177
rect 5163 29128 5164 29168
rect 5204 29128 5205 29168
rect 5163 29119 5205 29128
rect 5355 29168 5397 29177
rect 5355 29128 5356 29168
rect 5396 29128 5397 29168
rect 5355 29119 5397 29128
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 5739 29168 5781 29177
rect 5739 29128 5740 29168
rect 5780 29128 5781 29168
rect 5739 29119 5781 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 7171 29168 7229 29169
rect 7171 29128 7180 29168
rect 7220 29128 7229 29168
rect 7171 29127 7229 29128
rect 8035 29168 8093 29169
rect 8035 29128 8044 29168
rect 8084 29128 8093 29168
rect 8035 29127 8093 29128
rect 8707 29168 8765 29169
rect 8707 29128 8716 29168
rect 8756 29128 8765 29168
rect 8707 29127 8765 29128
rect 9099 29168 9141 29177
rect 9099 29128 9100 29168
rect 9140 29128 9141 29168
rect 9099 29119 9141 29128
rect 9955 29168 10013 29169
rect 9955 29128 9964 29168
rect 10004 29128 10013 29168
rect 9955 29127 10013 29128
rect 11299 29168 11357 29169
rect 11299 29128 11308 29168
rect 11348 29128 11357 29168
rect 11299 29127 11357 29128
rect 12163 29168 12221 29169
rect 12163 29128 12172 29168
rect 12212 29128 12221 29168
rect 12163 29127 12221 29128
rect 13987 29168 14045 29169
rect 13987 29128 13996 29168
rect 14036 29128 14045 29168
rect 13987 29127 14045 29128
rect 14283 29168 14325 29177
rect 14283 29128 14284 29168
rect 14324 29128 14325 29168
rect 14283 29119 14325 29128
rect 16099 29168 16157 29169
rect 16099 29128 16108 29168
rect 16148 29128 16157 29168
rect 16099 29127 16157 29128
rect 17731 29168 17789 29169
rect 17731 29128 17740 29168
rect 17780 29128 17789 29168
rect 17731 29127 17789 29128
rect 18595 29168 18653 29169
rect 18595 29128 18604 29168
rect 18644 29128 18653 29168
rect 18595 29127 18653 29128
rect 18987 29168 19029 29177
rect 18987 29128 18988 29168
rect 19028 29128 19029 29168
rect 18987 29119 19029 29128
rect 19179 29168 19221 29177
rect 19179 29128 19180 29168
rect 19220 29128 19221 29168
rect 19179 29119 19221 29128
rect 19843 29168 19901 29169
rect 19843 29128 19852 29168
rect 19892 29128 19901 29168
rect 19843 29127 19901 29128
rect 20043 29168 20085 29177
rect 20043 29128 20044 29168
rect 20084 29128 20085 29168
rect 20043 29119 20085 29128
rect 20235 29168 20277 29177
rect 20235 29128 20236 29168
rect 20276 29128 20277 29168
rect 20235 29119 20277 29128
rect 20323 29168 20381 29169
rect 20323 29128 20332 29168
rect 20372 29128 20381 29168
rect 20323 29127 20381 29128
rect 21667 29168 21725 29169
rect 21667 29128 21676 29168
rect 21716 29128 21725 29168
rect 21667 29127 21725 29128
rect 22531 29168 22589 29169
rect 22531 29128 22540 29168
rect 22580 29128 22589 29168
rect 22531 29127 22589 29128
rect 26283 29168 26325 29177
rect 26283 29128 26284 29168
rect 26324 29128 26325 29168
rect 26283 29119 26325 29128
rect 26379 29168 26421 29177
rect 26379 29128 26380 29168
rect 26420 29128 26421 29168
rect 26379 29119 26421 29128
rect 26475 29168 26517 29177
rect 26475 29128 26476 29168
rect 26516 29128 26517 29168
rect 26475 29119 26517 29128
rect 26571 29168 26613 29177
rect 26571 29128 26572 29168
rect 26612 29128 26613 29168
rect 26571 29119 26613 29128
rect 26763 29168 26805 29177
rect 26763 29128 26764 29168
rect 26804 29128 26805 29168
rect 26763 29119 26805 29128
rect 26955 29168 26997 29177
rect 26955 29128 26956 29168
rect 26996 29128 26997 29168
rect 26955 29119 26997 29128
rect 27043 29168 27101 29169
rect 27043 29128 27052 29168
rect 27092 29128 27101 29168
rect 27043 29127 27101 29128
rect 27243 29168 27285 29177
rect 27243 29128 27244 29168
rect 27284 29128 27285 29168
rect 27243 29119 27285 29128
rect 27435 29168 27477 29177
rect 27915 29170 27916 29210
rect 27956 29170 27957 29210
rect 35979 29212 35980 29252
rect 36020 29212 36021 29252
rect 35979 29203 36021 29212
rect 51627 29252 51669 29261
rect 51627 29212 51628 29252
rect 51668 29212 51669 29252
rect 51627 29203 51669 29212
rect 27435 29128 27436 29168
rect 27476 29128 27477 29168
rect 27435 29119 27477 29128
rect 27523 29168 27581 29169
rect 27523 29128 27532 29168
rect 27572 29128 27581 29168
rect 27915 29161 27957 29170
rect 28107 29168 28149 29177
rect 27523 29127 27581 29128
rect 28107 29128 28108 29168
rect 28148 29128 28149 29168
rect 28107 29119 28149 29128
rect 28195 29168 28253 29169
rect 28195 29128 28204 29168
rect 28244 29128 28253 29168
rect 28195 29127 28253 29128
rect 28395 29168 28437 29177
rect 28395 29128 28396 29168
rect 28436 29128 28437 29168
rect 28395 29119 28437 29128
rect 28483 29168 28541 29169
rect 28483 29128 28492 29168
rect 28532 29128 28541 29168
rect 28483 29127 28541 29128
rect 29067 29168 29109 29177
rect 29067 29128 29068 29168
rect 29108 29128 29109 29168
rect 29067 29119 29109 29128
rect 29259 29168 29301 29177
rect 29259 29128 29260 29168
rect 29300 29128 29301 29168
rect 29259 29119 29301 29128
rect 29347 29168 29405 29169
rect 29347 29128 29356 29168
rect 29396 29128 29405 29168
rect 29347 29127 29405 29128
rect 29835 29168 29877 29177
rect 29835 29128 29836 29168
rect 29876 29128 29877 29168
rect 29835 29119 29877 29128
rect 29923 29168 29981 29169
rect 29923 29128 29932 29168
rect 29972 29128 29981 29168
rect 29923 29127 29981 29128
rect 30115 29168 30173 29169
rect 30115 29128 30124 29168
rect 30164 29128 30173 29168
rect 30115 29127 30173 29128
rect 30219 29168 30261 29177
rect 30219 29128 30220 29168
rect 30260 29128 30261 29168
rect 30219 29119 30261 29128
rect 30411 29168 30453 29177
rect 30411 29128 30412 29168
rect 30452 29128 30453 29168
rect 30411 29119 30453 29128
rect 30603 29168 30645 29177
rect 30603 29128 30604 29168
rect 30644 29128 30645 29168
rect 30603 29119 30645 29128
rect 30699 29168 30741 29177
rect 30699 29128 30700 29168
rect 30740 29128 30741 29168
rect 30699 29119 30741 29128
rect 30795 29168 30837 29177
rect 30795 29128 30796 29168
rect 30836 29128 30837 29168
rect 30795 29119 30837 29128
rect 30891 29168 30933 29177
rect 30891 29128 30892 29168
rect 30932 29128 30933 29168
rect 30891 29119 30933 29128
rect 31075 29168 31133 29169
rect 31075 29128 31084 29168
rect 31124 29128 31133 29168
rect 31075 29127 31133 29128
rect 31947 29168 31989 29177
rect 31947 29128 31948 29168
rect 31988 29128 31989 29168
rect 31947 29119 31989 29128
rect 32611 29168 32669 29169
rect 32611 29128 32620 29168
rect 32660 29128 32669 29168
rect 32611 29127 32669 29128
rect 33283 29168 33341 29169
rect 33283 29128 33292 29168
rect 33332 29128 33341 29168
rect 33283 29127 33341 29128
rect 33483 29168 33525 29177
rect 33483 29128 33484 29168
rect 33524 29128 33525 29168
rect 33483 29119 33525 29128
rect 33675 29168 33717 29177
rect 33675 29128 33676 29168
rect 33716 29128 33717 29168
rect 33675 29119 33717 29128
rect 33763 29168 33821 29169
rect 33763 29128 33772 29168
rect 33812 29128 33821 29168
rect 33763 29127 33821 29128
rect 33955 29168 34013 29169
rect 33955 29128 33964 29168
rect 34004 29128 34013 29168
rect 33955 29127 34013 29128
rect 34827 29168 34869 29177
rect 34827 29128 34828 29168
rect 34868 29128 34869 29168
rect 34827 29119 34869 29128
rect 36355 29168 36413 29169
rect 36355 29128 36364 29168
rect 36404 29128 36413 29168
rect 36355 29127 36413 29128
rect 37219 29168 37277 29169
rect 37219 29128 37228 29168
rect 37268 29128 37277 29168
rect 37219 29127 37277 29128
rect 39811 29168 39869 29169
rect 39811 29128 39820 29168
rect 39860 29128 39869 29168
rect 39811 29127 39869 29128
rect 41643 29168 41685 29177
rect 41643 29128 41644 29168
rect 41684 29128 41685 29168
rect 41643 29119 41685 29128
rect 41827 29168 41885 29169
rect 41827 29128 41836 29168
rect 41876 29128 41885 29168
rect 41827 29127 41885 29128
rect 42891 29168 42933 29177
rect 42891 29128 42892 29168
rect 42932 29128 42933 29168
rect 42891 29119 42933 29128
rect 43267 29168 43325 29169
rect 43267 29128 43276 29168
rect 43316 29128 43325 29168
rect 43267 29127 43325 29128
rect 44139 29168 44181 29177
rect 44139 29128 44140 29168
rect 44180 29128 44181 29168
rect 44139 29119 44181 29128
rect 44611 29168 44669 29169
rect 44611 29128 44620 29168
rect 44660 29128 44669 29168
rect 44611 29127 44669 29128
rect 45859 29168 45917 29169
rect 45859 29128 45868 29168
rect 45908 29128 45917 29168
rect 45859 29127 45917 29128
rect 47107 29168 47165 29169
rect 47107 29128 47116 29168
rect 47156 29128 47165 29168
rect 47107 29127 47165 29128
rect 49027 29168 49085 29169
rect 49027 29128 49036 29168
rect 49076 29128 49085 29168
rect 49027 29127 49085 29128
rect 50371 29168 50429 29169
rect 50371 29128 50380 29168
rect 50420 29128 50429 29168
rect 50371 29127 50429 29128
rect 51235 29168 51293 29169
rect 51235 29128 51244 29168
rect 51284 29128 51293 29168
rect 51235 29127 51293 29128
rect 8619 29084 8661 29093
rect 8619 29044 8620 29084
rect 8660 29044 8661 29084
rect 8619 29035 8661 29044
rect 15435 29084 15477 29093
rect 15435 29044 15436 29084
rect 15476 29044 15477 29084
rect 15435 29035 15477 29044
rect 31755 29084 31797 29093
rect 31755 29044 31756 29084
rect 31796 29044 31797 29084
rect 31755 29035 31797 29044
rect 35779 29084 35837 29085
rect 35779 29044 35788 29084
rect 35828 29044 35837 29084
rect 35779 29043 35837 29044
rect 38955 29084 38997 29093
rect 38955 29044 38956 29084
rect 38996 29044 38997 29084
rect 38955 29035 38997 29044
rect 41443 29084 41501 29085
rect 41443 29044 41452 29084
rect 41492 29044 41501 29084
rect 41443 29043 41501 29044
rect 41739 29084 41781 29093
rect 41739 29044 41740 29084
rect 41780 29044 41781 29084
rect 41739 29035 41781 29044
rect 1803 29000 1845 29009
rect 1803 28960 1804 29000
rect 1844 28960 1845 29000
rect 1803 28951 1845 28960
rect 2763 29000 2805 29009
rect 2763 28960 2764 29000
rect 2804 28960 2805 29000
rect 2763 28951 2805 28960
rect 15243 29000 15285 29009
rect 15243 28960 15244 29000
rect 15284 28960 15285 29000
rect 15243 28951 15285 28960
rect 16587 29000 16629 29009
rect 16587 28960 16588 29000
rect 16628 28960 16629 29000
rect 16587 28951 16629 28960
rect 20043 29000 20085 29009
rect 20043 28960 20044 29000
rect 20084 28960 20085 29000
rect 20043 28951 20085 28960
rect 25419 29000 25461 29009
rect 25419 28960 25420 29000
rect 25460 28960 25461 29000
rect 25419 28951 25461 28960
rect 27243 29000 27285 29009
rect 27243 28960 27244 29000
rect 27284 28960 27285 29000
rect 27243 28951 27285 28960
rect 27915 29000 27957 29009
rect 27915 28960 27916 29000
rect 27956 28960 27957 29000
rect 27915 28951 27957 28960
rect 29067 29000 29109 29009
rect 29067 28960 29068 29000
rect 29108 28960 29109 29000
rect 29067 28951 29109 28960
rect 33003 29000 33045 29009
rect 33003 28960 33004 29000
rect 33044 28960 33045 29000
rect 33003 28951 33045 28960
rect 35403 29000 35445 29009
rect 35403 28960 35404 29000
rect 35444 28960 35445 29000
rect 35403 28951 35445 28960
rect 35595 29000 35637 29009
rect 35595 28960 35596 29000
rect 35636 28960 35637 29000
rect 35595 28951 35637 28960
rect 40875 29000 40917 29009
rect 40875 28960 40876 29000
rect 40916 28960 40917 29000
rect 40875 28951 40917 28960
rect 9291 28916 9333 28925
rect 9291 28876 9292 28916
rect 9332 28876 9333 28916
rect 9291 28867 9333 28876
rect 14659 28916 14717 28917
rect 14659 28876 14668 28916
rect 14708 28876 14717 28916
rect 14659 28875 14717 28876
rect 20515 28916 20573 28917
rect 20515 28876 20524 28916
rect 20564 28876 20573 28916
rect 20515 28875 20573 28876
rect 26763 28916 26805 28925
rect 26763 28876 26764 28916
rect 26804 28876 26805 28916
rect 26763 28867 26805 28876
rect 30411 28916 30453 28925
rect 30411 28876 30412 28916
rect 30452 28876 30453 28916
rect 30411 28867 30453 28876
rect 38371 28916 38429 28917
rect 38371 28876 38380 28916
rect 38420 28876 38429 28916
rect 38371 28875 38429 28876
rect 45771 28916 45813 28925
rect 45771 28876 45772 28916
rect 45812 28876 45813 28916
rect 45771 28867 45813 28876
rect 47787 28916 47829 28925
rect 47787 28876 47788 28916
rect 47828 28876 47829 28916
rect 47787 28867 47829 28876
rect 48355 28916 48413 28917
rect 48355 28876 48364 28916
rect 48404 28876 48413 28916
rect 48355 28875 48413 28876
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 3715 28580 3773 28581
rect 3715 28540 3724 28580
rect 3764 28540 3773 28580
rect 3715 28539 3773 28540
rect 20043 28580 20085 28589
rect 20043 28540 20044 28580
rect 20084 28540 20085 28580
rect 20043 28531 20085 28540
rect 27531 28580 27573 28589
rect 27531 28540 27532 28580
rect 27572 28540 27573 28580
rect 27531 28531 27573 28540
rect 31075 28580 31133 28581
rect 31075 28540 31084 28580
rect 31124 28540 31133 28580
rect 31075 28539 31133 28540
rect 34251 28580 34293 28589
rect 34251 28540 34252 28580
rect 34292 28540 34293 28580
rect 34251 28531 34293 28540
rect 39051 28580 39093 28589
rect 39051 28540 39052 28580
rect 39092 28540 39093 28580
rect 39051 28531 39093 28540
rect 39339 28580 39381 28589
rect 39339 28540 39340 28580
rect 39380 28540 39381 28580
rect 39339 28531 39381 28540
rect 47307 28580 47349 28589
rect 47307 28540 47308 28580
rect 47348 28540 47349 28580
rect 47307 28531 47349 28540
rect 6411 28496 6453 28505
rect 6411 28456 6412 28496
rect 6452 28456 6453 28496
rect 6411 28447 6453 28456
rect 8907 28496 8949 28505
rect 8907 28456 8908 28496
rect 8948 28456 8949 28496
rect 8907 28447 8949 28456
rect 11403 28496 11445 28505
rect 11403 28456 11404 28496
rect 11444 28456 11445 28496
rect 11403 28447 11445 28456
rect 16299 28496 16341 28505
rect 16299 28456 16300 28496
rect 16340 28456 16341 28496
rect 16299 28447 16341 28456
rect 19275 28496 19317 28505
rect 19275 28456 19276 28496
rect 19316 28456 19317 28496
rect 19275 28447 19317 28456
rect 22347 28496 22389 28505
rect 22347 28456 22348 28496
rect 22388 28456 22389 28496
rect 22347 28447 22389 28456
rect 35299 28496 35357 28497
rect 35299 28456 35308 28496
rect 35348 28456 35357 28496
rect 35299 28455 35357 28456
rect 36459 28496 36501 28505
rect 36459 28456 36460 28496
rect 36500 28456 36501 28496
rect 36459 28447 36501 28456
rect 42219 28496 42261 28505
rect 42219 28456 42220 28496
rect 42260 28456 42261 28496
rect 42219 28447 42261 28456
rect 47491 28496 47549 28497
rect 47491 28456 47500 28496
rect 47540 28456 47549 28496
rect 47491 28455 47549 28456
rect 50859 28496 50901 28505
rect 50859 28456 50860 28496
rect 50900 28456 50901 28496
rect 50859 28447 50901 28456
rect 51243 28496 51285 28505
rect 51243 28456 51244 28496
rect 51284 28456 51285 28496
rect 51243 28447 51285 28456
rect 41067 28412 41109 28421
rect 41067 28372 41068 28412
rect 41108 28372 41109 28412
rect 41067 28363 41109 28372
rect 45099 28412 45141 28421
rect 45099 28372 45100 28412
rect 45140 28372 45141 28412
rect 45099 28363 45141 28372
rect 44043 28342 44085 28351
rect 1699 28328 1757 28329
rect 1699 28288 1708 28328
rect 1748 28288 1757 28328
rect 1699 28287 1757 28288
rect 2563 28328 2621 28329
rect 2563 28288 2572 28328
rect 2612 28288 2621 28328
rect 2563 28287 2621 28288
rect 4011 28328 4053 28337
rect 4011 28288 4012 28328
rect 4052 28288 4053 28328
rect 4011 28279 4053 28288
rect 4203 28328 4245 28337
rect 4203 28288 4204 28328
rect 4244 28288 4245 28328
rect 4203 28279 4245 28288
rect 4291 28328 4349 28329
rect 4291 28288 4300 28328
rect 4340 28288 4349 28328
rect 4291 28287 4349 28288
rect 5155 28328 5213 28329
rect 5155 28288 5164 28328
rect 5204 28288 5213 28328
rect 5155 28287 5213 28288
rect 5347 28328 5405 28329
rect 5347 28288 5356 28328
rect 5396 28288 5405 28328
rect 5347 28287 5405 28288
rect 6603 28328 6645 28337
rect 6603 28288 6604 28328
rect 6644 28288 6645 28328
rect 6603 28279 6645 28288
rect 6699 28328 6741 28337
rect 6699 28288 6700 28328
rect 6740 28288 6741 28328
rect 6699 28279 6741 28288
rect 6795 28328 6837 28337
rect 6795 28288 6796 28328
rect 6836 28288 6837 28328
rect 6795 28279 6837 28288
rect 6891 28328 6933 28337
rect 6891 28288 6892 28328
rect 6932 28288 6933 28328
rect 6891 28279 6933 28288
rect 7083 28328 7125 28337
rect 7083 28288 7084 28328
rect 7124 28288 7125 28328
rect 7083 28279 7125 28288
rect 7275 28328 7317 28337
rect 7275 28288 7276 28328
rect 7316 28288 7317 28328
rect 7275 28279 7317 28288
rect 7363 28328 7421 28329
rect 7363 28288 7372 28328
rect 7412 28288 7421 28328
rect 7363 28287 7421 28288
rect 8227 28328 8285 28329
rect 8227 28288 8236 28328
rect 8276 28288 8285 28328
rect 8227 28287 8285 28288
rect 8715 28328 8757 28337
rect 8715 28288 8716 28328
rect 8756 28288 8757 28328
rect 8715 28279 8757 28288
rect 10147 28328 10205 28329
rect 10147 28288 10156 28328
rect 10196 28288 10205 28328
rect 10147 28287 10205 28288
rect 11883 28328 11925 28337
rect 11883 28288 11884 28328
rect 11924 28288 11925 28328
rect 11883 28279 11925 28288
rect 12067 28328 12125 28329
rect 12067 28288 12076 28328
rect 12116 28288 12125 28328
rect 12067 28287 12125 28288
rect 12267 28328 12309 28337
rect 12267 28288 12268 28328
rect 12308 28288 12309 28328
rect 12267 28279 12309 28288
rect 12451 28328 12509 28329
rect 12451 28288 12460 28328
rect 12500 28288 12509 28328
rect 12451 28287 12509 28288
rect 12643 28328 12701 28329
rect 12643 28288 12652 28328
rect 12692 28288 12701 28328
rect 12643 28287 12701 28288
rect 12747 28328 12789 28337
rect 12747 28288 12748 28328
rect 12788 28288 12789 28328
rect 12747 28279 12789 28288
rect 12939 28328 12981 28337
rect 12939 28288 12940 28328
rect 12980 28288 12981 28328
rect 12939 28279 12981 28288
rect 13131 28328 13173 28337
rect 13131 28288 13132 28328
rect 13172 28288 13173 28328
rect 13131 28279 13173 28288
rect 13795 28328 13853 28329
rect 13795 28288 13804 28328
rect 13844 28288 13853 28328
rect 13795 28287 13853 28288
rect 14083 28328 14141 28329
rect 14083 28288 14092 28328
rect 14132 28288 14141 28328
rect 14083 28287 14141 28288
rect 17923 28328 17981 28329
rect 17923 28288 17932 28328
rect 17972 28288 17981 28328
rect 17923 28287 17981 28288
rect 18699 28328 18741 28337
rect 18699 28288 18700 28328
rect 18740 28288 18741 28328
rect 18699 28279 18741 28288
rect 18795 28328 18837 28337
rect 18795 28288 18796 28328
rect 18836 28288 18837 28328
rect 18795 28279 18837 28288
rect 18891 28328 18933 28337
rect 18891 28288 18892 28328
rect 18932 28288 18933 28328
rect 18891 28279 18933 28288
rect 18987 28328 19029 28337
rect 18987 28288 18988 28328
rect 19028 28288 19029 28328
rect 18987 28279 19029 28288
rect 19363 28328 19421 28329
rect 19363 28288 19372 28328
rect 19412 28288 19421 28328
rect 19363 28287 19421 28288
rect 19563 28328 19605 28337
rect 19563 28288 19564 28328
rect 19604 28288 19605 28328
rect 19563 28279 19605 28288
rect 19659 28328 19701 28337
rect 19659 28288 19660 28328
rect 19700 28288 19701 28328
rect 19659 28279 19701 28288
rect 19755 28328 19797 28337
rect 19755 28288 19756 28328
rect 19796 28288 19797 28328
rect 19755 28279 19797 28288
rect 19851 28328 19893 28337
rect 19851 28288 19852 28328
rect 19892 28288 19893 28328
rect 19851 28279 19893 28288
rect 20043 28328 20085 28337
rect 20043 28288 20044 28328
rect 20084 28288 20085 28328
rect 20043 28279 20085 28288
rect 20235 28328 20277 28337
rect 20235 28288 20236 28328
rect 20276 28288 20277 28328
rect 20235 28279 20277 28288
rect 20323 28328 20381 28329
rect 20323 28288 20332 28328
rect 20372 28288 20381 28328
rect 20323 28287 20381 28288
rect 20523 28328 20565 28337
rect 20523 28288 20524 28328
rect 20564 28288 20565 28328
rect 20523 28279 20565 28288
rect 20619 28328 20661 28337
rect 20619 28288 20620 28328
rect 20660 28288 20661 28328
rect 20619 28279 20661 28288
rect 20715 28328 20757 28337
rect 20715 28288 20716 28328
rect 20756 28288 20757 28328
rect 20715 28279 20757 28288
rect 21091 28328 21149 28329
rect 21091 28288 21100 28328
rect 21140 28288 21149 28328
rect 21091 28287 21149 28288
rect 23395 28328 23453 28329
rect 23395 28288 23404 28328
rect 23444 28288 23453 28328
rect 23395 28287 23453 28288
rect 24355 28328 24413 28329
rect 24355 28288 24364 28328
rect 24404 28288 24413 28328
rect 24355 28287 24413 28288
rect 25315 28328 25373 28329
rect 25315 28288 25324 28328
rect 25364 28288 25373 28328
rect 25315 28287 25373 28288
rect 25987 28328 26045 28329
rect 25987 28288 25996 28328
rect 26036 28288 26045 28328
rect 25987 28287 26045 28288
rect 26475 28328 26517 28337
rect 26475 28288 26476 28328
rect 26516 28288 26517 28328
rect 26475 28279 26517 28288
rect 26571 28328 26613 28337
rect 26571 28288 26572 28328
rect 26612 28288 26613 28328
rect 26571 28279 26613 28288
rect 26667 28328 26709 28337
rect 26667 28288 26668 28328
rect 26708 28288 26709 28328
rect 26667 28279 26709 28288
rect 27723 28328 27765 28337
rect 27723 28288 27724 28328
rect 27764 28288 27765 28328
rect 27723 28279 27765 28288
rect 28491 28328 28533 28337
rect 28491 28288 28492 28328
rect 28532 28288 28533 28328
rect 28491 28279 28533 28288
rect 28587 28328 28629 28337
rect 28587 28288 28588 28328
rect 28628 28288 28629 28328
rect 28587 28279 28629 28288
rect 28771 28328 28829 28329
rect 28771 28288 28780 28328
rect 28820 28288 28829 28328
rect 28771 28287 28829 28288
rect 28875 28328 28917 28337
rect 28875 28288 28876 28328
rect 28916 28288 28917 28328
rect 28875 28279 28917 28288
rect 29067 28328 29109 28337
rect 29067 28288 29068 28328
rect 29108 28288 29109 28328
rect 29067 28279 29109 28288
rect 30603 28328 30645 28337
rect 30603 28288 30604 28328
rect 30644 28288 30645 28328
rect 30603 28279 30645 28288
rect 30699 28328 30741 28337
rect 30699 28288 30700 28328
rect 30740 28288 30741 28328
rect 30699 28279 30741 28288
rect 30795 28328 30837 28337
rect 30795 28288 30796 28328
rect 30836 28288 30837 28328
rect 30795 28279 30837 28288
rect 30891 28328 30933 28337
rect 30891 28288 30892 28328
rect 30932 28288 30933 28328
rect 30891 28279 30933 28288
rect 32227 28328 32285 28329
rect 32227 28288 32236 28328
rect 32276 28288 32285 28328
rect 32227 28287 32285 28288
rect 33091 28328 33149 28329
rect 33091 28288 33100 28328
rect 33140 28288 33149 28328
rect 33091 28287 33149 28288
rect 33483 28328 33525 28337
rect 33483 28288 33484 28328
rect 33524 28288 33525 28328
rect 33483 28279 33525 28288
rect 34339 28328 34397 28329
rect 34339 28288 34348 28328
rect 34388 28288 34397 28328
rect 34339 28287 34397 28288
rect 35691 28328 35733 28337
rect 35691 28288 35692 28328
rect 35732 28288 35733 28328
rect 35691 28279 35733 28288
rect 35971 28328 36029 28329
rect 35971 28288 35980 28328
rect 36020 28288 36029 28328
rect 35971 28287 36029 28288
rect 37131 28328 37173 28337
rect 37131 28288 37132 28328
rect 37172 28288 37173 28328
rect 37131 28279 37173 28288
rect 37227 28328 37269 28337
rect 37227 28288 37228 28328
rect 37268 28288 37269 28328
rect 37227 28279 37269 28288
rect 37323 28328 37365 28337
rect 37323 28288 37324 28328
rect 37364 28288 37365 28328
rect 37323 28279 37365 28288
rect 37419 28328 37461 28337
rect 40011 28333 40053 28342
rect 37419 28288 37420 28328
rect 37460 28288 37461 28328
rect 37419 28279 37461 28288
rect 38851 28328 38909 28329
rect 38851 28288 38860 28328
rect 38900 28288 38909 28328
rect 38851 28287 38909 28288
rect 39139 28328 39197 28329
rect 39139 28288 39148 28328
rect 39188 28288 39197 28328
rect 39139 28287 39197 28288
rect 39427 28328 39485 28329
rect 39427 28288 39436 28328
rect 39476 28288 39485 28328
rect 39427 28287 39485 28288
rect 40011 28293 40012 28333
rect 40052 28293 40053 28333
rect 40011 28284 40053 28293
rect 40483 28328 40541 28329
rect 40483 28288 40492 28328
rect 40532 28288 40541 28328
rect 40483 28287 40541 28288
rect 40971 28328 41013 28337
rect 40971 28288 40972 28328
rect 41012 28288 41013 28328
rect 40971 28279 41013 28288
rect 41451 28328 41493 28337
rect 41451 28288 41452 28328
rect 41492 28288 41493 28328
rect 41451 28279 41493 28288
rect 41547 28328 41589 28337
rect 41547 28288 41548 28328
rect 41588 28288 41589 28328
rect 41547 28279 41589 28288
rect 41923 28328 41981 28329
rect 41923 28288 41932 28328
rect 41972 28288 41981 28328
rect 41923 28287 41981 28288
rect 43171 28328 43229 28329
rect 43171 28288 43180 28328
rect 43220 28288 43229 28328
rect 43171 28287 43229 28288
rect 43371 28328 43413 28337
rect 43371 28288 43372 28328
rect 43412 28288 43413 28328
rect 43371 28279 43413 28288
rect 43467 28328 43509 28337
rect 43467 28288 43468 28328
rect 43508 28288 43509 28328
rect 43467 28279 43509 28288
rect 43563 28328 43605 28337
rect 43563 28288 43564 28328
rect 43604 28288 43605 28328
rect 43563 28279 43605 28288
rect 43659 28328 43701 28337
rect 43659 28288 43660 28328
rect 43700 28288 43701 28328
rect 44043 28302 44044 28342
rect 44084 28302 44085 28342
rect 44043 28293 44085 28302
rect 44515 28328 44573 28329
rect 43659 28279 43701 28288
rect 44515 28288 44524 28328
rect 44564 28288 44573 28328
rect 44515 28287 44573 28288
rect 45003 28328 45045 28337
rect 45003 28288 45004 28328
rect 45044 28288 45045 28328
rect 45003 28279 45045 28288
rect 45483 28328 45525 28337
rect 45483 28288 45484 28328
rect 45524 28288 45525 28328
rect 45483 28279 45525 28288
rect 45579 28328 45621 28337
rect 45579 28288 45580 28328
rect 45620 28288 45621 28328
rect 45579 28279 45621 28288
rect 46435 28328 46493 28329
rect 46435 28288 46444 28328
rect 46484 28288 46493 28328
rect 46435 28287 46493 28288
rect 46539 28328 46581 28337
rect 46539 28288 46540 28328
rect 46580 28288 46581 28328
rect 46539 28279 46581 28288
rect 46819 28328 46877 28329
rect 46819 28288 46828 28328
rect 46868 28288 46877 28328
rect 46819 28287 46877 28288
rect 47011 28328 47069 28329
rect 47011 28288 47020 28328
rect 47060 28288 47069 28328
rect 47011 28287 47069 28288
rect 47115 28328 47157 28337
rect 47115 28288 47116 28328
rect 47156 28288 47157 28328
rect 47115 28279 47157 28288
rect 47307 28328 47349 28337
rect 47307 28288 47308 28328
rect 47348 28288 47349 28328
rect 47307 28279 47349 28288
rect 48163 28328 48221 28329
rect 48163 28288 48172 28328
rect 48212 28288 48221 28328
rect 48163 28287 48221 28288
rect 48363 28328 48405 28337
rect 48363 28288 48364 28328
rect 48404 28288 48405 28328
rect 48363 28279 48405 28288
rect 48451 28328 48509 28329
rect 48451 28288 48460 28328
rect 48500 28288 48509 28328
rect 48451 28287 48509 28288
rect 48747 28328 48789 28337
rect 48747 28288 48748 28328
rect 48788 28288 48789 28328
rect 48747 28279 48789 28288
rect 48843 28328 48885 28337
rect 48843 28288 48844 28328
rect 48884 28288 48885 28328
rect 48843 28279 48885 28288
rect 48939 28328 48981 28337
rect 48939 28288 48940 28328
rect 48980 28288 48981 28328
rect 48939 28279 48981 28288
rect 49123 28328 49181 28329
rect 49123 28288 49132 28328
rect 49172 28288 49181 28328
rect 49123 28287 49181 28288
rect 50659 28328 50717 28329
rect 50659 28288 50668 28328
rect 50708 28288 50717 28328
rect 50659 28287 50717 28288
rect 1323 28244 1365 28253
rect 1323 28204 1324 28244
rect 1364 28204 1365 28244
rect 1323 28195 1365 28204
rect 4107 28244 4149 28253
rect 4107 28204 4108 28244
rect 4148 28204 4149 28244
rect 4107 28195 4149 28204
rect 7179 28244 7221 28253
rect 7179 28204 7180 28244
rect 7220 28204 7221 28244
rect 7179 28195 7221 28204
rect 11979 28244 12021 28253
rect 11979 28204 11980 28244
rect 12020 28204 12021 28244
rect 11979 28195 12021 28204
rect 12363 28244 12405 28253
rect 12363 28204 12364 28244
rect 12404 28204 12405 28244
rect 12363 28195 12405 28204
rect 17059 28244 17117 28245
rect 17059 28204 17068 28244
rect 17108 28204 17117 28244
rect 17059 28203 17117 28204
rect 21003 28244 21045 28253
rect 21003 28204 21004 28244
rect 21044 28204 21045 28244
rect 21003 28195 21045 28204
rect 28971 28244 29013 28253
rect 28971 28204 28972 28244
rect 29012 28204 29013 28244
rect 28971 28195 29013 28204
rect 35595 28244 35637 28253
rect 35595 28204 35596 28244
rect 35636 28204 35637 28244
rect 35595 28195 35637 28204
rect 49995 28244 50037 28253
rect 49995 28204 49996 28244
rect 50036 28204 50037 28244
rect 49995 28195 50037 28204
rect 4483 28160 4541 28161
rect 4483 28120 4492 28160
rect 4532 28120 4541 28160
rect 4483 28119 4541 28120
rect 6019 28160 6077 28161
rect 6019 28120 6028 28160
rect 6068 28120 6077 28160
rect 6019 28119 6077 28120
rect 7555 28160 7613 28161
rect 7555 28120 7564 28160
rect 7604 28120 7613 28160
rect 7555 28119 7613 28120
rect 10059 28160 10101 28169
rect 10059 28120 10060 28160
rect 10100 28120 10101 28160
rect 10059 28111 10101 28120
rect 12835 28160 12893 28161
rect 12835 28120 12844 28160
rect 12884 28120 12893 28160
rect 12835 28119 12893 28120
rect 14571 28160 14613 28169
rect 14571 28120 14572 28160
rect 14612 28120 14613 28160
rect 14571 28111 14613 28120
rect 20803 28160 20861 28161
rect 20803 28120 20812 28160
rect 20852 28120 20861 28160
rect 20803 28119 20861 28120
rect 22723 28160 22781 28161
rect 22723 28120 22732 28160
rect 22772 28120 22781 28160
rect 22723 28119 22781 28120
rect 26091 28160 26133 28169
rect 26091 28120 26092 28160
rect 26132 28120 26133 28160
rect 26091 28111 26133 28120
rect 26371 28160 26429 28161
rect 26371 28120 26380 28160
rect 26420 28120 26429 28160
rect 26371 28119 26429 28120
rect 28291 28160 28349 28161
rect 28291 28120 28300 28160
rect 28340 28120 28349 28160
rect 28291 28119 28349 28120
rect 38179 28160 38237 28161
rect 38179 28120 38188 28160
rect 38228 28120 38237 28160
rect 38179 28119 38237 28120
rect 39819 28160 39861 28169
rect 39819 28120 39820 28160
rect 39860 28120 39861 28160
rect 39819 28111 39861 28120
rect 43083 28160 43125 28169
rect 43083 28120 43084 28160
rect 43124 28120 43125 28160
rect 43083 28111 43125 28120
rect 43851 28160 43893 28169
rect 43851 28120 43852 28160
rect 43892 28120 43893 28160
rect 43851 28111 43893 28120
rect 46731 28160 46773 28169
rect 46731 28120 46732 28160
rect 46772 28120 46773 28160
rect 46731 28111 46773 28120
rect 48643 28160 48701 28161
rect 48643 28120 48652 28160
rect 48692 28120 48701 28160
rect 48643 28119 48701 28120
rect 49795 28160 49853 28161
rect 49795 28120 49804 28160
rect 49844 28120 49853 28160
rect 49795 28119 49853 28120
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 4683 27824 4725 27833
rect 4683 27784 4684 27824
rect 4724 27784 4725 27824
rect 4683 27775 4725 27784
rect 12171 27824 12213 27833
rect 12171 27784 12172 27824
rect 12212 27784 12213 27824
rect 12171 27775 12213 27784
rect 42891 27824 42933 27833
rect 42891 27784 42892 27824
rect 42932 27784 42933 27824
rect 42891 27775 42933 27784
rect 2667 27740 2709 27749
rect 2667 27700 2668 27740
rect 2708 27700 2709 27740
rect 2667 27691 2709 27700
rect 7467 27740 7509 27749
rect 7467 27700 7468 27740
rect 7508 27700 7509 27740
rect 7467 27691 7509 27700
rect 19851 27740 19893 27749
rect 19851 27700 19852 27740
rect 19892 27700 19893 27740
rect 19851 27691 19893 27700
rect 29739 27740 29781 27749
rect 29739 27700 29740 27740
rect 29780 27700 29781 27740
rect 29739 27691 29781 27700
rect 36363 27740 36405 27749
rect 36363 27700 36364 27740
rect 36404 27700 36405 27740
rect 36363 27691 36405 27700
rect 44427 27740 44469 27749
rect 44427 27700 44428 27740
rect 44468 27700 44469 27740
rect 44427 27691 44469 27700
rect 51627 27740 51669 27749
rect 51627 27700 51628 27740
rect 51668 27700 51669 27740
rect 51627 27691 51669 27700
rect 32150 27669 32192 27678
rect 2755 27656 2813 27657
rect 2755 27616 2764 27656
rect 2804 27616 2813 27656
rect 2755 27615 2813 27616
rect 3043 27656 3101 27657
rect 3043 27616 3052 27656
rect 3092 27616 3101 27656
rect 3043 27615 3101 27616
rect 3331 27656 3389 27657
rect 3331 27616 3340 27656
rect 3380 27616 3389 27656
rect 3331 27615 3389 27616
rect 3523 27656 3581 27657
rect 3523 27616 3532 27656
rect 3572 27616 3581 27656
rect 3523 27615 3581 27616
rect 3627 27656 3669 27665
rect 3627 27616 3628 27656
rect 3668 27616 3669 27656
rect 3627 27607 3669 27616
rect 3819 27656 3861 27665
rect 3819 27616 3820 27656
rect 3860 27616 3861 27656
rect 3819 27607 3861 27616
rect 4195 27656 4253 27657
rect 4195 27616 4204 27656
rect 4244 27616 4253 27656
rect 4195 27615 4253 27616
rect 5923 27656 5981 27657
rect 5923 27616 5932 27656
rect 5972 27616 5981 27656
rect 5923 27615 5981 27616
rect 6987 27656 7029 27665
rect 6987 27616 6988 27656
rect 7028 27616 7029 27656
rect 6987 27607 7029 27616
rect 7363 27656 7421 27657
rect 7363 27616 7372 27656
rect 7412 27616 7421 27656
rect 7363 27615 7421 27616
rect 7659 27656 7701 27665
rect 7659 27616 7660 27656
rect 7700 27616 7701 27656
rect 7659 27607 7701 27616
rect 7755 27656 7797 27665
rect 7755 27616 7756 27656
rect 7796 27616 7797 27656
rect 7755 27607 7797 27616
rect 7851 27656 7893 27665
rect 7851 27616 7852 27656
rect 7892 27616 7893 27656
rect 7851 27607 7893 27616
rect 7947 27656 7989 27665
rect 7947 27616 7948 27656
rect 7988 27616 7989 27656
rect 7947 27607 7989 27616
rect 8139 27656 8181 27665
rect 8139 27616 8140 27656
rect 8180 27616 8181 27656
rect 8139 27607 8181 27616
rect 8803 27656 8861 27657
rect 8803 27616 8812 27656
rect 8852 27616 8861 27656
rect 8803 27615 8861 27616
rect 9003 27656 9045 27665
rect 9003 27616 9004 27656
rect 9044 27616 9045 27656
rect 9003 27607 9045 27616
rect 9379 27656 9437 27657
rect 9379 27616 9388 27656
rect 9428 27616 9437 27656
rect 9379 27615 9437 27616
rect 10243 27656 10301 27657
rect 10243 27616 10252 27656
rect 10292 27616 10301 27656
rect 10243 27615 10301 27616
rect 11683 27656 11741 27657
rect 11683 27616 11692 27656
rect 11732 27616 11741 27656
rect 11683 27615 11741 27616
rect 12643 27656 12701 27657
rect 12643 27616 12652 27656
rect 12692 27616 12701 27656
rect 12643 27615 12701 27616
rect 13131 27656 13173 27665
rect 13131 27616 13132 27656
rect 13172 27616 13173 27656
rect 13131 27607 13173 27616
rect 13323 27656 13365 27665
rect 13323 27616 13324 27656
rect 13364 27616 13365 27656
rect 13323 27607 13365 27616
rect 13411 27656 13469 27657
rect 13411 27616 13420 27656
rect 13460 27616 13469 27656
rect 13411 27615 13469 27616
rect 13603 27656 13661 27657
rect 13603 27616 13612 27656
rect 13652 27616 13661 27656
rect 13603 27615 13661 27616
rect 13699 27656 13757 27657
rect 13699 27616 13708 27656
rect 13748 27616 13757 27656
rect 13699 27615 13757 27616
rect 13899 27656 13941 27665
rect 13899 27616 13900 27656
rect 13940 27616 13941 27656
rect 14142 27656 14200 27657
rect 13899 27607 13941 27616
rect 13987 27627 14045 27628
rect 13987 27587 13996 27627
rect 14036 27587 14045 27627
rect 14142 27616 14151 27656
rect 14191 27616 14200 27656
rect 14142 27615 14200 27616
rect 14755 27656 14813 27657
rect 14755 27616 14764 27656
rect 14804 27616 14813 27656
rect 14755 27615 14813 27616
rect 14851 27656 14909 27657
rect 14851 27616 14860 27656
rect 14900 27616 14909 27656
rect 14851 27615 14909 27616
rect 15051 27656 15093 27665
rect 15051 27616 15052 27656
rect 15092 27616 15093 27656
rect 15051 27607 15093 27616
rect 15147 27656 15189 27665
rect 15147 27616 15148 27656
rect 15188 27616 15189 27656
rect 16011 27656 16053 27665
rect 15147 27607 15189 27616
rect 15304 27641 15346 27650
rect 15304 27601 15305 27641
rect 15345 27601 15346 27641
rect 16011 27616 16012 27656
rect 16052 27616 16053 27656
rect 16011 27607 16053 27616
rect 16203 27656 16245 27665
rect 16203 27616 16204 27656
rect 16244 27616 16245 27656
rect 16203 27607 16245 27616
rect 16291 27656 16349 27657
rect 16291 27616 16300 27656
rect 16340 27616 16349 27656
rect 16291 27615 16349 27616
rect 17443 27656 17501 27657
rect 17443 27616 17452 27656
rect 17492 27616 17501 27656
rect 17443 27615 17501 27616
rect 18403 27656 18461 27657
rect 18403 27616 18412 27656
rect 18452 27616 18461 27656
rect 18403 27615 18461 27616
rect 19947 27656 19989 27665
rect 19947 27616 19948 27656
rect 19988 27616 19989 27656
rect 19947 27607 19989 27616
rect 20227 27656 20285 27657
rect 20227 27616 20236 27656
rect 20276 27616 20285 27656
rect 20227 27615 20285 27616
rect 20523 27656 20565 27665
rect 20523 27616 20524 27656
rect 20564 27616 20565 27656
rect 20523 27607 20565 27616
rect 20715 27656 20757 27665
rect 20715 27616 20716 27656
rect 20756 27616 20757 27656
rect 20715 27607 20757 27616
rect 20803 27656 20861 27657
rect 20803 27616 20812 27656
rect 20852 27616 20861 27656
rect 20803 27615 20861 27616
rect 21003 27656 21045 27665
rect 21003 27616 21004 27656
rect 21044 27616 21045 27656
rect 21003 27607 21045 27616
rect 21195 27656 21237 27665
rect 21195 27616 21196 27656
rect 21236 27616 21237 27656
rect 21195 27607 21237 27616
rect 21283 27656 21341 27657
rect 21283 27616 21292 27656
rect 21332 27616 21341 27656
rect 21283 27615 21341 27616
rect 21483 27656 21525 27665
rect 21483 27616 21484 27656
rect 21524 27616 21525 27656
rect 21483 27607 21525 27616
rect 21571 27656 21629 27657
rect 21571 27616 21580 27656
rect 21620 27616 21629 27656
rect 21571 27615 21629 27616
rect 21867 27656 21909 27665
rect 21867 27616 21868 27656
rect 21908 27616 21909 27656
rect 21867 27607 21909 27616
rect 22243 27656 22301 27657
rect 22243 27616 22252 27656
rect 22292 27616 22301 27656
rect 22243 27615 22301 27616
rect 23107 27656 23165 27657
rect 23107 27616 23116 27656
rect 23156 27616 23165 27656
rect 23107 27615 23165 27616
rect 24643 27656 24701 27657
rect 24643 27616 24652 27656
rect 24692 27616 24701 27656
rect 24835 27656 24893 27657
rect 24643 27615 24701 27616
rect 24747 27621 24789 27630
rect 15304 27592 15346 27601
rect 13987 27586 14045 27587
rect 24747 27581 24748 27621
rect 24788 27581 24789 27621
rect 24835 27616 24844 27656
rect 24884 27616 24893 27656
rect 24835 27615 24893 27616
rect 26283 27656 26325 27665
rect 26283 27616 26284 27656
rect 26324 27616 26325 27656
rect 26283 27607 26325 27616
rect 26755 27656 26813 27657
rect 26755 27616 26764 27656
rect 26804 27616 26813 27656
rect 26755 27615 26813 27616
rect 27715 27656 27773 27657
rect 27715 27616 27724 27656
rect 27764 27616 27773 27656
rect 27715 27615 27773 27616
rect 28011 27656 28053 27665
rect 28011 27616 28012 27656
rect 28052 27616 28053 27656
rect 28011 27607 28053 27616
rect 28107 27656 28149 27665
rect 28107 27616 28108 27656
rect 28148 27616 28149 27656
rect 28107 27607 28149 27616
rect 28491 27656 28533 27665
rect 28491 27616 28492 27656
rect 28532 27616 28533 27656
rect 28491 27607 28533 27616
rect 29059 27656 29117 27657
rect 29059 27616 29068 27656
rect 29108 27616 29117 27656
rect 29059 27615 29117 27616
rect 29547 27651 29589 27660
rect 29547 27611 29548 27651
rect 29588 27611 29589 27651
rect 29547 27602 29589 27611
rect 30507 27656 30549 27665
rect 30507 27616 30508 27656
rect 30548 27616 30549 27656
rect 30507 27607 30549 27616
rect 30699 27656 30741 27665
rect 30699 27616 30700 27656
rect 30740 27616 30741 27656
rect 30699 27607 30741 27616
rect 30787 27656 30845 27657
rect 30787 27616 30796 27656
rect 30836 27616 30845 27656
rect 30787 27615 30845 27616
rect 30987 27656 31029 27665
rect 30987 27616 30988 27656
rect 31028 27616 31029 27656
rect 30987 27607 31029 27616
rect 31179 27656 31221 27665
rect 31179 27616 31180 27656
rect 31220 27616 31221 27656
rect 31179 27607 31221 27616
rect 31267 27656 31325 27657
rect 31267 27616 31276 27656
rect 31316 27616 31325 27656
rect 31267 27615 31325 27616
rect 31467 27656 31509 27665
rect 31467 27616 31468 27656
rect 31508 27616 31509 27656
rect 31467 27607 31509 27616
rect 31563 27656 31605 27665
rect 31563 27616 31564 27656
rect 31604 27616 31605 27656
rect 31563 27607 31605 27616
rect 31659 27656 31701 27665
rect 31659 27616 31660 27656
rect 31700 27616 31701 27656
rect 31659 27607 31701 27616
rect 31755 27656 31797 27665
rect 31755 27616 31756 27656
rect 31796 27616 31797 27656
rect 31755 27607 31797 27616
rect 31947 27656 31989 27665
rect 31947 27616 31948 27656
rect 31988 27616 31989 27656
rect 32150 27629 32151 27669
rect 32191 27629 32192 27669
rect 32150 27620 32192 27629
rect 33283 27656 33341 27657
rect 31947 27607 31989 27616
rect 33283 27616 33292 27656
rect 33332 27616 33341 27656
rect 33283 27615 33341 27616
rect 34155 27656 34197 27665
rect 34155 27616 34156 27656
rect 34196 27616 34197 27656
rect 34155 27607 34197 27616
rect 34251 27656 34293 27665
rect 34251 27616 34252 27656
rect 34292 27616 34293 27656
rect 34251 27607 34293 27616
rect 34347 27656 34389 27665
rect 34347 27616 34348 27656
rect 34388 27616 34389 27656
rect 34347 27607 34389 27616
rect 34443 27656 34485 27665
rect 34443 27616 34444 27656
rect 34484 27616 34485 27656
rect 34443 27607 34485 27616
rect 35211 27656 35253 27665
rect 35211 27616 35212 27656
rect 35252 27616 35253 27656
rect 35211 27607 35253 27616
rect 36067 27656 36125 27657
rect 36067 27616 36076 27656
rect 36116 27616 36125 27656
rect 36067 27615 36125 27616
rect 36267 27656 36309 27665
rect 36267 27616 36268 27656
rect 36308 27616 36309 27656
rect 36267 27607 36309 27616
rect 36451 27656 36509 27657
rect 36451 27616 36460 27656
rect 36500 27616 36509 27656
rect 36451 27615 36509 27616
rect 37795 27656 37853 27657
rect 37795 27616 37804 27656
rect 37844 27616 37853 27656
rect 37795 27615 37853 27616
rect 38187 27656 38229 27665
rect 38187 27616 38188 27656
rect 38228 27616 38229 27656
rect 38187 27607 38229 27616
rect 38283 27656 38325 27665
rect 38283 27616 38284 27656
rect 38324 27616 38325 27656
rect 38283 27607 38325 27616
rect 38379 27656 38421 27665
rect 38379 27616 38380 27656
rect 38420 27616 38421 27656
rect 38379 27607 38421 27616
rect 38475 27656 38517 27665
rect 38475 27616 38476 27656
rect 38516 27616 38517 27656
rect 38475 27607 38517 27616
rect 38947 27656 39005 27657
rect 38947 27616 38956 27656
rect 38996 27616 39005 27656
rect 38947 27615 39005 27616
rect 39907 27656 39965 27657
rect 39907 27616 39916 27656
rect 39956 27616 39965 27656
rect 39907 27615 39965 27616
rect 40099 27656 40157 27657
rect 40099 27616 40108 27656
rect 40148 27616 40157 27656
rect 40099 27615 40157 27616
rect 42979 27656 43037 27657
rect 42979 27616 42988 27656
rect 43028 27616 43037 27656
rect 43275 27656 43317 27665
rect 42979 27615 43037 27616
rect 43171 27637 43229 27638
rect 43171 27597 43180 27637
rect 43220 27597 43229 27637
rect 43275 27616 43276 27656
rect 43316 27616 43317 27656
rect 43275 27607 43317 27616
rect 43467 27656 43509 27665
rect 43467 27616 43468 27656
rect 43508 27616 43509 27656
rect 43467 27607 43509 27616
rect 43659 27656 43701 27665
rect 43659 27616 43660 27656
rect 43700 27616 43701 27656
rect 43659 27607 43701 27616
rect 43755 27656 43797 27665
rect 43755 27616 43756 27656
rect 43796 27616 43797 27656
rect 43755 27607 43797 27616
rect 43851 27656 43893 27665
rect 43851 27616 43852 27656
rect 43892 27616 43893 27656
rect 43851 27607 43893 27616
rect 43947 27656 43989 27665
rect 43947 27616 43948 27656
rect 43988 27616 43989 27656
rect 43947 27607 43989 27616
rect 44331 27656 44373 27665
rect 44331 27616 44332 27656
rect 44372 27616 44373 27656
rect 44331 27607 44373 27616
rect 44515 27656 44573 27657
rect 44515 27616 44524 27656
rect 44564 27616 44573 27656
rect 44515 27615 44573 27616
rect 45099 27656 45141 27665
rect 45099 27616 45100 27656
rect 45140 27616 45141 27656
rect 45099 27607 45141 27616
rect 45195 27656 45237 27665
rect 45195 27616 45196 27656
rect 45236 27616 45237 27656
rect 45195 27607 45237 27616
rect 45291 27656 45333 27665
rect 45291 27616 45292 27656
rect 45332 27616 45333 27656
rect 45291 27607 45333 27616
rect 45387 27656 45429 27665
rect 45387 27616 45388 27656
rect 45428 27616 45429 27656
rect 45387 27607 45429 27616
rect 45963 27656 46005 27665
rect 45963 27616 45964 27656
rect 46004 27616 46005 27656
rect 45963 27607 46005 27616
rect 46155 27656 46197 27665
rect 46155 27616 46156 27656
rect 46196 27616 46197 27656
rect 46155 27607 46197 27616
rect 46243 27656 46301 27657
rect 46243 27616 46252 27656
rect 46292 27616 46301 27656
rect 46243 27615 46301 27616
rect 46915 27656 46973 27657
rect 46915 27616 46924 27656
rect 46964 27616 46973 27656
rect 46915 27615 46973 27616
rect 47203 27656 47261 27657
rect 47203 27616 47212 27656
rect 47252 27616 47261 27656
rect 47203 27615 47261 27616
rect 47499 27656 47541 27665
rect 47499 27616 47500 27656
rect 47540 27616 47541 27656
rect 47499 27607 47541 27616
rect 47595 27656 47637 27665
rect 47595 27616 47596 27656
rect 47636 27616 47637 27656
rect 47595 27607 47637 27616
rect 47691 27656 47733 27665
rect 47691 27616 47692 27656
rect 47732 27616 47733 27656
rect 47691 27607 47733 27616
rect 47787 27656 47829 27665
rect 47787 27616 47788 27656
rect 47828 27616 47829 27656
rect 47787 27607 47829 27616
rect 48171 27656 48213 27665
rect 48171 27616 48172 27656
rect 48212 27616 48213 27656
rect 48171 27607 48213 27616
rect 48267 27656 48309 27665
rect 48267 27616 48268 27656
rect 48308 27616 48309 27656
rect 48267 27607 48309 27616
rect 48363 27656 48405 27665
rect 48363 27616 48364 27656
rect 48404 27616 48405 27656
rect 48363 27607 48405 27616
rect 48459 27656 48501 27665
rect 48459 27616 48460 27656
rect 48500 27616 48501 27656
rect 48459 27607 48501 27616
rect 48643 27656 48701 27657
rect 48643 27616 48652 27656
rect 48692 27616 48701 27656
rect 48643 27615 48701 27616
rect 48747 27656 48789 27665
rect 48747 27616 48748 27656
rect 48788 27616 48789 27656
rect 48747 27607 48789 27616
rect 48939 27656 48981 27665
rect 48939 27616 48940 27656
rect 48980 27616 48981 27656
rect 48939 27607 48981 27616
rect 50371 27656 50429 27657
rect 50371 27616 50380 27656
rect 50420 27616 50429 27656
rect 50371 27615 50429 27616
rect 51235 27656 51293 27657
rect 51235 27616 51244 27656
rect 51284 27616 51293 27656
rect 51235 27615 51293 27616
rect 43171 27596 43229 27597
rect 5635 27572 5693 27573
rect 5635 27532 5644 27572
rect 5684 27532 5693 27572
rect 5635 27531 5693 27532
rect 19171 27572 19229 27573
rect 19171 27532 19180 27572
rect 19220 27532 19229 27572
rect 19171 27531 19229 27532
rect 24267 27572 24309 27581
rect 24747 27572 24789 27581
rect 25515 27572 25557 27581
rect 24267 27532 24268 27572
rect 24308 27532 24309 27572
rect 24267 27523 24309 27532
rect 25515 27532 25516 27572
rect 25556 27532 25557 27572
rect 25515 27523 25557 27532
rect 28587 27572 28629 27581
rect 28587 27532 28588 27572
rect 28628 27532 28629 27572
rect 28587 27523 28629 27532
rect 49227 27572 49269 27581
rect 49227 27532 49228 27572
rect 49268 27532 49269 27572
rect 49227 27523 49269 27532
rect 1707 27488 1749 27497
rect 1707 27448 1708 27488
rect 1748 27448 1749 27488
rect 1707 27439 1749 27448
rect 3243 27488 3285 27497
rect 3243 27448 3244 27488
rect 3284 27448 3285 27488
rect 3243 27439 3285 27448
rect 19555 27488 19613 27489
rect 19555 27448 19564 27488
rect 19604 27448 19613 27488
rect 19555 27447 19613 27448
rect 21003 27488 21045 27497
rect 21003 27448 21004 27488
rect 21044 27448 21045 27488
rect 21003 27439 21045 27448
rect 26091 27488 26133 27497
rect 26091 27448 26092 27488
rect 26132 27448 26133 27488
rect 26091 27439 26133 27448
rect 32043 27488 32085 27497
rect 32043 27448 32044 27488
rect 32084 27448 32085 27488
rect 32043 27439 32085 27448
rect 33099 27488 33141 27497
rect 33099 27448 33100 27488
rect 33140 27448 33141 27488
rect 33099 27439 33141 27448
rect 36939 27488 36981 27497
rect 36939 27448 36940 27488
rect 36980 27448 36981 27488
rect 36939 27439 36981 27448
rect 42219 27488 42261 27497
rect 42219 27448 42220 27488
rect 42260 27448 42261 27488
rect 42219 27439 42261 27448
rect 46443 27488 46485 27497
rect 46443 27448 46444 27488
rect 46484 27448 46485 27488
rect 46443 27439 46485 27448
rect 2955 27404 2997 27413
rect 2955 27364 2956 27404
rect 2996 27364 2997 27404
rect 2955 27355 2997 27364
rect 3819 27404 3861 27413
rect 3819 27364 3820 27404
rect 3860 27364 3861 27404
rect 3819 27355 3861 27364
rect 5451 27404 5493 27413
rect 5451 27364 5452 27404
rect 5492 27364 5493 27404
rect 5451 27355 5493 27364
rect 5835 27404 5877 27413
rect 5835 27364 5836 27404
rect 5876 27364 5877 27404
rect 5835 27355 5877 27364
rect 6795 27404 6837 27413
rect 6795 27364 6796 27404
rect 6836 27364 6837 27404
rect 6795 27355 6837 27364
rect 11395 27404 11453 27405
rect 11395 27364 11404 27404
rect 11444 27364 11453 27404
rect 11395 27363 11453 27364
rect 13131 27404 13173 27413
rect 13131 27364 13132 27404
rect 13172 27364 13173 27404
rect 13131 27355 13173 27364
rect 13611 27404 13653 27413
rect 13611 27364 13612 27404
rect 13652 27364 13653 27404
rect 13611 27355 13653 27364
rect 14763 27404 14805 27413
rect 14763 27364 14764 27404
rect 14804 27364 14805 27404
rect 14763 27355 14805 27364
rect 16011 27404 16053 27413
rect 16011 27364 16012 27404
rect 16052 27364 16053 27404
rect 16011 27355 16053 27364
rect 19371 27404 19413 27413
rect 19371 27364 19372 27404
rect 19412 27364 19413 27404
rect 19371 27355 19413 27364
rect 20523 27404 20565 27413
rect 20523 27364 20524 27404
rect 20564 27364 20565 27404
rect 20523 27355 20565 27364
rect 25131 27404 25173 27413
rect 25131 27364 25132 27404
rect 25172 27364 25173 27404
rect 25131 27355 25173 27364
rect 30507 27404 30549 27413
rect 30507 27364 30508 27404
rect 30548 27364 30549 27404
rect 30507 27355 30549 27364
rect 30987 27404 31029 27413
rect 30987 27364 30988 27404
rect 31028 27364 31029 27404
rect 30987 27355 31029 27364
rect 33955 27404 34013 27405
rect 33955 27364 33964 27404
rect 34004 27364 34013 27404
rect 33955 27363 34013 27364
rect 37707 27404 37749 27413
rect 37707 27364 37708 27404
rect 37748 27364 37749 27404
rect 37707 27355 37749 27364
rect 39619 27404 39677 27405
rect 39619 27364 39628 27404
rect 39668 27364 39677 27404
rect 39619 27363 39677 27364
rect 43467 27404 43509 27413
rect 43467 27364 43468 27404
rect 43508 27364 43509 27404
rect 43467 27355 43509 27364
rect 45963 27404 46005 27413
rect 45963 27364 45964 27404
rect 46004 27364 46005 27404
rect 45963 27355 46005 27364
rect 47019 27404 47061 27413
rect 47019 27364 47020 27404
rect 47060 27364 47061 27404
rect 47019 27355 47061 27364
rect 47307 27404 47349 27413
rect 47307 27364 47308 27404
rect 47348 27364 47349 27404
rect 47307 27355 47349 27364
rect 48939 27404 48981 27413
rect 48939 27364 48940 27404
rect 48980 27364 48981 27404
rect 48939 27355 48981 27364
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 3619 27068 3677 27069
rect 3619 27028 3628 27068
rect 3668 27028 3677 27068
rect 3619 27027 3677 27028
rect 4675 27068 4733 27069
rect 4675 27028 4684 27068
rect 4724 27028 4733 27068
rect 4675 27027 4733 27028
rect 7851 27068 7893 27077
rect 7851 27028 7852 27068
rect 7892 27028 7893 27068
rect 7851 27019 7893 27028
rect 9187 27068 9245 27069
rect 9187 27028 9196 27068
rect 9236 27028 9245 27068
rect 9187 27027 9245 27028
rect 11971 27068 12029 27069
rect 11971 27028 11980 27068
rect 12020 27028 12029 27068
rect 11971 27027 12029 27028
rect 13515 27068 13557 27077
rect 13515 27028 13516 27068
rect 13556 27028 13557 27068
rect 13515 27019 13557 27028
rect 14379 27068 14421 27077
rect 14379 27028 14380 27068
rect 14420 27028 14421 27068
rect 14379 27019 14421 27028
rect 15051 27068 15093 27077
rect 15051 27028 15052 27068
rect 15092 27028 15093 27068
rect 15051 27019 15093 27028
rect 21283 27068 21341 27069
rect 21283 27028 21292 27068
rect 21332 27028 21341 27068
rect 21283 27027 21341 27028
rect 27915 27068 27957 27077
rect 27915 27028 27916 27068
rect 27956 27028 27957 27068
rect 27915 27019 27957 27028
rect 31371 27068 31413 27077
rect 31371 27028 31372 27068
rect 31412 27028 31413 27068
rect 31371 27019 31413 27028
rect 31843 27068 31901 27069
rect 31843 27028 31852 27068
rect 31892 27028 31901 27068
rect 31843 27027 31901 27028
rect 32803 27068 32861 27069
rect 32803 27028 32812 27068
rect 32852 27028 32861 27068
rect 32803 27027 32861 27028
rect 38755 27068 38813 27069
rect 38755 27028 38764 27068
rect 38804 27028 38813 27068
rect 38755 27027 38813 27028
rect 39619 27068 39677 27069
rect 39619 27028 39628 27068
rect 39668 27028 39677 27068
rect 39619 27027 39677 27028
rect 47971 27068 48029 27069
rect 47971 27028 47980 27068
rect 48020 27028 48029 27068
rect 47971 27027 48029 27028
rect 48163 27068 48221 27069
rect 48163 27028 48172 27068
rect 48212 27028 48221 27068
rect 48163 27027 48221 27028
rect 49323 27068 49365 27077
rect 49323 27028 49324 27068
rect 49364 27028 49365 27068
rect 49323 27019 49365 27028
rect 10059 26984 10101 26993
rect 10059 26944 10060 26984
rect 10100 26944 10101 26984
rect 10059 26935 10101 26944
rect 18019 26984 18077 26985
rect 18019 26944 18028 26984
rect 18068 26944 18077 26984
rect 18019 26943 18077 26944
rect 19267 26984 19325 26985
rect 19267 26944 19276 26984
rect 19316 26944 19325 26984
rect 19267 26943 19325 26944
rect 22347 26984 22389 26993
rect 22347 26944 22348 26984
rect 22388 26944 22389 26984
rect 22347 26935 22389 26944
rect 24939 26984 24981 26993
rect 24939 26944 24940 26984
rect 24980 26944 24981 26984
rect 24939 26935 24981 26944
rect 26187 26984 26229 26993
rect 26187 26944 26188 26984
rect 26228 26944 26229 26984
rect 26187 26935 26229 26944
rect 44139 26900 44181 26909
rect 44139 26860 44140 26900
rect 44180 26860 44181 26900
rect 30411 26851 30453 26860
rect 44139 26851 44181 26860
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1603 26816 1661 26817
rect 1603 26776 1612 26816
rect 1652 26776 1661 26816
rect 1603 26775 1661 26776
rect 2467 26816 2525 26817
rect 2467 26776 2476 26816
rect 2516 26776 2525 26816
rect 2467 26775 2525 26776
rect 4483 26816 4541 26817
rect 4483 26776 4492 26816
rect 4532 26776 4541 26816
rect 4483 26775 4541 26776
rect 5827 26816 5885 26817
rect 5827 26776 5836 26816
rect 5876 26776 5885 26816
rect 5827 26775 5885 26776
rect 6691 26816 6749 26817
rect 6691 26776 6700 26816
rect 6740 26776 6749 26816
rect 6691 26775 6749 26776
rect 7083 26816 7125 26825
rect 7083 26776 7084 26816
rect 7124 26776 7125 26816
rect 7083 26767 7125 26776
rect 8427 26816 8469 26825
rect 8427 26776 8428 26816
rect 8468 26776 8469 26816
rect 8427 26767 8469 26776
rect 9859 26816 9917 26817
rect 9859 26776 9868 26816
rect 9908 26776 9917 26816
rect 9859 26775 9917 26776
rect 10531 26816 10589 26817
rect 10531 26776 10540 26816
rect 10580 26776 10589 26816
rect 10531 26775 10589 26776
rect 10723 26816 10781 26817
rect 10723 26776 10732 26816
rect 10772 26776 10781 26816
rect 10723 26775 10781 26776
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 11299 26816 11357 26817
rect 11299 26776 11308 26816
rect 11348 26776 11357 26816
rect 11299 26775 11357 26776
rect 11595 26816 11637 26825
rect 11595 26776 11596 26816
rect 11636 26776 11637 26816
rect 11595 26767 11637 26776
rect 12171 26816 12213 26825
rect 12171 26776 12172 26816
rect 12212 26776 12213 26816
rect 12171 26767 12213 26776
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12363 26816 12405 26825
rect 12363 26776 12364 26816
rect 12404 26776 12405 26816
rect 12363 26767 12405 26776
rect 12459 26816 12501 26825
rect 12459 26776 12460 26816
rect 12500 26776 12501 26816
rect 12459 26767 12501 26776
rect 13707 26816 13749 26825
rect 13707 26776 13708 26816
rect 13748 26776 13749 26816
rect 13707 26767 13749 26776
rect 14083 26816 14141 26817
rect 14083 26776 14092 26816
rect 14132 26776 14141 26816
rect 14083 26775 14141 26776
rect 14187 26816 14229 26825
rect 14187 26776 14188 26816
rect 14228 26776 14229 26816
rect 14187 26767 14229 26776
rect 14379 26816 14421 26825
rect 14379 26776 14380 26816
rect 14420 26776 14421 26816
rect 14379 26767 14421 26776
rect 14563 26816 14621 26817
rect 14563 26776 14572 26816
rect 14612 26776 14621 26816
rect 14563 26775 14621 26776
rect 14667 26816 14709 26825
rect 14667 26776 14668 26816
rect 14708 26776 14709 26816
rect 14667 26767 14709 26776
rect 14859 26816 14901 26825
rect 14859 26776 14860 26816
rect 14900 26776 14901 26816
rect 14859 26767 14901 26776
rect 15051 26816 15093 26825
rect 15051 26776 15052 26816
rect 15092 26776 15093 26816
rect 15051 26767 15093 26776
rect 15243 26816 15285 26825
rect 15243 26776 15244 26816
rect 15284 26776 15285 26816
rect 15243 26767 15285 26776
rect 15331 26816 15389 26817
rect 15331 26776 15340 26816
rect 15380 26776 15389 26816
rect 15331 26775 15389 26776
rect 16771 26816 16829 26817
rect 16771 26776 16780 26816
rect 16820 26776 16829 26816
rect 16771 26775 16829 26776
rect 16971 26816 17013 26825
rect 16971 26776 16972 26816
rect 17012 26776 17013 26816
rect 16971 26767 17013 26776
rect 17163 26816 17205 26825
rect 17163 26776 17164 26816
rect 17204 26776 17205 26816
rect 17163 26767 17205 26776
rect 17347 26816 17405 26817
rect 17347 26776 17356 26816
rect 17396 26776 17405 26816
rect 17347 26775 17405 26776
rect 17547 26816 17589 26825
rect 17547 26776 17548 26816
rect 17588 26776 17589 26816
rect 17547 26767 17589 26776
rect 17643 26816 17685 26825
rect 17643 26776 17644 26816
rect 17684 26776 17685 26816
rect 17643 26767 17685 26776
rect 17739 26816 17781 26825
rect 17739 26776 17740 26816
rect 17780 26776 17781 26816
rect 17739 26767 17781 26776
rect 18691 26816 18749 26817
rect 18691 26776 18700 26816
rect 18740 26776 18749 26816
rect 18691 26775 18749 26776
rect 19659 26816 19701 26825
rect 19659 26776 19660 26816
rect 19700 26776 19701 26816
rect 19659 26767 19701 26776
rect 19939 26816 19997 26817
rect 19939 26776 19948 26816
rect 19988 26776 19997 26816
rect 19939 26775 19997 26776
rect 20419 26816 20477 26817
rect 20419 26776 20428 26816
rect 20468 26776 20477 26816
rect 20419 26775 20477 26776
rect 21955 26816 22013 26817
rect 21955 26776 21964 26816
rect 22004 26776 22013 26816
rect 21955 26775 22013 26776
rect 24259 26816 24317 26817
rect 24259 26776 24268 26816
rect 24308 26776 24317 26816
rect 24259 26775 24317 26776
rect 24459 26816 24501 26825
rect 24459 26776 24460 26816
rect 24500 26776 24501 26816
rect 24459 26767 24501 26776
rect 24739 26816 24797 26817
rect 24739 26776 24748 26816
rect 24788 26776 24797 26816
rect 24739 26775 24797 26776
rect 27339 26816 27381 26825
rect 27339 26776 27340 26816
rect 27380 26776 27381 26816
rect 27339 26767 27381 26776
rect 28779 26816 28821 26825
rect 28779 26776 28780 26816
rect 28820 26776 28821 26816
rect 28779 26767 28821 26776
rect 28971 26816 29013 26825
rect 28971 26776 28972 26816
rect 29012 26776 29013 26816
rect 28971 26767 29013 26776
rect 29059 26816 29117 26817
rect 29059 26776 29068 26816
rect 29108 26776 29117 26816
rect 29059 26775 29117 26776
rect 29443 26816 29501 26817
rect 29443 26776 29452 26816
rect 29492 26776 29501 26816
rect 29443 26775 29501 26776
rect 29547 26816 29589 26825
rect 29547 26776 29548 26816
rect 29588 26776 29589 26816
rect 29547 26767 29589 26776
rect 29643 26816 29685 26825
rect 29643 26776 29644 26816
rect 29684 26776 29685 26816
rect 29643 26767 29685 26776
rect 30307 26816 30365 26817
rect 30307 26776 30316 26816
rect 30356 26776 30365 26816
rect 30411 26811 30412 26851
rect 30452 26811 30453 26851
rect 30411 26802 30453 26811
rect 30499 26816 30557 26817
rect 30307 26775 30365 26776
rect 30499 26776 30508 26816
rect 30548 26776 30557 26816
rect 30499 26775 30557 26776
rect 30891 26816 30933 26825
rect 30891 26776 30892 26816
rect 30932 26776 30933 26816
rect 30891 26767 30933 26776
rect 31083 26816 31125 26825
rect 31083 26776 31084 26816
rect 31124 26776 31125 26816
rect 31083 26767 31125 26776
rect 31171 26816 31229 26817
rect 31171 26776 31180 26816
rect 31220 26776 31229 26816
rect 31171 26775 31229 26776
rect 31371 26816 31413 26825
rect 31371 26776 31372 26816
rect 31412 26776 31413 26816
rect 31371 26767 31413 26776
rect 31563 26816 31605 26825
rect 31563 26776 31564 26816
rect 31604 26776 31605 26816
rect 31563 26767 31605 26776
rect 31651 26816 31709 26817
rect 31651 26776 31660 26816
rect 31700 26776 31709 26816
rect 31651 26775 31709 26776
rect 32139 26816 32181 26825
rect 32139 26776 32140 26816
rect 32180 26776 32181 26816
rect 32139 26767 32181 26776
rect 32235 26816 32277 26825
rect 32235 26776 32236 26816
rect 32276 26776 32277 26816
rect 32235 26767 32277 26776
rect 32515 26816 32573 26817
rect 32515 26776 32524 26816
rect 32564 26776 32573 26816
rect 32515 26775 32573 26776
rect 33955 26816 34013 26817
rect 33955 26776 33964 26816
rect 34004 26776 34013 26816
rect 33955 26775 34013 26776
rect 34819 26816 34877 26817
rect 34819 26776 34828 26816
rect 34868 26776 34877 26816
rect 34819 26775 34877 26776
rect 35499 26816 35541 26825
rect 35499 26776 35500 26816
rect 35540 26776 35541 26816
rect 35499 26767 35541 26776
rect 35595 26816 35637 26825
rect 35595 26776 35596 26816
rect 35636 26776 35637 26816
rect 35595 26767 35637 26776
rect 35691 26816 35733 26825
rect 35691 26776 35692 26816
rect 35732 26776 35733 26816
rect 35691 26767 35733 26776
rect 35883 26816 35925 26825
rect 35883 26776 35884 26816
rect 35924 26776 35925 26816
rect 35883 26767 35925 26776
rect 36075 26816 36117 26825
rect 36075 26776 36076 26816
rect 36116 26776 36117 26816
rect 36075 26767 36117 26776
rect 36163 26816 36221 26817
rect 36163 26776 36172 26816
rect 36212 26776 36221 26816
rect 36163 26775 36221 26776
rect 36739 26816 36797 26817
rect 36739 26776 36748 26816
rect 36788 26776 36797 26816
rect 36739 26775 36797 26776
rect 37603 26816 37661 26817
rect 37603 26776 37612 26816
rect 37652 26776 37661 26816
rect 37603 26775 37661 26776
rect 38947 26816 39005 26817
rect 38947 26776 38956 26816
rect 38996 26776 39005 26816
rect 38947 26775 39005 26776
rect 40299 26816 40341 26825
rect 40299 26776 40300 26816
rect 40340 26776 40341 26816
rect 40299 26767 40341 26776
rect 41739 26816 41781 26825
rect 41739 26776 41740 26816
rect 41780 26776 41781 26816
rect 41739 26767 41781 26776
rect 42115 26816 42173 26817
rect 42115 26776 42124 26816
rect 42164 26776 42173 26816
rect 42115 26775 42173 26776
rect 42979 26816 43037 26817
rect 42979 26776 42988 26816
rect 43028 26776 43037 26816
rect 42979 26775 43037 26776
rect 44995 26816 45053 26817
rect 44995 26776 45004 26816
rect 45044 26776 45053 26816
rect 44995 26775 45053 26776
rect 45579 26816 45621 26825
rect 45579 26776 45580 26816
rect 45620 26776 45621 26816
rect 45579 26767 45621 26776
rect 45955 26816 46013 26817
rect 45955 26776 45964 26816
rect 46004 26776 46013 26816
rect 45955 26775 46013 26776
rect 46819 26816 46877 26817
rect 46819 26776 46828 26816
rect 46868 26776 46877 26816
rect 46819 26775 46877 26776
rect 48835 26816 48893 26817
rect 48835 26776 48844 26816
rect 48884 26776 48893 26816
rect 48835 26775 48893 26776
rect 49027 26816 49085 26817
rect 49027 26776 49036 26816
rect 49076 26776 49085 26816
rect 49027 26775 49085 26776
rect 49131 26816 49173 26825
rect 49131 26776 49132 26816
rect 49172 26776 49173 26816
rect 49131 26767 49173 26776
rect 49323 26816 49365 26825
rect 49323 26776 49324 26816
rect 49364 26776 49365 26816
rect 49323 26767 49365 26776
rect 49611 26816 49653 26825
rect 49611 26776 49612 26816
rect 49652 26776 49653 26816
rect 49611 26767 49653 26776
rect 49987 26816 50045 26817
rect 49987 26776 49996 26816
rect 50036 26776 50045 26816
rect 49987 26775 50045 26776
rect 50851 26816 50909 26817
rect 50851 26776 50860 26816
rect 50900 26776 50909 26816
rect 50851 26775 50909 26776
rect 11691 26732 11733 26741
rect 11691 26692 11692 26732
rect 11732 26692 11733 26732
rect 11691 26683 11733 26692
rect 16875 26732 16917 26741
rect 16875 26692 16876 26732
rect 16916 26692 16917 26732
rect 16875 26683 16917 26692
rect 17259 26732 17301 26741
rect 17259 26692 17260 26732
rect 17300 26692 17301 26732
rect 17259 26683 17301 26692
rect 19563 26732 19605 26741
rect 19563 26692 19564 26732
rect 19604 26692 19605 26732
rect 19563 26683 19605 26692
rect 24363 26732 24405 26741
rect 24363 26692 24364 26732
rect 24404 26692 24405 26732
rect 24363 26683 24405 26692
rect 35211 26732 35253 26741
rect 35211 26692 35212 26732
rect 35252 26692 35253 26732
rect 35211 26683 35253 26692
rect 36363 26732 36405 26741
rect 36363 26692 36364 26732
rect 36404 26692 36405 26732
rect 36363 26683 36405 26692
rect 3811 26648 3869 26649
rect 3811 26608 3820 26648
rect 3860 26608 3869 26648
rect 3811 26607 3869 26608
rect 8043 26648 8085 26657
rect 8043 26608 8044 26648
rect 8084 26608 8085 26648
rect 8043 26599 8085 26608
rect 10443 26648 10485 26657
rect 10443 26608 10444 26648
rect 10484 26608 10485 26648
rect 10443 26599 10485 26608
rect 10915 26648 10973 26649
rect 10915 26608 10924 26648
rect 10964 26608 10973 26648
rect 10915 26607 10973 26608
rect 14755 26648 14813 26649
rect 14755 26608 14764 26648
rect 14804 26608 14813 26648
rect 14755 26607 14813 26608
rect 17827 26648 17885 26649
rect 17827 26608 17836 26648
rect 17876 26608 17885 26648
rect 17827 26607 17885 26608
rect 21091 26648 21149 26649
rect 21091 26608 21100 26648
rect 21140 26608 21149 26648
rect 21091 26607 21149 26608
rect 28867 26648 28925 26649
rect 28867 26608 28876 26648
rect 28916 26608 28925 26648
rect 28867 26607 28925 26608
rect 30027 26648 30069 26657
rect 30027 26608 30028 26648
rect 30068 26608 30069 26648
rect 30027 26599 30069 26608
rect 30979 26648 31037 26649
rect 30979 26608 30988 26648
rect 31028 26608 31037 26648
rect 30979 26607 31037 26608
rect 35395 26648 35453 26649
rect 35395 26608 35404 26648
rect 35444 26608 35453 26648
rect 35395 26607 35453 26608
rect 35971 26648 36029 26649
rect 35971 26608 35980 26648
rect 36020 26608 36029 26648
rect 35971 26607 36029 26608
rect 40683 26648 40725 26657
rect 40683 26608 40684 26648
rect 40724 26608 40725 26648
rect 40683 26599 40725 26608
rect 44323 26648 44381 26649
rect 44323 26608 44332 26648
rect 44372 26608 44381 26648
rect 44323 26607 44381 26608
rect 52003 26648 52061 26649
rect 52003 26608 52012 26648
rect 52052 26608 52061 26648
rect 52003 26607 52061 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 3619 26312 3677 26313
rect 3619 26272 3628 26312
rect 3668 26272 3677 26312
rect 3619 26271 3677 26272
rect 3811 26312 3869 26313
rect 3811 26272 3820 26312
rect 3860 26272 3869 26312
rect 3811 26271 3869 26272
rect 9187 26312 9245 26313
rect 9187 26272 9196 26312
rect 9236 26272 9245 26312
rect 9187 26271 9245 26272
rect 20619 26312 20661 26321
rect 20619 26272 20620 26312
rect 20660 26272 20661 26312
rect 20619 26263 20661 26272
rect 29635 26312 29693 26313
rect 29635 26272 29644 26312
rect 29684 26272 29693 26312
rect 29635 26271 29693 26272
rect 31755 26312 31797 26321
rect 31755 26272 31756 26312
rect 31796 26272 31797 26312
rect 31755 26263 31797 26272
rect 43555 26312 43613 26313
rect 43555 26272 43564 26312
rect 43604 26272 43613 26312
rect 43555 26271 43613 26272
rect 45675 26312 45717 26321
rect 45675 26272 45676 26312
rect 45716 26272 45717 26312
rect 45675 26263 45717 26272
rect 49803 26312 49845 26321
rect 49803 26272 49804 26312
rect 49844 26272 49845 26312
rect 49803 26263 49845 26272
rect 1227 26228 1269 26237
rect 1227 26188 1228 26228
rect 1268 26188 1269 26228
rect 1227 26179 1269 26188
rect 4395 26228 4437 26237
rect 4395 26188 4396 26228
rect 4436 26188 4437 26228
rect 4395 26179 4437 26188
rect 7851 26228 7893 26237
rect 7851 26188 7852 26228
rect 7892 26188 7893 26228
rect 7851 26179 7893 26188
rect 15147 26228 15189 26237
rect 15147 26188 15148 26228
rect 15188 26188 15189 26228
rect 15147 26179 15189 26188
rect 17163 26228 17205 26237
rect 17163 26188 17164 26228
rect 17204 26188 17205 26228
rect 17163 26179 17205 26188
rect 39147 26228 39189 26237
rect 39147 26188 39148 26228
rect 39188 26188 39189 26228
rect 39147 26179 39189 26188
rect 44235 26228 44277 26237
rect 44235 26188 44236 26228
rect 44276 26188 44277 26228
rect 44235 26179 44277 26188
rect 4011 26165 4053 26174
rect 1603 26144 1661 26145
rect 1603 26104 1612 26144
rect 1652 26104 1661 26144
rect 1603 26103 1661 26104
rect 2467 26144 2525 26145
rect 2467 26104 2476 26144
rect 2516 26104 2525 26144
rect 4011 26125 4012 26165
rect 4052 26125 4053 26165
rect 33859 26159 33917 26160
rect 4011 26116 4053 26125
rect 4107 26144 4149 26153
rect 2467 26103 2525 26104
rect 4107 26104 4108 26144
rect 4148 26104 4149 26144
rect 3907 26102 3965 26103
rect 3907 26062 3916 26102
rect 3956 26062 3965 26102
rect 4107 26095 4149 26104
rect 4299 26144 4341 26153
rect 4299 26104 4300 26144
rect 4340 26104 4341 26144
rect 4299 26095 4341 26104
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 4579 26144 4637 26145
rect 4579 26104 4588 26144
rect 4628 26104 4637 26144
rect 4579 26103 4637 26104
rect 4963 26144 5021 26145
rect 4963 26104 4972 26144
rect 5012 26104 5021 26144
rect 4963 26103 5021 26104
rect 5067 26144 5109 26153
rect 5067 26104 5068 26144
rect 5108 26104 5109 26144
rect 5067 26095 5109 26104
rect 5259 26144 5301 26153
rect 5259 26104 5260 26144
rect 5300 26104 5301 26144
rect 5259 26095 5301 26104
rect 6987 26144 7029 26153
rect 6987 26104 6988 26144
rect 7028 26104 7029 26144
rect 6987 26095 7029 26104
rect 7459 26144 7517 26145
rect 7459 26104 7468 26144
rect 7508 26104 7517 26144
rect 7459 26103 7517 26104
rect 7755 26144 7797 26153
rect 7755 26104 7756 26144
rect 7796 26104 7797 26144
rect 7755 26095 7797 26104
rect 9099 26144 9141 26153
rect 9099 26104 9100 26144
rect 9140 26104 9141 26144
rect 9099 26095 9141 26104
rect 9291 26144 9333 26153
rect 9291 26104 9292 26144
rect 9332 26104 9333 26144
rect 9291 26095 9333 26104
rect 9379 26144 9437 26145
rect 9379 26104 9388 26144
rect 9428 26104 9437 26144
rect 9379 26103 9437 26104
rect 10723 26144 10781 26145
rect 10723 26104 10732 26144
rect 10772 26104 10781 26144
rect 10723 26103 10781 26104
rect 10915 26144 10973 26145
rect 10915 26104 10924 26144
rect 10964 26104 10973 26144
rect 10915 26103 10973 26104
rect 11115 26144 11157 26153
rect 11115 26104 11116 26144
rect 11156 26104 11157 26144
rect 11115 26095 11157 26104
rect 11299 26144 11357 26145
rect 11299 26104 11308 26144
rect 11348 26104 11357 26144
rect 11299 26103 11357 26104
rect 12259 26144 12317 26145
rect 12259 26104 12268 26144
rect 12308 26104 12317 26144
rect 12259 26103 12317 26104
rect 12547 26144 12605 26145
rect 12547 26104 12556 26144
rect 12596 26104 12605 26144
rect 12547 26103 12605 26104
rect 12651 26144 12693 26153
rect 12651 26104 12652 26144
rect 12692 26104 12693 26144
rect 12651 26095 12693 26104
rect 12843 26144 12885 26153
rect 12843 26104 12844 26144
rect 12884 26104 12885 26144
rect 12843 26095 12885 26104
rect 13123 26144 13181 26145
rect 13123 26104 13132 26144
rect 13172 26104 13181 26144
rect 13123 26103 13181 26104
rect 13357 26137 13399 26146
rect 13357 26097 13358 26137
rect 13398 26097 13399 26137
rect 13357 26088 13399 26097
rect 13515 26144 13557 26153
rect 13515 26104 13516 26144
rect 13556 26104 13557 26144
rect 13515 26095 13557 26104
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13795 26144 13853 26145
rect 13795 26104 13804 26144
rect 13844 26104 13853 26144
rect 13795 26103 13853 26104
rect 13891 26144 13949 26145
rect 13891 26104 13900 26144
rect 13940 26104 13949 26144
rect 13891 26103 13949 26104
rect 14275 26144 14333 26145
rect 14275 26104 14284 26144
rect 14324 26104 14333 26144
rect 14275 26103 14333 26104
rect 14371 26144 14429 26145
rect 14371 26104 14380 26144
rect 14420 26104 14429 26144
rect 14371 26103 14429 26104
rect 14571 26144 14613 26153
rect 14571 26104 14572 26144
rect 14612 26104 14613 26144
rect 14571 26095 14613 26104
rect 14667 26144 14709 26153
rect 14667 26104 14668 26144
rect 14708 26104 14709 26144
rect 14667 26095 14709 26104
rect 14760 26144 14818 26145
rect 14760 26104 14769 26144
rect 14809 26104 14818 26144
rect 14760 26103 14818 26104
rect 15051 26144 15093 26153
rect 15051 26104 15052 26144
rect 15092 26104 15093 26144
rect 15051 26095 15093 26104
rect 15235 26144 15293 26145
rect 15235 26104 15244 26144
rect 15284 26104 15293 26144
rect 15235 26103 15293 26104
rect 15435 26144 15477 26153
rect 15435 26104 15436 26144
rect 15476 26104 15477 26144
rect 15435 26095 15477 26104
rect 15627 26144 15669 26153
rect 15627 26104 15628 26144
rect 15668 26104 15669 26144
rect 15627 26095 15669 26104
rect 15915 26144 15957 26153
rect 15915 26104 15916 26144
rect 15956 26104 15957 26144
rect 15915 26095 15957 26104
rect 16011 26144 16053 26153
rect 16011 26104 16012 26144
rect 16052 26104 16053 26144
rect 16011 26095 16053 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16107 26095 16149 26104
rect 16203 26144 16245 26153
rect 16203 26104 16204 26144
rect 16244 26104 16245 26144
rect 16203 26095 16245 26104
rect 16395 26144 16437 26153
rect 16395 26104 16396 26144
rect 16436 26104 16437 26144
rect 16395 26095 16437 26104
rect 16587 26144 16629 26153
rect 16587 26104 16588 26144
rect 16628 26104 16629 26144
rect 16587 26095 16629 26104
rect 16675 26144 16733 26145
rect 16675 26104 16684 26144
rect 16724 26104 16733 26144
rect 16675 26103 16733 26104
rect 17259 26144 17301 26153
rect 17259 26104 17260 26144
rect 17300 26104 17301 26144
rect 17259 26095 17301 26104
rect 17539 26144 17597 26145
rect 17539 26104 17548 26144
rect 17588 26104 17597 26144
rect 17539 26103 17597 26104
rect 18115 26144 18173 26145
rect 18115 26104 18124 26144
rect 18164 26104 18173 26144
rect 18115 26103 18173 26104
rect 18219 26144 18261 26153
rect 18219 26104 18220 26144
rect 18260 26104 18261 26144
rect 18219 26095 18261 26104
rect 18411 26144 18453 26153
rect 18411 26104 18412 26144
rect 18452 26104 18453 26144
rect 18411 26095 18453 26104
rect 18699 26144 18741 26153
rect 18699 26104 18700 26144
rect 18740 26104 18741 26144
rect 18699 26095 18741 26104
rect 18795 26144 18837 26153
rect 18795 26104 18796 26144
rect 18836 26104 18837 26144
rect 18795 26095 18837 26104
rect 18891 26144 18933 26153
rect 18891 26104 18892 26144
rect 18932 26104 18933 26144
rect 18891 26095 18933 26104
rect 18987 26144 19029 26153
rect 18987 26104 18988 26144
rect 19028 26104 19029 26144
rect 18987 26095 19029 26104
rect 19179 26144 19221 26153
rect 19179 26104 19180 26144
rect 19220 26104 19221 26144
rect 19179 26095 19221 26104
rect 19275 26144 19317 26153
rect 19275 26104 19276 26144
rect 19316 26104 19317 26144
rect 19275 26095 19317 26104
rect 19467 26144 19509 26153
rect 19467 26104 19468 26144
rect 19508 26104 19509 26144
rect 19363 26102 19421 26103
rect 3907 26061 3965 26062
rect 9667 26060 9725 26061
rect 9667 26020 9676 26060
rect 9716 26020 9725 26060
rect 9667 26019 9725 26020
rect 11019 26060 11061 26069
rect 19363 26062 19372 26102
rect 19412 26062 19421 26102
rect 19467 26095 19509 26104
rect 19651 26144 19709 26145
rect 19651 26104 19660 26144
rect 19700 26104 19709 26144
rect 19651 26103 19709 26104
rect 20515 26144 20573 26145
rect 20515 26104 20524 26144
rect 20564 26104 20573 26144
rect 20515 26103 20573 26104
rect 20907 26144 20949 26153
rect 20907 26104 20908 26144
rect 20948 26104 20949 26144
rect 20907 26095 20949 26104
rect 22051 26144 22109 26145
rect 22051 26104 22060 26144
rect 22100 26104 22109 26144
rect 22051 26103 22109 26104
rect 22915 26144 22973 26145
rect 22915 26104 22924 26144
rect 22964 26104 22973 26144
rect 22915 26103 22973 26104
rect 23307 26144 23349 26153
rect 23307 26104 23308 26144
rect 23348 26104 23349 26144
rect 23307 26095 23349 26104
rect 23691 26144 23733 26153
rect 23691 26104 23692 26144
rect 23732 26104 23733 26144
rect 23691 26095 23733 26104
rect 23787 26144 23829 26153
rect 23787 26104 23788 26144
rect 23828 26104 23829 26144
rect 23787 26095 23829 26104
rect 23883 26144 23925 26153
rect 23883 26104 23884 26144
rect 23924 26104 23925 26144
rect 23883 26095 23925 26104
rect 23979 26144 24021 26153
rect 23979 26104 23980 26144
rect 24020 26104 24021 26144
rect 23979 26095 24021 26104
rect 25123 26144 25181 26145
rect 25123 26104 25132 26144
rect 25172 26104 25181 26144
rect 25123 26103 25181 26104
rect 25795 26144 25853 26145
rect 25795 26104 25804 26144
rect 25844 26104 25853 26144
rect 25795 26103 25853 26104
rect 25899 26139 25941 26148
rect 25899 26099 25900 26139
rect 25940 26099 25941 26139
rect 25987 26144 26045 26145
rect 25987 26104 25996 26144
rect 26036 26104 26045 26144
rect 25987 26103 26045 26104
rect 26947 26144 27005 26145
rect 26947 26104 26956 26144
rect 26996 26104 27005 26144
rect 26947 26103 27005 26104
rect 27523 26144 27581 26145
rect 27523 26104 27532 26144
rect 27572 26104 27581 26144
rect 27523 26103 27581 26104
rect 27627 26139 27669 26148
rect 25899 26090 25941 26099
rect 27627 26099 27628 26139
rect 27668 26099 27669 26139
rect 27715 26144 27773 26145
rect 27715 26104 27724 26144
rect 27764 26104 27773 26144
rect 27715 26103 27773 26104
rect 28387 26144 28445 26145
rect 28387 26104 28396 26144
rect 28436 26104 28445 26144
rect 28387 26103 28445 26104
rect 29347 26144 29405 26145
rect 29347 26104 29356 26144
rect 29396 26104 29405 26144
rect 29347 26103 29405 26104
rect 29547 26144 29589 26153
rect 29547 26104 29548 26144
rect 29588 26104 29589 26144
rect 27627 26090 27669 26099
rect 29547 26095 29589 26104
rect 29739 26144 29781 26153
rect 29739 26104 29740 26144
rect 29780 26104 29781 26144
rect 29739 26095 29781 26104
rect 29827 26144 29885 26145
rect 29827 26104 29836 26144
rect 29876 26104 29885 26144
rect 29827 26103 29885 26104
rect 30883 26144 30941 26145
rect 30883 26104 30892 26144
rect 30932 26104 30941 26144
rect 31075 26144 31133 26145
rect 30883 26103 30941 26104
rect 30987 26109 31029 26118
rect 30987 26069 30988 26109
rect 31028 26069 31029 26109
rect 31075 26104 31084 26144
rect 31124 26104 31133 26144
rect 31075 26103 31133 26104
rect 32139 26144 32181 26153
rect 32139 26104 32140 26144
rect 32180 26104 32181 26144
rect 32139 26095 32181 26104
rect 33667 26144 33725 26145
rect 33667 26104 33676 26144
rect 33716 26104 33725 26144
rect 33859 26119 33868 26159
rect 33908 26119 33917 26159
rect 33859 26118 33917 26119
rect 33963 26144 34005 26153
rect 33667 26103 33725 26104
rect 33963 26104 33964 26144
rect 34004 26104 34005 26144
rect 33963 26095 34005 26104
rect 34155 26144 34197 26153
rect 34155 26104 34156 26144
rect 34196 26104 34197 26144
rect 34155 26095 34197 26104
rect 35971 26144 36029 26145
rect 35971 26104 35980 26144
rect 36020 26104 36029 26144
rect 35971 26103 36029 26104
rect 39339 26139 39381 26148
rect 39339 26099 39340 26139
rect 39380 26099 39381 26139
rect 39811 26144 39869 26145
rect 39811 26104 39820 26144
rect 39860 26104 39869 26144
rect 39811 26103 39869 26104
rect 40299 26144 40341 26153
rect 40299 26104 40300 26144
rect 40340 26104 40341 26144
rect 39339 26090 39381 26099
rect 40299 26095 40341 26104
rect 40395 26144 40437 26153
rect 40395 26104 40396 26144
rect 40436 26104 40437 26144
rect 40395 26095 40437 26104
rect 40779 26144 40821 26153
rect 40779 26104 40780 26144
rect 40820 26104 40821 26144
rect 40779 26095 40821 26104
rect 40875 26144 40917 26153
rect 40875 26104 40876 26144
rect 40916 26104 40917 26144
rect 40875 26095 40917 26104
rect 42219 26144 42261 26153
rect 42219 26104 42220 26144
rect 42260 26104 42261 26144
rect 42219 26095 42261 26104
rect 42315 26144 42357 26153
rect 42315 26104 42316 26144
rect 42356 26104 42357 26144
rect 42315 26095 42357 26104
rect 42411 26144 42453 26153
rect 42411 26104 42412 26144
rect 42452 26104 42453 26144
rect 42411 26095 42453 26104
rect 42507 26144 42549 26153
rect 42507 26104 42508 26144
rect 42548 26104 42549 26144
rect 42507 26095 42549 26104
rect 42795 26144 42837 26153
rect 42795 26104 42796 26144
rect 42836 26104 42837 26144
rect 42795 26095 42837 26104
rect 42883 26144 42941 26145
rect 42883 26104 42892 26144
rect 42932 26104 42941 26144
rect 42883 26103 42941 26104
rect 43075 26144 43133 26145
rect 43075 26104 43084 26144
rect 43124 26104 43133 26144
rect 43075 26103 43133 26104
rect 43179 26144 43221 26153
rect 43179 26104 43180 26144
rect 43220 26104 43221 26144
rect 43179 26095 43221 26104
rect 43371 26144 43413 26153
rect 43371 26104 43372 26144
rect 43412 26104 43413 26144
rect 43371 26095 43413 26104
rect 43659 26144 43701 26153
rect 43659 26104 43660 26144
rect 43700 26104 43701 26144
rect 43659 26095 43701 26104
rect 43755 26144 43797 26153
rect 43755 26104 43756 26144
rect 43796 26104 43797 26144
rect 43755 26095 43797 26104
rect 43851 26144 43893 26153
rect 43851 26104 43852 26144
rect 43892 26104 43893 26144
rect 43851 26095 43893 26104
rect 44331 26144 44373 26153
rect 44331 26104 44332 26144
rect 44372 26104 44373 26144
rect 44331 26095 44373 26104
rect 44427 26144 44469 26153
rect 44427 26104 44428 26144
rect 44468 26104 44469 26144
rect 44427 26095 44469 26104
rect 44523 26144 44565 26153
rect 44523 26104 44524 26144
rect 44564 26104 44565 26144
rect 44523 26095 44565 26104
rect 44715 26144 44757 26153
rect 44715 26104 44716 26144
rect 44756 26104 44757 26144
rect 44715 26095 44757 26104
rect 44899 26144 44957 26145
rect 44899 26104 44908 26144
rect 44948 26104 44957 26144
rect 44899 26103 44957 26104
rect 46051 26144 46109 26145
rect 46051 26104 46060 26144
rect 46100 26104 46109 26144
rect 46051 26103 46109 26104
rect 46155 26144 46197 26153
rect 46155 26104 46156 26144
rect 46196 26104 46197 26144
rect 46155 26095 46197 26104
rect 46347 26144 46389 26153
rect 46347 26104 46348 26144
rect 46388 26104 46389 26144
rect 46347 26095 46389 26104
rect 47203 26144 47261 26145
rect 47203 26104 47212 26144
rect 47252 26104 47261 26144
rect 47203 26103 47261 26104
rect 47403 26144 47445 26153
rect 47403 26104 47404 26144
rect 47444 26104 47445 26144
rect 47403 26095 47445 26104
rect 47499 26144 47541 26153
rect 47499 26104 47500 26144
rect 47540 26104 47541 26144
rect 47499 26095 47541 26104
rect 47595 26144 47637 26153
rect 47595 26104 47596 26144
rect 47636 26104 47637 26144
rect 47595 26095 47637 26104
rect 47691 26144 47733 26153
rect 47691 26104 47692 26144
rect 47732 26104 47733 26144
rect 47691 26095 47733 26104
rect 47883 26144 47925 26153
rect 47883 26104 47884 26144
rect 47924 26104 47925 26144
rect 47883 26095 47925 26104
rect 48075 26144 48117 26153
rect 48075 26104 48076 26144
rect 48116 26104 48117 26144
rect 48075 26095 48117 26104
rect 48163 26144 48221 26145
rect 48163 26104 48172 26144
rect 48212 26104 48221 26144
rect 48163 26103 48221 26104
rect 48931 26144 48989 26145
rect 48931 26104 48940 26144
rect 48980 26104 48989 26144
rect 48931 26103 48989 26104
rect 49891 26144 49949 26145
rect 49891 26104 49900 26144
rect 49940 26104 49949 26144
rect 49891 26103 49949 26104
rect 50755 26144 50813 26145
rect 50755 26104 50764 26144
rect 50804 26104 50813 26144
rect 50755 26103 50813 26104
rect 50955 26144 50997 26153
rect 50955 26104 50956 26144
rect 50996 26104 50997 26144
rect 50955 26095 50997 26104
rect 51619 26144 51677 26145
rect 51619 26104 51628 26144
rect 51668 26104 51677 26144
rect 51619 26103 51677 26104
rect 19363 26061 19421 26062
rect 11019 26020 11020 26060
rect 11060 26020 11061 26060
rect 11019 26011 11061 26020
rect 24267 26060 24309 26069
rect 30987 26060 31029 26069
rect 45859 26060 45917 26061
rect 24267 26020 24268 26060
rect 24308 26020 24309 26060
rect 24267 26011 24309 26020
rect 45859 26020 45868 26060
rect 45908 26020 45917 26060
rect 45859 26019 45917 26020
rect 1035 25976 1077 25985
rect 1035 25936 1036 25976
rect 1076 25936 1077 25976
rect 1035 25927 1077 25936
rect 5259 25976 5301 25985
rect 5259 25936 5260 25976
rect 5300 25936 5301 25976
rect 5259 25927 5301 25936
rect 5643 25976 5685 25985
rect 5643 25936 5644 25976
rect 5684 25936 5685 25976
rect 5643 25927 5685 25936
rect 6411 25976 6453 25985
rect 6411 25936 6412 25976
rect 6452 25936 6453 25976
rect 6411 25927 6453 25936
rect 8907 25976 8949 25985
rect 8907 25936 8908 25976
rect 8948 25936 8949 25976
rect 8907 25927 8949 25936
rect 12843 25976 12885 25985
rect 12843 25936 12844 25976
rect 12884 25936 12885 25976
rect 12843 25927 12885 25936
rect 16867 25976 16925 25977
rect 16867 25936 16876 25976
rect 16916 25936 16925 25976
rect 16867 25935 16925 25936
rect 18411 25976 18453 25985
rect 18411 25936 18412 25976
rect 18452 25936 18453 25976
rect 18411 25927 18453 25936
rect 29067 25976 29109 25985
rect 29067 25936 29068 25976
rect 29108 25936 29109 25976
rect 29067 25927 29109 25936
rect 34155 25976 34197 25985
rect 34155 25936 34156 25976
rect 34196 25936 34197 25976
rect 34155 25927 34197 25936
rect 36843 25976 36885 25985
rect 36843 25936 36844 25976
rect 36884 25936 36885 25976
rect 36843 25927 36885 25936
rect 44811 25976 44853 25985
rect 44811 25936 44812 25976
rect 44852 25936 44853 25976
rect 44811 25927 44853 25936
rect 45291 25976 45333 25985
rect 45291 25936 45292 25976
rect 45332 25936 45333 25976
rect 45291 25927 45333 25936
rect 48747 25976 48789 25985
rect 48747 25936 48748 25976
rect 48788 25936 48789 25976
rect 48747 25927 48789 25936
rect 8131 25892 8189 25893
rect 8131 25852 8140 25892
rect 8180 25852 8189 25892
rect 8131 25851 8189 25852
rect 10051 25892 10109 25893
rect 10051 25852 10060 25892
rect 10100 25852 10109 25892
rect 10051 25851 10109 25852
rect 13035 25892 13077 25901
rect 13035 25852 13036 25892
rect 13076 25852 13077 25892
rect 13035 25843 13077 25852
rect 13899 25892 13941 25901
rect 13899 25852 13900 25892
rect 13940 25852 13941 25892
rect 13899 25843 13941 25852
rect 14283 25892 14325 25901
rect 14283 25852 14284 25892
rect 14324 25852 14325 25892
rect 14283 25843 14325 25852
rect 15435 25892 15477 25901
rect 15435 25852 15436 25892
rect 15476 25852 15477 25892
rect 15435 25843 15477 25852
rect 16395 25892 16437 25901
rect 16395 25852 16396 25892
rect 16436 25852 16437 25892
rect 16395 25843 16437 25852
rect 20323 25892 20381 25893
rect 20323 25852 20332 25892
rect 20372 25852 20381 25892
rect 20323 25851 20381 25852
rect 25515 25892 25557 25901
rect 25515 25852 25516 25892
rect 25556 25852 25557 25892
rect 25515 25843 25557 25852
rect 26275 25892 26333 25893
rect 26275 25852 26284 25892
rect 26324 25852 26333 25892
rect 26275 25851 26333 25852
rect 27243 25892 27285 25901
rect 27243 25852 27244 25892
rect 27284 25852 27285 25892
rect 27243 25843 27285 25852
rect 30603 25892 30645 25901
rect 30603 25852 30604 25892
rect 30644 25852 30645 25892
rect 30603 25843 30645 25852
rect 33579 25892 33621 25901
rect 33579 25852 33580 25892
rect 33620 25852 33621 25892
rect 33579 25843 33621 25852
rect 36643 25892 36701 25893
rect 36643 25852 36652 25892
rect 36692 25852 36701 25892
rect 36643 25851 36701 25852
rect 43371 25892 43413 25901
rect 43371 25852 43372 25892
rect 43412 25852 43413 25892
rect 43371 25843 43413 25852
rect 46347 25892 46389 25901
rect 46347 25852 46348 25892
rect 46388 25852 46389 25892
rect 46347 25843 46389 25852
rect 46531 25892 46589 25893
rect 46531 25852 46540 25892
rect 46580 25852 46589 25892
rect 46531 25851 46589 25852
rect 47883 25892 47925 25901
rect 47883 25852 47884 25892
rect 47924 25852 47925 25892
rect 47883 25843 47925 25852
rect 49603 25892 49661 25893
rect 49603 25852 49612 25892
rect 49652 25852 49661 25892
rect 49603 25851 49661 25852
rect 50083 25892 50141 25893
rect 50083 25852 50092 25892
rect 50132 25852 50141 25892
rect 50083 25851 50141 25852
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 11491 25556 11549 25557
rect 11491 25516 11500 25556
rect 11540 25516 11549 25556
rect 11491 25515 11549 25516
rect 13131 25556 13173 25565
rect 13131 25516 13132 25556
rect 13172 25516 13173 25556
rect 13131 25507 13173 25516
rect 15051 25556 15093 25565
rect 15051 25516 15052 25556
rect 15092 25516 15093 25556
rect 15051 25507 15093 25516
rect 17451 25556 17493 25565
rect 17451 25516 17452 25556
rect 17492 25516 17493 25556
rect 17451 25507 17493 25516
rect 17931 25556 17973 25565
rect 17931 25516 17932 25556
rect 17972 25516 17973 25556
rect 17931 25507 17973 25516
rect 19363 25556 19421 25557
rect 19363 25516 19372 25556
rect 19412 25516 19421 25556
rect 19363 25515 19421 25516
rect 24555 25556 24597 25565
rect 24555 25516 24556 25556
rect 24596 25516 24597 25556
rect 24555 25507 24597 25516
rect 31659 25556 31701 25565
rect 31659 25516 31660 25556
rect 31700 25516 31701 25556
rect 31659 25507 31701 25516
rect 39627 25556 39669 25565
rect 39627 25516 39628 25556
rect 39668 25516 39669 25556
rect 39627 25507 39669 25516
rect 41251 25556 41309 25557
rect 41251 25516 41260 25556
rect 41300 25516 41309 25556
rect 41251 25515 41309 25516
rect 42411 25556 42453 25565
rect 42411 25516 42412 25556
rect 42452 25516 42453 25556
rect 42411 25507 42453 25516
rect 47203 25556 47261 25557
rect 47203 25516 47212 25556
rect 47252 25516 47261 25556
rect 47203 25515 47261 25516
rect 51139 25556 51197 25557
rect 51139 25516 51148 25556
rect 51188 25516 51197 25556
rect 51139 25515 51197 25516
rect 1611 25472 1653 25481
rect 1611 25432 1612 25472
rect 1652 25432 1653 25472
rect 1611 25423 1653 25432
rect 6699 25472 6741 25481
rect 6699 25432 6700 25472
rect 6740 25432 6741 25472
rect 6699 25423 6741 25432
rect 27531 25472 27573 25481
rect 27531 25432 27532 25472
rect 27572 25432 27573 25472
rect 27531 25423 27573 25432
rect 28203 25472 28245 25481
rect 28203 25432 28204 25472
rect 28244 25432 28245 25472
rect 28203 25423 28245 25432
rect 29835 25472 29877 25481
rect 29835 25432 29836 25472
rect 29876 25432 29877 25472
rect 29835 25423 29877 25432
rect 32523 25472 32565 25481
rect 32523 25432 32524 25472
rect 32564 25432 32565 25472
rect 32523 25423 32565 25432
rect 33003 25472 33045 25481
rect 33003 25432 33004 25472
rect 33044 25432 33045 25472
rect 33003 25423 33045 25432
rect 44331 25472 44373 25481
rect 44331 25432 44332 25472
rect 44372 25432 44373 25472
rect 44331 25423 44373 25432
rect 22731 25388 22773 25397
rect 22731 25348 22732 25388
rect 22772 25348 22773 25388
rect 22731 25339 22773 25348
rect 38475 25388 38517 25397
rect 38475 25348 38476 25388
rect 38516 25348 38517 25388
rect 38475 25339 38517 25348
rect 3435 25304 3477 25313
rect 3435 25264 3436 25304
rect 3476 25264 3477 25304
rect 3435 25255 3477 25264
rect 3531 25304 3573 25313
rect 3531 25264 3532 25304
rect 3572 25264 3573 25304
rect 3531 25255 3573 25264
rect 3627 25304 3669 25313
rect 3627 25264 3628 25304
rect 3668 25264 3669 25304
rect 3627 25255 3669 25264
rect 3819 25304 3861 25313
rect 3819 25264 3820 25304
rect 3860 25264 3861 25304
rect 3819 25255 3861 25264
rect 3915 25304 3957 25313
rect 3915 25264 3916 25304
rect 3956 25264 3957 25304
rect 3915 25255 3957 25264
rect 4011 25304 4053 25313
rect 4011 25264 4012 25304
rect 4052 25264 4053 25304
rect 4011 25255 4053 25264
rect 4107 25304 4149 25313
rect 4107 25264 4108 25304
rect 4148 25264 4149 25304
rect 4107 25255 4149 25264
rect 4291 25304 4349 25305
rect 4291 25264 4300 25304
rect 4340 25264 4349 25304
rect 4291 25263 4349 25264
rect 4971 25304 5013 25313
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 4971 25255 5013 25264
rect 5827 25304 5885 25305
rect 5827 25264 5836 25304
rect 5876 25264 5885 25304
rect 5827 25263 5885 25264
rect 6979 25304 7037 25305
rect 6979 25264 6988 25304
rect 7028 25264 7037 25304
rect 6979 25263 7037 25264
rect 7843 25304 7901 25305
rect 7843 25264 7852 25304
rect 7892 25264 7901 25304
rect 7843 25263 7901 25264
rect 8715 25304 8757 25313
rect 8715 25264 8716 25304
rect 8756 25264 8757 25304
rect 8715 25255 8757 25264
rect 9099 25304 9141 25313
rect 9099 25264 9100 25304
rect 9140 25264 9141 25304
rect 9099 25255 9141 25264
rect 9475 25304 9533 25305
rect 9475 25264 9484 25304
rect 9524 25264 9533 25304
rect 9475 25263 9533 25264
rect 10339 25304 10397 25305
rect 10339 25264 10348 25304
rect 10388 25264 10397 25304
rect 10339 25263 10397 25264
rect 11683 25304 11741 25305
rect 11683 25264 11692 25304
rect 11732 25264 11741 25304
rect 11683 25263 11741 25264
rect 12939 25304 12981 25313
rect 12939 25264 12940 25304
rect 12980 25264 12981 25304
rect 12939 25255 12981 25264
rect 13795 25304 13853 25305
rect 13795 25264 13804 25304
rect 13844 25264 13853 25304
rect 13795 25263 13853 25264
rect 13995 25304 14037 25313
rect 13995 25264 13996 25304
rect 14036 25264 14037 25304
rect 13995 25255 14037 25264
rect 14091 25304 14133 25313
rect 14091 25264 14092 25304
rect 14132 25264 14133 25304
rect 14091 25255 14133 25264
rect 14187 25304 14229 25313
rect 14187 25264 14188 25304
rect 14228 25264 14229 25304
rect 14187 25255 14229 25264
rect 14283 25304 14325 25313
rect 14283 25264 14284 25304
rect 14324 25264 14325 25304
rect 14283 25255 14325 25264
rect 14659 25304 14717 25305
rect 14659 25264 14668 25304
rect 14708 25264 14717 25304
rect 14659 25263 14717 25264
rect 14763 25304 14805 25313
rect 14763 25264 14764 25304
rect 14804 25264 14805 25304
rect 14763 25255 14805 25264
rect 15235 25304 15293 25305
rect 15235 25264 15244 25304
rect 15284 25264 15293 25304
rect 15235 25263 15293 25264
rect 16107 25304 16149 25313
rect 16107 25264 16108 25304
rect 16148 25264 16149 25304
rect 16107 25255 16149 25264
rect 17155 25304 17213 25305
rect 17155 25264 17164 25304
rect 17204 25264 17213 25304
rect 17155 25263 17213 25264
rect 17259 25304 17301 25313
rect 17259 25264 17260 25304
rect 17300 25264 17301 25304
rect 17259 25255 17301 25264
rect 17451 25304 17493 25313
rect 17451 25264 17452 25304
rect 17492 25264 17493 25304
rect 17451 25255 17493 25264
rect 17635 25304 17693 25305
rect 17635 25264 17644 25304
rect 17684 25264 17693 25304
rect 17635 25263 17693 25264
rect 17739 25304 17781 25313
rect 17739 25264 17740 25304
rect 17780 25264 17781 25304
rect 17739 25255 17781 25264
rect 17931 25304 17973 25313
rect 17931 25264 17932 25304
rect 17972 25264 17973 25304
rect 17931 25255 17973 25264
rect 19171 25304 19229 25305
rect 19171 25264 19180 25304
rect 19220 25264 19229 25304
rect 19171 25263 19229 25264
rect 20515 25304 20573 25305
rect 20515 25264 20524 25304
rect 20564 25264 20573 25304
rect 20515 25263 20573 25264
rect 21379 25304 21437 25305
rect 21379 25264 21388 25304
rect 21428 25264 21437 25304
rect 21379 25263 21437 25264
rect 21771 25304 21813 25313
rect 21771 25264 21772 25304
rect 21812 25264 21813 25304
rect 21771 25255 21813 25264
rect 23587 25304 23645 25305
rect 23587 25264 23596 25304
rect 23636 25264 23645 25304
rect 23587 25263 23645 25264
rect 24835 25304 24893 25305
rect 24835 25264 24844 25304
rect 24884 25264 24893 25304
rect 24835 25263 24893 25264
rect 25131 25304 25173 25313
rect 25131 25264 25132 25304
rect 25172 25264 25173 25304
rect 25131 25255 25173 25264
rect 25507 25304 25565 25305
rect 25507 25264 25516 25304
rect 25556 25264 25565 25304
rect 25507 25263 25565 25264
rect 26371 25304 26429 25305
rect 26371 25264 26380 25304
rect 26420 25264 26429 25304
rect 26371 25263 26429 25264
rect 27907 25304 27965 25305
rect 27907 25264 27916 25304
rect 27956 25264 27965 25304
rect 27907 25263 27965 25264
rect 31171 25304 31229 25305
rect 31171 25264 31180 25304
rect 31220 25264 31229 25304
rect 31171 25263 31229 25264
rect 32707 25304 32765 25305
rect 32707 25264 32716 25304
rect 32756 25264 32765 25304
rect 32707 25263 32765 25264
rect 32811 25304 32853 25313
rect 32811 25264 32812 25304
rect 32852 25264 32853 25304
rect 32811 25255 32853 25264
rect 33003 25304 33045 25313
rect 33003 25264 33004 25304
rect 33044 25264 33045 25304
rect 33003 25255 33045 25264
rect 33859 25304 33917 25305
rect 33859 25264 33868 25304
rect 33908 25264 33917 25304
rect 33859 25263 33917 25264
rect 34059 25304 34101 25313
rect 34059 25264 34060 25304
rect 34100 25264 34101 25304
rect 34059 25255 34101 25264
rect 34155 25304 34197 25313
rect 34155 25264 34156 25304
rect 34196 25264 34197 25304
rect 34155 25255 34197 25264
rect 34251 25304 34293 25313
rect 34251 25264 34252 25304
rect 34292 25264 34293 25304
rect 34251 25255 34293 25264
rect 34347 25304 34389 25313
rect 34347 25264 34348 25304
rect 34388 25264 34389 25304
rect 34347 25255 34389 25264
rect 34731 25304 34773 25313
rect 34731 25264 34732 25304
rect 34772 25264 34773 25304
rect 34731 25255 34773 25264
rect 34827 25304 34869 25313
rect 34827 25264 34828 25304
rect 34868 25264 34869 25304
rect 34827 25255 34869 25264
rect 34923 25304 34965 25313
rect 34923 25264 34924 25304
rect 34964 25264 34965 25304
rect 34923 25255 34965 25264
rect 35203 25304 35261 25305
rect 35203 25264 35212 25304
rect 35252 25264 35261 25304
rect 35203 25263 35261 25264
rect 36075 25304 36117 25313
rect 36075 25264 36076 25304
rect 36116 25264 36117 25304
rect 36075 25255 36117 25264
rect 36451 25304 36509 25305
rect 36451 25264 36460 25304
rect 36500 25264 36509 25304
rect 36451 25263 36509 25264
rect 37315 25304 37373 25305
rect 37315 25264 37324 25304
rect 37364 25264 37373 25304
rect 39051 25304 39093 25313
rect 37315 25263 37373 25264
rect 38942 25293 38984 25302
rect 38942 25253 38943 25293
rect 38983 25253 38984 25293
rect 39051 25264 39052 25304
rect 39092 25264 39093 25304
rect 39051 25255 39093 25264
rect 39331 25304 39389 25305
rect 39331 25264 39340 25304
rect 39380 25264 39389 25304
rect 39331 25263 39389 25264
rect 40291 25304 40349 25305
rect 40291 25264 40300 25304
rect 40340 25264 40349 25304
rect 40291 25263 40349 25264
rect 40491 25304 40533 25313
rect 40491 25264 40492 25304
rect 40532 25264 40533 25304
rect 40491 25255 40533 25264
rect 40587 25304 40629 25313
rect 40587 25264 40588 25304
rect 40628 25264 40629 25304
rect 40587 25255 40629 25264
rect 41643 25304 41685 25313
rect 41643 25264 41644 25304
rect 41684 25264 41685 25304
rect 41643 25255 41685 25264
rect 41923 25304 41981 25305
rect 41923 25264 41932 25304
rect 41972 25264 41981 25304
rect 41923 25263 41981 25264
rect 42315 25304 42357 25313
rect 42315 25264 42316 25304
rect 42356 25264 42357 25304
rect 42315 25255 42357 25264
rect 42499 25304 42557 25305
rect 42499 25264 42508 25304
rect 42548 25264 42557 25304
rect 42499 25263 42557 25264
rect 43363 25304 43421 25305
rect 43363 25264 43372 25304
rect 43412 25264 43421 25304
rect 43363 25263 43421 25264
rect 43755 25304 43797 25313
rect 43755 25264 43756 25304
rect 43796 25264 43797 25304
rect 43755 25255 43797 25264
rect 43851 25304 43893 25313
rect 43851 25264 43852 25304
rect 43892 25264 43893 25304
rect 43851 25255 43893 25264
rect 43947 25304 43989 25313
rect 43947 25264 43948 25304
rect 43988 25264 43989 25304
rect 43947 25255 43989 25264
rect 44043 25304 44085 25313
rect 44043 25264 44044 25304
rect 44084 25264 44085 25304
rect 44043 25255 44085 25264
rect 44331 25304 44373 25313
rect 44331 25264 44332 25304
rect 44372 25264 44373 25304
rect 44331 25255 44373 25264
rect 44523 25304 44565 25313
rect 44523 25264 44524 25304
rect 44564 25264 44565 25304
rect 44523 25255 44565 25264
rect 44611 25304 44669 25305
rect 44611 25264 44620 25304
rect 44660 25264 44669 25304
rect 44611 25263 44669 25264
rect 44811 25304 44853 25313
rect 44811 25264 44812 25304
rect 44852 25264 44853 25304
rect 44811 25255 44853 25264
rect 45187 25304 45245 25305
rect 45187 25264 45196 25304
rect 45236 25264 45245 25304
rect 45187 25263 45245 25264
rect 46051 25304 46109 25305
rect 46051 25264 46060 25304
rect 46100 25264 46109 25304
rect 46051 25263 46109 25264
rect 47403 25304 47445 25313
rect 47403 25264 47404 25304
rect 47444 25264 47445 25304
rect 47403 25255 47445 25264
rect 47499 25304 47541 25313
rect 47499 25264 47500 25304
rect 47540 25264 47541 25304
rect 47499 25255 47541 25264
rect 47595 25304 47637 25313
rect 47595 25264 47596 25304
rect 47636 25264 47637 25304
rect 47595 25255 47637 25264
rect 47875 25304 47933 25305
rect 47875 25264 47884 25304
rect 47924 25264 47933 25304
rect 47875 25263 47933 25264
rect 49123 25304 49181 25305
rect 49123 25264 49132 25304
rect 49172 25264 49181 25304
rect 49123 25263 49181 25264
rect 49987 25304 50045 25305
rect 49987 25264 49996 25304
rect 50036 25264 50045 25304
rect 49987 25263 50045 25264
rect 38942 25244 38984 25253
rect 12363 25220 12405 25229
rect 12363 25180 12364 25220
rect 12404 25180 12405 25220
rect 12363 25171 12405 25180
rect 35019 25220 35061 25229
rect 35019 25180 35020 25220
rect 35060 25180 35061 25220
rect 35019 25171 35061 25180
rect 41547 25220 41589 25229
rect 41547 25180 41548 25220
rect 41588 25180 41589 25220
rect 41547 25171 41589 25180
rect 47691 25220 47733 25229
rect 47691 25180 47692 25220
rect 47732 25180 47733 25220
rect 47691 25171 47733 25180
rect 48555 25220 48597 25229
rect 48555 25180 48556 25220
rect 48596 25180 48597 25220
rect 48555 25171 48597 25180
rect 48747 25220 48789 25229
rect 48747 25180 48748 25220
rect 48788 25180 48789 25220
rect 48747 25171 48789 25180
rect 3331 25136 3389 25137
rect 3331 25096 3340 25136
rect 3380 25096 3389 25136
rect 3331 25095 3389 25096
rect 5155 25136 5213 25137
rect 5155 25096 5164 25136
rect 5204 25096 5213 25136
rect 5155 25095 5213 25096
rect 14571 25132 14613 25141
rect 14571 25092 14572 25132
rect 14612 25092 14613 25132
rect 14571 25083 14613 25092
rect 19083 25136 19125 25145
rect 19083 25096 19084 25136
rect 19124 25096 19125 25136
rect 19083 25087 19125 25096
rect 33187 25136 33245 25137
rect 33187 25096 33196 25136
rect 33236 25096 33245 25136
rect 33187 25095 33245 25096
rect 35875 25136 35933 25137
rect 35875 25096 35884 25136
rect 35924 25096 35933 25136
rect 35875 25095 35933 25096
rect 40771 25136 40829 25137
rect 40771 25096 40780 25136
rect 40820 25096 40829 25136
rect 40771 25095 40829 25096
rect 42691 25136 42749 25137
rect 42691 25096 42700 25136
rect 42740 25096 42749 25136
rect 42691 25095 42749 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 28107 24858 28149 24867
rect 28107 24818 28108 24858
rect 28148 24818 28149 24858
rect 28107 24809 28149 24818
rect 13315 24800 13373 24801
rect 13315 24760 13324 24800
rect 13364 24760 13373 24800
rect 13315 24759 13373 24760
rect 16195 24800 16253 24801
rect 16195 24760 16204 24800
rect 16244 24760 16253 24800
rect 16195 24759 16253 24760
rect 16867 24800 16925 24801
rect 16867 24760 16876 24800
rect 16916 24760 16925 24800
rect 16867 24759 16925 24760
rect 19075 24800 19133 24801
rect 19075 24760 19084 24800
rect 19124 24760 19133 24800
rect 19075 24759 19133 24760
rect 21571 24800 21629 24801
rect 21571 24760 21580 24800
rect 21620 24760 21629 24800
rect 21571 24759 21629 24760
rect 25803 24800 25845 24809
rect 25803 24760 25804 24800
rect 25844 24760 25845 24800
rect 25803 24751 25845 24760
rect 28387 24800 28445 24801
rect 28387 24760 28396 24800
rect 28436 24760 28445 24800
rect 28387 24759 28445 24760
rect 31747 24800 31805 24801
rect 31747 24760 31756 24800
rect 31796 24760 31805 24800
rect 31747 24759 31805 24760
rect 35203 24800 35261 24801
rect 35203 24760 35212 24800
rect 35252 24760 35261 24800
rect 35203 24759 35261 24760
rect 35683 24800 35741 24801
rect 35683 24760 35692 24800
rect 35732 24760 35741 24800
rect 35683 24759 35741 24760
rect 39819 24800 39861 24809
rect 39819 24760 39820 24800
rect 39860 24760 39861 24800
rect 39819 24751 39861 24760
rect 44131 24800 44189 24801
rect 44131 24760 44140 24800
rect 44180 24760 44189 24800
rect 44131 24759 44189 24760
rect 44611 24800 44669 24801
rect 44611 24760 44620 24800
rect 44660 24760 44669 24800
rect 44611 24759 44669 24760
rect 45475 24800 45533 24801
rect 45475 24760 45484 24800
rect 45524 24760 45533 24800
rect 45475 24759 45533 24760
rect 46339 24800 46397 24801
rect 46339 24760 46348 24800
rect 46388 24760 46397 24800
rect 46339 24759 46397 24760
rect 46531 24800 46589 24801
rect 46531 24760 46540 24800
rect 46580 24760 46589 24800
rect 46531 24759 46589 24760
rect 5067 24716 5109 24725
rect 5067 24676 5068 24716
rect 5108 24676 5109 24716
rect 5067 24667 5109 24676
rect 10347 24716 10389 24725
rect 10347 24676 10348 24716
rect 10388 24676 10389 24716
rect 10347 24667 10389 24676
rect 10827 24716 10869 24725
rect 10827 24676 10828 24716
rect 10868 24676 10869 24716
rect 10827 24667 10869 24676
rect 12651 24716 12693 24725
rect 12651 24676 12652 24716
rect 12692 24676 12693 24716
rect 12651 24667 12693 24676
rect 32811 24716 32853 24725
rect 32811 24676 32812 24716
rect 32852 24676 32853 24716
rect 32811 24667 32853 24676
rect 38475 24716 38517 24725
rect 38475 24676 38476 24716
rect 38516 24676 38517 24716
rect 38475 24667 38517 24676
rect 48939 24716 48981 24725
rect 48939 24676 48940 24716
rect 48980 24676 48981 24716
rect 48939 24667 48981 24676
rect 14379 24653 14421 24662
rect 1131 24632 1173 24641
rect 1131 24592 1132 24632
rect 1172 24592 1173 24632
rect 1131 24583 1173 24592
rect 1507 24632 1565 24633
rect 1507 24592 1516 24632
rect 1556 24592 1565 24632
rect 1507 24591 1565 24592
rect 2371 24632 2429 24633
rect 2371 24592 2380 24632
rect 2420 24592 2429 24632
rect 2371 24591 2429 24592
rect 4195 24632 4253 24633
rect 4195 24592 4204 24632
rect 4244 24592 4253 24632
rect 4195 24591 4253 24592
rect 4491 24632 4533 24641
rect 4491 24592 4492 24632
rect 4532 24592 4533 24632
rect 4491 24583 4533 24592
rect 4587 24632 4629 24641
rect 4587 24592 4588 24632
rect 4628 24592 4629 24632
rect 4587 24583 4629 24592
rect 5443 24632 5501 24633
rect 5443 24592 5452 24632
rect 5492 24592 5501 24632
rect 5443 24591 5501 24592
rect 6307 24632 6365 24633
rect 6307 24592 6316 24632
rect 6356 24592 6365 24632
rect 6307 24591 6365 24592
rect 7747 24632 7805 24633
rect 7747 24592 7756 24632
rect 7796 24592 7805 24632
rect 7747 24591 7805 24592
rect 8043 24632 8085 24641
rect 8043 24592 8044 24632
rect 8084 24592 8085 24632
rect 8043 24583 8085 24592
rect 8139 24632 8181 24641
rect 8139 24592 8140 24632
rect 8180 24592 8181 24632
rect 8139 24583 8181 24592
rect 9283 24632 9341 24633
rect 9283 24592 9292 24632
rect 9332 24592 9341 24632
rect 9283 24591 9341 24592
rect 10251 24632 10293 24641
rect 10251 24592 10252 24632
rect 10292 24592 10293 24632
rect 10251 24583 10293 24592
rect 10435 24632 10493 24633
rect 10435 24592 10444 24632
rect 10484 24592 10493 24632
rect 10435 24591 10493 24592
rect 10627 24632 10685 24633
rect 10627 24592 10636 24632
rect 10676 24592 10685 24632
rect 10627 24591 10685 24592
rect 10731 24632 10773 24641
rect 10731 24592 10732 24632
rect 10772 24592 10773 24632
rect 10731 24583 10773 24592
rect 10923 24632 10965 24641
rect 10923 24592 10924 24632
rect 10964 24592 10965 24632
rect 10923 24583 10965 24592
rect 11779 24632 11837 24633
rect 11779 24592 11788 24632
rect 11828 24592 11837 24632
rect 11779 24591 11837 24592
rect 12259 24632 12317 24633
rect 12259 24592 12268 24632
rect 12308 24592 12317 24632
rect 12259 24591 12317 24592
rect 12555 24632 12597 24641
rect 12555 24592 12556 24632
rect 12596 24592 12597 24632
rect 12555 24583 12597 24592
rect 13123 24632 13181 24633
rect 13123 24592 13132 24632
rect 13172 24592 13181 24632
rect 13123 24591 13181 24592
rect 13227 24632 13269 24641
rect 13227 24592 13228 24632
rect 13268 24592 13269 24632
rect 13227 24583 13269 24592
rect 13419 24632 13461 24641
rect 13419 24592 13420 24632
rect 13460 24592 13461 24632
rect 13419 24583 13461 24592
rect 13603 24632 13661 24633
rect 13603 24592 13612 24632
rect 13652 24592 13661 24632
rect 13603 24591 13661 24592
rect 13707 24632 13749 24641
rect 13707 24592 13708 24632
rect 13748 24592 13749 24632
rect 13707 24583 13749 24592
rect 13899 24632 13941 24641
rect 13899 24592 13900 24632
rect 13940 24592 13941 24632
rect 13899 24583 13941 24592
rect 14091 24632 14133 24641
rect 14091 24592 14092 24632
rect 14132 24592 14133 24632
rect 14091 24583 14133 24592
rect 14187 24632 14229 24641
rect 14187 24592 14188 24632
rect 14228 24592 14229 24632
rect 14187 24583 14229 24592
rect 14283 24632 14325 24641
rect 14283 24592 14284 24632
rect 14324 24592 14325 24632
rect 14379 24613 14380 24653
rect 14420 24613 14421 24653
rect 14379 24604 14421 24613
rect 14763 24632 14805 24641
rect 14283 24583 14325 24592
rect 14763 24592 14764 24632
rect 14804 24592 14805 24632
rect 14763 24583 14805 24592
rect 14859 24632 14901 24641
rect 14859 24592 14860 24632
rect 14900 24592 14901 24632
rect 14859 24583 14901 24592
rect 14955 24632 14997 24641
rect 14955 24592 14956 24632
rect 14996 24592 14997 24632
rect 14955 24583 14997 24592
rect 15051 24632 15093 24641
rect 15051 24592 15052 24632
rect 15092 24592 15093 24632
rect 15051 24583 15093 24592
rect 15243 24632 15285 24641
rect 15243 24592 15244 24632
rect 15284 24592 15285 24632
rect 15243 24583 15285 24592
rect 15531 24632 15573 24641
rect 15531 24592 15532 24632
rect 15572 24592 15573 24632
rect 15531 24583 15573 24592
rect 15723 24632 15765 24641
rect 15723 24592 15724 24632
rect 15764 24592 15765 24632
rect 15723 24583 15765 24592
rect 15819 24632 15861 24641
rect 15819 24592 15820 24632
rect 15860 24592 15861 24632
rect 15819 24583 15861 24592
rect 15915 24632 15957 24641
rect 15915 24592 15916 24632
rect 15956 24592 15957 24632
rect 15915 24583 15957 24592
rect 16011 24632 16053 24641
rect 16011 24592 16012 24632
rect 16052 24592 16053 24632
rect 16011 24583 16053 24592
rect 16299 24632 16341 24641
rect 16299 24592 16300 24632
rect 16340 24592 16341 24632
rect 16299 24583 16341 24592
rect 16395 24632 16437 24641
rect 16395 24592 16396 24632
rect 16436 24592 16437 24632
rect 16395 24583 16437 24592
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 16491 24583 16533 24592
rect 16675 24632 16733 24633
rect 16675 24592 16684 24632
rect 16724 24592 16733 24632
rect 16675 24591 16733 24592
rect 16779 24632 16821 24641
rect 16779 24592 16780 24632
rect 16820 24592 16821 24632
rect 16779 24583 16821 24592
rect 16971 24632 17013 24641
rect 16971 24592 16972 24632
rect 17012 24592 17013 24632
rect 16971 24583 17013 24592
rect 17451 24632 17493 24641
rect 17451 24592 17452 24632
rect 17492 24592 17493 24632
rect 17451 24583 17493 24592
rect 17547 24632 17589 24641
rect 17547 24592 17548 24632
rect 17588 24592 17589 24632
rect 17547 24583 17589 24592
rect 17827 24632 17885 24633
rect 17827 24592 17836 24632
rect 17876 24592 17885 24632
rect 17827 24591 17885 24592
rect 18603 24632 18645 24641
rect 18603 24592 18604 24632
rect 18644 24592 18645 24632
rect 18603 24583 18645 24592
rect 18795 24632 18837 24641
rect 18795 24592 18796 24632
rect 18836 24592 18837 24632
rect 18795 24583 18837 24592
rect 18883 24632 18941 24633
rect 18883 24592 18892 24632
rect 18932 24592 18941 24632
rect 18883 24591 18941 24592
rect 19747 24632 19805 24633
rect 19747 24592 19756 24632
rect 19796 24592 19805 24632
rect 19747 24591 19805 24592
rect 19939 24632 19997 24633
rect 19939 24592 19948 24632
rect 19988 24592 19997 24632
rect 19939 24591 19997 24592
rect 22243 24632 22301 24633
rect 22243 24592 22252 24632
rect 22292 24592 22301 24632
rect 22243 24591 22301 24592
rect 22435 24632 22493 24633
rect 22435 24592 22444 24632
rect 22484 24592 22493 24632
rect 22435 24591 22493 24592
rect 23307 24632 23349 24641
rect 23307 24592 23308 24632
rect 23348 24592 23349 24632
rect 23307 24583 23349 24592
rect 25707 24632 25749 24641
rect 25707 24592 25708 24632
rect 25748 24592 25749 24632
rect 25707 24583 25749 24592
rect 25899 24632 25941 24641
rect 25899 24592 25900 24632
rect 25940 24592 25941 24632
rect 25899 24583 25941 24592
rect 27915 24632 27957 24641
rect 27915 24592 27916 24632
rect 27956 24592 27957 24632
rect 27915 24583 27957 24592
rect 28003 24632 28061 24633
rect 28003 24592 28012 24632
rect 28052 24592 28061 24632
rect 28003 24591 28061 24592
rect 28299 24632 28341 24641
rect 28299 24592 28300 24632
rect 28340 24592 28341 24632
rect 28299 24583 28341 24592
rect 28491 24632 28533 24641
rect 28491 24592 28492 24632
rect 28532 24592 28533 24632
rect 28491 24583 28533 24592
rect 28579 24632 28637 24633
rect 28579 24592 28588 24632
rect 28628 24592 28637 24632
rect 28579 24591 28637 24592
rect 29355 24632 29397 24641
rect 29355 24592 29356 24632
rect 29396 24592 29397 24632
rect 29355 24583 29397 24592
rect 29731 24632 29789 24633
rect 29731 24592 29740 24632
rect 29780 24592 29789 24632
rect 29731 24591 29789 24592
rect 30595 24632 30653 24633
rect 30595 24592 30604 24632
rect 30644 24592 30653 24632
rect 30595 24591 30653 24592
rect 33187 24632 33245 24633
rect 33187 24592 33196 24632
rect 33236 24592 33245 24632
rect 33187 24591 33245 24592
rect 34051 24632 34109 24633
rect 34051 24592 34060 24632
rect 34100 24592 34109 24632
rect 34051 24591 34109 24592
rect 35595 24632 35637 24641
rect 35595 24592 35596 24632
rect 35636 24592 35637 24632
rect 35595 24583 35637 24592
rect 35787 24632 35829 24641
rect 35787 24592 35788 24632
rect 35828 24592 35829 24632
rect 35787 24583 35829 24592
rect 35875 24632 35933 24633
rect 35875 24592 35884 24632
rect 35924 24592 35933 24632
rect 35875 24591 35933 24592
rect 36067 24632 36125 24633
rect 36067 24592 36076 24632
rect 36116 24592 36125 24632
rect 36067 24591 36125 24592
rect 36747 24632 36789 24641
rect 36747 24592 36748 24632
rect 36788 24592 36789 24632
rect 36747 24583 36789 24592
rect 36843 24632 36885 24641
rect 36843 24592 36844 24632
rect 36884 24592 36885 24632
rect 36843 24583 36885 24592
rect 37795 24632 37853 24633
rect 37795 24592 37804 24632
rect 37844 24592 37853 24632
rect 37795 24591 37853 24592
rect 38283 24627 38325 24636
rect 38283 24587 38284 24627
rect 38324 24587 38325 24627
rect 38283 24578 38325 24587
rect 40011 24627 40053 24636
rect 40011 24587 40012 24627
rect 40052 24587 40053 24627
rect 40483 24632 40541 24633
rect 40483 24592 40492 24632
rect 40532 24592 40541 24632
rect 40483 24591 40541 24592
rect 41451 24632 41493 24641
rect 41451 24592 41452 24632
rect 41492 24592 41493 24632
rect 40011 24578 40053 24587
rect 41451 24583 41493 24592
rect 41547 24632 41589 24641
rect 41547 24592 41548 24632
rect 41588 24592 41589 24632
rect 41547 24583 41589 24592
rect 43371 24632 43413 24641
rect 43371 24592 43372 24632
rect 43412 24592 43413 24632
rect 43371 24583 43413 24592
rect 43851 24632 43893 24641
rect 43851 24592 43852 24632
rect 43892 24592 43893 24632
rect 43851 24583 43893 24592
rect 43947 24632 43989 24641
rect 43947 24592 43948 24632
rect 43988 24592 43989 24632
rect 43947 24583 43989 24592
rect 44043 24632 44085 24641
rect 44043 24592 44044 24632
rect 44084 24592 44085 24632
rect 44043 24583 44085 24592
rect 44331 24632 44373 24641
rect 44331 24592 44332 24632
rect 44372 24592 44373 24632
rect 44331 24583 44373 24592
rect 44427 24632 44469 24641
rect 44427 24592 44428 24632
rect 44468 24592 44469 24632
rect 44427 24583 44469 24592
rect 44523 24632 44565 24641
rect 44523 24592 44524 24632
rect 44564 24592 44565 24632
rect 44523 24583 44565 24592
rect 44803 24632 44861 24633
rect 44803 24592 44812 24632
rect 44852 24592 44861 24632
rect 44803 24591 44861 24592
rect 45667 24632 45725 24633
rect 45667 24592 45676 24632
rect 45716 24592 45725 24632
rect 45667 24591 45725 24592
rect 47203 24632 47261 24633
rect 47203 24592 47212 24632
rect 47252 24592 47261 24632
rect 47203 24591 47261 24592
rect 47403 24632 47445 24641
rect 47403 24592 47404 24632
rect 47444 24592 47445 24632
rect 47403 24583 47445 24592
rect 47499 24632 47541 24641
rect 47499 24592 47500 24632
rect 47540 24592 47541 24632
rect 47499 24583 47541 24592
rect 47595 24632 47637 24641
rect 47595 24592 47596 24632
rect 47636 24592 47637 24632
rect 47595 24583 47637 24592
rect 47691 24632 47733 24641
rect 47691 24592 47692 24632
rect 47732 24592 47733 24632
rect 47691 24583 47733 24592
rect 47979 24632 48021 24641
rect 47979 24592 47980 24632
rect 48020 24592 48021 24632
rect 47979 24583 48021 24592
rect 48171 24632 48213 24641
rect 48171 24592 48172 24632
rect 48212 24592 48213 24632
rect 48171 24583 48213 24592
rect 48259 24632 48317 24633
rect 48259 24592 48268 24632
rect 48308 24592 48317 24632
rect 48259 24591 48317 24592
rect 48459 24632 48501 24641
rect 48459 24592 48460 24632
rect 48500 24592 48501 24632
rect 48459 24583 48501 24592
rect 48651 24632 48693 24641
rect 48651 24592 48652 24632
rect 48692 24592 48693 24632
rect 48651 24583 48693 24592
rect 48739 24632 48797 24633
rect 48739 24592 48748 24632
rect 48788 24592 48797 24632
rect 48739 24591 48797 24592
rect 49027 24632 49085 24633
rect 49027 24592 49036 24632
rect 49076 24592 49085 24632
rect 49027 24591 49085 24592
rect 49419 24632 49461 24641
rect 49419 24592 49420 24632
rect 49460 24592 49461 24632
rect 49419 24583 49461 24592
rect 49795 24632 49853 24633
rect 49795 24592 49804 24632
rect 49844 24592 49853 24632
rect 49795 24591 49853 24592
rect 50659 24632 50717 24633
rect 50659 24592 50668 24632
rect 50708 24592 50717 24632
rect 50659 24591 50717 24592
rect 51819 24632 51861 24641
rect 51819 24592 51820 24632
rect 51860 24592 51861 24632
rect 51819 24583 51861 24592
rect 3531 24548 3573 24557
rect 3531 24508 3532 24548
rect 3572 24508 3573 24548
rect 3531 24499 3573 24508
rect 36171 24548 36213 24557
rect 36171 24508 36172 24548
rect 36212 24508 36213 24548
rect 36171 24499 36213 24508
rect 37227 24548 37269 24557
rect 37227 24508 37228 24548
rect 37268 24508 37269 24548
rect 37227 24499 37269 24508
rect 37323 24548 37365 24557
rect 37323 24508 37324 24548
rect 37364 24508 37365 24548
rect 37323 24499 37365 24508
rect 40971 24548 41013 24557
rect 40971 24508 40972 24548
rect 41012 24508 41013 24548
rect 40971 24499 41013 24508
rect 41067 24548 41109 24557
rect 41067 24508 41068 24548
rect 41108 24508 41109 24548
rect 41067 24499 41109 24508
rect 8419 24464 8477 24465
rect 8419 24424 8428 24464
rect 8468 24424 8477 24464
rect 8419 24423 8477 24424
rect 10059 24464 10101 24473
rect 10059 24424 10060 24464
rect 10100 24424 10101 24464
rect 10059 24415 10101 24424
rect 15531 24464 15573 24473
rect 15531 24424 15532 24464
rect 15572 24424 15573 24464
rect 15531 24415 15573 24424
rect 17155 24464 17213 24465
rect 17155 24424 17164 24464
rect 17204 24424 17213 24464
rect 17155 24423 17213 24424
rect 18603 24464 18645 24473
rect 18603 24424 18604 24464
rect 18644 24424 18645 24464
rect 18603 24415 18645 24424
rect 20811 24464 20853 24473
rect 20811 24424 20812 24464
rect 20852 24424 20853 24464
rect 20811 24415 20853 24424
rect 21387 24464 21429 24473
rect 21387 24424 21388 24464
rect 21428 24424 21429 24464
rect 21387 24415 21429 24424
rect 27627 24464 27669 24473
rect 27627 24424 27628 24464
rect 27668 24424 27669 24464
rect 27627 24415 27669 24424
rect 38859 24464 38901 24473
rect 38859 24424 38860 24464
rect 38900 24424 38901 24464
rect 38859 24415 38901 24424
rect 42315 24464 42357 24473
rect 42315 24424 42316 24464
rect 42356 24424 42357 24464
rect 42315 24415 42357 24424
rect 48459 24464 48501 24473
rect 48459 24424 48460 24464
rect 48500 24424 48501 24464
rect 48459 24415 48501 24424
rect 4867 24380 4925 24381
rect 4867 24340 4876 24380
rect 4916 24340 4925 24380
rect 4867 24339 4925 24340
rect 7459 24380 7517 24381
rect 7459 24340 7468 24380
rect 7508 24340 7517 24380
rect 7459 24339 7517 24340
rect 8611 24380 8669 24381
rect 8611 24340 8620 24380
rect 8660 24340 8669 24380
rect 8611 24339 8669 24340
rect 11107 24380 11165 24381
rect 11107 24340 11116 24380
rect 11156 24340 11165 24380
rect 11107 24339 11165 24340
rect 12931 24380 12989 24381
rect 12931 24340 12940 24380
rect 12980 24340 12989 24380
rect 12931 24339 12989 24340
rect 13899 24380 13941 24389
rect 13899 24340 13900 24380
rect 13940 24340 13941 24380
rect 13899 24331 13941 24340
rect 20611 24380 20669 24381
rect 20611 24340 20620 24380
rect 20660 24340 20669 24380
rect 20611 24339 20669 24340
rect 22731 24380 22773 24389
rect 22731 24340 22732 24380
rect 22772 24340 22773 24380
rect 22731 24331 22773 24340
rect 42987 24380 43029 24389
rect 42987 24340 42988 24380
rect 43028 24340 43029 24380
rect 42987 24331 43029 24340
rect 45475 24380 45533 24381
rect 45475 24340 45484 24380
rect 45524 24340 45533 24380
rect 45475 24339 45533 24340
rect 46339 24380 46397 24381
rect 46339 24340 46348 24380
rect 46388 24340 46397 24380
rect 46339 24339 46397 24340
rect 46531 24380 46589 24381
rect 46531 24340 46540 24380
rect 46580 24340 46589 24380
rect 46531 24339 46589 24340
rect 47979 24380 48021 24389
rect 47979 24340 47980 24380
rect 48020 24340 48021 24380
rect 47979 24331 48021 24340
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 12451 24044 12509 24045
rect 12451 24004 12460 24044
rect 12500 24004 12509 24044
rect 12451 24003 12509 24004
rect 19563 24044 19605 24053
rect 19563 24004 19564 24044
rect 19604 24004 19605 24044
rect 19563 23995 19605 24004
rect 22435 24044 22493 24045
rect 22435 24004 22444 24044
rect 22484 24004 22493 24044
rect 22435 24003 22493 24004
rect 29451 24044 29493 24053
rect 29451 24004 29452 24044
rect 29492 24004 29493 24044
rect 29451 23995 29493 24004
rect 37131 24044 37173 24053
rect 37131 24004 37132 24044
rect 37172 24004 37173 24044
rect 37131 23995 37173 24004
rect 45099 24044 45141 24053
rect 45099 24004 45100 24044
rect 45140 24004 45141 24044
rect 45099 23995 45141 24004
rect 47587 24044 47645 24045
rect 47587 24004 47596 24044
rect 47636 24004 47645 24044
rect 47587 24003 47645 24004
rect 1707 23960 1749 23969
rect 1707 23920 1708 23960
rect 1748 23920 1749 23960
rect 1707 23911 1749 23920
rect 3523 23960 3581 23961
rect 3523 23920 3532 23960
rect 3572 23920 3581 23960
rect 3523 23919 3581 23920
rect 4971 23960 5013 23969
rect 4971 23920 4972 23960
rect 5012 23920 5013 23960
rect 4971 23911 5013 23920
rect 6315 23960 6357 23969
rect 6315 23920 6316 23960
rect 6356 23920 6357 23960
rect 6315 23911 6357 23920
rect 13603 23960 13661 23961
rect 13603 23920 13612 23960
rect 13652 23920 13661 23960
rect 13603 23919 13661 23920
rect 16395 23960 16437 23969
rect 16395 23920 16396 23960
rect 16436 23920 16437 23960
rect 16395 23911 16437 23920
rect 17931 23960 17973 23969
rect 17931 23920 17932 23960
rect 17972 23920 17973 23960
rect 17931 23911 17973 23920
rect 23395 23960 23453 23961
rect 23395 23920 23404 23960
rect 23444 23920 23453 23960
rect 23395 23919 23453 23920
rect 32427 23960 32469 23969
rect 32427 23920 32428 23960
rect 32468 23920 32469 23960
rect 32427 23911 32469 23920
rect 44323 23960 44381 23961
rect 44323 23920 44332 23960
rect 44372 23920 44381 23960
rect 44323 23919 44381 23920
rect 45867 23960 45909 23969
rect 45867 23920 45868 23960
rect 45908 23920 45909 23960
rect 45867 23911 45909 23920
rect 49515 23960 49557 23969
rect 49515 23920 49516 23960
rect 49556 23920 49557 23960
rect 49515 23911 49557 23920
rect 49899 23960 49941 23969
rect 49899 23920 49900 23960
rect 49940 23920 49941 23960
rect 49899 23911 49941 23920
rect 27723 23876 27765 23885
rect 27723 23836 27724 23876
rect 27764 23836 27765 23876
rect 27723 23827 27765 23836
rect 34347 23876 34389 23885
rect 34347 23836 34348 23876
rect 34388 23836 34389 23876
rect 34347 23827 34389 23836
rect 34627 23876 34685 23877
rect 34627 23836 34636 23876
rect 34676 23836 34685 23876
rect 34627 23835 34685 23836
rect 2283 23792 2325 23801
rect 2283 23752 2284 23792
rect 2324 23752 2325 23792
rect 2283 23743 2325 23752
rect 2371 23792 2429 23793
rect 2371 23752 2380 23792
rect 2420 23752 2429 23792
rect 2371 23751 2429 23752
rect 2563 23792 2621 23793
rect 2563 23752 2572 23792
rect 2612 23752 2621 23792
rect 2563 23751 2621 23752
rect 2667 23792 2709 23801
rect 2667 23752 2668 23792
rect 2708 23752 2709 23792
rect 2667 23743 2709 23752
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3051 23743 3093 23752
rect 3243 23792 3285 23801
rect 3243 23752 3244 23792
rect 3284 23752 3285 23792
rect 3243 23743 3285 23752
rect 3331 23792 3389 23793
rect 3331 23752 3340 23792
rect 3380 23752 3389 23792
rect 3331 23751 3389 23752
rect 4195 23792 4253 23793
rect 4195 23752 4204 23792
rect 4244 23752 4253 23792
rect 4195 23751 4253 23752
rect 4491 23792 4533 23801
rect 4491 23752 4492 23792
rect 4532 23752 4533 23792
rect 4491 23743 4533 23752
rect 4587 23792 4629 23801
rect 4587 23752 4588 23792
rect 4628 23752 4629 23792
rect 4587 23743 4629 23752
rect 4683 23792 4725 23801
rect 4683 23752 4684 23792
rect 4724 23752 4725 23792
rect 4683 23743 4725 23752
rect 4867 23792 4925 23793
rect 4867 23752 4876 23792
rect 4916 23752 4925 23792
rect 4867 23751 4925 23752
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 5259 23792 5301 23801
rect 5259 23752 5260 23792
rect 5300 23752 5301 23792
rect 5259 23743 5301 23752
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 5451 23792 5493 23801
rect 5451 23752 5452 23792
rect 5492 23752 5493 23792
rect 5451 23743 5493 23752
rect 5643 23792 5685 23801
rect 5643 23752 5644 23792
rect 5684 23752 5685 23792
rect 5643 23743 5685 23752
rect 5739 23792 5781 23801
rect 5739 23752 5740 23792
rect 5780 23752 5781 23792
rect 5739 23743 5781 23752
rect 5835 23792 5877 23801
rect 5835 23752 5836 23792
rect 5876 23752 5877 23792
rect 5835 23743 5877 23752
rect 6499 23792 6557 23793
rect 6499 23752 6508 23792
rect 6548 23752 6557 23792
rect 6499 23751 6557 23752
rect 7747 23792 7805 23793
rect 7747 23752 7756 23792
rect 7796 23752 7805 23792
rect 7747 23751 7805 23752
rect 8611 23792 8669 23793
rect 8611 23752 8620 23792
rect 8660 23752 8669 23792
rect 8611 23751 8669 23752
rect 10059 23792 10101 23801
rect 10059 23752 10060 23792
rect 10100 23752 10101 23792
rect 10059 23743 10101 23752
rect 10435 23792 10493 23793
rect 10435 23752 10444 23792
rect 10484 23752 10493 23792
rect 10435 23751 10493 23752
rect 11299 23792 11357 23793
rect 11299 23752 11308 23792
rect 11348 23752 11357 23792
rect 11299 23751 11357 23752
rect 12643 23792 12701 23793
rect 12643 23752 12652 23792
rect 12692 23752 12701 23792
rect 12643 23751 12701 23752
rect 12931 23792 12989 23793
rect 12931 23752 12940 23792
rect 12980 23752 12989 23792
rect 12931 23751 12989 23752
rect 14467 23792 14525 23793
rect 14467 23752 14476 23792
rect 14516 23752 14525 23792
rect 14467 23751 14525 23752
rect 14667 23792 14709 23801
rect 14667 23752 14668 23792
rect 14708 23752 14709 23792
rect 14667 23743 14709 23752
rect 14851 23792 14909 23793
rect 14851 23752 14860 23792
rect 14900 23752 14909 23792
rect 14851 23751 14909 23752
rect 15147 23792 15189 23801
rect 15147 23752 15148 23792
rect 15188 23752 15189 23792
rect 15147 23743 15189 23752
rect 15243 23792 15285 23801
rect 15243 23752 15244 23792
rect 15284 23752 15285 23792
rect 15243 23743 15285 23752
rect 15339 23792 15381 23801
rect 15339 23752 15340 23792
rect 15380 23752 15381 23792
rect 15339 23743 15381 23752
rect 15627 23792 15669 23801
rect 15627 23752 15628 23792
rect 15668 23752 15669 23792
rect 15627 23743 15669 23752
rect 15723 23792 15765 23801
rect 15723 23752 15724 23792
rect 15764 23752 15765 23792
rect 15723 23743 15765 23752
rect 16099 23792 16157 23793
rect 16099 23752 16108 23792
rect 16148 23752 16157 23792
rect 16099 23751 16157 23752
rect 16203 23792 16245 23801
rect 16203 23752 16204 23792
rect 16244 23752 16245 23792
rect 16203 23743 16245 23752
rect 16395 23792 16437 23801
rect 16395 23752 16396 23792
rect 16436 23752 16437 23792
rect 16395 23743 16437 23752
rect 16587 23792 16629 23801
rect 16587 23752 16588 23792
rect 16628 23752 16629 23792
rect 16587 23743 16629 23752
rect 16683 23792 16725 23801
rect 16683 23752 16684 23792
rect 16724 23752 16725 23792
rect 16683 23743 16725 23752
rect 16779 23792 16821 23801
rect 16779 23752 16780 23792
rect 16820 23752 16821 23792
rect 16779 23743 16821 23752
rect 17059 23792 17117 23793
rect 17059 23752 17068 23792
rect 17108 23752 17117 23792
rect 17059 23751 17117 23752
rect 19083 23792 19125 23801
rect 19083 23752 19084 23792
rect 19124 23752 19125 23792
rect 19083 23743 19125 23752
rect 19179 23792 19221 23801
rect 19179 23752 19180 23792
rect 19220 23752 19221 23792
rect 19179 23743 19221 23752
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 19371 23792 19413 23801
rect 19371 23752 19372 23792
rect 19412 23752 19413 23792
rect 19371 23743 19413 23752
rect 19563 23792 19605 23801
rect 19563 23752 19564 23792
rect 19604 23752 19605 23792
rect 19563 23743 19605 23752
rect 19755 23792 19797 23801
rect 19755 23752 19756 23792
rect 19796 23752 19797 23792
rect 19755 23743 19797 23752
rect 19843 23792 19901 23793
rect 19843 23752 19852 23792
rect 19892 23752 19901 23792
rect 19843 23751 19901 23752
rect 20043 23792 20085 23801
rect 20043 23752 20044 23792
rect 20084 23752 20085 23792
rect 20043 23743 20085 23752
rect 20419 23792 20477 23793
rect 20419 23752 20428 23792
rect 20468 23752 20477 23792
rect 20419 23751 20477 23752
rect 21283 23792 21341 23793
rect 21283 23752 21292 23792
rect 21332 23752 21341 23792
rect 21283 23751 21341 23752
rect 22627 23792 22685 23793
rect 22627 23752 22636 23792
rect 22676 23752 22685 23792
rect 22627 23751 22685 23752
rect 22731 23792 22773 23801
rect 22731 23752 22732 23792
rect 22772 23752 22773 23792
rect 22731 23743 22773 23752
rect 22915 23792 22973 23793
rect 22915 23752 22924 23792
rect 22964 23752 22973 23792
rect 22915 23751 22973 23752
rect 23403 23792 23445 23801
rect 23403 23752 23404 23792
rect 23444 23752 23445 23792
rect 23403 23743 23445 23752
rect 23499 23792 23541 23801
rect 23499 23752 23500 23792
rect 23540 23752 23541 23792
rect 23499 23743 23541 23752
rect 23683 23792 23741 23793
rect 23683 23752 23692 23792
rect 23732 23752 23741 23792
rect 23683 23751 23741 23752
rect 23883 23792 23925 23801
rect 23883 23752 23884 23792
rect 23924 23752 23925 23792
rect 23883 23743 23925 23752
rect 24651 23792 24693 23801
rect 24651 23752 24652 23792
rect 24692 23752 24693 23792
rect 24651 23743 24693 23752
rect 24843 23792 24885 23801
rect 24843 23752 24844 23792
rect 24884 23752 24885 23792
rect 24843 23743 24885 23752
rect 25027 23792 25085 23793
rect 25027 23752 25036 23792
rect 25076 23752 25085 23792
rect 25027 23751 25085 23752
rect 25227 23792 25269 23801
rect 25227 23752 25228 23792
rect 25268 23752 25269 23792
rect 25227 23743 25269 23752
rect 25315 23792 25373 23793
rect 25315 23752 25324 23792
rect 25364 23752 25373 23792
rect 25315 23751 25373 23752
rect 25707 23792 25749 23801
rect 25707 23752 25708 23792
rect 25748 23752 25749 23792
rect 25707 23743 25749 23752
rect 25803 23792 25845 23801
rect 25803 23752 25804 23792
rect 25844 23752 25845 23792
rect 25803 23743 25845 23752
rect 25987 23792 26045 23793
rect 25987 23752 25996 23792
rect 26036 23752 26045 23792
rect 25987 23751 26045 23752
rect 26091 23792 26133 23801
rect 26091 23752 26092 23792
rect 26132 23752 26133 23792
rect 26091 23743 26133 23752
rect 26275 23792 26333 23793
rect 26275 23752 26284 23792
rect 26324 23752 26333 23792
rect 26275 23751 26333 23752
rect 26475 23792 26517 23801
rect 26475 23752 26476 23792
rect 26516 23752 26517 23792
rect 26475 23743 26517 23752
rect 26659 23792 26717 23793
rect 26659 23752 26668 23792
rect 26708 23752 26717 23792
rect 26659 23751 26717 23752
rect 27139 23792 27197 23793
rect 27139 23752 27148 23792
rect 27188 23752 27197 23792
rect 27139 23751 27197 23752
rect 27243 23792 27285 23801
rect 27243 23752 27244 23792
rect 27284 23752 27285 23792
rect 27243 23743 27285 23752
rect 27435 23792 27477 23801
rect 27435 23752 27436 23792
rect 27476 23752 27477 23792
rect 27435 23743 27477 23752
rect 27627 23792 27669 23801
rect 27627 23752 27628 23792
rect 27668 23752 27669 23792
rect 27627 23743 27669 23752
rect 27811 23792 27869 23793
rect 27811 23752 27820 23792
rect 27860 23752 27869 23792
rect 27811 23751 27869 23752
rect 28099 23792 28157 23793
rect 28099 23752 28108 23792
rect 28148 23752 28157 23792
rect 28099 23751 28157 23752
rect 28491 23792 28533 23801
rect 28491 23752 28492 23792
rect 28532 23752 28533 23792
rect 28491 23743 28533 23752
rect 28587 23792 28629 23801
rect 28587 23752 28588 23792
rect 28628 23752 28629 23792
rect 28587 23743 28629 23752
rect 28683 23792 28725 23801
rect 28683 23752 28684 23792
rect 28724 23752 28725 23792
rect 28683 23743 28725 23752
rect 28779 23792 28821 23801
rect 28779 23752 28780 23792
rect 28820 23752 28821 23792
rect 28779 23743 28821 23752
rect 29067 23792 29109 23801
rect 29067 23752 29068 23792
rect 29108 23752 29109 23792
rect 29067 23743 29109 23752
rect 29163 23792 29205 23801
rect 29163 23752 29164 23792
rect 29204 23752 29205 23792
rect 29163 23743 29205 23752
rect 29259 23792 29301 23801
rect 29259 23752 29260 23792
rect 29300 23752 29301 23792
rect 29259 23743 29301 23752
rect 29451 23792 29493 23801
rect 29451 23752 29452 23792
rect 29492 23752 29493 23792
rect 29451 23743 29493 23752
rect 29643 23792 29685 23801
rect 29643 23752 29644 23792
rect 29684 23752 29685 23792
rect 29643 23743 29685 23752
rect 29731 23792 29789 23793
rect 29731 23752 29740 23792
rect 29780 23752 29789 23792
rect 29731 23751 29789 23752
rect 30787 23792 30845 23793
rect 30787 23752 30796 23792
rect 30836 23752 30845 23792
rect 30787 23751 30845 23752
rect 31083 23792 31125 23801
rect 31083 23752 31084 23792
rect 31124 23752 31125 23792
rect 31083 23743 31125 23752
rect 31179 23792 31221 23801
rect 31179 23752 31180 23792
rect 31220 23752 31221 23792
rect 31179 23743 31221 23752
rect 31275 23792 31317 23801
rect 31275 23752 31276 23792
rect 31316 23752 31317 23792
rect 31275 23743 31317 23752
rect 33091 23792 33149 23793
rect 33091 23752 33100 23792
rect 33140 23752 33149 23792
rect 33091 23751 33149 23752
rect 33475 23792 33533 23793
rect 33475 23752 33484 23792
rect 33524 23752 33533 23792
rect 33475 23751 33533 23752
rect 35683 23792 35741 23793
rect 35683 23752 35692 23792
rect 35732 23752 35741 23792
rect 35683 23751 35741 23752
rect 36747 23792 36789 23801
rect 36747 23752 36748 23792
rect 36788 23752 36789 23792
rect 36747 23743 36789 23752
rect 37219 23792 37277 23793
rect 37219 23752 37228 23792
rect 37268 23752 37277 23792
rect 37219 23751 37277 23752
rect 37411 23792 37469 23793
rect 37411 23752 37420 23792
rect 37460 23752 37469 23792
rect 37411 23751 37469 23752
rect 37515 23792 37557 23801
rect 37515 23752 37516 23792
rect 37556 23752 37557 23792
rect 37515 23743 37557 23752
rect 37707 23792 37749 23801
rect 37707 23752 37708 23792
rect 37748 23752 37749 23792
rect 37707 23743 37749 23752
rect 37899 23792 37941 23801
rect 37899 23752 37900 23792
rect 37940 23752 37941 23792
rect 37899 23743 37941 23752
rect 37995 23792 38037 23801
rect 37995 23752 37996 23792
rect 38036 23752 38037 23792
rect 37995 23743 38037 23752
rect 38091 23792 38133 23801
rect 38091 23752 38092 23792
rect 38132 23752 38133 23792
rect 38091 23743 38133 23752
rect 38187 23792 38229 23801
rect 38187 23752 38188 23792
rect 38228 23752 38229 23792
rect 38187 23743 38229 23752
rect 38755 23792 38813 23793
rect 38755 23752 38764 23792
rect 38804 23752 38813 23792
rect 38755 23751 38813 23752
rect 39619 23792 39677 23793
rect 39619 23752 39628 23792
rect 39668 23752 39677 23792
rect 39619 23751 39677 23752
rect 41731 23792 41789 23793
rect 41731 23752 41740 23792
rect 41780 23752 41789 23792
rect 41731 23751 41789 23752
rect 41931 23792 41973 23801
rect 41931 23752 41932 23792
rect 41972 23752 41973 23792
rect 41931 23743 41973 23752
rect 42307 23792 42365 23793
rect 42307 23752 42316 23792
rect 42356 23752 42365 23792
rect 42307 23751 42365 23752
rect 43171 23792 43229 23793
rect 43171 23752 43180 23792
rect 43220 23752 43229 23792
rect 43171 23751 43229 23752
rect 44611 23792 44669 23793
rect 44611 23752 44620 23792
rect 44660 23752 44669 23792
rect 44611 23751 44669 23752
rect 45763 23792 45821 23793
rect 45763 23752 45772 23792
rect 45812 23752 45821 23792
rect 45763 23751 45821 23752
rect 46155 23792 46197 23801
rect 46155 23752 46156 23792
rect 46196 23752 46197 23792
rect 46155 23743 46197 23752
rect 46923 23792 46965 23801
rect 46923 23752 46924 23792
rect 46964 23752 46965 23792
rect 46923 23743 46965 23752
rect 48259 23792 48317 23793
rect 48259 23752 48268 23792
rect 48308 23752 48317 23792
rect 48259 23751 48317 23752
rect 48451 23792 48509 23793
rect 48451 23752 48460 23792
rect 48500 23752 48509 23792
rect 48451 23751 48509 23752
rect 2763 23708 2805 23717
rect 2763 23668 2764 23708
rect 2804 23668 2805 23708
rect 2763 23659 2805 23668
rect 5931 23708 5973 23717
rect 5931 23668 5932 23708
rect 5972 23668 5973 23708
rect 5931 23659 5973 23668
rect 7179 23708 7221 23717
rect 7179 23668 7180 23708
rect 7220 23668 7221 23708
rect 7179 23659 7221 23668
rect 7371 23708 7413 23717
rect 7371 23668 7372 23708
rect 7412 23668 7413 23708
rect 7371 23659 7413 23668
rect 14763 23708 14805 23717
rect 14763 23668 14764 23708
rect 14804 23668 14805 23708
rect 14763 23659 14805 23668
rect 15051 23708 15093 23717
rect 15051 23668 15052 23708
rect 15092 23668 15093 23708
rect 15051 23659 15093 23668
rect 23299 23708 23357 23709
rect 23299 23668 23308 23708
rect 23348 23668 23357 23708
rect 23299 23667 23357 23668
rect 23787 23708 23829 23717
rect 23787 23668 23788 23708
rect 23828 23668 23829 23708
rect 23787 23659 23829 23668
rect 26571 23708 26613 23717
rect 26571 23668 26572 23708
rect 26612 23668 26613 23708
rect 26571 23659 26613 23668
rect 35971 23708 36029 23709
rect 35971 23668 35980 23708
rect 36020 23668 36029 23708
rect 35971 23667 36029 23668
rect 38379 23708 38421 23717
rect 38379 23668 38380 23708
rect 38420 23668 38421 23708
rect 38379 23659 38421 23668
rect 3139 23624 3197 23625
rect 3139 23584 3148 23624
rect 3188 23584 3197 23624
rect 3139 23583 3197 23584
rect 4387 23624 4445 23625
rect 4387 23584 4396 23624
rect 4436 23584 4445 23624
rect 4387 23583 4445 23584
rect 9763 23624 9821 23625
rect 9763 23584 9772 23624
rect 9812 23584 9821 23624
rect 9763 23583 9821 23584
rect 12747 23624 12789 23633
rect 12747 23584 12748 23624
rect 12788 23584 12789 23624
rect 12747 23575 12789 23584
rect 13795 23624 13853 23625
rect 13795 23584 13804 23624
rect 13844 23584 13853 23624
rect 13795 23583 13853 23584
rect 15907 23624 15965 23625
rect 15907 23584 15916 23624
rect 15956 23584 15965 23624
rect 15907 23583 15965 23584
rect 16867 23624 16925 23625
rect 16867 23584 16876 23624
rect 16916 23584 16925 23624
rect 16867 23583 16925 23584
rect 17731 23624 17789 23625
rect 17731 23584 17740 23624
rect 17780 23584 17789 23624
rect 17731 23583 17789 23584
rect 22923 23624 22965 23633
rect 22923 23584 22924 23624
rect 22964 23584 22965 23624
rect 22923 23575 22965 23584
rect 23115 23624 23157 23633
rect 23115 23584 23116 23624
rect 23156 23584 23157 23624
rect 23115 23575 23157 23584
rect 23203 23624 23261 23625
rect 23203 23584 23212 23624
rect 23252 23584 23261 23624
rect 23203 23583 23261 23584
rect 24747 23624 24789 23633
rect 24747 23584 24748 23624
rect 24788 23584 24789 23624
rect 24747 23575 24789 23584
rect 25035 23624 25077 23633
rect 25035 23584 25036 23624
rect 25076 23584 25077 23624
rect 25035 23575 25077 23584
rect 25507 23624 25565 23625
rect 25507 23584 25516 23624
rect 25556 23584 25565 23624
rect 25507 23583 25565 23584
rect 26283 23624 26325 23633
rect 26283 23584 26284 23624
rect 26324 23584 26325 23624
rect 26283 23575 26325 23584
rect 27331 23624 27389 23625
rect 27331 23584 27340 23624
rect 27380 23584 27389 23624
rect 27331 23583 27389 23584
rect 28003 23624 28061 23625
rect 28003 23584 28012 23624
rect 28052 23584 28061 23624
rect 28003 23583 28061 23584
rect 28291 23624 28349 23625
rect 28291 23584 28300 23624
rect 28340 23584 28349 23624
rect 28291 23583 28349 23584
rect 28963 23624 29021 23625
rect 28963 23584 28972 23624
rect 29012 23584 29021 23624
rect 28963 23583 29021 23584
rect 30891 23624 30933 23633
rect 30891 23584 30892 23624
rect 30932 23584 30933 23624
rect 30891 23575 30933 23584
rect 31363 23624 31421 23625
rect 31363 23584 31372 23624
rect 31412 23584 31421 23624
rect 31363 23583 31421 23584
rect 34827 23624 34869 23633
rect 34827 23584 34828 23624
rect 34868 23584 34869 23624
rect 34827 23575 34869 23584
rect 35011 23624 35069 23625
rect 35011 23584 35020 23624
rect 35060 23584 35069 23624
rect 35011 23583 35069 23584
rect 37131 23624 37173 23633
rect 37131 23584 37132 23624
rect 37172 23584 37173 23624
rect 37131 23575 37173 23584
rect 37603 23624 37661 23625
rect 37603 23584 37612 23624
rect 37652 23584 37661 23624
rect 37603 23583 37661 23584
rect 40771 23624 40829 23625
rect 40771 23584 40780 23624
rect 40820 23584 40829 23624
rect 40771 23583 40829 23584
rect 41059 23624 41117 23625
rect 41059 23584 41068 23624
rect 41108 23584 41117 23624
rect 41059 23583 41117 23584
rect 47587 23624 47645 23625
rect 47587 23584 47596 23624
rect 47636 23584 47645 23624
rect 47587 23583 47645 23584
rect 49123 23624 49181 23625
rect 49123 23584 49132 23624
rect 49172 23584 49181 23624
rect 49123 23583 49181 23584
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 3619 23288 3677 23289
rect 3619 23248 3628 23288
rect 3668 23248 3677 23288
rect 3619 23247 3677 23248
rect 6027 23288 6069 23297
rect 6027 23248 6028 23288
rect 6068 23248 6069 23288
rect 6027 23239 6069 23248
rect 7171 23288 7229 23289
rect 7171 23248 7180 23288
rect 7220 23248 7229 23288
rect 7171 23247 7229 23248
rect 11115 23288 11157 23297
rect 11115 23248 11116 23288
rect 11156 23248 11157 23288
rect 11115 23239 11157 23248
rect 12067 23288 12125 23289
rect 12067 23248 12076 23288
rect 12116 23248 12125 23288
rect 12067 23247 12125 23248
rect 16003 23288 16061 23289
rect 16003 23248 16012 23288
rect 16052 23248 16061 23288
rect 16003 23247 16061 23248
rect 19747 23288 19805 23289
rect 19747 23248 19756 23288
rect 19796 23248 19805 23288
rect 19747 23247 19805 23248
rect 25891 23288 25949 23289
rect 25891 23248 25900 23288
rect 25940 23248 25949 23288
rect 25891 23247 25949 23248
rect 28779 23288 28821 23297
rect 28779 23248 28780 23288
rect 28820 23248 28821 23288
rect 28779 23239 28821 23248
rect 29067 23288 29109 23297
rect 29067 23248 29068 23288
rect 29108 23248 29109 23288
rect 29067 23239 29109 23248
rect 30891 23288 30933 23297
rect 30891 23248 30892 23288
rect 30932 23248 30933 23288
rect 30891 23239 30933 23248
rect 36547 23288 36605 23289
rect 36547 23248 36556 23288
rect 36596 23248 36605 23288
rect 36547 23247 36605 23248
rect 37123 23288 37181 23289
rect 37123 23248 37132 23288
rect 37172 23248 37181 23288
rect 37123 23247 37181 23248
rect 38371 23288 38429 23289
rect 38371 23248 38380 23288
rect 38420 23248 38429 23288
rect 38371 23247 38429 23248
rect 43075 23288 43133 23289
rect 43075 23248 43084 23288
rect 43124 23248 43133 23288
rect 43075 23247 43133 23248
rect 1227 23204 1269 23213
rect 1227 23164 1228 23204
rect 1268 23164 1269 23204
rect 1227 23155 1269 23164
rect 7467 23204 7509 23213
rect 7467 23164 7468 23204
rect 7508 23164 7509 23204
rect 7467 23155 7509 23164
rect 13611 23204 13653 23213
rect 13611 23164 13612 23204
rect 13652 23164 13653 23204
rect 13611 23155 13653 23164
rect 17355 23204 17397 23213
rect 17355 23164 17356 23204
rect 17396 23164 17397 23204
rect 17355 23155 17397 23164
rect 26283 23204 26325 23213
rect 26283 23164 26284 23204
rect 26324 23164 26325 23204
rect 26283 23155 26325 23164
rect 29547 23204 29589 23213
rect 29547 23164 29548 23204
rect 29588 23164 29589 23204
rect 29547 23155 29589 23164
rect 35787 23204 35829 23213
rect 35787 23164 35788 23204
rect 35828 23164 35829 23204
rect 35787 23155 35829 23164
rect 47403 23204 47445 23213
rect 47403 23164 47404 23204
rect 47444 23164 47445 23204
rect 47403 23155 47445 23164
rect 1603 23120 1661 23121
rect 1603 23080 1612 23120
rect 1652 23080 1661 23120
rect 1603 23079 1661 23080
rect 2467 23120 2525 23121
rect 2467 23080 2476 23120
rect 2516 23080 2525 23120
rect 2467 23079 2525 23080
rect 3915 23120 3957 23129
rect 3915 23080 3916 23120
rect 3956 23080 3957 23120
rect 3915 23071 3957 23080
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4195 23120 4253 23121
rect 4195 23080 4204 23120
rect 4244 23080 4253 23120
rect 4195 23079 4253 23080
rect 4483 23120 4541 23121
rect 4483 23080 4492 23120
rect 4532 23080 4541 23120
rect 4483 23079 4541 23080
rect 4779 23120 4821 23129
rect 4779 23080 4780 23120
rect 4820 23080 4821 23120
rect 4779 23071 4821 23080
rect 4875 23120 4917 23129
rect 4875 23080 4876 23120
rect 4916 23080 4917 23120
rect 4875 23071 4917 23080
rect 5451 23120 5493 23129
rect 5451 23080 5452 23120
rect 5492 23080 5493 23120
rect 5451 23071 5493 23080
rect 5539 23120 5597 23121
rect 5539 23080 5548 23120
rect 5588 23080 5597 23120
rect 5539 23079 5597 23080
rect 5731 23120 5789 23121
rect 5731 23080 5740 23120
rect 5780 23080 5789 23120
rect 5731 23079 5789 23080
rect 6115 23120 6173 23121
rect 6115 23080 6124 23120
rect 6164 23080 6173 23120
rect 6115 23079 6173 23080
rect 6699 23120 6741 23129
rect 6699 23080 6700 23120
rect 6740 23080 6741 23120
rect 6699 23071 6741 23080
rect 6787 23120 6845 23121
rect 6787 23080 6796 23120
rect 6836 23080 6845 23120
rect 6787 23079 6845 23080
rect 6979 23120 7037 23121
rect 6979 23080 6988 23120
rect 7028 23080 7037 23120
rect 6979 23079 7037 23080
rect 7083 23120 7125 23129
rect 7083 23080 7084 23120
rect 7124 23080 7125 23120
rect 7083 23071 7125 23080
rect 7275 23120 7317 23129
rect 7275 23080 7276 23120
rect 7316 23080 7317 23120
rect 7275 23071 7317 23080
rect 8131 23120 8189 23121
rect 8131 23080 8140 23120
rect 8180 23080 8189 23120
rect 8131 23079 8189 23080
rect 8331 23120 8373 23129
rect 8331 23080 8332 23120
rect 8372 23080 8373 23120
rect 8331 23071 8373 23080
rect 8427 23120 8469 23129
rect 8427 23080 8428 23120
rect 8468 23080 8469 23120
rect 8427 23071 8469 23080
rect 8523 23120 8565 23129
rect 8523 23080 8524 23120
rect 8564 23080 8565 23120
rect 8523 23071 8565 23080
rect 8619 23120 8661 23129
rect 8619 23080 8620 23120
rect 8660 23080 8661 23120
rect 8619 23071 8661 23080
rect 9195 23120 9237 23129
rect 9195 23080 9196 23120
rect 9236 23080 9237 23120
rect 9195 23071 9237 23080
rect 9291 23120 9333 23129
rect 9291 23080 9292 23120
rect 9332 23080 9333 23120
rect 9291 23071 9333 23080
rect 9387 23120 9429 23129
rect 9387 23080 9388 23120
rect 9428 23080 9429 23120
rect 9387 23071 9429 23080
rect 9483 23120 9525 23129
rect 9483 23080 9484 23120
rect 9524 23080 9525 23120
rect 9483 23071 9525 23080
rect 9675 23120 9717 23129
rect 9675 23080 9676 23120
rect 9716 23080 9717 23120
rect 9675 23071 9717 23080
rect 9867 23120 9909 23129
rect 9867 23080 9868 23120
rect 9908 23080 9909 23120
rect 9867 23071 9909 23080
rect 9955 23120 10013 23121
rect 9955 23080 9964 23120
rect 10004 23080 10013 23120
rect 9955 23079 10013 23080
rect 11203 23120 11261 23121
rect 11203 23080 11212 23120
rect 11252 23080 11261 23120
rect 11203 23079 11261 23080
rect 11395 23120 11453 23121
rect 11395 23080 11404 23120
rect 11444 23080 11453 23120
rect 11395 23079 11453 23080
rect 12259 23120 12317 23121
rect 12259 23080 12268 23120
rect 12308 23080 12317 23120
rect 12259 23079 12317 23080
rect 12363 23120 12405 23129
rect 12363 23080 12364 23120
rect 12404 23080 12405 23120
rect 12363 23071 12405 23080
rect 12555 23120 12597 23129
rect 12555 23080 12556 23120
rect 12596 23080 12597 23120
rect 12555 23071 12597 23080
rect 12739 23120 12797 23121
rect 12739 23080 12748 23120
rect 12788 23080 12797 23120
rect 12739 23079 12797 23080
rect 13987 23120 14045 23121
rect 13987 23080 13996 23120
rect 14036 23080 14045 23120
rect 13987 23079 14045 23080
rect 14851 23120 14909 23121
rect 14851 23080 14860 23120
rect 14900 23080 14909 23120
rect 14851 23079 14909 23080
rect 16291 23120 16349 23121
rect 16291 23080 16300 23120
rect 16340 23080 16349 23120
rect 16291 23079 16349 23080
rect 17731 23120 17789 23121
rect 17731 23080 17740 23120
rect 17780 23080 17789 23120
rect 17731 23079 17789 23080
rect 18595 23120 18653 23121
rect 18595 23080 18604 23120
rect 18644 23080 18653 23120
rect 18595 23079 18653 23080
rect 20611 23120 20669 23121
rect 20611 23080 20620 23120
rect 20660 23080 20669 23120
rect 20611 23079 20669 23080
rect 23115 23120 23157 23129
rect 23115 23080 23116 23120
rect 23156 23080 23157 23120
rect 23115 23071 23157 23080
rect 23403 23127 23445 23136
rect 23403 23087 23404 23127
rect 23444 23087 23445 23127
rect 23403 23078 23445 23087
rect 23691 23120 23733 23129
rect 23691 23080 23692 23120
rect 23732 23080 23733 23120
rect 23691 23071 23733 23080
rect 23787 23120 23829 23129
rect 23787 23080 23788 23120
rect 23828 23080 23829 23120
rect 23787 23071 23829 23080
rect 23883 23120 23925 23129
rect 23883 23080 23884 23120
rect 23924 23080 23925 23120
rect 23883 23071 23925 23080
rect 23979 23120 24021 23129
rect 23979 23080 23980 23120
rect 24020 23080 24021 23120
rect 23979 23071 24021 23080
rect 24363 23120 24405 23129
rect 24363 23080 24364 23120
rect 24404 23080 24405 23120
rect 24363 23071 24405 23080
rect 24451 23120 24509 23121
rect 24451 23080 24460 23120
rect 24500 23080 24509 23120
rect 24451 23079 24509 23080
rect 25027 23120 25085 23121
rect 25027 23080 25036 23120
rect 25076 23080 25085 23120
rect 25027 23079 25085 23080
rect 25419 23120 25461 23129
rect 25419 23080 25420 23120
rect 25460 23080 25461 23120
rect 25419 23071 25461 23080
rect 25611 23120 25653 23129
rect 25611 23080 25612 23120
rect 25652 23080 25653 23120
rect 25611 23071 25653 23080
rect 25707 23120 25749 23129
rect 25707 23080 25708 23120
rect 25748 23080 25749 23120
rect 25707 23071 25749 23080
rect 25803 23120 25845 23129
rect 25803 23080 25804 23120
rect 25844 23080 25845 23120
rect 25803 23071 25845 23080
rect 26083 23120 26141 23121
rect 26083 23080 26092 23120
rect 26132 23080 26141 23120
rect 26083 23079 26141 23080
rect 26187 23120 26229 23129
rect 26187 23080 26188 23120
rect 26228 23080 26229 23120
rect 26187 23071 26229 23080
rect 26379 23120 26421 23129
rect 26379 23080 26380 23120
rect 26420 23080 26421 23120
rect 26379 23071 26421 23080
rect 26571 23120 26613 23129
rect 26571 23080 26572 23120
rect 26612 23080 26613 23120
rect 26571 23071 26613 23080
rect 26667 23120 26709 23129
rect 26667 23080 26668 23120
rect 26708 23080 26709 23120
rect 26667 23071 26709 23080
rect 26763 23120 26805 23129
rect 26763 23080 26764 23120
rect 26804 23080 26805 23120
rect 26763 23071 26805 23080
rect 26859 23120 26901 23129
rect 26859 23080 26860 23120
rect 26900 23080 26901 23120
rect 26859 23071 26901 23080
rect 27043 23120 27101 23121
rect 27043 23080 27052 23120
rect 27092 23080 27101 23120
rect 27043 23079 27101 23080
rect 27243 23120 27285 23129
rect 27243 23080 27244 23120
rect 27284 23080 27285 23120
rect 27243 23071 27285 23080
rect 27331 23120 27389 23121
rect 27331 23080 27340 23120
rect 27380 23080 27389 23120
rect 27331 23079 27389 23080
rect 27723 23120 27765 23129
rect 27723 23080 27724 23120
rect 27764 23080 27765 23120
rect 27723 23071 27765 23080
rect 27811 23120 27869 23121
rect 27811 23080 27820 23120
rect 27860 23080 27869 23120
rect 27811 23079 27869 23080
rect 28291 23120 28349 23121
rect 28291 23080 28300 23120
rect 28340 23080 28349 23120
rect 28291 23079 28349 23080
rect 28491 23120 28533 23129
rect 28491 23080 28492 23120
rect 28532 23080 28533 23120
rect 28491 23071 28533 23080
rect 28579 23120 28637 23121
rect 28579 23080 28588 23120
rect 28628 23080 28637 23120
rect 28579 23079 28637 23080
rect 28971 23120 29013 23129
rect 28971 23080 28972 23120
rect 29012 23080 29013 23120
rect 28971 23071 29013 23080
rect 29163 23120 29205 23129
rect 29163 23080 29164 23120
rect 29204 23080 29205 23120
rect 29163 23071 29205 23080
rect 29443 23120 29501 23121
rect 29443 23080 29452 23120
rect 29492 23080 29501 23120
rect 29443 23079 29501 23080
rect 29643 23120 29685 23129
rect 29643 23080 29644 23120
rect 29684 23080 29685 23120
rect 29643 23071 29685 23080
rect 30403 23120 30461 23121
rect 30403 23080 30412 23120
rect 30452 23080 30461 23120
rect 30403 23079 30461 23080
rect 31563 23120 31605 23129
rect 31563 23080 31564 23120
rect 31604 23080 31605 23120
rect 31563 23071 31605 23080
rect 31755 23120 31797 23129
rect 31755 23080 31756 23120
rect 31796 23080 31797 23120
rect 31755 23071 31797 23080
rect 31843 23120 31901 23121
rect 31843 23080 31852 23120
rect 31892 23080 31901 23120
rect 31843 23079 31901 23080
rect 32899 23120 32957 23121
rect 32899 23080 32908 23120
rect 32948 23080 32957 23120
rect 32899 23079 32957 23080
rect 33579 23120 33621 23129
rect 33579 23080 33580 23120
rect 33620 23080 33621 23120
rect 33579 23071 33621 23080
rect 33859 23120 33917 23121
rect 33859 23080 33868 23120
rect 33908 23080 33917 23120
rect 33859 23079 33917 23080
rect 35019 23120 35061 23129
rect 35019 23080 35020 23120
rect 35060 23080 35061 23120
rect 35019 23071 35061 23080
rect 35115 23120 35157 23129
rect 35115 23080 35116 23120
rect 35156 23080 35157 23120
rect 35115 23071 35157 23080
rect 35211 23120 35253 23129
rect 35211 23080 35212 23120
rect 35252 23080 35253 23120
rect 35211 23071 35253 23080
rect 35307 23120 35349 23129
rect 35307 23080 35308 23120
rect 35348 23080 35349 23120
rect 35307 23071 35349 23080
rect 35883 23120 35925 23129
rect 35883 23080 35884 23120
rect 35924 23080 35925 23120
rect 35883 23071 35925 23080
rect 36163 23120 36221 23121
rect 36163 23080 36172 23120
rect 36212 23080 36221 23120
rect 36163 23079 36221 23080
rect 36459 23120 36501 23129
rect 36459 23080 36460 23120
rect 36500 23080 36501 23120
rect 36459 23071 36501 23080
rect 36651 23120 36693 23129
rect 36651 23080 36652 23120
rect 36692 23080 36693 23120
rect 36651 23071 36693 23080
rect 36739 23120 36797 23121
rect 36739 23080 36748 23120
rect 36788 23080 36797 23120
rect 36739 23079 36797 23080
rect 37795 23120 37853 23121
rect 37795 23080 37804 23120
rect 37844 23080 37853 23120
rect 37795 23079 37853 23080
rect 39043 23120 39101 23121
rect 39043 23080 39052 23120
rect 39092 23080 39101 23120
rect 39043 23079 39101 23080
rect 39331 23120 39389 23121
rect 39331 23080 39340 23120
rect 39380 23080 39389 23120
rect 39331 23079 39389 23080
rect 40291 23120 40349 23121
rect 40291 23080 40300 23120
rect 40340 23080 40349 23120
rect 40291 23079 40349 23080
rect 40579 23120 40637 23121
rect 40579 23080 40588 23120
rect 40628 23080 40637 23120
rect 40579 23079 40637 23080
rect 40683 23120 40725 23129
rect 40683 23080 40684 23120
rect 40724 23080 40725 23120
rect 40683 23071 40725 23080
rect 41251 23120 41309 23121
rect 41251 23080 41260 23120
rect 41300 23080 41309 23120
rect 41251 23079 41309 23080
rect 41355 23120 41397 23129
rect 41355 23080 41356 23120
rect 41396 23080 41397 23120
rect 41355 23071 41397 23080
rect 41547 23120 41589 23129
rect 41547 23080 41548 23120
rect 41588 23080 41589 23120
rect 41547 23071 41589 23080
rect 41739 23120 41781 23129
rect 41739 23080 41740 23120
rect 41780 23080 41781 23120
rect 41739 23071 41781 23080
rect 41835 23120 41877 23129
rect 41835 23080 41836 23120
rect 41876 23080 41877 23120
rect 41835 23071 41877 23080
rect 41931 23120 41973 23129
rect 41931 23080 41932 23120
rect 41972 23080 41973 23120
rect 41931 23071 41973 23080
rect 42027 23120 42069 23129
rect 42027 23080 42028 23120
rect 42068 23080 42069 23120
rect 42027 23071 42069 23080
rect 42211 23120 42269 23121
rect 42211 23080 42220 23120
rect 42260 23080 42269 23120
rect 42211 23079 42269 23080
rect 43747 23120 43805 23121
rect 43747 23080 43756 23120
rect 43796 23080 43805 23120
rect 43747 23079 43805 23080
rect 44803 23120 44861 23121
rect 44803 23080 44812 23120
rect 44852 23080 44861 23120
rect 44803 23079 44861 23080
rect 46147 23120 46205 23121
rect 46147 23080 46156 23120
rect 46196 23080 46205 23120
rect 46147 23079 46205 23080
rect 47011 23120 47069 23121
rect 47011 23080 47020 23120
rect 47060 23080 47069 23120
rect 47011 23079 47069 23080
rect 48643 23120 48701 23121
rect 48643 23080 48652 23120
rect 48692 23080 48701 23120
rect 48643 23079 48701 23080
rect 49891 23120 49949 23121
rect 49891 23080 49900 23120
rect 49940 23080 49949 23120
rect 49891 23079 49949 23080
rect 50755 23120 50813 23121
rect 50755 23080 50764 23120
rect 50804 23080 50813 23120
rect 50755 23079 50813 23080
rect 51147 23120 51189 23129
rect 51147 23080 51148 23120
rect 51188 23080 51189 23120
rect 51147 23071 51189 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 24739 23036 24797 23037
rect 24739 22996 24748 23036
rect 24788 22996 24797 23036
rect 24739 22995 24797 22996
rect 25131 23036 25173 23045
rect 25131 22996 25132 23036
rect 25172 22996 25173 23036
rect 25131 22987 25173 22996
rect 25323 23036 25365 23045
rect 25323 22996 25324 23036
rect 25364 22996 25365 23036
rect 25323 22987 25365 22996
rect 28099 23036 28157 23037
rect 28099 22996 28108 23036
rect 28148 22996 28157 23036
rect 28099 22995 28157 22996
rect 30115 23036 30173 23037
rect 30115 22996 30124 23036
rect 30164 22996 30173 23036
rect 30115 22995 30173 22996
rect 37987 23036 38045 23037
rect 37987 22996 37996 23036
rect 38036 22996 38045 23036
rect 37987 22995 38045 22996
rect 44139 23036 44181 23045
rect 44139 22996 44140 23036
rect 44180 22996 44181 23036
rect 44139 22987 44181 22996
rect 5155 22952 5213 22953
rect 5155 22912 5164 22952
rect 5204 22912 5213 22952
rect 5155 22911 5213 22912
rect 10347 22952 10389 22961
rect 10347 22912 10348 22952
rect 10388 22912 10389 22952
rect 10347 22903 10389 22912
rect 12555 22952 12597 22961
rect 12555 22912 12556 22952
rect 12596 22912 12597 22952
rect 12555 22903 12597 22912
rect 23403 22952 23445 22961
rect 23403 22912 23404 22952
rect 23444 22912 23445 22952
rect 23403 22903 23445 22912
rect 25227 22952 25269 22961
rect 25227 22912 25228 22952
rect 25268 22912 25269 22952
rect 25227 22903 25269 22912
rect 29931 22952 29973 22961
rect 29931 22912 29932 22952
rect 29972 22912 29973 22952
rect 29931 22903 29973 22912
rect 32043 22952 32085 22961
rect 32043 22912 32044 22952
rect 32084 22912 32085 22952
rect 32043 22903 32085 22912
rect 34155 22952 34197 22961
rect 34155 22912 34156 22952
rect 34196 22912 34197 22952
rect 34155 22903 34197 22912
rect 39627 22952 39669 22961
rect 39627 22912 39628 22952
rect 39668 22912 39669 22952
rect 39627 22903 39669 22912
rect 41067 22952 41109 22961
rect 41067 22912 41068 22952
rect 41108 22912 41109 22952
rect 41067 22903 41109 22912
rect 41547 22952 41589 22961
rect 41547 22912 41548 22952
rect 41588 22912 41589 22952
rect 41547 22903 41589 22912
rect 44995 22952 45053 22953
rect 44995 22912 45004 22952
rect 45044 22912 45053 22952
rect 44995 22911 45053 22912
rect 47595 22952 47637 22961
rect 47595 22912 47596 22952
rect 47636 22912 47637 22952
rect 47595 22903 47637 22912
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 3915 22868 3957 22877
rect 3915 22828 3916 22868
rect 3956 22828 3957 22868
rect 3915 22819 3957 22828
rect 5835 22868 5877 22877
rect 5835 22828 5836 22868
rect 5876 22828 5877 22868
rect 5835 22819 5877 22828
rect 9675 22868 9717 22877
rect 9675 22828 9676 22868
rect 9716 22828 9717 22868
rect 9675 22819 9717 22828
rect 13411 22868 13469 22869
rect 13411 22828 13420 22868
rect 13460 22828 13469 22868
rect 13411 22827 13469 22828
rect 16963 22868 17021 22869
rect 16963 22828 16972 22868
rect 17012 22828 17021 22868
rect 16963 22827 17021 22828
rect 19939 22868 19997 22869
rect 19939 22828 19948 22868
rect 19988 22828 19997 22868
rect 19939 22827 19997 22828
rect 24651 22868 24693 22877
rect 24651 22828 24652 22868
rect 24692 22828 24693 22868
rect 24651 22819 24693 22828
rect 27051 22868 27093 22877
rect 27051 22828 27052 22868
rect 27092 22828 27093 22868
rect 27051 22819 27093 22828
rect 31563 22868 31605 22877
rect 31563 22828 31564 22868
rect 31604 22828 31605 22868
rect 31563 22819 31605 22828
rect 35491 22868 35549 22869
rect 35491 22828 35500 22868
rect 35540 22828 35549 22868
rect 35491 22827 35549 22828
rect 37123 22868 37181 22869
rect 37123 22828 37132 22868
rect 37172 22828 37181 22868
rect 37123 22827 37181 22828
rect 40011 22868 40053 22877
rect 40011 22828 40012 22868
rect 40052 22828 40053 22868
rect 40011 22819 40053 22828
rect 42883 22868 42941 22869
rect 42883 22828 42892 22868
rect 42932 22828 42941 22868
rect 42883 22827 42941 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 4963 22532 5021 22533
rect 4963 22492 4972 22532
rect 5012 22492 5021 22532
rect 4963 22491 5021 22492
rect 5643 22532 5685 22541
rect 5643 22492 5644 22532
rect 5684 22492 5685 22532
rect 5643 22483 5685 22492
rect 8707 22532 8765 22533
rect 8707 22492 8716 22532
rect 8756 22492 8765 22532
rect 8707 22491 8765 22492
rect 11299 22532 11357 22533
rect 11299 22492 11308 22532
rect 11348 22492 11357 22532
rect 11299 22491 11357 22492
rect 12747 22532 12789 22541
rect 12747 22492 12748 22532
rect 12788 22492 12789 22532
rect 12747 22483 12789 22492
rect 14859 22532 14901 22541
rect 14859 22492 14860 22532
rect 14900 22492 14901 22532
rect 14859 22483 14901 22492
rect 19275 22532 19317 22541
rect 19275 22492 19276 22532
rect 19316 22492 19317 22532
rect 19275 22483 19317 22492
rect 20043 22532 20085 22541
rect 20043 22492 20044 22532
rect 20084 22492 20085 22532
rect 20043 22483 20085 22492
rect 23787 22532 23829 22541
rect 23787 22492 23788 22532
rect 23828 22492 23829 22532
rect 23787 22483 23829 22492
rect 24459 22532 24501 22541
rect 24459 22492 24460 22532
rect 24500 22492 24501 22532
rect 24459 22483 24501 22492
rect 26083 22532 26141 22533
rect 26083 22492 26092 22532
rect 26132 22492 26141 22532
rect 26083 22491 26141 22492
rect 30699 22532 30741 22541
rect 30699 22492 30700 22532
rect 30740 22492 30741 22532
rect 30699 22483 30741 22492
rect 33955 22532 34013 22533
rect 33955 22492 33964 22532
rect 34004 22492 34013 22532
rect 33955 22491 34013 22492
rect 36835 22532 36893 22533
rect 36835 22492 36844 22532
rect 36884 22492 36893 22532
rect 36835 22491 36893 22492
rect 40683 22532 40725 22541
rect 40683 22492 40684 22532
rect 40724 22492 40725 22532
rect 40683 22483 40725 22492
rect 44715 22532 44757 22541
rect 44715 22492 44716 22532
rect 44756 22492 44757 22532
rect 44715 22483 44757 22492
rect 45763 22532 45821 22533
rect 45763 22492 45772 22532
rect 45812 22492 45821 22532
rect 45763 22491 45821 22492
rect 49131 22532 49173 22541
rect 49131 22492 49132 22532
rect 49172 22492 49173 22532
rect 49131 22483 49173 22492
rect 7083 22448 7125 22457
rect 7083 22408 7084 22448
rect 7124 22408 7125 22448
rect 7083 22399 7125 22408
rect 13995 22448 14037 22457
rect 13995 22408 13996 22448
rect 14036 22408 14037 22448
rect 13995 22399 14037 22408
rect 15723 22448 15765 22457
rect 15723 22408 15724 22448
rect 15764 22408 15765 22448
rect 15723 22399 15765 22408
rect 18507 22448 18549 22457
rect 18507 22408 18508 22448
rect 18548 22408 18549 22448
rect 18507 22399 18549 22408
rect 21675 22448 21717 22457
rect 21675 22408 21676 22448
rect 21716 22408 21717 22448
rect 21675 22399 21717 22408
rect 24651 22448 24693 22457
rect 24651 22408 24652 22448
rect 24692 22408 24693 22448
rect 24651 22399 24693 22408
rect 37323 22448 37365 22457
rect 37323 22408 37324 22448
rect 37364 22408 37365 22448
rect 37323 22399 37365 22408
rect 46155 22448 46197 22457
rect 46155 22408 46156 22448
rect 46196 22408 46197 22448
rect 46155 22399 46197 22408
rect 3627 22364 3669 22373
rect 3627 22324 3628 22364
rect 3668 22324 3669 22364
rect 3627 22315 3669 22324
rect 8235 22364 8277 22373
rect 8235 22324 8236 22364
rect 8276 22324 8277 22364
rect 8235 22315 8277 22324
rect 29163 22364 29205 22373
rect 29163 22324 29164 22364
rect 29204 22324 29205 22364
rect 29163 22315 29205 22324
rect 1227 22280 1269 22289
rect 1227 22240 1228 22280
rect 1268 22240 1269 22280
rect 1227 22231 1269 22240
rect 1603 22280 1661 22281
rect 1603 22240 1612 22280
rect 1652 22240 1661 22280
rect 1603 22239 1661 22240
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2467 22239 2525 22240
rect 3915 22280 3957 22289
rect 3915 22240 3916 22280
rect 3956 22240 3957 22280
rect 3915 22231 3957 22240
rect 4011 22280 4053 22289
rect 4011 22240 4012 22280
rect 4052 22240 4053 22280
rect 4011 22231 4053 22240
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 4291 22280 4349 22281
rect 4291 22240 4300 22280
rect 4340 22240 4349 22280
rect 4291 22239 4349 22240
rect 5155 22280 5213 22281
rect 5155 22240 5164 22280
rect 5204 22240 5213 22280
rect 5155 22239 5213 22240
rect 6027 22280 6069 22289
rect 6027 22240 6028 22280
rect 6068 22240 6069 22280
rect 6027 22231 6069 22240
rect 6411 22280 6453 22289
rect 6411 22240 6412 22280
rect 6452 22240 6453 22280
rect 6411 22231 6453 22240
rect 6507 22280 6549 22289
rect 6507 22240 6508 22280
rect 6548 22240 6549 22280
rect 6507 22231 6549 22240
rect 6603 22280 6645 22289
rect 6603 22240 6604 22280
rect 6644 22240 6645 22280
rect 6603 22231 6645 22240
rect 7363 22280 7421 22281
rect 7363 22240 7372 22280
rect 7412 22240 7421 22280
rect 7363 22239 7421 22240
rect 9379 22280 9437 22281
rect 9379 22240 9388 22280
rect 9428 22240 9437 22280
rect 9379 22239 9437 22240
rect 9571 22280 9629 22281
rect 9571 22240 9580 22280
rect 9620 22240 9629 22280
rect 9571 22239 9629 22240
rect 10627 22280 10685 22281
rect 10627 22240 10636 22280
rect 10676 22240 10685 22280
rect 10627 22239 10685 22240
rect 10923 22280 10965 22289
rect 10923 22240 10924 22280
rect 10964 22240 10965 22280
rect 10923 22231 10965 22240
rect 11019 22280 11061 22289
rect 11019 22240 11020 22280
rect 11060 22240 11061 22280
rect 11019 22231 11061 22240
rect 12067 22280 12125 22281
rect 12067 22240 12076 22280
rect 12116 22240 12125 22280
rect 12067 22239 12125 22240
rect 12939 22280 12981 22289
rect 12939 22240 12940 22280
rect 12980 22240 12981 22280
rect 12939 22231 12981 22240
rect 13515 22280 13557 22289
rect 13515 22240 13516 22280
rect 13556 22240 13557 22280
rect 13515 22231 13557 22240
rect 13611 22280 13653 22289
rect 13611 22240 13612 22280
rect 13652 22240 13653 22280
rect 13611 22231 13653 22240
rect 13707 22280 13749 22289
rect 13707 22240 13708 22280
rect 13748 22240 13749 22280
rect 13707 22231 13749 22240
rect 13803 22280 13845 22289
rect 13803 22240 13804 22280
rect 13844 22240 13845 22280
rect 13803 22231 13845 22240
rect 14563 22280 14621 22281
rect 14563 22240 14572 22280
rect 14612 22240 14621 22280
rect 14563 22239 14621 22240
rect 15523 22280 15581 22281
rect 15523 22240 15532 22280
rect 15572 22240 15581 22280
rect 15523 22239 15581 22240
rect 16099 22280 16157 22281
rect 16099 22240 16108 22280
rect 16148 22240 16157 22280
rect 16099 22239 16157 22240
rect 17155 22280 17213 22281
rect 17155 22240 17164 22280
rect 17204 22240 17213 22280
rect 17155 22239 17213 22240
rect 18123 22280 18165 22289
rect 18123 22240 18124 22280
rect 18164 22240 18165 22280
rect 18123 22231 18165 22240
rect 18219 22280 18261 22289
rect 18219 22240 18220 22280
rect 18260 22240 18261 22280
rect 18219 22231 18261 22240
rect 18315 22280 18357 22289
rect 18315 22240 18316 22280
rect 18356 22240 18357 22280
rect 18315 22231 18357 22240
rect 18883 22280 18941 22281
rect 18883 22240 18892 22280
rect 18932 22240 18941 22280
rect 18883 22239 18941 22240
rect 19171 22280 19229 22281
rect 19171 22240 19180 22280
rect 19220 22240 19229 22280
rect 19171 22239 19229 22240
rect 19939 22280 19997 22281
rect 19939 22240 19948 22280
rect 19988 22240 19997 22280
rect 19939 22239 19997 22240
rect 23115 22280 23157 22289
rect 23115 22240 23116 22280
rect 23156 22240 23157 22280
rect 23115 22231 23157 22240
rect 23299 22280 23357 22281
rect 23299 22240 23308 22280
rect 23348 22240 23357 22280
rect 23299 22239 23357 22240
rect 23491 22280 23549 22281
rect 23491 22240 23500 22280
rect 23540 22240 23549 22280
rect 23491 22239 23549 22240
rect 23595 22280 23637 22289
rect 23595 22240 23596 22280
rect 23636 22240 23637 22280
rect 23595 22231 23637 22240
rect 23787 22280 23829 22289
rect 23787 22240 23788 22280
rect 23828 22240 23829 22280
rect 23787 22231 23829 22240
rect 23979 22280 24021 22289
rect 23979 22240 23980 22280
rect 24020 22240 24021 22280
rect 23979 22231 24021 22240
rect 24171 22280 24213 22289
rect 24171 22240 24172 22280
rect 24212 22240 24213 22280
rect 24171 22231 24213 22240
rect 24259 22280 24317 22281
rect 24259 22240 24268 22280
rect 24308 22240 24317 22280
rect 24259 22239 24317 22240
rect 24651 22280 24693 22289
rect 24651 22240 24652 22280
rect 24692 22240 24693 22280
rect 24651 22231 24693 22240
rect 24939 22280 24981 22289
rect 24939 22240 24940 22280
rect 24980 22240 24981 22280
rect 24939 22231 24981 22240
rect 25035 22280 25077 22289
rect 25035 22240 25036 22280
rect 25076 22240 25077 22280
rect 25035 22231 25077 22240
rect 25411 22280 25469 22281
rect 25411 22240 25420 22280
rect 25460 22240 25469 22280
rect 25411 22239 25469 22240
rect 27235 22280 27293 22281
rect 27235 22240 27244 22280
rect 27284 22240 27293 22280
rect 27235 22239 27293 22240
rect 27427 22280 27485 22281
rect 27427 22240 27436 22280
rect 27476 22240 27485 22280
rect 27427 22239 27485 22240
rect 28587 22280 28629 22289
rect 28587 22240 28588 22280
rect 28628 22240 28629 22280
rect 28587 22231 28629 22240
rect 28683 22280 28725 22289
rect 28683 22240 28684 22280
rect 28724 22240 28725 22280
rect 28683 22231 28725 22240
rect 28779 22280 28821 22289
rect 28779 22240 28780 22280
rect 28820 22240 28821 22280
rect 28779 22231 28821 22240
rect 28875 22280 28917 22289
rect 28875 22240 28876 22280
rect 28916 22240 28917 22280
rect 28875 22231 28917 22240
rect 29931 22280 29973 22289
rect 29931 22240 29932 22280
rect 29972 22240 29973 22280
rect 29931 22231 29973 22240
rect 30403 22280 30461 22281
rect 30403 22240 30412 22280
rect 30452 22240 30461 22280
rect 30403 22239 30461 22240
rect 31563 22280 31605 22289
rect 31563 22240 31564 22280
rect 31604 22240 31605 22280
rect 31563 22231 31605 22240
rect 31939 22280 31997 22281
rect 31939 22240 31948 22280
rect 31988 22240 31997 22280
rect 31939 22239 31997 22240
rect 32803 22280 32861 22281
rect 32803 22240 32812 22280
rect 32852 22240 32861 22280
rect 32803 22239 32861 22240
rect 34443 22280 34485 22289
rect 34443 22240 34444 22280
rect 34484 22240 34485 22280
rect 34443 22231 34485 22240
rect 34819 22280 34877 22281
rect 34819 22240 34828 22280
rect 34868 22240 34877 22280
rect 34819 22239 34877 22240
rect 35683 22280 35741 22281
rect 35683 22240 35692 22280
rect 35732 22240 35741 22280
rect 35683 22239 35741 22240
rect 37507 22280 37565 22281
rect 37507 22240 37516 22280
rect 37556 22240 37565 22280
rect 37507 22239 37565 22240
rect 38571 22280 38613 22289
rect 38571 22240 38572 22280
rect 38612 22240 38613 22280
rect 38571 22231 38613 22240
rect 38667 22280 38709 22289
rect 38667 22240 38668 22280
rect 38708 22240 38709 22280
rect 38667 22231 38709 22240
rect 38763 22280 38805 22289
rect 38763 22240 38764 22280
rect 38804 22240 38805 22280
rect 38763 22231 38805 22240
rect 38947 22280 39005 22281
rect 38947 22240 38956 22280
rect 38996 22240 39005 22280
rect 38947 22239 39005 22240
rect 39051 22280 39093 22289
rect 39051 22240 39052 22280
rect 39092 22240 39093 22280
rect 39051 22231 39093 22240
rect 39243 22280 39285 22289
rect 39243 22240 39244 22280
rect 39284 22240 39285 22280
rect 39243 22231 39285 22240
rect 40099 22280 40157 22281
rect 40099 22240 40108 22280
rect 40148 22240 40157 22280
rect 40099 22239 40157 22240
rect 40387 22280 40445 22281
rect 40387 22240 40396 22280
rect 40436 22240 40445 22280
rect 40387 22239 40445 22240
rect 41347 22280 41405 22281
rect 41347 22240 41356 22280
rect 41396 22240 41405 22280
rect 41347 22239 41405 22240
rect 41643 22280 41685 22289
rect 41643 22240 41644 22280
rect 41684 22240 41685 22280
rect 41643 22231 41685 22240
rect 41739 22280 41781 22289
rect 41739 22240 41740 22280
rect 41780 22240 41781 22280
rect 41739 22231 41781 22240
rect 41835 22280 41877 22289
rect 41835 22240 41836 22280
rect 41876 22240 41877 22280
rect 41835 22231 41877 22240
rect 42027 22280 42069 22289
rect 42027 22240 42028 22280
rect 42068 22240 42069 22280
rect 42027 22231 42069 22240
rect 42115 22280 42173 22281
rect 42115 22240 42124 22280
rect 42164 22240 42173 22280
rect 42115 22239 42173 22240
rect 42315 22280 42357 22289
rect 42315 22240 42316 22280
rect 42356 22240 42357 22280
rect 42315 22231 42357 22240
rect 42691 22280 42749 22281
rect 42691 22240 42700 22280
rect 42740 22240 42749 22280
rect 42691 22239 42749 22240
rect 43555 22280 43613 22281
rect 43555 22240 43564 22280
rect 43604 22240 43613 22280
rect 43555 22239 43613 22240
rect 45091 22280 45149 22281
rect 45091 22240 45100 22280
rect 45140 22240 45149 22280
rect 45091 22239 45149 22240
rect 46731 22280 46773 22289
rect 46731 22240 46732 22280
rect 46772 22240 46773 22280
rect 46731 22231 46773 22240
rect 47107 22280 47165 22281
rect 47107 22240 47116 22280
rect 47156 22240 47165 22280
rect 47107 22239 47165 22240
rect 47971 22280 48029 22281
rect 47971 22240 47980 22280
rect 48020 22240 48029 22280
rect 47971 22239 48029 22240
rect 23211 22196 23253 22205
rect 23211 22156 23212 22196
rect 23252 22156 23253 22196
rect 23211 22147 23253 22156
rect 643 22112 701 22113
rect 643 22072 652 22112
rect 692 22072 701 22112
rect 643 22071 701 22072
rect 3811 22112 3869 22113
rect 3811 22072 3820 22112
rect 3860 22072 3869 22112
rect 3811 22071 3869 22072
rect 6691 22112 6749 22113
rect 6691 22072 6700 22112
rect 6740 22072 6749 22112
rect 6691 22071 6749 22072
rect 10243 22112 10301 22113
rect 10243 22072 10252 22112
rect 10292 22072 10301 22112
rect 10243 22071 10301 22072
rect 16771 22112 16829 22113
rect 16771 22072 16780 22112
rect 16820 22072 16829 22112
rect 16771 22071 16829 22072
rect 17827 22112 17885 22113
rect 17827 22072 17836 22112
rect 17876 22072 17885 22112
rect 17827 22071 17885 22072
rect 18019 22112 18077 22113
rect 18019 22072 18028 22112
rect 18068 22072 18077 22112
rect 18019 22071 18077 22072
rect 18987 22112 19029 22121
rect 18987 22072 18988 22112
rect 19028 22072 19029 22112
rect 18987 22063 19029 22072
rect 24067 22112 24125 22113
rect 24067 22072 24076 22112
rect 24116 22072 24125 22112
rect 24067 22071 24125 22072
rect 25219 22112 25277 22113
rect 25219 22072 25228 22112
rect 25268 22072 25277 22112
rect 25219 22071 25277 22072
rect 26083 22112 26141 22113
rect 26083 22072 26092 22112
rect 26132 22072 26141 22112
rect 26083 22071 26141 22072
rect 26563 22112 26621 22113
rect 26563 22072 26572 22112
rect 26612 22072 26621 22112
rect 26563 22071 26621 22072
rect 28099 22112 28157 22113
rect 28099 22072 28108 22112
rect 28148 22072 28157 22112
rect 28099 22071 28157 22072
rect 30891 22112 30933 22121
rect 30891 22072 30892 22112
rect 30932 22072 30933 22112
rect 30891 22063 30933 22072
rect 38179 22112 38237 22113
rect 38179 22072 38188 22112
rect 38228 22072 38237 22112
rect 38179 22071 38237 22072
rect 38467 22112 38525 22113
rect 38467 22072 38476 22112
rect 38516 22072 38525 22112
rect 38467 22071 38525 22072
rect 39139 22112 39197 22113
rect 39139 22072 39148 22112
rect 39188 22072 39197 22112
rect 39139 22071 39197 22072
rect 39427 22112 39485 22113
rect 39427 22072 39436 22112
rect 39476 22072 39485 22112
rect 39427 22071 39485 22072
rect 41539 22112 41597 22113
rect 41539 22072 41548 22112
rect 41588 22072 41597 22112
rect 41539 22071 41597 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 4963 21776 5021 21777
rect 4963 21736 4972 21776
rect 5012 21736 5021 21776
rect 4963 21735 5021 21736
rect 8995 21776 9053 21777
rect 8995 21736 9004 21776
rect 9044 21736 9053 21776
rect 8995 21735 9053 21736
rect 9187 21776 9245 21777
rect 9187 21736 9196 21776
rect 9236 21736 9245 21776
rect 9187 21735 9245 21736
rect 15427 21776 15485 21777
rect 15427 21736 15436 21776
rect 15476 21736 15485 21776
rect 15427 21735 15485 21736
rect 16491 21776 16533 21785
rect 16491 21736 16492 21776
rect 16532 21736 16533 21776
rect 16491 21727 16533 21736
rect 19651 21776 19709 21777
rect 19651 21736 19660 21776
rect 19700 21736 19709 21776
rect 19651 21735 19709 21736
rect 25707 21776 25749 21785
rect 25707 21736 25708 21776
rect 25748 21736 25749 21776
rect 25707 21727 25749 21736
rect 27331 21776 27389 21777
rect 27331 21736 27340 21776
rect 27380 21736 27389 21776
rect 27331 21735 27389 21736
rect 30595 21776 30653 21777
rect 30595 21736 30604 21776
rect 30644 21736 30653 21776
rect 30595 21735 30653 21736
rect 36267 21776 36309 21785
rect 36267 21736 36268 21776
rect 36308 21736 36309 21776
rect 36267 21727 36309 21736
rect 36931 21776 36989 21777
rect 36931 21736 36940 21776
rect 36980 21736 36989 21776
rect 36931 21735 36989 21736
rect 45283 21776 45341 21777
rect 45283 21736 45292 21776
rect 45332 21736 45341 21776
rect 45283 21735 45341 21736
rect 2763 21692 2805 21701
rect 2763 21652 2764 21692
rect 2804 21652 2805 21692
rect 2763 21643 2805 21652
rect 11595 21692 11637 21701
rect 11595 21652 11596 21692
rect 11636 21652 11637 21692
rect 11595 21643 11637 21652
rect 13035 21692 13077 21701
rect 13035 21652 13036 21692
rect 13076 21652 13077 21692
rect 13035 21643 13077 21652
rect 17259 21692 17301 21701
rect 17259 21652 17260 21692
rect 17300 21652 17301 21692
rect 17259 21643 17301 21652
rect 25323 21692 25365 21701
rect 25323 21652 25324 21692
rect 25364 21652 25365 21692
rect 25323 21643 25365 21652
rect 28203 21692 28245 21701
rect 28203 21652 28204 21692
rect 28244 21652 28245 21692
rect 28203 21643 28245 21652
rect 39339 21692 39381 21701
rect 39339 21652 39340 21692
rect 39380 21652 39381 21692
rect 39339 21643 39381 21652
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 2859 21608 2901 21617
rect 2859 21568 2860 21608
rect 2900 21568 2901 21608
rect 2859 21559 2901 21568
rect 2947 21608 3005 21609
rect 2947 21568 2956 21608
rect 2996 21568 3005 21608
rect 2947 21567 3005 21568
rect 3139 21608 3197 21609
rect 3139 21568 3148 21608
rect 3188 21568 3197 21608
rect 3139 21567 3197 21568
rect 4099 21608 4157 21609
rect 4099 21568 4108 21608
rect 4148 21568 4157 21608
rect 4099 21567 4157 21568
rect 4491 21608 4533 21617
rect 4491 21568 4492 21608
rect 4532 21568 4533 21608
rect 4491 21559 4533 21568
rect 4683 21608 4725 21617
rect 4683 21568 4684 21608
rect 4724 21568 4725 21608
rect 4683 21559 4725 21568
rect 4771 21608 4829 21609
rect 4771 21568 4780 21608
rect 4820 21568 4829 21608
rect 4771 21567 4829 21568
rect 5067 21608 5109 21617
rect 5067 21568 5068 21608
rect 5108 21568 5109 21608
rect 5067 21559 5109 21568
rect 5163 21608 5205 21617
rect 5163 21568 5164 21608
rect 5204 21568 5205 21608
rect 5163 21559 5205 21568
rect 5259 21608 5301 21617
rect 5259 21568 5260 21608
rect 5300 21568 5301 21608
rect 5259 21559 5301 21568
rect 5539 21608 5597 21609
rect 5539 21568 5548 21608
rect 5588 21568 5597 21608
rect 5539 21567 5597 21568
rect 5731 21608 5789 21609
rect 5731 21568 5740 21608
rect 5780 21568 5789 21608
rect 5731 21567 5789 21568
rect 6411 21608 6453 21617
rect 6411 21568 6412 21608
rect 6452 21568 6453 21608
rect 6411 21559 6453 21568
rect 6603 21608 6645 21617
rect 6603 21568 6604 21608
rect 6644 21568 6645 21608
rect 6603 21559 6645 21568
rect 6979 21608 7037 21609
rect 6979 21568 6988 21608
rect 7028 21568 7037 21608
rect 6979 21567 7037 21568
rect 7843 21608 7901 21609
rect 7843 21568 7852 21608
rect 7892 21568 7901 21608
rect 7843 21567 7901 21568
rect 10339 21608 10397 21609
rect 10339 21568 10348 21608
rect 10388 21568 10397 21608
rect 10339 21567 10397 21568
rect 11203 21608 11261 21609
rect 11203 21568 11212 21608
rect 11252 21568 11261 21608
rect 11203 21567 11261 21568
rect 13411 21608 13469 21609
rect 13411 21568 13420 21608
rect 13460 21568 13469 21608
rect 13411 21567 13469 21568
rect 14275 21608 14333 21609
rect 14275 21568 14284 21608
rect 14324 21568 14333 21608
rect 14275 21567 14333 21568
rect 15627 21608 15669 21617
rect 15627 21568 15628 21608
rect 15668 21568 15669 21608
rect 15627 21559 15669 21568
rect 15715 21608 15773 21609
rect 15715 21568 15724 21608
rect 15764 21568 15773 21608
rect 15715 21567 15773 21568
rect 16875 21608 16917 21617
rect 16875 21568 16876 21608
rect 16916 21568 16917 21608
rect 16875 21559 16917 21568
rect 17635 21608 17693 21609
rect 17635 21568 17644 21608
rect 17684 21568 17693 21608
rect 17635 21567 17693 21568
rect 18499 21608 18557 21609
rect 18499 21568 18508 21608
rect 18548 21568 18557 21608
rect 18499 21567 18557 21568
rect 21195 21608 21237 21617
rect 21195 21568 21196 21608
rect 21236 21568 21237 21608
rect 21195 21559 21237 21568
rect 21571 21608 21629 21609
rect 21571 21568 21580 21608
rect 21620 21568 21629 21608
rect 21571 21567 21629 21568
rect 22435 21608 22493 21609
rect 22435 21568 22444 21608
rect 22484 21568 22493 21608
rect 22435 21567 22493 21568
rect 23683 21608 23741 21609
rect 23683 21568 23692 21608
rect 23732 21568 23741 21608
rect 23683 21567 23741 21568
rect 24355 21608 24413 21609
rect 24355 21568 24364 21608
rect 24404 21568 24413 21608
rect 24355 21567 24413 21568
rect 24459 21608 24501 21617
rect 24459 21568 24460 21608
rect 24500 21568 24501 21608
rect 24459 21559 24501 21568
rect 25227 21608 25269 21617
rect 25227 21568 25228 21608
rect 25268 21568 25269 21608
rect 25227 21559 25269 21568
rect 25411 21608 25469 21609
rect 25411 21568 25420 21608
rect 25460 21568 25469 21608
rect 25411 21567 25469 21568
rect 25611 21608 25653 21617
rect 25611 21568 25612 21608
rect 25652 21568 25653 21608
rect 25611 21559 25653 21568
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 25803 21559 25845 21568
rect 26083 21608 26141 21609
rect 26083 21568 26092 21608
rect 26132 21568 26141 21608
rect 26083 21567 26141 21568
rect 27043 21608 27101 21609
rect 27043 21568 27052 21608
rect 27092 21568 27101 21608
rect 27043 21567 27101 21568
rect 27531 21608 27573 21617
rect 27531 21568 27532 21608
rect 27572 21568 27573 21608
rect 27531 21559 27573 21568
rect 27627 21608 27669 21617
rect 27627 21568 27628 21608
rect 27668 21568 27669 21608
rect 27627 21559 27669 21568
rect 28579 21608 28637 21609
rect 28579 21568 28588 21608
rect 28628 21568 28637 21608
rect 28579 21567 28637 21568
rect 29443 21608 29501 21609
rect 29443 21568 29452 21608
rect 29492 21568 29501 21608
rect 29443 21567 29501 21568
rect 35779 21608 35837 21609
rect 35779 21568 35788 21608
rect 35828 21568 35837 21608
rect 35779 21567 35837 21568
rect 38083 21608 38141 21609
rect 38083 21568 38092 21608
rect 38132 21568 38141 21608
rect 38083 21567 38141 21568
rect 38947 21608 39005 21609
rect 38947 21568 38956 21608
rect 38996 21568 39005 21608
rect 38947 21567 39005 21568
rect 40291 21608 40349 21609
rect 40291 21568 40300 21608
rect 40340 21568 40349 21608
rect 40291 21567 40349 21568
rect 41155 21608 41213 21609
rect 41155 21568 41164 21608
rect 41204 21568 41213 21608
rect 41155 21567 41213 21568
rect 41443 21608 41501 21609
rect 41443 21568 41452 21608
rect 41492 21568 41501 21608
rect 41443 21567 41501 21568
rect 41635 21608 41693 21609
rect 41635 21568 41644 21608
rect 41684 21568 41693 21608
rect 41635 21567 41693 21568
rect 41739 21608 41781 21617
rect 41739 21568 41740 21608
rect 41780 21568 41781 21608
rect 41739 21559 41781 21568
rect 41931 21608 41973 21617
rect 41931 21568 41932 21608
rect 41972 21568 41973 21608
rect 41931 21559 41973 21568
rect 42115 21608 42173 21609
rect 42115 21568 42124 21608
rect 42164 21568 42173 21608
rect 42115 21567 42173 21568
rect 43267 21608 43325 21609
rect 43267 21568 43276 21608
rect 43316 21568 43325 21608
rect 43267 21567 43325 21568
rect 44427 21608 44469 21617
rect 44427 21568 44428 21608
rect 44468 21568 44469 21608
rect 44427 21559 44469 21568
rect 44515 21608 44573 21609
rect 44515 21568 44524 21608
rect 44564 21568 44573 21608
rect 44515 21567 44573 21568
rect 44715 21608 44757 21617
rect 44715 21568 44716 21608
rect 44756 21568 44757 21608
rect 44715 21559 44757 21568
rect 44811 21608 44853 21617
rect 44811 21568 44812 21608
rect 44852 21568 44853 21608
rect 44811 21559 44853 21568
rect 44907 21608 44949 21617
rect 44907 21568 44908 21608
rect 44948 21568 44949 21608
rect 44907 21559 44949 21568
rect 45003 21608 45045 21617
rect 45003 21568 45004 21608
rect 45044 21568 45045 21608
rect 45003 21559 45045 21568
rect 45195 21608 45237 21617
rect 45195 21568 45196 21608
rect 45236 21568 45237 21608
rect 45195 21559 45237 21568
rect 45387 21608 45429 21617
rect 45387 21568 45388 21608
rect 45428 21568 45429 21608
rect 45387 21559 45429 21568
rect 45475 21608 45533 21609
rect 45475 21568 45484 21608
rect 45524 21568 45533 21608
rect 45475 21567 45533 21568
rect 24835 21524 24893 21525
rect 24835 21484 24844 21524
rect 24884 21484 24893 21524
rect 24835 21483 24893 21484
rect 1707 21440 1749 21449
rect 1707 21400 1708 21440
rect 1748 21400 1749 21440
rect 1707 21391 1749 21400
rect 2187 21440 2229 21449
rect 2187 21400 2188 21440
rect 2228 21400 2229 21440
rect 2187 21391 2229 21400
rect 4491 21440 4533 21449
rect 4491 21400 4492 21440
rect 4532 21400 4533 21440
rect 4491 21391 4533 21400
rect 5451 21440 5493 21449
rect 5451 21400 5452 21440
rect 5492 21400 5493 21440
rect 5451 21391 5493 21400
rect 11787 21440 11829 21449
rect 11787 21400 11788 21440
rect 11828 21400 11829 21440
rect 11787 21391 11829 21400
rect 24171 21440 24213 21449
rect 24171 21400 24172 21440
rect 24212 21400 24213 21440
rect 24171 21391 24213 21400
rect 25035 21440 25077 21449
rect 25035 21400 25036 21440
rect 25076 21400 25077 21440
rect 25035 21391 25077 21400
rect 28011 21440 28053 21449
rect 28011 21400 28012 21440
rect 28052 21400 28053 21440
rect 28011 21391 28053 21400
rect 34923 21440 34965 21449
rect 34923 21400 34924 21440
rect 34964 21400 34965 21440
rect 34923 21391 34965 21400
rect 41931 21440 41973 21449
rect 41931 21400 41932 21440
rect 41972 21400 41973 21440
rect 41931 21391 41973 21400
rect 43563 21440 43605 21449
rect 43563 21400 43564 21440
rect 43604 21400 43605 21440
rect 43563 21391 43605 21400
rect 39619 21356 39677 21357
rect 39619 21316 39628 21356
rect 39668 21316 39677 21356
rect 39619 21315 39677 21316
rect 40483 21356 40541 21357
rect 40483 21316 40492 21356
rect 40532 21316 40541 21356
rect 40483 21315 40541 21316
rect 41355 21356 41397 21365
rect 41355 21316 41356 21356
rect 41396 21316 41397 21356
rect 41355 21307 41397 21316
rect 42787 21356 42845 21357
rect 42787 21316 42796 21356
rect 42836 21316 42845 21356
rect 42787 21315 42845 21316
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 4099 21020 4157 21021
rect 4099 20980 4108 21020
rect 4148 20980 4157 21020
rect 4099 20979 4157 20980
rect 5923 21020 5981 21021
rect 5923 20980 5932 21020
rect 5972 20980 5981 21020
rect 5923 20979 5981 20980
rect 6211 21020 6269 21021
rect 6211 20980 6220 21020
rect 6260 20980 6269 21020
rect 6211 20979 6269 20980
rect 11683 21020 11741 21021
rect 11683 20980 11692 21020
rect 11732 20980 11741 21020
rect 11683 20979 11741 20980
rect 16971 21020 17013 21029
rect 16971 20980 16972 21020
rect 17012 20980 17013 21020
rect 16971 20971 17013 20980
rect 33771 21020 33813 21029
rect 33771 20980 33772 21020
rect 33812 20980 33813 21020
rect 33771 20971 33813 20980
rect 37227 21020 37269 21029
rect 37227 20980 37228 21020
rect 37268 20980 37269 21020
rect 37227 20971 37269 20980
rect 37803 21020 37845 21029
rect 37803 20980 37804 21020
rect 37844 20980 37845 21020
rect 37803 20971 37845 20980
rect 38955 21020 38997 21029
rect 38955 20980 38956 21020
rect 38996 20980 38997 21020
rect 38955 20971 38997 20980
rect 44619 21020 44661 21029
rect 44619 20980 44620 21020
rect 44660 20980 44661 21020
rect 44619 20971 44661 20980
rect 16107 20936 16149 20945
rect 16107 20896 16108 20936
rect 16148 20896 16149 20936
rect 16107 20887 16149 20896
rect 25035 20936 25077 20945
rect 25035 20896 25036 20936
rect 25076 20896 25077 20936
rect 25035 20887 25077 20896
rect 27627 20936 27669 20945
rect 27627 20896 27628 20936
rect 27668 20896 27669 20936
rect 27627 20887 27669 20896
rect 29067 20936 29109 20945
rect 29067 20896 29068 20936
rect 29108 20896 29109 20936
rect 29067 20887 29109 20896
rect 34827 20936 34869 20945
rect 34827 20896 34828 20936
rect 34868 20896 34869 20936
rect 34827 20887 34869 20896
rect 13227 20852 13269 20861
rect 13227 20812 13228 20852
rect 13268 20812 13269 20852
rect 13227 20803 13269 20812
rect 17259 20852 17301 20861
rect 17259 20812 17260 20852
rect 17300 20812 17301 20852
rect 17259 20803 17301 20812
rect 21291 20852 21333 20861
rect 21291 20812 21292 20852
rect 21332 20812 21333 20852
rect 21291 20803 21333 20812
rect 25707 20852 25749 20861
rect 25707 20812 25708 20852
rect 25748 20812 25749 20852
rect 25707 20803 25749 20812
rect 41643 20852 41685 20861
rect 41643 20812 41644 20852
rect 41684 20812 41685 20852
rect 41643 20803 41685 20812
rect 20131 20779 20189 20780
rect 1707 20768 1749 20777
rect 1707 20728 1708 20768
rect 1748 20728 1749 20768
rect 1707 20719 1749 20728
rect 2083 20768 2141 20769
rect 2083 20728 2092 20768
rect 2132 20728 2141 20768
rect 2083 20727 2141 20728
rect 2947 20768 3005 20769
rect 2947 20728 2956 20768
rect 2996 20728 3005 20768
rect 2947 20727 3005 20728
rect 5059 20768 5117 20769
rect 5059 20728 5068 20768
rect 5108 20728 5117 20768
rect 5059 20727 5117 20728
rect 5251 20768 5309 20769
rect 5251 20728 5260 20768
rect 5300 20728 5309 20768
rect 5251 20727 5309 20728
rect 6883 20768 6941 20769
rect 6883 20728 6892 20768
rect 6932 20728 6941 20768
rect 6883 20727 6941 20728
rect 7363 20768 7421 20769
rect 7363 20728 7372 20768
rect 7412 20728 7421 20768
rect 7363 20727 7421 20728
rect 8803 20768 8861 20769
rect 8803 20728 8812 20768
rect 8852 20728 8861 20768
rect 8803 20727 8861 20728
rect 8995 20768 9053 20769
rect 8995 20728 9004 20768
rect 9044 20728 9053 20768
rect 8995 20727 9053 20728
rect 9283 20768 9341 20769
rect 9283 20728 9292 20768
rect 9332 20728 9341 20768
rect 9283 20727 9341 20728
rect 9579 20768 9621 20777
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 9675 20768 9717 20777
rect 9675 20728 9676 20768
rect 9716 20728 9717 20768
rect 9675 20719 9717 20728
rect 9771 20768 9813 20777
rect 9771 20728 9772 20768
rect 9812 20728 9813 20768
rect 9771 20719 9813 20728
rect 9867 20768 9909 20777
rect 9867 20728 9868 20768
rect 9908 20728 9909 20768
rect 9867 20719 9909 20728
rect 10347 20768 10389 20777
rect 10347 20728 10348 20768
rect 10388 20728 10389 20768
rect 10347 20719 10389 20728
rect 10539 20768 10581 20777
rect 10539 20728 10540 20768
rect 10580 20728 10581 20768
rect 10539 20719 10581 20728
rect 10627 20768 10685 20769
rect 10627 20728 10636 20768
rect 10676 20728 10685 20768
rect 10627 20727 10685 20728
rect 11491 20768 11549 20769
rect 11491 20728 11500 20768
rect 11540 20728 11549 20768
rect 11491 20727 11549 20728
rect 12075 20768 12117 20777
rect 12075 20728 12076 20768
rect 12116 20728 12117 20768
rect 12075 20719 12117 20728
rect 12355 20768 12413 20769
rect 12355 20728 12364 20768
rect 12404 20728 12413 20768
rect 12355 20727 12413 20728
rect 13995 20768 14037 20777
rect 13995 20728 13996 20768
rect 14036 20728 14037 20768
rect 13995 20719 14037 20728
rect 15147 20768 15189 20777
rect 15147 20728 15148 20768
rect 15188 20728 15189 20768
rect 15147 20719 15189 20728
rect 15339 20768 15381 20777
rect 15339 20728 15340 20768
rect 15380 20728 15381 20768
rect 15339 20719 15381 20728
rect 15427 20768 15485 20769
rect 15427 20728 15436 20768
rect 15476 20728 15485 20768
rect 15427 20727 15485 20728
rect 15627 20768 15669 20777
rect 15627 20728 15628 20768
rect 15668 20728 15669 20768
rect 15627 20719 15669 20728
rect 15723 20768 15765 20777
rect 15723 20728 15724 20768
rect 15764 20728 15765 20768
rect 15723 20719 15765 20728
rect 15819 20768 15861 20777
rect 15819 20728 15820 20768
rect 15860 20728 15861 20768
rect 15819 20719 15861 20728
rect 15915 20768 15957 20777
rect 15915 20728 15916 20768
rect 15956 20728 15957 20768
rect 15915 20719 15957 20728
rect 16675 20768 16733 20769
rect 16675 20728 16684 20768
rect 16724 20728 16733 20768
rect 16675 20727 16733 20728
rect 16779 20768 16821 20777
rect 16779 20728 16780 20768
rect 16820 20728 16821 20768
rect 16779 20719 16821 20728
rect 16971 20768 17013 20777
rect 16971 20728 16972 20768
rect 17012 20728 17013 20768
rect 16971 20719 17013 20728
rect 18115 20768 18173 20769
rect 18115 20728 18124 20768
rect 18164 20728 18173 20768
rect 18115 20727 18173 20728
rect 19267 20768 19325 20769
rect 19267 20728 19276 20768
rect 19316 20728 19325 20768
rect 20131 20739 20140 20779
rect 20180 20739 20189 20779
rect 20131 20738 20189 20739
rect 22147 20768 22205 20769
rect 19267 20727 19325 20728
rect 22147 20728 22156 20768
rect 22196 20728 22205 20768
rect 22147 20727 22205 20728
rect 22347 20768 22389 20777
rect 22347 20728 22348 20768
rect 22388 20728 22389 20768
rect 22347 20719 22389 20728
rect 22443 20768 22485 20777
rect 22443 20728 22444 20768
rect 22484 20728 22485 20768
rect 22443 20719 22485 20728
rect 22539 20768 22581 20777
rect 22539 20728 22540 20768
rect 22580 20728 22581 20768
rect 22539 20719 22581 20728
rect 24459 20768 24501 20777
rect 24459 20728 24460 20768
rect 24500 20728 24501 20768
rect 24459 20719 24501 20728
rect 26563 20768 26621 20769
rect 26563 20728 26572 20768
rect 26612 20728 26621 20768
rect 26563 20727 26621 20728
rect 26947 20768 27005 20769
rect 26947 20728 26956 20768
rect 26996 20728 27005 20768
rect 26947 20727 27005 20728
rect 33283 20768 33341 20769
rect 33283 20728 33292 20768
rect 33332 20728 33341 20768
rect 33283 20727 33341 20728
rect 35403 20768 35445 20777
rect 35403 20728 35404 20768
rect 35444 20728 35445 20768
rect 35403 20719 35445 20728
rect 35499 20768 35541 20777
rect 35499 20728 35500 20768
rect 35540 20728 35541 20768
rect 35499 20719 35541 20728
rect 35595 20768 35637 20777
rect 35595 20728 35596 20768
rect 35636 20728 35637 20768
rect 35595 20719 35637 20728
rect 37123 20768 37181 20769
rect 37123 20728 37132 20768
rect 37172 20728 37181 20768
rect 37123 20727 37181 20728
rect 37891 20768 37949 20769
rect 37891 20728 37900 20768
rect 37940 20728 37949 20768
rect 37891 20727 37949 20728
rect 39043 20768 39101 20769
rect 39043 20728 39052 20768
rect 39092 20728 39101 20768
rect 39043 20727 39101 20728
rect 39243 20768 39285 20777
rect 39243 20728 39244 20768
rect 39284 20728 39285 20768
rect 39243 20719 39285 20728
rect 39619 20768 39677 20769
rect 39619 20728 39628 20768
rect 39668 20728 39677 20768
rect 39619 20727 39677 20728
rect 40483 20768 40541 20769
rect 40483 20728 40492 20768
rect 40532 20728 40541 20768
rect 40483 20727 40541 20728
rect 42219 20768 42261 20777
rect 42219 20728 42220 20768
rect 42260 20728 42261 20768
rect 42219 20719 42261 20728
rect 42595 20768 42653 20769
rect 42595 20728 42604 20768
rect 42644 20728 42653 20768
rect 42595 20727 42653 20728
rect 43459 20768 43517 20769
rect 43459 20728 43468 20768
rect 43508 20728 43517 20768
rect 43459 20727 43517 20728
rect 10827 20684 10869 20693
rect 10827 20644 10828 20684
rect 10868 20644 10869 20684
rect 10827 20635 10869 20644
rect 11979 20684 12021 20693
rect 11979 20644 11980 20684
rect 12020 20644 12021 20684
rect 11979 20635 12021 20644
rect 18891 20684 18933 20693
rect 18891 20644 18892 20684
rect 18932 20644 18933 20684
rect 18891 20635 18933 20644
rect 643 20600 701 20601
rect 643 20560 652 20600
rect 692 20560 701 20600
rect 643 20559 701 20560
rect 4387 20600 4445 20601
rect 4387 20560 4396 20600
rect 4436 20560 4445 20600
rect 4387 20559 4445 20560
rect 7851 20600 7893 20609
rect 7851 20560 7852 20600
rect 7892 20560 7893 20600
rect 7851 20551 7893 20560
rect 9195 20600 9237 20609
rect 9195 20560 9196 20600
rect 9236 20560 9237 20600
rect 9195 20551 9237 20560
rect 10435 20600 10493 20601
rect 10435 20560 10444 20600
rect 10484 20560 10493 20600
rect 10435 20559 10493 20560
rect 15235 20600 15293 20601
rect 15235 20560 15244 20600
rect 15284 20560 15293 20600
rect 15235 20559 15293 20560
rect 21475 20600 21533 20601
rect 21475 20560 21484 20600
rect 21524 20560 21533 20600
rect 21475 20559 21533 20560
rect 22627 20600 22685 20601
rect 22627 20560 22636 20600
rect 22676 20560 22685 20600
rect 22627 20559 22685 20560
rect 33771 20600 33813 20609
rect 33771 20560 33772 20600
rect 33812 20560 33813 20600
rect 33771 20551 33813 20560
rect 35299 20600 35357 20601
rect 35299 20560 35308 20600
rect 35348 20560 35357 20600
rect 35299 20559 35357 20560
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 21099 20322 21141 20331
rect 21099 20282 21100 20322
rect 21140 20282 21141 20322
rect 21099 20273 21141 20282
rect 643 20264 701 20265
rect 643 20224 652 20264
rect 692 20224 701 20264
rect 643 20223 701 20224
rect 6499 20264 6557 20265
rect 6499 20224 6508 20264
rect 6548 20224 6557 20264
rect 6499 20223 6557 20224
rect 21763 20264 21821 20265
rect 21763 20224 21772 20264
rect 21812 20224 21821 20264
rect 21763 20223 21821 20224
rect 21955 20264 22013 20265
rect 21955 20224 21964 20264
rect 22004 20224 22013 20264
rect 21955 20223 22013 20224
rect 4107 20180 4149 20189
rect 4107 20140 4108 20180
rect 4148 20140 4149 20180
rect 4107 20131 4149 20140
rect 15627 20180 15669 20189
rect 15627 20140 15628 20180
rect 15668 20140 15669 20180
rect 15627 20131 15669 20140
rect 19755 20180 19797 20189
rect 19755 20140 19756 20180
rect 19796 20140 19797 20180
rect 19755 20131 19797 20140
rect 21475 20180 21533 20181
rect 21475 20140 21484 20180
rect 21524 20140 21533 20180
rect 21475 20139 21533 20140
rect 26667 20180 26709 20189
rect 26667 20140 26668 20180
rect 26708 20140 26709 20180
rect 26667 20131 26709 20140
rect 39723 20180 39765 20189
rect 39723 20140 39724 20180
rect 39764 20140 39765 20180
rect 39723 20131 39765 20140
rect 4483 20096 4541 20097
rect 4483 20056 4492 20096
rect 4532 20056 4541 20096
rect 4483 20055 4541 20056
rect 5347 20096 5405 20097
rect 5347 20056 5356 20096
rect 5396 20056 5405 20096
rect 5347 20055 5405 20056
rect 6795 20096 6837 20105
rect 6795 20056 6796 20096
rect 6836 20056 6837 20096
rect 6795 20047 6837 20056
rect 6987 20096 7029 20105
rect 6987 20056 6988 20096
rect 7028 20056 7029 20096
rect 6987 20047 7029 20056
rect 7075 20096 7133 20097
rect 7075 20056 7084 20096
rect 7124 20056 7133 20096
rect 7075 20055 7133 20056
rect 7651 20096 7709 20097
rect 7651 20056 7660 20096
rect 7700 20056 7709 20096
rect 7651 20055 7709 20056
rect 9291 20096 9333 20105
rect 9291 20056 9292 20096
rect 9332 20056 9333 20096
rect 9291 20047 9333 20056
rect 10147 20096 10205 20097
rect 10147 20056 10156 20096
rect 10196 20056 10205 20096
rect 10147 20055 10205 20056
rect 10443 20096 10485 20105
rect 10443 20056 10444 20096
rect 10484 20056 10485 20096
rect 10443 20047 10485 20056
rect 10819 20096 10877 20097
rect 10819 20056 10828 20096
rect 10868 20056 10877 20096
rect 10819 20055 10877 20056
rect 11683 20096 11741 20097
rect 11683 20056 11692 20096
rect 11732 20056 11741 20096
rect 11683 20055 11741 20056
rect 12931 20096 12989 20097
rect 12931 20056 12940 20096
rect 12980 20056 12989 20096
rect 12931 20055 12989 20056
rect 15427 20096 15485 20097
rect 15427 20056 15436 20096
rect 15476 20056 15485 20096
rect 15427 20055 15485 20056
rect 16291 20096 16349 20097
rect 16291 20056 16300 20096
rect 16340 20056 16349 20096
rect 16291 20055 16349 20056
rect 16683 20096 16725 20105
rect 16683 20056 16684 20096
rect 16724 20056 16725 20096
rect 16683 20047 16725 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19371 20096 19413 20105
rect 19371 20056 19372 20096
rect 19412 20056 19413 20096
rect 19371 20047 19413 20056
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19563 20096 19605 20105
rect 19563 20056 19564 20096
rect 19604 20056 19605 20096
rect 19563 20047 19605 20056
rect 20419 20096 20477 20097
rect 20419 20056 20428 20096
rect 20468 20056 20477 20096
rect 20419 20055 20477 20056
rect 20907 20096 20949 20105
rect 20907 20056 20908 20096
rect 20948 20056 20949 20096
rect 20907 20047 20949 20056
rect 20995 20096 21053 20097
rect 20995 20056 21004 20096
rect 21044 20056 21053 20096
rect 20995 20055 21053 20056
rect 21667 20096 21725 20097
rect 21667 20056 21676 20096
rect 21716 20056 21725 20096
rect 21667 20055 21725 20056
rect 22155 20096 22197 20105
rect 22155 20056 22156 20096
rect 22196 20056 22197 20096
rect 22155 20047 22197 20056
rect 22251 20096 22293 20105
rect 22251 20056 22252 20096
rect 22292 20056 22293 20096
rect 22251 20047 22293 20056
rect 23299 20096 23357 20097
rect 23299 20056 23308 20096
rect 23348 20056 23357 20096
rect 23299 20055 23357 20056
rect 24075 20096 24117 20105
rect 24075 20056 24076 20096
rect 24116 20056 24117 20096
rect 24075 20047 24117 20056
rect 24259 20096 24317 20097
rect 24259 20056 24268 20096
rect 24308 20056 24317 20096
rect 24259 20055 24317 20056
rect 24843 20096 24885 20105
rect 24843 20056 24844 20096
rect 24884 20056 24885 20096
rect 25411 20104 25469 20105
rect 25411 20064 25420 20104
rect 25460 20064 25469 20104
rect 25411 20063 25469 20064
rect 25803 20096 25845 20105
rect 24843 20047 24885 20056
rect 25803 20056 25804 20096
rect 25844 20056 25845 20096
rect 25803 20047 25845 20056
rect 26083 20096 26141 20097
rect 26083 20056 26092 20096
rect 26132 20056 26141 20096
rect 26083 20055 26141 20056
rect 26275 20096 26333 20097
rect 26275 20056 26284 20096
rect 26324 20056 26333 20096
rect 26275 20055 26333 20056
rect 26571 20096 26613 20105
rect 26571 20056 26572 20096
rect 26612 20056 26613 20096
rect 26571 20047 26613 20056
rect 26755 20096 26813 20097
rect 26755 20056 26764 20096
rect 26804 20056 26813 20096
rect 26755 20055 26813 20056
rect 26947 20096 27005 20097
rect 26947 20056 26956 20096
rect 26996 20056 27005 20096
rect 26947 20055 27005 20056
rect 27907 20096 27965 20097
rect 27907 20056 27916 20096
rect 27956 20056 27965 20096
rect 27907 20055 27965 20056
rect 28587 20096 28629 20105
rect 28587 20056 28588 20096
rect 28628 20056 28629 20096
rect 28587 20047 28629 20056
rect 28963 20096 29021 20097
rect 28963 20056 28972 20096
rect 29012 20056 29021 20096
rect 28963 20055 29021 20056
rect 29827 20096 29885 20097
rect 29827 20056 29836 20096
rect 29876 20056 29885 20096
rect 29827 20055 29885 20056
rect 31467 20096 31509 20105
rect 31467 20056 31468 20096
rect 31508 20056 31509 20096
rect 31467 20047 31509 20056
rect 31843 20096 31901 20097
rect 31843 20056 31852 20096
rect 31892 20056 31901 20096
rect 31843 20055 31901 20056
rect 32323 20096 32381 20097
rect 32323 20056 32332 20096
rect 32372 20056 32381 20096
rect 32323 20055 32381 20056
rect 33283 20096 33341 20097
rect 33283 20056 33292 20096
rect 33332 20056 33341 20096
rect 33283 20055 33341 20056
rect 34347 20096 34389 20105
rect 34347 20056 34348 20096
rect 34388 20056 34389 20096
rect 34347 20047 34389 20056
rect 34723 20096 34781 20097
rect 34723 20056 34732 20096
rect 34772 20056 34781 20096
rect 34723 20055 34781 20056
rect 35587 20096 35645 20097
rect 35587 20056 35596 20096
rect 35636 20056 35645 20096
rect 35587 20055 35645 20056
rect 36835 20096 36893 20097
rect 36835 20056 36844 20096
rect 36884 20056 36893 20096
rect 36835 20055 36893 20056
rect 39819 20096 39861 20105
rect 39819 20056 39820 20096
rect 39860 20056 39861 20096
rect 39819 20047 39861 20056
rect 39915 20096 39957 20105
rect 39915 20056 39916 20096
rect 39956 20056 39957 20096
rect 39915 20047 39957 20056
rect 40011 20096 40053 20105
rect 40011 20056 40012 20096
rect 40052 20056 40053 20096
rect 40011 20047 40053 20056
rect 40203 20096 40245 20105
rect 40203 20056 40204 20096
rect 40244 20056 40245 20096
rect 40203 20047 40245 20056
rect 40395 20096 40437 20105
rect 40395 20056 40396 20096
rect 40436 20056 40437 20096
rect 40395 20047 40437 20056
rect 40483 20096 40541 20097
rect 40483 20056 40492 20096
rect 40532 20056 40541 20096
rect 40483 20055 40541 20056
rect 33571 20012 33629 20013
rect 33571 19972 33580 20012
rect 33620 19972 33629 20012
rect 33571 19971 33629 19972
rect 6795 19928 6837 19937
rect 6795 19888 6796 19928
rect 6836 19888 6837 19928
rect 6795 19879 6837 19888
rect 13227 19928 13269 19937
rect 13227 19888 13228 19928
rect 13268 19888 13269 19928
rect 13227 19879 13269 19888
rect 16875 19928 16917 19937
rect 16875 19888 16876 19928
rect 16916 19888 16917 19928
rect 16875 19879 16917 19888
rect 18507 19928 18549 19937
rect 18507 19888 18508 19928
rect 18548 19888 18549 19928
rect 18507 19879 18549 19888
rect 19083 19928 19125 19937
rect 19083 19888 19084 19928
rect 19124 19888 19125 19928
rect 19083 19879 19125 19888
rect 20619 19928 20661 19937
rect 20619 19888 20620 19928
rect 20660 19888 20661 19928
rect 20619 19879 20661 19888
rect 23499 19928 23541 19937
rect 23499 19888 23500 19928
rect 23540 19888 23541 19928
rect 23499 19879 23541 19888
rect 24843 19928 24885 19937
rect 24843 19888 24844 19928
rect 24884 19888 24885 19928
rect 24843 19879 24885 19888
rect 26283 19928 26325 19937
rect 26283 19888 26284 19928
rect 26324 19888 26325 19928
rect 26283 19879 26325 19888
rect 28395 19928 28437 19937
rect 28395 19888 28396 19928
rect 28436 19888 28437 19928
rect 28395 19879 28437 19888
rect 37899 19928 37941 19937
rect 37899 19888 37900 19928
rect 37940 19888 37941 19928
rect 37899 19879 37941 19888
rect 39531 19928 39573 19937
rect 39531 19888 39532 19928
rect 39572 19888 39573 19928
rect 39531 19879 39573 19888
rect 40203 19928 40245 19937
rect 40203 19888 40204 19928
rect 40244 19888 40245 19928
rect 40203 19879 40245 19888
rect 42795 19928 42837 19937
rect 42795 19888 42796 19928
rect 42836 19888 42837 19928
rect 42795 19879 42837 19888
rect 7947 19844 7989 19853
rect 7947 19804 7948 19844
rect 7988 19804 7989 19844
rect 7947 19795 7989 19804
rect 14755 19844 14813 19845
rect 14755 19804 14764 19844
rect 14804 19804 14813 19844
rect 14755 19803 14813 19804
rect 22627 19844 22685 19845
rect 22627 19804 22636 19844
rect 22676 19804 22685 19844
rect 22627 19803 22685 19804
rect 24171 19844 24213 19853
rect 24171 19804 24172 19844
rect 24212 19804 24213 19844
rect 24171 19795 24213 19804
rect 25035 19844 25077 19853
rect 25035 19804 25036 19844
rect 25076 19804 25077 19844
rect 25035 19795 25077 19804
rect 25323 19844 25365 19853
rect 25323 19804 25324 19844
rect 25364 19804 25365 19844
rect 25323 19795 25365 19804
rect 30979 19844 31037 19845
rect 30979 19804 30988 19844
rect 31028 19804 31037 19844
rect 30979 19803 31037 19804
rect 31947 19844 31989 19853
rect 31947 19804 31948 19844
rect 31988 19804 31989 19844
rect 31947 19795 31989 19804
rect 33771 19844 33813 19853
rect 33771 19804 33772 19844
rect 33812 19804 33813 19844
rect 33771 19795 33813 19804
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 5355 19508 5397 19517
rect 5355 19468 5356 19508
rect 5396 19468 5397 19508
rect 5355 19459 5397 19468
rect 10347 19508 10389 19517
rect 10347 19468 10348 19508
rect 10388 19468 10389 19508
rect 10347 19459 10389 19468
rect 14851 19508 14909 19509
rect 14851 19468 14860 19508
rect 14900 19468 14909 19508
rect 14851 19467 14909 19468
rect 17443 19508 17501 19509
rect 17443 19468 17452 19508
rect 17492 19468 17501 19508
rect 17443 19467 17501 19468
rect 20811 19508 20853 19517
rect 20811 19468 20812 19508
rect 20852 19468 20853 19508
rect 20811 19459 20853 19468
rect 34915 19508 34973 19509
rect 34915 19468 34924 19508
rect 34964 19468 34973 19508
rect 34915 19467 34973 19468
rect 1995 19424 2037 19433
rect 1995 19384 1996 19424
rect 2036 19384 2037 19424
rect 1995 19375 2037 19384
rect 3723 19424 3765 19433
rect 3723 19384 3724 19424
rect 3764 19384 3765 19424
rect 3723 19375 3765 19384
rect 5835 19424 5877 19433
rect 5835 19384 5836 19424
rect 5876 19384 5877 19424
rect 5835 19375 5877 19384
rect 36363 19424 36405 19433
rect 36363 19384 36364 19424
rect 36404 19384 36405 19424
rect 36363 19375 36405 19384
rect 8907 19340 8949 19349
rect 8907 19300 8908 19340
rect 8948 19300 8949 19340
rect 8907 19291 8949 19300
rect 35107 19340 35165 19341
rect 35107 19300 35116 19340
rect 35156 19300 35165 19340
rect 35107 19299 35165 19300
rect 3915 19256 3957 19265
rect 3915 19216 3916 19256
rect 3956 19216 3957 19256
rect 3915 19207 3957 19216
rect 4011 19256 4053 19265
rect 4011 19216 4012 19256
rect 4052 19216 4053 19256
rect 4011 19207 4053 19216
rect 4203 19256 4245 19265
rect 4203 19216 4204 19256
rect 4244 19216 4245 19256
rect 4203 19207 4245 19216
rect 4483 19256 4541 19257
rect 4483 19216 4492 19256
rect 4532 19216 4541 19256
rect 4483 19215 4541 19216
rect 5443 19256 5501 19257
rect 5443 19216 5452 19256
rect 5492 19216 5501 19256
rect 5443 19215 5501 19216
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6219 19256 6261 19265
rect 6219 19216 6220 19256
rect 6260 19216 6261 19256
rect 6219 19207 6261 19216
rect 6883 19256 6941 19257
rect 6883 19216 6892 19256
rect 6932 19216 6941 19256
rect 6883 19215 6941 19216
rect 7747 19256 7805 19257
rect 7747 19216 7756 19256
rect 7796 19216 7805 19256
rect 7747 19215 7805 19216
rect 10435 19256 10493 19257
rect 10435 19216 10444 19256
rect 10484 19216 10493 19256
rect 10435 19215 10493 19216
rect 10635 19256 10677 19265
rect 10635 19216 10636 19256
rect 10676 19216 10677 19256
rect 10635 19207 10677 19216
rect 11299 19256 11357 19257
rect 11299 19216 11308 19256
rect 11348 19216 11357 19256
rect 11299 19215 11357 19216
rect 11683 19256 11741 19257
rect 11683 19216 11692 19256
rect 11732 19216 11741 19256
rect 11683 19215 11741 19216
rect 11787 19256 11829 19265
rect 11787 19216 11788 19256
rect 11828 19216 11829 19256
rect 11787 19207 11829 19216
rect 11971 19256 12029 19257
rect 11971 19216 11980 19256
rect 12020 19216 12029 19256
rect 11971 19215 12029 19216
rect 12075 19256 12117 19265
rect 12075 19216 12076 19256
rect 12116 19216 12117 19256
rect 12075 19207 12117 19216
rect 12267 19256 12309 19265
rect 12267 19216 12268 19256
rect 12308 19216 12309 19256
rect 12267 19207 12309 19216
rect 12835 19256 12893 19257
rect 12835 19216 12844 19256
rect 12884 19216 12893 19256
rect 12835 19215 12893 19216
rect 13699 19256 13757 19257
rect 13699 19216 13708 19256
rect 13748 19216 13757 19256
rect 13699 19215 13757 19216
rect 15051 19256 15093 19265
rect 15051 19216 15052 19256
rect 15092 19216 15093 19256
rect 15051 19207 15093 19216
rect 15427 19256 15485 19257
rect 15427 19216 15436 19256
rect 15476 19216 15485 19256
rect 15427 19215 15485 19216
rect 16291 19256 16349 19257
rect 16291 19216 16300 19256
rect 16340 19216 16349 19256
rect 16291 19215 16349 19216
rect 17643 19256 17685 19265
rect 17643 19216 17644 19256
rect 17684 19216 17685 19256
rect 17643 19207 17685 19216
rect 17931 19256 17973 19265
rect 17931 19216 17932 19256
rect 17972 19216 17973 19256
rect 17931 19207 17973 19216
rect 18499 19256 18557 19257
rect 18499 19216 18508 19256
rect 18548 19216 18557 19256
rect 18499 19215 18557 19216
rect 19363 19256 19421 19257
rect 19363 19216 19372 19256
rect 19412 19216 19421 19256
rect 19363 19215 19421 19216
rect 20707 19256 20765 19257
rect 20707 19216 20716 19256
rect 20756 19216 20765 19256
rect 20707 19215 20765 19216
rect 20995 19256 21053 19257
rect 20995 19216 21004 19256
rect 21044 19216 21053 19256
rect 20995 19215 21053 19216
rect 22155 19256 22197 19265
rect 22155 19216 22156 19256
rect 22196 19216 22197 19256
rect 22155 19207 22197 19216
rect 22531 19256 22589 19257
rect 22531 19216 22540 19256
rect 22580 19216 22589 19256
rect 22531 19215 22589 19216
rect 23395 19256 23453 19257
rect 23395 19216 23404 19256
rect 23444 19216 23453 19256
rect 23395 19215 23453 19216
rect 24555 19256 24597 19265
rect 24555 19216 24556 19256
rect 24596 19216 24597 19256
rect 24555 19207 24597 19216
rect 25603 19256 25661 19257
rect 25603 19216 25612 19256
rect 25652 19216 25661 19256
rect 25603 19215 25661 19216
rect 25795 19256 25853 19257
rect 25795 19216 25804 19256
rect 25844 19216 25853 19256
rect 25795 19215 25853 19216
rect 26083 19256 26141 19257
rect 26083 19216 26092 19256
rect 26132 19216 26141 19256
rect 26083 19215 26141 19216
rect 26659 19256 26717 19257
rect 26659 19216 26668 19256
rect 26708 19216 26717 19256
rect 26659 19215 26717 19216
rect 28011 19256 28053 19265
rect 28011 19216 28012 19256
rect 28052 19216 28053 19256
rect 28011 19207 28053 19216
rect 28107 19256 28149 19265
rect 28107 19216 28108 19256
rect 28148 19216 28149 19256
rect 28107 19207 28149 19216
rect 28203 19256 28245 19265
rect 28203 19216 28204 19256
rect 28244 19216 28245 19256
rect 28203 19207 28245 19216
rect 28299 19256 28341 19265
rect 28299 19216 28300 19256
rect 28340 19216 28341 19256
rect 28299 19207 28341 19216
rect 28675 19256 28733 19257
rect 28675 19216 28684 19256
rect 28724 19216 28733 19256
rect 28675 19215 28733 19216
rect 29163 19256 29205 19265
rect 29163 19216 29164 19256
rect 29204 19216 29205 19256
rect 29163 19207 29205 19216
rect 29259 19256 29301 19265
rect 29259 19216 29260 19256
rect 29300 19216 29301 19256
rect 29259 19207 29301 19216
rect 29355 19256 29397 19265
rect 29355 19216 29356 19256
rect 29396 19216 29397 19256
rect 29355 19207 29397 19216
rect 29547 19256 29589 19265
rect 29547 19216 29548 19256
rect 29588 19216 29589 19256
rect 29547 19207 29589 19216
rect 29923 19256 29981 19257
rect 29923 19216 29932 19256
rect 29972 19216 29981 19256
rect 29923 19215 29981 19216
rect 30787 19256 30845 19257
rect 30787 19216 30796 19256
rect 30836 19216 30845 19256
rect 30787 19215 30845 19216
rect 31947 19256 31989 19265
rect 31947 19216 31948 19256
rect 31988 19216 31989 19256
rect 31947 19207 31989 19216
rect 33195 19256 33237 19265
rect 33195 19216 33196 19256
rect 33236 19216 33237 19256
rect 33195 19207 33237 19216
rect 33867 19256 33909 19265
rect 33867 19216 33868 19256
rect 33908 19216 33909 19256
rect 33867 19207 33909 19216
rect 33963 19256 34005 19265
rect 33963 19216 33964 19256
rect 34004 19216 34005 19256
rect 33963 19207 34005 19216
rect 34059 19256 34101 19265
rect 34059 19216 34060 19256
rect 34100 19216 34101 19256
rect 34059 19207 34101 19216
rect 34243 19256 34301 19257
rect 34243 19216 34252 19256
rect 34292 19216 34301 19256
rect 34243 19215 34301 19216
rect 35299 19256 35357 19257
rect 35299 19216 35308 19256
rect 35348 19216 35357 19256
rect 35299 19215 35357 19216
rect 35395 19256 35453 19257
rect 35395 19216 35404 19256
rect 35444 19216 35453 19256
rect 35395 19215 35453 19216
rect 36939 19256 36981 19265
rect 36939 19216 36940 19256
rect 36980 19216 36981 19256
rect 36939 19207 36981 19216
rect 37323 19256 37365 19265
rect 37323 19216 37324 19256
rect 37364 19216 37365 19256
rect 37323 19207 37365 19216
rect 37699 19256 37757 19257
rect 37699 19216 37708 19256
rect 37748 19216 37757 19256
rect 37699 19215 37757 19216
rect 38563 19256 38621 19257
rect 38563 19216 38572 19256
rect 38612 19216 38621 19256
rect 38563 19215 38621 19216
rect 39723 19256 39765 19265
rect 39723 19216 39724 19256
rect 39764 19216 39765 19256
rect 39723 19207 39765 19216
rect 40675 19256 40733 19257
rect 40675 19216 40684 19256
rect 40724 19216 40733 19256
rect 40675 19215 40733 19216
rect 6507 19172 6549 19181
rect 6507 19132 6508 19172
rect 6548 19132 6549 19172
rect 6507 19123 6549 19132
rect 12459 19172 12501 19181
rect 12459 19132 12460 19172
rect 12500 19132 12501 19172
rect 12459 19123 12501 19132
rect 18123 19172 18165 19181
rect 18123 19132 18124 19172
rect 18164 19132 18165 19172
rect 18123 19123 18165 19132
rect 32419 19172 32477 19173
rect 32419 19132 32428 19172
rect 32468 19132 32477 19172
rect 32419 19131 32477 19132
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 4107 19088 4149 19097
rect 4107 19048 4108 19088
rect 4148 19048 4149 19088
rect 4107 19039 4149 19048
rect 5155 19088 5213 19089
rect 5155 19048 5164 19088
rect 5204 19048 5213 19088
rect 5155 19047 5213 19048
rect 6307 19088 6365 19089
rect 6307 19048 6316 19088
rect 6356 19048 6365 19088
rect 6307 19047 6365 19048
rect 12163 19088 12221 19089
rect 12163 19048 12172 19088
rect 12212 19048 12221 19088
rect 12163 19047 12221 19048
rect 17835 19088 17877 19097
rect 17835 19048 17836 19088
rect 17876 19048 17877 19088
rect 17835 19039 17877 19048
rect 20515 19088 20573 19089
rect 20515 19048 20524 19088
rect 20564 19048 20573 19088
rect 20515 19047 20573 19048
rect 21667 19088 21725 19089
rect 21667 19048 21676 19088
rect 21716 19048 21725 19088
rect 21667 19047 21725 19048
rect 25899 19088 25941 19097
rect 25899 19048 25900 19088
rect 25940 19048 25941 19088
rect 25899 19039 25941 19048
rect 27147 19088 27189 19097
rect 27147 19048 27148 19088
rect 27188 19048 27189 19088
rect 27147 19039 27189 19048
rect 27811 19088 27869 19089
rect 27811 19048 27820 19088
rect 27860 19048 27869 19088
rect 27811 19047 27869 19048
rect 28779 19088 28821 19097
rect 28779 19048 28780 19088
rect 28820 19048 28821 19088
rect 28779 19039 28821 19048
rect 29059 19088 29117 19089
rect 29059 19048 29068 19088
rect 29108 19048 29117 19088
rect 29059 19047 29117 19048
rect 33763 19088 33821 19089
rect 33763 19048 33772 19088
rect 33812 19048 33821 19088
rect 33763 19047 33821 19048
rect 40003 19088 40061 19089
rect 40003 19048 40012 19088
rect 40052 19048 40061 19088
rect 40003 19047 40061 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 31843 18794 31901 18795
rect 643 18752 701 18753
rect 643 18712 652 18752
rect 692 18712 701 18752
rect 643 18711 701 18712
rect 3715 18752 3773 18753
rect 3715 18712 3724 18752
rect 3764 18712 3773 18752
rect 3715 18711 3773 18712
rect 4579 18752 4637 18753
rect 4579 18712 4588 18752
rect 4628 18712 4637 18752
rect 4579 18711 4637 18712
rect 4771 18752 4829 18753
rect 4771 18712 4780 18752
rect 4820 18712 4829 18752
rect 4771 18711 4829 18712
rect 6787 18752 6845 18753
rect 6787 18712 6796 18752
rect 6836 18712 6845 18752
rect 6787 18711 6845 18712
rect 11587 18752 11645 18753
rect 11587 18712 11596 18752
rect 11636 18712 11645 18752
rect 11587 18711 11645 18712
rect 12451 18752 12509 18753
rect 12451 18712 12460 18752
rect 12500 18712 12509 18752
rect 12451 18711 12509 18712
rect 13315 18752 13373 18753
rect 13315 18712 13324 18752
rect 13364 18712 13373 18752
rect 13315 18711 13373 18712
rect 14947 18752 15005 18753
rect 14947 18712 14956 18752
rect 14996 18712 15005 18752
rect 14947 18711 15005 18712
rect 16395 18752 16437 18761
rect 16395 18712 16396 18752
rect 16436 18712 16437 18752
rect 16395 18703 16437 18712
rect 19555 18752 19613 18753
rect 19555 18712 19564 18752
rect 19604 18712 19613 18752
rect 19555 18711 19613 18712
rect 20523 18752 20565 18761
rect 20523 18712 20524 18752
rect 20564 18712 20565 18752
rect 20523 18703 20565 18712
rect 22051 18752 22109 18753
rect 22051 18712 22060 18752
rect 22100 18712 22109 18752
rect 22051 18711 22109 18712
rect 24739 18752 24797 18753
rect 24739 18712 24748 18752
rect 24788 18712 24797 18752
rect 24739 18711 24797 18712
rect 26667 18752 26709 18761
rect 31843 18754 31852 18794
rect 31892 18754 31901 18794
rect 31843 18753 31901 18754
rect 26667 18712 26668 18752
rect 26708 18712 26709 18752
rect 26667 18703 26709 18712
rect 35403 18752 35445 18761
rect 35403 18712 35404 18752
rect 35444 18712 35445 18752
rect 35403 18703 35445 18712
rect 36355 18752 36413 18753
rect 36355 18712 36364 18752
rect 36404 18712 36413 18752
rect 36355 18711 36413 18712
rect 1323 18668 1365 18677
rect 1323 18628 1324 18668
rect 1364 18628 1365 18668
rect 1323 18619 1365 18628
rect 23115 18668 23157 18677
rect 23115 18628 23116 18668
rect 23156 18628 23157 18668
rect 23115 18619 23157 18628
rect 1699 18584 1757 18585
rect 1699 18544 1708 18584
rect 1748 18544 1757 18584
rect 1699 18543 1757 18544
rect 2563 18584 2621 18585
rect 2563 18544 2572 18584
rect 2612 18544 2621 18584
rect 2563 18543 2621 18544
rect 3907 18584 3965 18585
rect 3907 18544 3916 18584
rect 3956 18544 3965 18584
rect 3907 18543 3965 18544
rect 4867 18584 4925 18585
rect 4867 18544 4876 18584
rect 4916 18544 4925 18584
rect 4867 18543 4925 18544
rect 6595 18584 6653 18585
rect 6595 18544 6604 18584
rect 6644 18544 6653 18584
rect 6595 18543 6653 18544
rect 7459 18584 7517 18585
rect 7459 18544 7468 18584
rect 7508 18544 7517 18584
rect 7459 18543 7517 18544
rect 7659 18584 7701 18593
rect 7659 18544 7660 18584
rect 7700 18544 7701 18584
rect 7659 18535 7701 18544
rect 7851 18584 7893 18593
rect 7851 18544 7852 18584
rect 7892 18544 7893 18584
rect 7851 18535 7893 18544
rect 7939 18584 7997 18585
rect 7939 18544 7948 18584
rect 7988 18544 7997 18584
rect 7939 18543 7997 18544
rect 10251 18584 10293 18593
rect 10251 18544 10252 18584
rect 10292 18544 10293 18584
rect 10251 18535 10293 18544
rect 10347 18584 10389 18593
rect 10347 18544 10348 18584
rect 10388 18544 10389 18584
rect 10347 18535 10389 18544
rect 10443 18584 10485 18593
rect 10443 18544 10444 18584
rect 10484 18544 10485 18584
rect 10443 18535 10485 18544
rect 10539 18584 10581 18593
rect 10539 18544 10540 18584
rect 10580 18544 10581 18584
rect 10539 18535 10581 18544
rect 10819 18584 10877 18585
rect 10819 18544 10828 18584
rect 10868 18544 10877 18584
rect 10819 18543 10877 18544
rect 11115 18584 11157 18593
rect 11115 18544 11116 18584
rect 11156 18544 11157 18584
rect 11115 18535 11157 18544
rect 11211 18584 11253 18593
rect 11211 18544 11212 18584
rect 11252 18544 11253 18584
rect 11211 18535 11253 18544
rect 11307 18584 11349 18593
rect 11307 18544 11308 18584
rect 11348 18544 11349 18584
rect 11307 18535 11349 18544
rect 11403 18584 11445 18593
rect 11403 18544 11404 18584
rect 11444 18544 11445 18584
rect 11403 18535 11445 18544
rect 12259 18584 12317 18585
rect 12259 18544 12268 18584
rect 12308 18544 12317 18584
rect 12259 18543 12317 18544
rect 13123 18584 13181 18585
rect 13123 18544 13132 18584
rect 13172 18544 13181 18584
rect 13123 18543 13181 18544
rect 13987 18584 14045 18585
rect 13987 18544 13996 18584
rect 14036 18544 14045 18584
rect 13987 18543 14045 18544
rect 15051 18584 15093 18593
rect 15051 18544 15052 18584
rect 15092 18544 15093 18584
rect 15051 18535 15093 18544
rect 15147 18584 15189 18593
rect 15147 18544 15148 18584
rect 15188 18544 15189 18584
rect 15147 18535 15189 18544
rect 15243 18584 15285 18593
rect 15243 18544 15244 18584
rect 15284 18544 15285 18584
rect 15243 18535 15285 18544
rect 15427 18584 15485 18585
rect 15427 18544 15436 18584
rect 15476 18544 15485 18584
rect 15427 18543 15485 18544
rect 16107 18584 16149 18593
rect 16107 18544 16108 18584
rect 16148 18544 16149 18584
rect 16107 18535 16149 18544
rect 16291 18584 16349 18585
rect 16291 18544 16300 18584
rect 16340 18544 16349 18584
rect 16291 18543 16349 18544
rect 20227 18584 20285 18585
rect 20227 18544 20236 18584
rect 20276 18544 20285 18584
rect 20227 18543 20285 18544
rect 20611 18584 20669 18585
rect 20611 18544 20620 18584
rect 20660 18544 20669 18584
rect 20611 18543 20669 18544
rect 20803 18584 20861 18585
rect 20803 18544 20812 18584
rect 20852 18544 20861 18584
rect 20803 18543 20861 18544
rect 21195 18584 21237 18593
rect 21195 18544 21196 18584
rect 21236 18544 21237 18584
rect 21195 18535 21237 18544
rect 21379 18584 21437 18585
rect 21379 18544 21388 18584
rect 21428 18544 21437 18584
rect 21379 18543 21437 18544
rect 22243 18584 22301 18585
rect 22243 18544 22252 18584
rect 22292 18544 22301 18584
rect 22243 18543 22301 18544
rect 22635 18584 22677 18593
rect 22635 18544 22636 18584
rect 22676 18544 22677 18584
rect 22635 18535 22677 18544
rect 23211 18584 23253 18593
rect 23211 18544 23212 18584
rect 23252 18544 23253 18584
rect 23211 18535 23253 18544
rect 23307 18584 23349 18593
rect 23307 18544 23308 18584
rect 23348 18544 23349 18584
rect 23307 18535 23349 18544
rect 23403 18584 23445 18593
rect 23403 18544 23404 18584
rect 23444 18544 23445 18584
rect 23403 18535 23445 18544
rect 23595 18584 23637 18593
rect 23595 18544 23596 18584
rect 23636 18544 23637 18584
rect 23595 18535 23637 18544
rect 23691 18584 23733 18593
rect 23691 18544 23692 18584
rect 23732 18544 23733 18584
rect 23691 18535 23733 18544
rect 23787 18584 23829 18593
rect 23787 18544 23788 18584
rect 23828 18544 23829 18584
rect 23787 18535 23829 18544
rect 23883 18584 23925 18593
rect 23883 18544 23884 18584
rect 23924 18544 23925 18584
rect 23883 18535 23925 18544
rect 24067 18584 24125 18585
rect 24067 18544 24076 18584
rect 24116 18544 24125 18584
rect 24067 18543 24125 18544
rect 25131 18584 25173 18593
rect 25131 18544 25132 18584
rect 25172 18544 25173 18584
rect 25131 18535 25173 18544
rect 26667 18584 26709 18593
rect 26667 18544 26668 18584
rect 26708 18544 26709 18584
rect 26667 18535 26709 18544
rect 26755 18584 26813 18585
rect 26755 18544 26764 18584
rect 26804 18544 26813 18584
rect 26755 18543 26813 18544
rect 27147 18584 27189 18593
rect 27147 18544 27148 18584
rect 27188 18544 27189 18584
rect 27147 18535 27189 18544
rect 27523 18584 27581 18585
rect 27523 18544 27532 18584
rect 27572 18544 27581 18584
rect 27523 18543 27581 18544
rect 28387 18584 28445 18585
rect 28387 18544 28396 18584
rect 28436 18544 28445 18584
rect 28387 18543 28445 18544
rect 29547 18584 29589 18593
rect 29547 18544 29548 18584
rect 29588 18544 29589 18584
rect 29547 18535 29589 18544
rect 29827 18584 29885 18585
rect 29827 18544 29836 18584
rect 29876 18544 29885 18584
rect 29827 18543 29885 18544
rect 31363 18584 31421 18585
rect 31363 18544 31372 18584
rect 31412 18544 31421 18584
rect 31363 18543 31421 18544
rect 31651 18584 31709 18585
rect 31651 18544 31660 18584
rect 31700 18544 31709 18584
rect 31651 18543 31709 18544
rect 31843 18584 31901 18585
rect 31843 18544 31852 18584
rect 31892 18544 31901 18584
rect 31843 18543 31901 18544
rect 32227 18584 32285 18585
rect 32227 18544 32236 18584
rect 32276 18544 32285 18584
rect 32227 18543 32285 18544
rect 33099 18584 33141 18593
rect 33099 18544 33100 18584
rect 33140 18544 33141 18584
rect 33099 18535 33141 18544
rect 33571 18584 33629 18585
rect 33571 18544 33580 18584
rect 33620 18544 33629 18584
rect 33571 18543 33629 18544
rect 33675 18584 33717 18593
rect 33675 18544 33676 18584
rect 33716 18544 33717 18584
rect 33675 18535 33717 18544
rect 33867 18584 33909 18593
rect 33867 18544 33868 18584
rect 33908 18544 33909 18584
rect 33867 18535 33909 18544
rect 34251 18584 34293 18593
rect 34251 18544 34252 18584
rect 34292 18544 34293 18584
rect 34251 18535 34293 18544
rect 34339 18584 34397 18585
rect 34339 18544 34348 18584
rect 34388 18544 34397 18584
rect 34339 18543 34397 18544
rect 35019 18584 35061 18593
rect 35019 18544 35020 18584
rect 35060 18544 35061 18584
rect 35019 18535 35061 18544
rect 35107 18584 35165 18585
rect 35107 18544 35116 18584
rect 35156 18544 35165 18584
rect 35107 18543 35165 18544
rect 35678 18584 35736 18585
rect 35678 18544 35687 18584
rect 35727 18544 35736 18584
rect 35678 18543 35736 18544
rect 35787 18584 35829 18593
rect 35787 18544 35788 18584
rect 35828 18544 35829 18584
rect 35787 18535 35829 18544
rect 35883 18584 35925 18593
rect 35883 18544 35884 18584
rect 35924 18544 35925 18584
rect 35883 18535 35925 18544
rect 36067 18584 36125 18585
rect 36067 18544 36076 18584
rect 36116 18544 36125 18584
rect 36067 18543 36125 18544
rect 36163 18584 36221 18585
rect 36163 18544 36172 18584
rect 36212 18544 36221 18584
rect 36163 18543 36221 18544
rect 37027 18584 37085 18585
rect 37027 18544 37036 18584
rect 37076 18544 37085 18584
rect 37027 18543 37085 18544
rect 37227 18584 37269 18593
rect 37227 18544 37228 18584
rect 37268 18544 37269 18584
rect 37227 18535 37269 18544
rect 37323 18584 37365 18593
rect 37323 18544 37324 18584
rect 37364 18544 37365 18584
rect 37323 18535 37365 18544
rect 37419 18584 37461 18593
rect 37419 18544 37420 18584
rect 37460 18544 37461 18584
rect 37419 18535 37461 18544
rect 37515 18584 37557 18593
rect 37515 18544 37516 18584
rect 37556 18544 37557 18584
rect 37515 18535 37557 18544
rect 37891 18584 37949 18585
rect 37891 18544 37900 18584
rect 37940 18544 37949 18584
rect 37891 18543 37949 18544
rect 38851 18584 38909 18585
rect 38851 18544 38860 18584
rect 38900 18544 38909 18584
rect 38851 18543 38909 18544
rect 39235 18584 39293 18585
rect 39235 18544 39244 18584
rect 39284 18544 39293 18584
rect 39235 18543 39293 18544
rect 40483 18584 40541 18585
rect 40483 18544 40492 18584
rect 40532 18544 40541 18584
rect 40483 18543 40541 18544
rect 41443 18584 41501 18585
rect 41443 18544 41452 18584
rect 41492 18544 41501 18584
rect 41443 18543 41501 18544
rect 20907 18500 20949 18509
rect 20907 18460 20908 18500
rect 20948 18460 20949 18500
rect 20907 18451 20949 18460
rect 21099 18500 21141 18509
rect 21099 18460 21100 18500
rect 21140 18460 21141 18500
rect 21099 18451 21141 18460
rect 22347 18500 22389 18509
rect 22347 18460 22348 18500
rect 22388 18460 22389 18500
rect 22347 18451 22389 18460
rect 22539 18500 22581 18509
rect 22539 18460 22540 18500
rect 22580 18460 22581 18500
rect 22539 18451 22581 18460
rect 26571 18500 26613 18509
rect 26571 18460 26572 18500
rect 26612 18460 26613 18500
rect 26571 18451 26613 18460
rect 34627 18500 34685 18501
rect 34627 18460 34636 18500
rect 34676 18460 34685 18500
rect 34627 18459 34685 18460
rect 5739 18416 5781 18425
rect 5739 18376 5740 18416
rect 5780 18376 5781 18416
rect 5739 18367 5781 18376
rect 7659 18416 7701 18425
rect 7659 18376 7660 18416
rect 7700 18376 7701 18416
rect 7659 18367 7701 18376
rect 9387 18416 9429 18425
rect 9387 18376 9388 18416
rect 9428 18376 9429 18416
rect 9387 18367 9429 18376
rect 14187 18416 14229 18425
rect 14187 18376 14188 18416
rect 14228 18376 14229 18416
rect 14187 18367 14229 18376
rect 18219 18416 18261 18425
rect 18219 18376 18220 18416
rect 18260 18376 18261 18416
rect 18219 18367 18261 18376
rect 21003 18416 21045 18425
rect 21003 18376 21004 18416
rect 21044 18376 21045 18416
rect 21003 18367 21045 18376
rect 22443 18416 22485 18425
rect 22443 18376 22444 18416
rect 22484 18376 22485 18416
rect 22443 18367 22485 18376
rect 25707 18416 25749 18425
rect 25707 18376 25708 18416
rect 25748 18376 25749 18416
rect 25707 18367 25749 18376
rect 26475 18416 26517 18425
rect 26475 18376 26476 18416
rect 26516 18376 26517 18416
rect 26475 18367 26517 18376
rect 33867 18416 33909 18425
rect 33867 18376 33868 18416
rect 33908 18376 33909 18416
rect 33867 18367 33909 18376
rect 4579 18332 4637 18333
rect 4579 18292 4588 18332
rect 4628 18292 4637 18332
rect 4579 18291 4637 18292
rect 5059 18332 5117 18333
rect 5059 18292 5068 18332
rect 5108 18292 5117 18332
rect 5059 18291 5117 18292
rect 5923 18332 5981 18333
rect 5923 18292 5932 18332
rect 5972 18292 5981 18332
rect 5923 18291 5981 18292
rect 10923 18332 10965 18341
rect 10923 18292 10924 18332
rect 10964 18292 10965 18332
rect 10923 18283 10965 18292
rect 24739 18332 24797 18333
rect 24739 18292 24748 18332
rect 24788 18292 24797 18332
rect 24739 18291 24797 18292
rect 30499 18332 30557 18333
rect 30499 18292 30508 18332
rect 30548 18292 30557 18332
rect 30499 18291 30557 18292
rect 30691 18332 30749 18333
rect 30691 18292 30700 18332
rect 30740 18292 30749 18332
rect 30691 18291 30749 18292
rect 36171 18332 36213 18341
rect 36171 18292 36172 18332
rect 36212 18292 36213 18332
rect 36171 18283 36213 18292
rect 39915 18332 39957 18341
rect 39915 18292 39916 18332
rect 39956 18292 39957 18332
rect 39915 18283 39957 18292
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 3907 17996 3965 17997
rect 3907 17956 3916 17996
rect 3956 17956 3965 17996
rect 3907 17955 3965 17956
rect 11299 17996 11357 17997
rect 11299 17956 11308 17996
rect 11348 17956 11357 17996
rect 11299 17955 11357 17956
rect 14955 17996 14997 18005
rect 14955 17956 14956 17996
rect 14996 17956 14997 17996
rect 14955 17947 14997 17956
rect 20139 17996 20181 18005
rect 20139 17956 20140 17996
rect 20180 17956 20181 17996
rect 20139 17947 20181 17956
rect 24363 17996 24405 18005
rect 24363 17956 24364 17996
rect 24404 17956 24405 17996
rect 24363 17947 24405 17956
rect 26091 17996 26133 18005
rect 26091 17956 26092 17996
rect 26132 17956 26133 17996
rect 26091 17947 26133 17956
rect 28963 17996 29021 17997
rect 28963 17956 28972 17996
rect 29012 17956 29021 17996
rect 28963 17955 29021 17956
rect 29827 17996 29885 17997
rect 29827 17956 29836 17996
rect 29876 17956 29885 17996
rect 29827 17955 29885 17956
rect 30315 17996 30357 18005
rect 30315 17956 30316 17996
rect 30356 17956 30357 17996
rect 30315 17947 30357 17956
rect 34155 17996 34197 18005
rect 34155 17956 34156 17996
rect 34196 17956 34197 17996
rect 34155 17947 34197 17956
rect 34635 17996 34677 18005
rect 34635 17956 34636 17996
rect 34676 17956 34677 17996
rect 34635 17947 34677 17956
rect 1323 17912 1365 17921
rect 1323 17872 1324 17912
rect 1364 17872 1365 17912
rect 1323 17863 1365 17872
rect 4683 17912 4725 17921
rect 4683 17872 4684 17912
rect 4724 17872 4725 17912
rect 4683 17863 4725 17872
rect 8715 17912 8757 17921
rect 8715 17872 8716 17912
rect 8756 17872 8757 17912
rect 8715 17863 8757 17872
rect 27243 17912 27285 17921
rect 27243 17872 27244 17912
rect 27284 17872 27285 17912
rect 27243 17863 27285 17872
rect 27915 17912 27957 17921
rect 27915 17872 27916 17912
rect 27956 17872 27957 17912
rect 27915 17863 27957 17872
rect 37707 17912 37749 17921
rect 37707 17872 37708 17912
rect 37748 17872 37749 17912
rect 37707 17863 37749 17872
rect 31747 17828 31805 17829
rect 31747 17788 31756 17828
rect 31796 17788 31805 17828
rect 31747 17787 31805 17788
rect 36651 17828 36693 17837
rect 36651 17788 36652 17828
rect 36692 17788 36693 17828
rect 36651 17779 36693 17788
rect 24904 17759 24946 17768
rect 1891 17744 1949 17745
rect 1891 17704 1900 17744
rect 1940 17704 1949 17744
rect 1891 17703 1949 17704
rect 2755 17744 2813 17745
rect 2755 17704 2764 17744
rect 2804 17704 2813 17744
rect 2755 17703 2813 17704
rect 4387 17744 4445 17745
rect 4387 17704 4396 17744
rect 4436 17704 4445 17744
rect 4387 17703 4445 17704
rect 4491 17744 4533 17753
rect 4491 17704 4492 17744
rect 4532 17704 4533 17744
rect 4491 17695 4533 17704
rect 4675 17744 4733 17745
rect 4675 17704 4684 17744
rect 4724 17704 4733 17744
rect 4675 17703 4733 17704
rect 4867 17744 4925 17745
rect 4867 17704 4876 17744
rect 4916 17704 4925 17744
rect 4867 17703 4925 17704
rect 5739 17744 5781 17753
rect 5739 17704 5740 17744
rect 5780 17704 5781 17744
rect 5739 17695 5781 17704
rect 6115 17744 6173 17745
rect 6115 17704 6124 17744
rect 6164 17704 6173 17744
rect 6115 17703 6173 17704
rect 6979 17744 7037 17745
rect 6979 17704 6988 17744
rect 7028 17704 7037 17744
rect 6979 17703 7037 17704
rect 8419 17744 8477 17745
rect 8419 17704 8428 17744
rect 8468 17704 8477 17744
rect 8419 17703 8477 17704
rect 8523 17744 8565 17753
rect 8523 17704 8524 17744
rect 8564 17704 8565 17744
rect 8523 17695 8565 17704
rect 8715 17744 8757 17753
rect 8715 17704 8716 17744
rect 8756 17704 8757 17744
rect 8715 17695 8757 17704
rect 8907 17744 8949 17753
rect 8907 17704 8908 17744
rect 8948 17704 8949 17744
rect 8907 17695 8949 17704
rect 9283 17744 9341 17745
rect 9283 17704 9292 17744
rect 9332 17704 9341 17744
rect 9283 17703 9341 17704
rect 10147 17744 10205 17745
rect 10147 17704 10156 17744
rect 10196 17704 10205 17744
rect 10147 17703 10205 17704
rect 11683 17744 11741 17745
rect 11683 17704 11692 17744
rect 11732 17704 11741 17744
rect 11683 17703 11741 17704
rect 12363 17744 12405 17753
rect 12363 17704 12364 17744
rect 12404 17704 12405 17744
rect 12363 17695 12405 17704
rect 12555 17744 12597 17753
rect 12555 17704 12556 17744
rect 12596 17704 12597 17744
rect 12555 17695 12597 17704
rect 12931 17744 12989 17745
rect 12931 17704 12940 17744
rect 12980 17704 12989 17744
rect 12931 17703 12989 17704
rect 13795 17744 13853 17745
rect 13795 17704 13804 17744
rect 13844 17704 13853 17744
rect 13795 17703 13853 17704
rect 15907 17744 15965 17745
rect 15907 17704 15916 17744
rect 15956 17704 15965 17744
rect 15907 17703 15965 17704
rect 17739 17744 17781 17753
rect 17739 17704 17740 17744
rect 17780 17704 17781 17744
rect 17739 17695 17781 17704
rect 18115 17744 18173 17745
rect 18115 17704 18124 17744
rect 18164 17704 18173 17744
rect 18115 17703 18173 17704
rect 18979 17744 19037 17745
rect 18979 17704 18988 17744
rect 19028 17704 19037 17744
rect 18979 17703 19037 17704
rect 20811 17744 20853 17753
rect 20811 17704 20812 17744
rect 20852 17704 20853 17744
rect 20811 17695 20853 17704
rect 21475 17744 21533 17745
rect 21475 17704 21484 17744
rect 21524 17704 21533 17744
rect 21475 17703 21533 17704
rect 21667 17744 21725 17745
rect 21667 17704 21676 17744
rect 21716 17704 21725 17744
rect 21667 17703 21725 17704
rect 22539 17744 22581 17753
rect 22539 17704 22540 17744
rect 22580 17704 22581 17744
rect 22539 17695 22581 17704
rect 22915 17744 22973 17745
rect 22915 17704 22924 17744
rect 22964 17704 22973 17744
rect 22915 17703 22973 17704
rect 23019 17744 23061 17753
rect 23019 17704 23020 17744
rect 23060 17704 23061 17744
rect 23019 17695 23061 17704
rect 23211 17744 23253 17753
rect 23211 17704 23212 17744
rect 23252 17704 23253 17744
rect 23211 17695 23253 17704
rect 23395 17744 23453 17745
rect 23395 17704 23404 17744
rect 23444 17704 23453 17744
rect 23395 17703 23453 17704
rect 23499 17744 23541 17753
rect 23499 17704 23500 17744
rect 23540 17704 23541 17744
rect 23499 17695 23541 17704
rect 23691 17744 23733 17753
rect 23691 17704 23692 17744
rect 23732 17704 23733 17744
rect 23691 17695 23733 17704
rect 23883 17744 23925 17753
rect 23883 17704 23884 17744
rect 23924 17704 23925 17744
rect 23883 17695 23925 17704
rect 24075 17744 24117 17753
rect 24075 17704 24076 17744
rect 24116 17704 24117 17744
rect 24075 17695 24117 17704
rect 24163 17744 24221 17745
rect 24163 17704 24172 17744
rect 24212 17704 24221 17744
rect 24163 17703 24221 17704
rect 24355 17744 24413 17745
rect 24355 17704 24364 17744
rect 24404 17704 24413 17744
rect 24355 17703 24413 17704
rect 24451 17744 24509 17745
rect 24451 17704 24460 17744
rect 24500 17704 24509 17744
rect 24451 17703 24509 17704
rect 24651 17744 24693 17753
rect 24651 17704 24652 17744
rect 24692 17704 24693 17744
rect 24651 17695 24693 17704
rect 24747 17744 24789 17753
rect 24747 17704 24748 17744
rect 24788 17704 24789 17744
rect 24904 17719 24905 17759
rect 24945 17719 24946 17759
rect 24904 17710 24946 17719
rect 26091 17744 26133 17753
rect 24747 17695 24789 17704
rect 26091 17704 26092 17744
rect 26132 17704 26133 17744
rect 26091 17695 26133 17704
rect 26283 17744 26325 17753
rect 26283 17704 26284 17744
rect 26324 17704 26325 17744
rect 26283 17695 26325 17704
rect 26563 17744 26621 17745
rect 26563 17704 26572 17744
rect 26612 17704 26621 17744
rect 26563 17703 26621 17704
rect 27435 17744 27477 17753
rect 27435 17704 27436 17744
rect 27476 17704 27477 17744
rect 27435 17695 27477 17704
rect 27619 17744 27677 17745
rect 27619 17704 27628 17744
rect 27668 17704 27677 17744
rect 27619 17703 27677 17704
rect 27915 17744 27957 17753
rect 27915 17704 27916 17744
rect 27956 17704 27957 17744
rect 27915 17695 27957 17704
rect 28291 17744 28349 17745
rect 28291 17704 28300 17744
rect 28340 17704 28349 17744
rect 28291 17703 28349 17704
rect 29155 17744 29213 17745
rect 29155 17704 29164 17744
rect 29204 17704 29213 17744
rect 29155 17703 29213 17704
rect 30979 17744 31037 17745
rect 30979 17704 30988 17744
rect 31028 17704 31037 17744
rect 30979 17703 31037 17704
rect 31363 17744 31421 17745
rect 31363 17704 31372 17744
rect 31412 17704 31421 17744
rect 31363 17703 31421 17704
rect 31555 17744 31613 17745
rect 31555 17704 31564 17744
rect 31604 17704 31613 17744
rect 31555 17703 31613 17704
rect 31843 17744 31901 17745
rect 31843 17704 31852 17744
rect 31892 17704 31901 17744
rect 31843 17703 31901 17704
rect 33195 17744 33237 17753
rect 33195 17704 33196 17744
rect 33236 17704 33237 17744
rect 33195 17695 33237 17704
rect 34155 17744 34197 17753
rect 34155 17704 34156 17744
rect 34196 17704 34197 17744
rect 34155 17695 34197 17704
rect 34347 17744 34389 17753
rect 34347 17704 34348 17744
rect 34388 17704 34389 17744
rect 34347 17695 34389 17704
rect 34435 17744 34493 17745
rect 34435 17704 34444 17744
rect 34484 17704 34493 17744
rect 34435 17703 34493 17704
rect 34627 17744 34685 17745
rect 34627 17704 34636 17744
rect 34676 17704 34685 17744
rect 34627 17703 34685 17704
rect 34723 17744 34781 17745
rect 34723 17704 34732 17744
rect 34772 17704 34781 17744
rect 34723 17703 34781 17704
rect 34923 17744 34965 17753
rect 34923 17704 34924 17744
rect 34964 17704 34965 17744
rect 34923 17695 34965 17704
rect 35019 17744 35061 17753
rect 35019 17704 35020 17744
rect 35060 17704 35061 17744
rect 35019 17695 35061 17704
rect 35112 17744 35170 17745
rect 35112 17704 35121 17744
rect 35161 17704 35170 17744
rect 35112 17703 35170 17704
rect 35403 17744 35445 17753
rect 35403 17704 35404 17744
rect 35444 17704 35445 17744
rect 35403 17695 35445 17704
rect 35499 17744 35541 17753
rect 35499 17704 35500 17744
rect 35540 17704 35541 17744
rect 35499 17695 35541 17704
rect 35595 17744 35637 17753
rect 35595 17704 35596 17744
rect 35636 17704 35637 17744
rect 35595 17695 35637 17704
rect 35691 17744 35733 17753
rect 35691 17704 35692 17744
rect 35732 17704 35733 17744
rect 35691 17695 35733 17704
rect 36555 17744 36597 17753
rect 36555 17704 36556 17744
rect 36596 17704 36597 17744
rect 36555 17695 36597 17704
rect 36747 17744 36789 17753
rect 36747 17704 36748 17744
rect 36788 17704 36789 17744
rect 36747 17695 36789 17704
rect 37035 17744 37077 17753
rect 37035 17704 37036 17744
rect 37076 17704 37077 17744
rect 37227 17744 37269 17753
rect 37035 17695 37077 17704
rect 37131 17723 37173 17732
rect 37131 17683 37132 17723
rect 37172 17683 37173 17723
rect 37227 17704 37228 17744
rect 37268 17704 37269 17744
rect 37227 17695 37269 17704
rect 37411 17744 37469 17745
rect 37411 17704 37420 17744
rect 37460 17704 37469 17744
rect 37411 17703 37469 17704
rect 37515 17744 37557 17753
rect 37515 17704 37516 17744
rect 37556 17704 37557 17744
rect 37515 17695 37557 17704
rect 37707 17744 37749 17753
rect 37707 17704 37708 17744
rect 37748 17704 37749 17744
rect 37707 17695 37749 17704
rect 37891 17744 37949 17745
rect 37891 17704 37900 17744
rect 37940 17704 37949 17744
rect 37891 17703 37949 17704
rect 38763 17744 38805 17753
rect 38763 17704 38764 17744
rect 38804 17704 38805 17744
rect 38763 17695 38805 17704
rect 39139 17744 39197 17745
rect 39139 17704 39148 17744
rect 39188 17704 39197 17744
rect 39139 17703 39197 17704
rect 40003 17744 40061 17745
rect 40003 17704 40012 17744
rect 40052 17704 40061 17744
rect 40003 17703 40061 17704
rect 41251 17744 41309 17745
rect 41251 17704 41260 17744
rect 41300 17704 41309 17744
rect 41251 17703 41309 17704
rect 37131 17674 37173 17683
rect 1515 17660 1557 17669
rect 1515 17620 1516 17660
rect 1556 17620 1557 17660
rect 1515 17611 1557 17620
rect 16771 17660 16829 17661
rect 16771 17620 16780 17660
rect 16820 17620 16829 17660
rect 16771 17619 16829 17620
rect 23115 17660 23157 17669
rect 23115 17620 23116 17660
rect 23156 17620 23157 17660
rect 23115 17611 23157 17620
rect 23595 17660 23637 17669
rect 23595 17620 23596 17660
rect 23636 17620 23637 17660
rect 23595 17611 23637 17620
rect 23979 17660 24021 17669
rect 23979 17620 23980 17660
rect 24020 17620 24021 17660
rect 23979 17611 24021 17620
rect 26755 17660 26813 17661
rect 26755 17620 26764 17660
rect 26804 17620 26813 17660
rect 26755 17619 26813 17620
rect 27531 17660 27573 17669
rect 27531 17620 27532 17660
rect 27572 17620 27573 17660
rect 27531 17611 27573 17620
rect 32419 17660 32477 17661
rect 32419 17620 32428 17660
rect 32468 17620 32477 17660
rect 32419 17619 32477 17620
rect 36939 17660 36981 17669
rect 36939 17620 36940 17660
rect 36980 17620 36981 17660
rect 36939 17611 36981 17620
rect 643 17576 701 17577
rect 643 17536 652 17576
rect 692 17536 701 17576
rect 643 17535 701 17536
rect 5539 17576 5597 17577
rect 5539 17536 5548 17576
rect 5588 17536 5597 17576
rect 5539 17535 5597 17536
rect 8131 17576 8189 17577
rect 8131 17536 8140 17576
rect 8180 17536 8189 17576
rect 8131 17535 8189 17536
rect 26467 17576 26525 17577
rect 26467 17536 26476 17576
rect 26516 17536 26525 17576
rect 26467 17535 26525 17536
rect 28107 17576 28149 17585
rect 28107 17536 28108 17576
rect 28148 17536 28149 17576
rect 28107 17527 28149 17536
rect 38563 17576 38621 17577
rect 38563 17536 38572 17576
rect 38612 17536 38621 17576
rect 38563 17535 38621 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 27723 17298 27765 17307
rect 27723 17258 27724 17298
rect 27764 17258 27765 17298
rect 27723 17249 27765 17258
rect 643 17240 701 17241
rect 643 17200 652 17240
rect 692 17200 701 17240
rect 643 17199 701 17200
rect 3723 17240 3765 17249
rect 3723 17200 3724 17240
rect 3764 17200 3765 17240
rect 3723 17191 3765 17200
rect 4387 17240 4445 17241
rect 4387 17200 4396 17240
rect 4436 17200 4445 17240
rect 4387 17199 4445 17200
rect 5835 17240 5877 17249
rect 5835 17200 5836 17240
rect 5876 17200 5877 17240
rect 5835 17191 5877 17200
rect 20803 17240 20861 17241
rect 20803 17200 20812 17240
rect 20852 17200 20861 17240
rect 20803 17199 20861 17200
rect 21867 17240 21909 17249
rect 21867 17200 21868 17240
rect 21908 17200 21909 17240
rect 21867 17191 21909 17200
rect 23395 17240 23453 17241
rect 23395 17200 23404 17240
rect 23444 17200 23453 17240
rect 23395 17199 23453 17200
rect 24163 17240 24221 17241
rect 24163 17200 24172 17240
rect 24212 17200 24221 17240
rect 24163 17199 24221 17200
rect 24643 17240 24701 17241
rect 24643 17200 24652 17240
rect 24692 17200 24701 17240
rect 24643 17199 24701 17200
rect 25411 17240 25469 17241
rect 25411 17200 25420 17240
rect 25460 17200 25469 17240
rect 25411 17199 25469 17200
rect 26563 17240 26621 17241
rect 26563 17200 26572 17240
rect 26612 17200 26621 17240
rect 26563 17199 26621 17200
rect 36643 17240 36701 17241
rect 36643 17200 36652 17240
rect 36692 17200 36701 17240
rect 36643 17199 36701 17200
rect 38275 17240 38333 17241
rect 38275 17200 38284 17240
rect 38324 17200 38333 17240
rect 38275 17199 38333 17200
rect 39147 17240 39189 17249
rect 39147 17200 39148 17240
rect 39188 17200 39189 17240
rect 39147 17191 39189 17200
rect 4099 17156 4157 17157
rect 4099 17116 4108 17156
rect 4148 17116 4157 17156
rect 4099 17115 4157 17116
rect 19371 17156 19413 17165
rect 19371 17116 19372 17156
rect 19412 17116 19413 17156
rect 19371 17107 19413 17116
rect 35019 17156 35061 17165
rect 35019 17116 35020 17156
rect 35060 17116 35061 17156
rect 35019 17107 35061 17116
rect 3243 17072 3285 17081
rect 3243 17032 3244 17072
rect 3284 17032 3285 17072
rect 3243 17023 3285 17032
rect 3435 17072 3477 17081
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3627 17072 3669 17081
rect 3627 17032 3628 17072
rect 3668 17032 3669 17072
rect 3627 17023 3669 17032
rect 3819 17072 3861 17081
rect 3819 17032 3820 17072
rect 3860 17032 3861 17072
rect 3819 17023 3861 17032
rect 3915 17072 3957 17081
rect 3915 17032 3916 17072
rect 3956 17032 3957 17072
rect 3915 17023 3957 17032
rect 4291 17072 4349 17073
rect 4291 17032 4300 17072
rect 4340 17032 4349 17072
rect 4291 17031 4349 17032
rect 4683 17072 4725 17081
rect 4683 17032 4684 17072
rect 4724 17032 4725 17072
rect 4683 17023 4725 17032
rect 4779 17072 4821 17081
rect 4779 17032 4780 17072
rect 4820 17032 4821 17072
rect 4779 17023 4821 17032
rect 4875 17072 4917 17081
rect 4875 17032 4876 17072
rect 4916 17032 4917 17072
rect 4875 17023 4917 17032
rect 4971 17072 5013 17081
rect 4971 17032 4972 17072
rect 5012 17032 5013 17072
rect 4971 17023 5013 17032
rect 5643 17072 5685 17081
rect 5643 17032 5644 17072
rect 5684 17032 5685 17072
rect 5643 17023 5685 17032
rect 5739 17072 5781 17081
rect 5739 17032 5740 17072
rect 5780 17032 5781 17072
rect 5739 17023 5781 17032
rect 5931 17072 5973 17081
rect 5931 17032 5932 17072
rect 5972 17032 5973 17072
rect 5931 17023 5973 17032
rect 6115 17072 6173 17073
rect 6115 17032 6124 17072
rect 6164 17032 6173 17072
rect 6115 17031 6173 17032
rect 6795 17072 6837 17081
rect 6795 17032 6796 17072
rect 6836 17032 6837 17072
rect 6795 17023 6837 17032
rect 7651 17072 7709 17073
rect 7651 17032 7660 17072
rect 7700 17032 7709 17072
rect 7651 17031 7709 17032
rect 7851 17072 7893 17081
rect 7851 17032 7852 17072
rect 7892 17032 7893 17072
rect 7851 17023 7893 17032
rect 7947 17072 7989 17081
rect 7947 17032 7948 17072
rect 7988 17032 7989 17072
rect 7947 17023 7989 17032
rect 8043 17072 8085 17081
rect 8043 17032 8044 17072
rect 8084 17032 8085 17072
rect 8043 17023 8085 17032
rect 8139 17072 8181 17081
rect 8139 17032 8140 17072
rect 8180 17032 8181 17072
rect 8139 17023 8181 17032
rect 8323 17072 8381 17073
rect 8323 17032 8332 17072
rect 8372 17032 8381 17072
rect 8323 17031 8381 17032
rect 8523 17072 8565 17081
rect 8523 17032 8524 17072
rect 8564 17032 8565 17072
rect 8523 17023 8565 17032
rect 11203 17072 11261 17073
rect 11203 17032 11212 17072
rect 11252 17032 11261 17072
rect 11203 17031 11261 17032
rect 11595 17072 11637 17081
rect 11595 17032 11596 17072
rect 11636 17032 11637 17072
rect 11595 17023 11637 17032
rect 12451 17072 12509 17073
rect 12451 17032 12460 17072
rect 12500 17032 12509 17072
rect 12451 17031 12509 17032
rect 12643 17072 12701 17073
rect 12643 17032 12652 17072
rect 12692 17032 12701 17072
rect 12643 17031 12701 17032
rect 13603 17072 13661 17073
rect 13603 17032 13612 17072
rect 13652 17032 13661 17072
rect 13603 17031 13661 17032
rect 15235 17072 15293 17073
rect 15235 17032 15244 17072
rect 15284 17032 15293 17072
rect 15235 17031 15293 17032
rect 15427 17072 15485 17073
rect 15427 17032 15436 17072
rect 15476 17032 15485 17072
rect 15427 17031 15485 17032
rect 16675 17072 16733 17073
rect 16675 17032 16684 17072
rect 16724 17032 16733 17072
rect 16675 17031 16733 17032
rect 17539 17072 17597 17073
rect 17539 17032 17548 17072
rect 17588 17032 17597 17072
rect 17539 17031 17597 17032
rect 17931 17072 17973 17081
rect 17931 17032 17932 17072
rect 17972 17032 17973 17072
rect 17931 17023 17973 17032
rect 18307 17072 18365 17073
rect 18307 17032 18316 17072
rect 18356 17032 18365 17072
rect 18307 17031 18365 17032
rect 20035 17072 20093 17073
rect 20035 17032 20044 17072
rect 20084 17032 20093 17072
rect 20035 17031 20093 17032
rect 20331 17072 20373 17081
rect 20331 17032 20332 17072
rect 20372 17032 20373 17072
rect 20331 17023 20373 17032
rect 20523 17072 20565 17081
rect 20523 17032 20524 17072
rect 20564 17032 20565 17072
rect 20523 17023 20565 17032
rect 20611 17072 20669 17073
rect 20611 17032 20620 17072
rect 20660 17032 20669 17072
rect 20611 17031 20669 17032
rect 20907 17072 20949 17081
rect 20907 17032 20908 17072
rect 20948 17032 20949 17072
rect 20907 17023 20949 17032
rect 21003 17072 21045 17081
rect 21003 17032 21004 17072
rect 21044 17032 21045 17072
rect 21003 17023 21045 17032
rect 21099 17072 21141 17081
rect 21099 17032 21100 17072
rect 21140 17032 21141 17072
rect 21099 17023 21141 17032
rect 21483 17072 21525 17081
rect 21483 17032 21484 17072
rect 21524 17032 21525 17072
rect 21483 17023 21525 17032
rect 22531 17072 22589 17073
rect 22531 17032 22540 17072
rect 22580 17032 22589 17072
rect 22531 17031 22589 17032
rect 23499 17072 23541 17081
rect 23499 17032 23500 17072
rect 23540 17032 23541 17072
rect 23499 17023 23541 17032
rect 23595 17072 23637 17081
rect 23595 17032 23596 17072
rect 23636 17032 23637 17072
rect 23595 17023 23637 17032
rect 23691 17072 23733 17081
rect 23691 17032 23692 17072
rect 23732 17032 23733 17072
rect 23691 17023 23733 17032
rect 23883 17072 23925 17081
rect 23883 17032 23884 17072
rect 23924 17032 23925 17072
rect 23883 17023 23925 17032
rect 23979 17072 24021 17081
rect 23979 17032 23980 17072
rect 24020 17032 24021 17072
rect 23979 17023 24021 17032
rect 24075 17072 24117 17081
rect 24075 17032 24076 17072
rect 24116 17032 24117 17072
rect 24075 17023 24117 17032
rect 24363 17072 24405 17081
rect 24363 17032 24364 17072
rect 24404 17032 24405 17072
rect 24363 17023 24405 17032
rect 24459 17072 24501 17081
rect 24459 17032 24460 17072
rect 24500 17032 24501 17072
rect 24459 17023 24501 17032
rect 24555 17072 24597 17081
rect 24555 17032 24556 17072
rect 24596 17032 24597 17072
rect 24555 17023 24597 17032
rect 25219 17072 25277 17073
rect 25219 17032 25228 17072
rect 25268 17032 25277 17072
rect 25219 17031 25277 17032
rect 25323 17072 25365 17081
rect 25323 17032 25324 17072
rect 25364 17032 25365 17072
rect 25323 17023 25365 17032
rect 25515 17072 25557 17081
rect 25515 17032 25516 17072
rect 25556 17032 25557 17072
rect 25515 17023 25557 17032
rect 26475 17072 26517 17081
rect 26475 17032 26476 17072
rect 26516 17032 26517 17072
rect 26475 17023 26517 17032
rect 26667 17072 26709 17081
rect 26667 17032 26668 17072
rect 26708 17032 26709 17072
rect 26667 17023 26709 17032
rect 26755 17072 26813 17073
rect 26755 17032 26764 17072
rect 26804 17032 26813 17072
rect 26755 17031 26813 17032
rect 27235 17072 27293 17073
rect 27235 17032 27244 17072
rect 27284 17032 27293 17072
rect 27235 17031 27293 17032
rect 27331 17072 27389 17073
rect 27331 17032 27340 17072
rect 27380 17032 27389 17072
rect 27331 17031 27389 17032
rect 27915 17072 27957 17081
rect 27915 17032 27916 17072
rect 27956 17032 27957 17072
rect 27811 17030 27869 17031
rect 3339 16988 3381 16997
rect 27811 16990 27820 17030
rect 27860 16990 27869 17030
rect 27915 17023 27957 17032
rect 28766 17072 28824 17073
rect 28766 17032 28775 17072
rect 28815 17032 28824 17072
rect 28766 17031 28824 17032
rect 28875 17072 28917 17081
rect 28875 17032 28876 17072
rect 28916 17032 28917 17072
rect 28875 17023 28917 17032
rect 28971 17072 29013 17081
rect 28971 17032 28972 17072
rect 29012 17032 29013 17072
rect 28971 17023 29013 17032
rect 29155 17072 29213 17073
rect 29155 17032 29164 17072
rect 29204 17032 29213 17072
rect 29155 17031 29213 17032
rect 29251 17072 29309 17073
rect 29251 17032 29260 17072
rect 29300 17032 29309 17072
rect 29251 17031 29309 17032
rect 30403 17072 30461 17073
rect 30403 17032 30412 17072
rect 30452 17032 30461 17072
rect 30403 17031 30461 17032
rect 31171 17072 31229 17073
rect 31171 17032 31180 17072
rect 31220 17032 31229 17072
rect 31171 17031 31229 17032
rect 31363 17072 31421 17073
rect 31363 17032 31372 17072
rect 31412 17032 31421 17072
rect 31363 17031 31421 17032
rect 31651 17072 31709 17073
rect 31651 17032 31660 17072
rect 31700 17032 31709 17072
rect 31651 17031 31709 17032
rect 31947 17072 31989 17081
rect 31947 17032 31948 17072
rect 31988 17032 31989 17072
rect 31947 17023 31989 17032
rect 32043 17072 32085 17081
rect 32043 17032 32044 17072
rect 32084 17032 32085 17072
rect 32043 17023 32085 17032
rect 32139 17072 32181 17081
rect 32139 17032 32140 17072
rect 32180 17032 32181 17072
rect 32139 17023 32181 17032
rect 32235 17072 32277 17081
rect 32235 17032 32236 17072
rect 32276 17032 32277 17072
rect 32235 17023 32277 17032
rect 33379 17072 33437 17073
rect 33379 17032 33388 17072
rect 33428 17032 33437 17072
rect 33379 17031 33437 17032
rect 33763 17072 33821 17073
rect 33763 17032 33772 17072
rect 33812 17032 33821 17072
rect 33763 17031 33821 17032
rect 34923 17072 34965 17081
rect 34923 17032 34924 17072
rect 34964 17032 34965 17072
rect 34923 17023 34965 17032
rect 35107 17072 35165 17073
rect 35107 17032 35116 17072
rect 35156 17032 35165 17072
rect 35107 17031 35165 17032
rect 35875 17072 35933 17073
rect 35875 17032 35884 17072
rect 35924 17032 35933 17072
rect 35875 17031 35933 17032
rect 36075 17072 36117 17081
rect 36075 17032 36076 17072
rect 36116 17032 36117 17072
rect 36075 17023 36117 17032
rect 36299 17072 36357 17073
rect 36299 17032 36308 17072
rect 36348 17032 36357 17072
rect 36299 17031 36357 17032
rect 36459 17072 36501 17081
rect 36459 17032 36460 17072
rect 36500 17032 36501 17072
rect 36459 17023 36501 17032
rect 36555 17072 36597 17081
rect 36555 17032 36556 17072
rect 36596 17032 36597 17072
rect 36555 17023 36597 17032
rect 36739 17072 36797 17073
rect 36739 17032 36748 17072
rect 36788 17032 36797 17072
rect 36739 17031 36797 17032
rect 36835 17072 36893 17073
rect 36835 17032 36844 17072
rect 36884 17032 36893 17072
rect 36835 17031 36893 17032
rect 37064 17072 37122 17073
rect 37064 17032 37073 17072
rect 37113 17032 37122 17072
rect 37064 17031 37122 17032
rect 37227 17072 37269 17081
rect 37227 17032 37228 17072
rect 37268 17032 37269 17072
rect 37603 17072 37661 17073
rect 37227 17023 37269 17032
rect 37323 17057 37365 17066
rect 37323 17017 37324 17057
rect 37364 17017 37365 17057
rect 37323 17008 37365 17017
rect 37515 17057 37557 17066
rect 37515 17017 37516 17057
rect 37556 17017 37557 17057
rect 37603 17032 37612 17072
rect 37652 17032 37661 17072
rect 37603 17031 37661 17032
rect 38187 17072 38229 17081
rect 38187 17032 38188 17072
rect 38228 17032 38229 17072
rect 38187 17023 38229 17032
rect 38379 17072 38421 17081
rect 38379 17032 38380 17072
rect 38420 17032 38421 17072
rect 38379 17023 38421 17032
rect 38467 17072 38525 17073
rect 38467 17032 38476 17072
rect 38516 17032 38525 17072
rect 38467 17031 38525 17032
rect 39619 17072 39677 17073
rect 39619 17032 39628 17072
rect 39668 17032 39677 17072
rect 39619 17031 39677 17032
rect 39915 17072 39957 17081
rect 39915 17032 39916 17072
rect 39956 17032 39957 17072
rect 39915 17023 39957 17032
rect 40291 17072 40349 17073
rect 40291 17032 40300 17072
rect 40340 17032 40349 17072
rect 40291 17031 40349 17032
rect 41155 17072 41213 17073
rect 41155 17032 41164 17072
rect 41204 17032 41213 17072
rect 41155 17031 41213 17032
rect 37515 17008 37557 17017
rect 27811 16989 27869 16990
rect 3339 16948 3340 16988
rect 3380 16948 3381 16988
rect 3339 16939 3381 16948
rect 29547 16988 29589 16997
rect 29547 16948 29548 16988
rect 29588 16948 29589 16988
rect 29547 16939 29589 16948
rect 31555 16988 31613 16989
rect 31555 16948 31564 16988
rect 31604 16948 31613 16988
rect 31555 16947 31613 16948
rect 37987 16988 38045 16989
rect 37987 16948 37996 16988
rect 38036 16948 38045 16988
rect 37987 16947 38045 16948
rect 9867 16904 9909 16913
rect 9867 16864 9868 16904
rect 9908 16864 9909 16904
rect 9867 16855 9909 16864
rect 14379 16904 14421 16913
rect 14379 16864 14380 16904
rect 14420 16864 14421 16904
rect 14379 16855 14421 16864
rect 20331 16904 20373 16913
rect 20331 16864 20332 16904
rect 20372 16864 20373 16904
rect 20331 16855 20373 16864
rect 34443 16904 34485 16913
rect 34443 16864 34444 16904
rect 34484 16864 34485 16904
rect 34443 16855 34485 16864
rect 5155 16820 5213 16821
rect 5155 16780 5164 16820
rect 5204 16780 5213 16820
rect 5155 16779 5213 16780
rect 6979 16820 7037 16821
rect 6979 16780 6988 16820
rect 7028 16780 7037 16820
rect 6979 16779 7037 16780
rect 8427 16820 8469 16829
rect 8427 16780 8428 16820
rect 8468 16780 8469 16820
rect 8427 16771 8469 16780
rect 10531 16820 10589 16821
rect 10531 16780 10540 16820
rect 10580 16780 10589 16820
rect 10531 16779 10589 16780
rect 14563 16820 14621 16821
rect 14563 16780 14572 16820
rect 14612 16780 14621 16820
rect 14563 16779 14621 16780
rect 18979 16820 19037 16821
rect 18979 16780 18988 16820
rect 19028 16780 19037 16820
rect 18979 16779 19037 16780
rect 21675 16820 21717 16829
rect 21675 16780 21676 16820
rect 21716 16780 21717 16820
rect 21675 16771 21717 16780
rect 23203 16820 23261 16821
rect 23203 16780 23212 16820
rect 23252 16780 23261 16820
rect 23203 16779 23261 16780
rect 27435 16820 27477 16829
rect 27435 16780 27436 16820
rect 27476 16780 27477 16820
rect 27435 16771 27477 16780
rect 28203 16820 28245 16829
rect 28203 16780 28204 16820
rect 28244 16780 28245 16820
rect 28203 16771 28245 16780
rect 29259 16820 29301 16829
rect 29259 16780 29260 16820
rect 29300 16780 29301 16820
rect 29259 16771 29301 16780
rect 32907 16820 32949 16829
rect 32907 16780 32908 16820
rect 32948 16780 32949 16820
rect 32907 16771 32949 16780
rect 34059 16820 34101 16829
rect 34059 16780 34060 16820
rect 34100 16780 34101 16820
rect 34059 16771 34101 16780
rect 35979 16820 36021 16829
rect 35979 16780 35980 16820
rect 36020 16780 36021 16820
rect 35979 16771 36021 16780
rect 37611 16820 37653 16829
rect 37611 16780 37612 16820
rect 37652 16780 37653 16820
rect 37611 16771 37653 16780
rect 39147 16820 39189 16829
rect 39147 16780 39148 16820
rect 39188 16780 39189 16820
rect 39147 16771 39189 16780
rect 42315 16820 42357 16829
rect 42315 16780 42316 16820
rect 42356 16780 42357 16820
rect 42315 16771 42357 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 6411 16484 6453 16493
rect 6411 16444 6412 16484
rect 6452 16444 6453 16484
rect 6411 16435 6453 16444
rect 8139 16484 8181 16493
rect 8139 16444 8140 16484
rect 8180 16444 8181 16484
rect 8139 16435 8181 16444
rect 8427 16484 8469 16493
rect 8427 16444 8428 16484
rect 8468 16444 8469 16484
rect 8427 16435 8469 16444
rect 11779 16484 11837 16485
rect 11779 16444 11788 16484
rect 11828 16444 11837 16484
rect 11779 16443 11837 16444
rect 15627 16484 15669 16493
rect 15627 16444 15628 16484
rect 15668 16444 15669 16484
rect 15627 16435 15669 16444
rect 26667 16484 26709 16493
rect 26667 16444 26668 16484
rect 26708 16444 26709 16484
rect 26667 16435 26709 16444
rect 1419 16400 1461 16409
rect 1419 16360 1420 16400
rect 1460 16360 1461 16400
rect 1419 16351 1461 16360
rect 5451 16400 5493 16409
rect 5451 16360 5452 16400
rect 5492 16360 5493 16400
rect 5451 16351 5493 16360
rect 12075 16400 12117 16409
rect 12075 16360 12076 16400
rect 12116 16360 12117 16400
rect 12075 16351 12117 16360
rect 13035 16400 13077 16409
rect 13035 16360 13036 16400
rect 13076 16360 13077 16400
rect 13035 16351 13077 16360
rect 16491 16400 16533 16409
rect 16491 16360 16492 16400
rect 16532 16360 16533 16400
rect 16491 16351 16533 16360
rect 20331 16400 20373 16409
rect 20331 16360 20332 16400
rect 20372 16360 20373 16400
rect 20331 16351 20373 16360
rect 21387 16400 21429 16409
rect 21387 16360 21388 16400
rect 21428 16360 21429 16400
rect 21387 16351 21429 16360
rect 21963 16400 22005 16409
rect 21963 16360 21964 16400
rect 22004 16360 22005 16400
rect 21963 16351 22005 16360
rect 22155 16400 22197 16409
rect 22155 16360 22156 16400
rect 22196 16360 22197 16400
rect 22155 16351 22197 16360
rect 37035 16400 37077 16409
rect 37035 16360 37036 16400
rect 37076 16360 37077 16400
rect 37035 16351 37077 16360
rect 38475 16400 38517 16409
rect 38475 16360 38476 16400
rect 38516 16360 38517 16400
rect 38475 16351 38517 16360
rect 39427 16400 39485 16401
rect 39427 16360 39436 16400
rect 39476 16360 39485 16400
rect 39427 16359 39485 16360
rect 41163 16400 41205 16409
rect 41163 16360 41164 16400
rect 41204 16360 41205 16400
rect 41163 16351 41205 16360
rect 6603 16316 6645 16325
rect 6603 16276 6604 16316
rect 6644 16276 6645 16316
rect 6603 16267 6645 16276
rect 20235 16316 20277 16325
rect 20235 16276 20236 16316
rect 20276 16276 20277 16316
rect 20235 16267 20277 16276
rect 20427 16316 20469 16325
rect 20427 16276 20428 16316
rect 20468 16276 20469 16316
rect 20427 16267 20469 16276
rect 21291 16316 21333 16325
rect 21291 16276 21292 16316
rect 21332 16276 21333 16316
rect 21291 16267 21333 16276
rect 21483 16316 21525 16325
rect 21483 16276 21484 16316
rect 21524 16276 21525 16316
rect 21483 16267 21525 16276
rect 27715 16316 27773 16317
rect 27715 16276 27724 16316
rect 27764 16276 27773 16316
rect 27715 16275 27773 16276
rect 3051 16232 3093 16241
rect 3051 16192 3052 16232
rect 3092 16192 3093 16232
rect 3051 16183 3093 16192
rect 3243 16232 3285 16241
rect 3243 16192 3244 16232
rect 3284 16192 3285 16232
rect 3243 16183 3285 16192
rect 3435 16232 3477 16241
rect 3435 16192 3436 16232
rect 3476 16192 3477 16232
rect 3435 16183 3477 16192
rect 3627 16232 3669 16241
rect 3627 16192 3628 16232
rect 3668 16192 3669 16232
rect 3627 16183 3669 16192
rect 3723 16232 3765 16241
rect 3723 16192 3724 16232
rect 3764 16192 3765 16232
rect 3723 16183 3765 16192
rect 4011 16232 4053 16241
rect 4011 16192 4012 16232
rect 4052 16192 4053 16232
rect 4011 16183 4053 16192
rect 4675 16232 4733 16233
rect 4675 16192 4684 16232
rect 4724 16192 4733 16232
rect 4675 16191 4733 16192
rect 4971 16232 5013 16241
rect 4971 16192 4972 16232
rect 5012 16192 5013 16232
rect 4971 16183 5013 16192
rect 5163 16232 5205 16241
rect 5163 16192 5164 16232
rect 5204 16192 5205 16232
rect 5163 16183 5205 16192
rect 5451 16232 5493 16241
rect 5451 16192 5452 16232
rect 5492 16192 5493 16232
rect 5451 16183 5493 16192
rect 5643 16232 5685 16241
rect 5643 16192 5644 16232
rect 5684 16192 5685 16232
rect 5643 16183 5685 16192
rect 5731 16232 5789 16233
rect 5731 16192 5740 16232
rect 5780 16192 5789 16232
rect 5731 16191 5789 16192
rect 5931 16232 5973 16241
rect 5931 16192 5932 16232
rect 5972 16192 5973 16232
rect 5931 16183 5973 16192
rect 6123 16232 6165 16241
rect 6123 16192 6124 16232
rect 6164 16192 6165 16232
rect 6123 16183 6165 16192
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 7083 16232 7125 16241
rect 7083 16192 7084 16232
rect 7124 16192 7125 16232
rect 7083 16183 7125 16192
rect 7171 16232 7229 16233
rect 7171 16192 7180 16232
rect 7220 16192 7229 16232
rect 7171 16191 7229 16192
rect 7563 16232 7605 16241
rect 7563 16192 7564 16232
rect 7604 16192 7605 16232
rect 7563 16183 7605 16192
rect 7843 16232 7901 16233
rect 7843 16192 7852 16232
rect 7892 16192 7901 16232
rect 7843 16191 7901 16192
rect 7947 16232 7989 16241
rect 7947 16192 7948 16232
rect 7988 16192 7989 16232
rect 7947 16183 7989 16192
rect 8131 16232 8189 16233
rect 8131 16192 8140 16232
rect 8180 16192 8189 16232
rect 8131 16191 8189 16192
rect 8323 16232 8381 16233
rect 8323 16192 8332 16232
rect 8372 16192 8381 16232
rect 8323 16191 8381 16192
rect 8515 16232 8573 16233
rect 8515 16192 8524 16232
rect 8564 16192 8573 16232
rect 8515 16191 8573 16192
rect 9387 16232 9429 16241
rect 9387 16192 9388 16232
rect 9428 16192 9429 16232
rect 9387 16183 9429 16192
rect 9763 16232 9821 16233
rect 9763 16192 9772 16232
rect 9812 16192 9821 16232
rect 9763 16191 9821 16192
rect 10627 16232 10685 16233
rect 10627 16192 10636 16232
rect 10676 16192 10685 16232
rect 10627 16191 10685 16192
rect 12075 16232 12117 16241
rect 12075 16192 12076 16232
rect 12116 16192 12117 16232
rect 12075 16183 12117 16192
rect 12267 16232 12309 16241
rect 12267 16192 12268 16232
rect 12308 16192 12309 16232
rect 12267 16183 12309 16192
rect 12355 16232 12413 16233
rect 12355 16192 12364 16232
rect 12404 16192 12413 16232
rect 12355 16191 12413 16192
rect 13219 16232 13277 16233
rect 13219 16192 13228 16232
rect 13268 16192 13277 16232
rect 13219 16191 13277 16192
rect 14091 16232 14133 16241
rect 14091 16192 14092 16232
rect 14132 16192 14133 16232
rect 14091 16183 14133 16192
rect 15331 16232 15389 16233
rect 15331 16192 15340 16232
rect 15380 16192 15389 16232
rect 15331 16191 15389 16192
rect 16491 16232 16533 16241
rect 16491 16192 16492 16232
rect 16532 16192 16533 16232
rect 16491 16183 16533 16192
rect 16683 16232 16725 16241
rect 16683 16192 16684 16232
rect 16724 16192 16725 16232
rect 16683 16183 16725 16192
rect 18595 16232 18653 16233
rect 18595 16192 18604 16232
rect 18644 16192 18653 16232
rect 18595 16191 18653 16192
rect 18883 16232 18941 16233
rect 18883 16192 18892 16232
rect 18932 16192 18941 16232
rect 18883 16191 18941 16192
rect 19363 16232 19421 16233
rect 19363 16192 19372 16232
rect 19412 16192 19421 16232
rect 19363 16191 19421 16192
rect 19651 16232 19709 16233
rect 19651 16192 19660 16232
rect 19700 16192 19709 16232
rect 19651 16191 19709 16192
rect 20523 16232 20565 16241
rect 20523 16192 20524 16232
rect 20564 16192 20565 16232
rect 20131 16190 20189 16191
rect 3147 16148 3189 16157
rect 20131 16150 20140 16190
rect 20180 16150 20189 16190
rect 20523 16183 20565 16192
rect 20715 16232 20757 16241
rect 20715 16192 20716 16232
rect 20756 16192 20757 16232
rect 20715 16183 20757 16192
rect 20811 16232 20853 16241
rect 20811 16192 20812 16232
rect 20852 16192 20853 16232
rect 20811 16183 20853 16192
rect 20907 16232 20949 16241
rect 20907 16192 20908 16232
rect 20948 16192 20949 16232
rect 20907 16183 20949 16192
rect 21003 16232 21045 16241
rect 21003 16192 21004 16232
rect 21044 16192 21045 16232
rect 21003 16183 21045 16192
rect 21195 16232 21237 16241
rect 21195 16192 21196 16232
rect 21236 16192 21237 16232
rect 21195 16183 21237 16192
rect 21571 16232 21629 16233
rect 21571 16192 21580 16232
rect 21620 16192 21629 16232
rect 21571 16191 21629 16192
rect 21963 16232 22005 16241
rect 21963 16192 21964 16232
rect 22004 16192 22005 16232
rect 21963 16183 22005 16192
rect 22339 16232 22397 16233
rect 22339 16192 22348 16232
rect 22388 16192 22397 16232
rect 22339 16191 22397 16192
rect 22443 16232 22485 16241
rect 22443 16192 22444 16232
rect 22484 16192 22485 16232
rect 22443 16183 22485 16192
rect 22635 16232 22677 16241
rect 22635 16192 22636 16232
rect 22676 16192 22677 16232
rect 22635 16183 22677 16192
rect 22827 16232 22869 16241
rect 22827 16192 22828 16232
rect 22868 16192 22869 16232
rect 22827 16183 22869 16192
rect 22923 16232 22965 16241
rect 22923 16192 22924 16232
rect 22964 16192 22965 16232
rect 22923 16183 22965 16192
rect 23395 16232 23453 16233
rect 23395 16192 23404 16232
rect 23444 16192 23453 16232
rect 23395 16191 23453 16192
rect 24355 16232 24413 16233
rect 24355 16192 24364 16232
rect 24404 16192 24413 16232
rect 24355 16191 24413 16192
rect 24739 16232 24797 16233
rect 24739 16192 24748 16232
rect 24788 16192 24797 16232
rect 24739 16191 24797 16192
rect 26187 16232 26229 16241
rect 26187 16192 26188 16232
rect 26228 16192 26229 16232
rect 26187 16183 26229 16192
rect 26283 16232 26325 16241
rect 26283 16192 26284 16232
rect 26324 16192 26325 16232
rect 26283 16183 26325 16192
rect 26379 16232 26421 16241
rect 26379 16192 26380 16232
rect 26420 16192 26421 16232
rect 26379 16183 26421 16192
rect 26475 16232 26517 16241
rect 26475 16192 26476 16232
rect 26516 16192 26517 16232
rect 26475 16183 26517 16192
rect 26667 16232 26709 16241
rect 26667 16192 26668 16232
rect 26708 16192 26709 16232
rect 26667 16183 26709 16192
rect 26859 16232 26901 16241
rect 26859 16192 26860 16232
rect 26900 16192 26901 16232
rect 26859 16183 26901 16192
rect 26947 16232 27005 16233
rect 26947 16192 26956 16232
rect 26996 16192 27005 16232
rect 26947 16191 27005 16192
rect 27427 16232 27485 16233
rect 27427 16192 27436 16232
rect 27476 16192 27485 16232
rect 27427 16191 27485 16192
rect 27523 16232 27581 16233
rect 27523 16192 27532 16232
rect 27572 16192 27581 16232
rect 27523 16191 27581 16192
rect 27907 16232 27965 16233
rect 27907 16192 27916 16232
rect 27956 16192 27965 16232
rect 27907 16191 27965 16192
rect 28011 16232 28053 16241
rect 28011 16192 28012 16232
rect 28052 16192 28053 16232
rect 28011 16183 28053 16192
rect 28195 16232 28253 16233
rect 28195 16192 28204 16232
rect 28244 16192 28253 16232
rect 28195 16191 28253 16192
rect 28387 16232 28445 16233
rect 28387 16192 28396 16232
rect 28436 16192 28445 16232
rect 28387 16191 28445 16192
rect 28491 16232 28533 16241
rect 28491 16192 28492 16232
rect 28532 16192 28533 16232
rect 28491 16183 28533 16192
rect 28675 16232 28733 16233
rect 28675 16192 28684 16232
rect 28724 16192 28733 16232
rect 28675 16191 28733 16192
rect 28963 16232 29021 16233
rect 28963 16192 28972 16232
rect 29012 16192 29021 16232
rect 28963 16191 29021 16192
rect 29067 16232 29109 16241
rect 29067 16192 29068 16232
rect 29108 16192 29109 16232
rect 29067 16183 29109 16192
rect 29259 16232 29301 16241
rect 29259 16192 29260 16232
rect 29300 16192 29301 16232
rect 29259 16183 29301 16192
rect 29931 16232 29973 16241
rect 29931 16192 29932 16232
rect 29972 16192 29973 16232
rect 29931 16183 29973 16192
rect 30027 16232 30069 16241
rect 30027 16192 30028 16232
rect 30068 16192 30069 16232
rect 30027 16183 30069 16192
rect 30123 16232 30165 16241
rect 30123 16192 30124 16232
rect 30164 16192 30165 16232
rect 30123 16183 30165 16192
rect 30507 16232 30549 16241
rect 30507 16192 30508 16232
rect 30548 16192 30549 16232
rect 30507 16183 30549 16192
rect 32427 16232 32469 16241
rect 32427 16192 32428 16232
rect 32468 16192 32469 16232
rect 32427 16183 32469 16192
rect 32803 16232 32861 16233
rect 32803 16192 32812 16232
rect 32852 16192 32861 16232
rect 32803 16191 32861 16192
rect 32907 16232 32949 16241
rect 32907 16192 32908 16232
rect 32948 16192 32949 16232
rect 32907 16183 32949 16192
rect 33099 16232 33141 16241
rect 33099 16192 33100 16232
rect 33140 16192 33141 16232
rect 33099 16183 33141 16192
rect 33283 16232 33341 16233
rect 33283 16192 33292 16232
rect 33332 16192 33341 16232
rect 33283 16191 33341 16192
rect 33483 16232 33525 16241
rect 33483 16192 33484 16232
rect 33524 16192 33525 16232
rect 33483 16183 33525 16192
rect 33571 16232 33629 16233
rect 33571 16192 33580 16232
rect 33620 16192 33629 16232
rect 33571 16191 33629 16192
rect 33763 16232 33821 16233
rect 33763 16192 33772 16232
rect 33812 16192 33821 16232
rect 33763 16191 33821 16192
rect 33963 16232 34005 16241
rect 33963 16192 33964 16232
rect 34004 16192 34005 16232
rect 33963 16183 34005 16192
rect 34051 16232 34109 16233
rect 34051 16192 34060 16232
rect 34100 16192 34109 16232
rect 34051 16191 34109 16192
rect 34627 16232 34685 16233
rect 34627 16192 34636 16232
rect 34676 16192 34685 16232
rect 34627 16191 34685 16192
rect 35587 16232 35645 16233
rect 35587 16192 35596 16232
rect 35636 16192 35645 16232
rect 35587 16191 35645 16192
rect 35787 16232 35829 16241
rect 35787 16192 35788 16232
rect 35828 16192 35829 16232
rect 35787 16183 35829 16192
rect 35979 16232 36021 16241
rect 35979 16192 35980 16232
rect 36020 16192 36021 16232
rect 35979 16183 36021 16192
rect 36067 16232 36125 16233
rect 36067 16192 36076 16232
rect 36116 16192 36125 16232
rect 36067 16191 36125 16192
rect 36267 16232 36309 16241
rect 36267 16192 36268 16232
rect 36308 16192 36309 16232
rect 36267 16183 36309 16192
rect 36363 16232 36405 16241
rect 36363 16192 36364 16232
rect 36404 16192 36405 16232
rect 36363 16183 36405 16192
rect 36459 16232 36501 16241
rect 36459 16192 36460 16232
rect 36500 16192 36501 16232
rect 36459 16183 36501 16192
rect 36555 16232 36597 16241
rect 36555 16192 36556 16232
rect 36596 16192 36597 16232
rect 36555 16183 36597 16192
rect 36939 16232 36981 16241
rect 36939 16192 36940 16232
rect 36980 16192 36981 16232
rect 36939 16183 36981 16192
rect 37123 16232 37181 16233
rect 37123 16192 37132 16232
rect 37172 16192 37181 16232
rect 37123 16191 37181 16192
rect 37323 16232 37365 16241
rect 37323 16192 37324 16232
rect 37364 16192 37365 16232
rect 37323 16183 37365 16192
rect 37419 16232 37461 16241
rect 37419 16192 37420 16232
rect 37460 16192 37461 16232
rect 37419 16183 37461 16192
rect 37515 16232 37557 16241
rect 37515 16192 37516 16232
rect 37556 16192 37557 16232
rect 37515 16183 37557 16192
rect 37611 16232 37653 16241
rect 37611 16192 37612 16232
rect 37652 16192 37653 16232
rect 37611 16183 37653 16192
rect 38083 16232 38141 16233
rect 38083 16192 38092 16232
rect 38132 16192 38141 16232
rect 38083 16191 38141 16192
rect 38187 16232 38229 16241
rect 38187 16192 38188 16232
rect 38228 16192 38229 16232
rect 38187 16183 38229 16192
rect 38947 16232 39005 16233
rect 38947 16192 38956 16232
rect 38996 16192 39005 16232
rect 38947 16191 39005 16192
rect 39147 16232 39189 16241
rect 39147 16192 39148 16232
rect 39188 16192 39189 16232
rect 39147 16183 39189 16192
rect 39235 16232 39293 16233
rect 39235 16192 39244 16232
rect 39284 16192 39293 16232
rect 39235 16191 39293 16192
rect 40099 16232 40157 16233
rect 40099 16192 40108 16232
rect 40148 16192 40157 16232
rect 40099 16191 40157 16192
rect 40299 16232 40341 16241
rect 40299 16192 40300 16232
rect 40340 16192 40341 16232
rect 40299 16183 40341 16192
rect 40963 16232 41021 16233
rect 40963 16192 40972 16232
rect 41012 16192 41021 16232
rect 40963 16191 41021 16192
rect 20131 16149 20189 16150
rect 3147 16108 3148 16148
rect 3188 16108 3189 16148
rect 3147 16099 3189 16108
rect 16195 16148 16253 16149
rect 16195 16108 16204 16148
rect 16244 16108 16253 16148
rect 16195 16107 16253 16108
rect 19075 16148 19133 16149
rect 19075 16108 19084 16148
rect 19124 16108 19133 16148
rect 19075 16107 19133 16108
rect 19843 16148 19901 16149
rect 19843 16108 19852 16148
rect 19892 16108 19901 16148
rect 19843 16107 19901 16108
rect 24547 16148 24605 16149
rect 24547 16108 24556 16148
rect 24596 16108 24605 16148
rect 24547 16107 24605 16108
rect 29163 16148 29205 16157
rect 29163 16108 29164 16148
rect 29204 16108 29205 16148
rect 29163 16099 29205 16108
rect 31651 16148 31709 16149
rect 31651 16108 31660 16148
rect 31700 16108 31709 16148
rect 31651 16107 31709 16108
rect 33003 16148 33045 16157
rect 33003 16108 33004 16148
rect 33044 16108 33045 16148
rect 33003 16099 33045 16108
rect 35883 16148 35925 16157
rect 35883 16108 35884 16148
rect 35924 16108 35925 16148
rect 35883 16099 35925 16108
rect 643 16064 701 16065
rect 643 16024 652 16064
rect 692 16024 701 16064
rect 643 16023 701 16024
rect 3531 16064 3573 16073
rect 3531 16024 3532 16064
rect 3572 16024 3573 16064
rect 3531 16015 3573 16024
rect 5067 16064 5109 16073
rect 5067 16024 5068 16064
rect 5108 16024 5109 16064
rect 5067 16015 5109 16024
rect 6027 16064 6069 16073
rect 6027 16024 6028 16064
rect 6068 16024 6069 16064
rect 6027 16015 6069 16024
rect 22531 16064 22589 16065
rect 22531 16024 22540 16064
rect 22580 16024 22589 16064
rect 22531 16023 22589 16024
rect 23107 16064 23165 16065
rect 23107 16024 23116 16064
rect 23156 16024 23165 16064
rect 23107 16023 23165 16024
rect 24835 16064 24893 16065
rect 24835 16024 24844 16064
rect 24884 16024 24893 16064
rect 24835 16023 24893 16024
rect 28203 16064 28245 16073
rect 28203 16024 28204 16064
rect 28244 16024 28245 16064
rect 28203 16015 28245 16024
rect 28683 16064 28725 16073
rect 28683 16024 28684 16064
rect 28724 16024 28725 16064
rect 28683 16015 28725 16024
rect 29827 16064 29885 16065
rect 29827 16024 29836 16064
rect 29876 16024 29885 16064
rect 29827 16023 29885 16024
rect 30891 16064 30933 16073
rect 30891 16024 30892 16064
rect 30932 16024 30933 16064
rect 30891 16015 30933 16024
rect 33291 16064 33333 16073
rect 33291 16024 33292 16064
rect 33332 16024 33333 16064
rect 33291 16015 33333 16024
rect 33771 16064 33813 16073
rect 33771 16024 33772 16064
rect 33812 16024 33813 16064
rect 33771 16015 33813 16024
rect 37995 16060 38037 16069
rect 37995 16020 37996 16060
rect 38036 16020 38037 16060
rect 37995 16011 38037 16020
rect 38955 16064 38997 16073
rect 38955 16024 38956 16064
rect 38996 16024 38997 16064
rect 38955 16015 38997 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 21675 15759 21717 15768
rect 7659 15732 7701 15741
rect 3811 15728 3869 15729
rect 3811 15688 3820 15728
rect 3860 15688 3869 15728
rect 3811 15687 3869 15688
rect 4099 15728 4157 15729
rect 4099 15688 4108 15728
rect 4148 15688 4157 15728
rect 4099 15687 4157 15688
rect 7659 15692 7660 15732
rect 7700 15692 7701 15732
rect 7659 15683 7701 15692
rect 8235 15728 8277 15737
rect 8235 15688 8236 15728
rect 8276 15688 8277 15728
rect 8235 15679 8277 15688
rect 11683 15728 11741 15729
rect 11683 15688 11692 15728
rect 11732 15688 11741 15728
rect 11683 15687 11741 15688
rect 19363 15728 19421 15729
rect 19363 15688 19372 15728
rect 19412 15688 19421 15728
rect 19363 15687 19421 15688
rect 19843 15728 19901 15729
rect 19843 15688 19852 15728
rect 19892 15688 19901 15728
rect 19843 15687 19901 15688
rect 20323 15728 20381 15729
rect 20323 15688 20332 15728
rect 20372 15688 20381 15728
rect 21675 15719 21676 15759
rect 21716 15719 21717 15759
rect 21675 15710 21717 15719
rect 23587 15728 23645 15729
rect 20323 15687 20381 15688
rect 23587 15688 23596 15728
rect 23636 15688 23645 15728
rect 23587 15687 23645 15688
rect 23875 15728 23933 15729
rect 23875 15688 23884 15728
rect 23924 15688 23933 15728
rect 23875 15687 23933 15688
rect 25611 15728 25653 15737
rect 25611 15688 25612 15728
rect 25652 15688 25653 15728
rect 25611 15679 25653 15688
rect 27435 15728 27477 15737
rect 27435 15688 27436 15728
rect 27476 15688 27477 15728
rect 27435 15679 27477 15688
rect 27907 15728 27965 15729
rect 27907 15688 27916 15728
rect 27956 15688 27965 15728
rect 27907 15687 27965 15688
rect 30507 15728 30549 15737
rect 33867 15732 33909 15741
rect 30507 15688 30508 15728
rect 30548 15688 30549 15728
rect 30507 15679 30549 15688
rect 32707 15728 32765 15729
rect 32707 15688 32716 15728
rect 32756 15688 32765 15728
rect 32707 15687 32765 15688
rect 33867 15692 33868 15732
rect 33908 15692 33909 15732
rect 33867 15683 33909 15692
rect 35779 15728 35837 15729
rect 35779 15688 35788 15728
rect 35828 15688 35837 15728
rect 35779 15687 35837 15688
rect 36843 15728 36885 15737
rect 36843 15688 36844 15728
rect 36884 15688 36885 15728
rect 36843 15679 36885 15688
rect 38667 15728 38709 15737
rect 38667 15688 38668 15728
rect 38708 15688 38709 15728
rect 38667 15679 38709 15688
rect 19075 15644 19133 15645
rect 19075 15604 19084 15644
rect 19124 15604 19133 15644
rect 19075 15603 19133 15604
rect 19555 15644 19613 15645
rect 19555 15604 19564 15644
rect 19604 15604 19613 15644
rect 19555 15603 19613 15604
rect 21003 15644 21045 15653
rect 21003 15604 21004 15644
rect 21044 15604 21045 15644
rect 21003 15595 21045 15604
rect 25899 15644 25941 15653
rect 25899 15604 25900 15644
rect 25940 15604 25941 15644
rect 25899 15595 25941 15604
rect 939 15560 981 15569
rect 939 15520 940 15560
rect 980 15520 981 15560
rect 939 15511 981 15520
rect 1315 15560 1373 15561
rect 1315 15520 1324 15560
rect 1364 15520 1373 15560
rect 1315 15519 1373 15520
rect 2179 15560 2237 15561
rect 2179 15520 2188 15560
rect 2228 15520 2237 15560
rect 2179 15519 2237 15520
rect 4003 15560 4061 15561
rect 4003 15520 4012 15560
rect 4052 15520 4061 15560
rect 4003 15519 4061 15520
rect 4291 15560 4349 15561
rect 4291 15520 4300 15560
rect 4340 15520 4349 15560
rect 4291 15519 4349 15520
rect 4395 15560 4437 15569
rect 4395 15520 4396 15560
rect 4436 15520 4437 15560
rect 4395 15511 4437 15520
rect 4579 15560 4637 15561
rect 4579 15520 4588 15560
rect 4628 15520 4637 15560
rect 4579 15519 4637 15520
rect 4771 15560 4829 15561
rect 4771 15520 4780 15560
rect 4820 15520 4829 15560
rect 4771 15519 4829 15520
rect 6307 15560 6365 15561
rect 6307 15520 6316 15560
rect 6356 15520 6365 15560
rect 6307 15519 6365 15520
rect 6499 15560 6557 15561
rect 6499 15520 6508 15560
rect 6548 15520 6557 15560
rect 6499 15519 6557 15520
rect 6603 15560 6645 15569
rect 6603 15520 6604 15560
rect 6644 15520 6645 15560
rect 6603 15511 6645 15520
rect 7467 15560 7509 15569
rect 7467 15520 7468 15560
rect 7508 15520 7509 15560
rect 7467 15511 7509 15520
rect 7555 15560 7613 15561
rect 7555 15520 7564 15560
rect 7604 15520 7613 15560
rect 7555 15519 7613 15520
rect 7843 15560 7901 15561
rect 7843 15520 7852 15560
rect 7892 15520 7901 15560
rect 7843 15519 7901 15520
rect 8139 15560 8181 15569
rect 8139 15520 8140 15560
rect 8180 15520 8181 15560
rect 8139 15511 8181 15520
rect 8331 15560 8373 15569
rect 8331 15520 8332 15560
rect 8372 15520 8373 15560
rect 8331 15511 8373 15520
rect 8523 15560 8565 15569
rect 8523 15520 8524 15560
rect 8564 15520 8565 15560
rect 8523 15511 8565 15520
rect 8715 15560 8757 15569
rect 8715 15520 8716 15560
rect 8756 15520 8757 15560
rect 8715 15511 8757 15520
rect 8811 15560 8853 15569
rect 8811 15520 8812 15560
rect 8852 15520 8853 15560
rect 8811 15511 8853 15520
rect 9091 15560 9149 15561
rect 9091 15520 9100 15560
rect 9140 15520 9149 15560
rect 9091 15519 9149 15520
rect 9291 15560 9333 15569
rect 9291 15520 9292 15560
rect 9332 15520 9333 15560
rect 9291 15511 9333 15520
rect 9667 15560 9725 15561
rect 9667 15520 9676 15560
rect 9716 15520 9725 15560
rect 9667 15519 9725 15520
rect 10531 15560 10589 15561
rect 10531 15520 10540 15560
rect 10580 15520 10589 15560
rect 10531 15519 10589 15520
rect 12939 15560 12981 15569
rect 12939 15520 12940 15560
rect 12980 15520 12981 15560
rect 12939 15511 12981 15520
rect 13315 15560 13373 15561
rect 13315 15520 13324 15560
rect 13364 15520 13373 15560
rect 13315 15519 13373 15520
rect 14179 15560 14237 15561
rect 14179 15520 14188 15560
rect 14228 15520 14237 15560
rect 14179 15519 14237 15520
rect 15427 15560 15485 15561
rect 15427 15520 15436 15560
rect 15476 15520 15485 15560
rect 15427 15519 15485 15520
rect 16291 15560 16349 15561
rect 16291 15520 16300 15560
rect 16340 15520 16349 15560
rect 16291 15519 16349 15520
rect 16683 15560 16725 15569
rect 16683 15520 16684 15560
rect 16724 15520 16725 15560
rect 16683 15511 16725 15520
rect 16771 15560 16829 15561
rect 16771 15520 16780 15560
rect 16820 15520 16829 15560
rect 16771 15519 16829 15520
rect 18595 15560 18653 15561
rect 18595 15520 18604 15560
rect 18644 15520 18653 15560
rect 18595 15519 18653 15520
rect 18699 15560 18741 15569
rect 18699 15520 18700 15560
rect 18740 15520 18741 15560
rect 18699 15511 18741 15520
rect 18891 15560 18933 15569
rect 18891 15520 18892 15560
rect 18932 15520 18933 15560
rect 18891 15511 18933 15520
rect 19267 15560 19325 15561
rect 19267 15520 19276 15560
rect 19316 15520 19325 15560
rect 19267 15519 19325 15520
rect 19747 15560 19805 15561
rect 19747 15520 19756 15560
rect 19796 15520 19805 15560
rect 19747 15519 19805 15520
rect 20043 15560 20085 15569
rect 20043 15520 20044 15560
rect 20084 15520 20085 15560
rect 20043 15511 20085 15520
rect 20139 15560 20181 15569
rect 20139 15520 20140 15560
rect 20180 15520 20181 15560
rect 20139 15511 20181 15520
rect 20235 15560 20277 15569
rect 20235 15520 20236 15560
rect 20276 15520 20277 15560
rect 20235 15511 20277 15520
rect 20715 15560 20757 15569
rect 20715 15520 20716 15560
rect 20756 15520 20757 15560
rect 20715 15511 20757 15520
rect 20811 15560 20853 15569
rect 20811 15520 20812 15560
rect 20852 15520 20853 15560
rect 20811 15511 20853 15520
rect 20907 15560 20949 15569
rect 20907 15520 20908 15560
rect 20948 15520 20949 15560
rect 20907 15511 20949 15520
rect 21483 15560 21525 15569
rect 21483 15520 21484 15560
rect 21524 15520 21525 15560
rect 21483 15511 21525 15520
rect 21867 15560 21909 15569
rect 21867 15520 21868 15560
rect 21908 15520 21909 15560
rect 21571 15518 21629 15519
rect 6699 15476 6741 15485
rect 6699 15436 6700 15476
rect 6740 15436 6741 15476
rect 6699 15427 6741 15436
rect 7947 15476 7989 15485
rect 21571 15478 21580 15518
rect 21620 15478 21629 15518
rect 21867 15511 21909 15520
rect 22059 15560 22101 15569
rect 22059 15520 22060 15560
rect 22100 15520 22101 15560
rect 22059 15511 22101 15520
rect 22243 15560 22301 15561
rect 22243 15520 22252 15560
rect 22292 15520 22301 15560
rect 22243 15519 22301 15520
rect 22443 15560 22485 15569
rect 22443 15520 22444 15560
rect 22484 15520 22485 15560
rect 22443 15511 22485 15520
rect 22531 15560 22589 15561
rect 22531 15520 22540 15560
rect 22580 15520 22589 15560
rect 22531 15519 22589 15520
rect 22731 15560 22773 15569
rect 22731 15520 22732 15560
rect 22772 15520 22773 15560
rect 22731 15511 22773 15520
rect 23107 15560 23165 15561
rect 23107 15520 23116 15560
rect 23156 15520 23165 15560
rect 23107 15519 23165 15520
rect 23779 15560 23837 15561
rect 23779 15520 23788 15560
rect 23828 15520 23837 15560
rect 23779 15519 23837 15520
rect 24067 15560 24125 15561
rect 24067 15520 24076 15560
rect 24116 15520 24125 15560
rect 24067 15519 24125 15520
rect 24267 15560 24309 15569
rect 24267 15520 24268 15560
rect 24308 15520 24309 15560
rect 24267 15511 24309 15520
rect 24739 15560 24797 15561
rect 24739 15520 24748 15560
rect 24788 15520 24797 15560
rect 24739 15519 24797 15520
rect 25131 15560 25173 15569
rect 25131 15520 25132 15560
rect 25172 15520 25173 15560
rect 25131 15511 25173 15520
rect 25315 15560 25373 15561
rect 25315 15520 25324 15560
rect 25364 15520 25373 15560
rect 25315 15519 25373 15520
rect 25419 15560 25461 15569
rect 25419 15520 25420 15560
rect 25460 15520 25461 15560
rect 25419 15511 25461 15520
rect 25603 15560 25661 15561
rect 25603 15520 25612 15560
rect 25652 15520 25661 15560
rect 25603 15519 25661 15520
rect 26091 15560 26133 15569
rect 26091 15520 26092 15560
rect 26132 15520 26133 15560
rect 26091 15511 26133 15520
rect 27627 15560 27669 15569
rect 27627 15520 27628 15560
rect 27668 15520 27669 15560
rect 27627 15511 27669 15520
rect 28011 15560 28053 15569
rect 28011 15520 28012 15560
rect 28052 15520 28053 15560
rect 28011 15511 28053 15520
rect 28107 15560 28149 15569
rect 28107 15520 28108 15560
rect 28148 15520 28149 15560
rect 28107 15511 28149 15520
rect 28203 15560 28245 15569
rect 28203 15520 28204 15560
rect 28244 15520 28245 15560
rect 28203 15511 28245 15520
rect 28387 15560 28445 15561
rect 28387 15520 28396 15560
rect 28436 15520 28445 15560
rect 28387 15519 28445 15520
rect 29259 15560 29301 15569
rect 29259 15520 29260 15560
rect 29300 15520 29301 15560
rect 29259 15511 29301 15520
rect 29355 15560 29397 15569
rect 29355 15520 29356 15560
rect 29396 15520 29397 15560
rect 29355 15511 29397 15520
rect 29451 15560 29493 15569
rect 29451 15520 29452 15560
rect 29492 15520 29493 15560
rect 29451 15511 29493 15520
rect 29547 15560 29589 15569
rect 29547 15520 29548 15560
rect 29588 15520 29589 15560
rect 29547 15511 29589 15520
rect 29739 15560 29781 15569
rect 29739 15520 29740 15560
rect 29780 15520 29781 15560
rect 29739 15511 29781 15520
rect 29931 15560 29973 15569
rect 29931 15520 29932 15560
rect 29972 15520 29973 15560
rect 29931 15511 29973 15520
rect 30027 15560 30069 15569
rect 30027 15520 30028 15560
rect 30068 15520 30069 15560
rect 30027 15511 30069 15520
rect 30595 15560 30653 15561
rect 30595 15520 30604 15560
rect 30644 15520 30653 15560
rect 30595 15519 30653 15520
rect 31555 15560 31613 15561
rect 31555 15520 31564 15560
rect 31604 15520 31613 15560
rect 31555 15519 31613 15520
rect 31651 15560 31709 15561
rect 31651 15520 31660 15560
rect 31700 15520 31709 15560
rect 31651 15519 31709 15520
rect 31851 15560 31893 15569
rect 31851 15520 31852 15560
rect 31892 15520 31893 15560
rect 32040 15560 32098 15561
rect 31851 15511 31893 15520
rect 31939 15531 31997 15532
rect 31939 15491 31948 15531
rect 31988 15491 31997 15531
rect 32040 15520 32049 15560
rect 32089 15520 32098 15560
rect 32040 15519 32098 15520
rect 32414 15560 32472 15561
rect 32414 15520 32423 15560
rect 32463 15520 32472 15560
rect 32414 15519 32472 15520
rect 32523 15560 32565 15569
rect 32523 15520 32524 15560
rect 32564 15520 32565 15560
rect 32523 15511 32565 15520
rect 32619 15560 32661 15569
rect 32619 15520 32620 15560
rect 32660 15520 32661 15560
rect 32619 15511 32661 15520
rect 32803 15560 32861 15561
rect 32803 15520 32812 15560
rect 32852 15520 32861 15560
rect 32803 15519 32861 15520
rect 32899 15560 32957 15561
rect 32899 15520 32908 15560
rect 32948 15520 32957 15560
rect 32899 15519 32957 15520
rect 33675 15560 33717 15569
rect 33675 15520 33676 15560
rect 33716 15520 33717 15560
rect 33675 15511 33717 15520
rect 33763 15560 33821 15561
rect 33763 15520 33772 15560
rect 33812 15520 33821 15560
rect 33763 15519 33821 15520
rect 34339 15560 34397 15561
rect 34339 15520 34348 15560
rect 34388 15520 34397 15560
rect 34339 15519 34397 15520
rect 34435 15560 34493 15561
rect 34435 15520 34444 15560
rect 34484 15520 34493 15560
rect 34435 15519 34493 15520
rect 34819 15560 34877 15561
rect 34819 15520 34828 15560
rect 34868 15520 34877 15560
rect 34819 15519 34877 15520
rect 34923 15560 34965 15569
rect 34923 15520 34924 15560
rect 34964 15520 34965 15560
rect 34923 15511 34965 15520
rect 35019 15560 35061 15569
rect 35019 15520 35020 15560
rect 35060 15520 35061 15560
rect 35019 15511 35061 15520
rect 35403 15560 35445 15569
rect 35403 15520 35404 15560
rect 35444 15520 35445 15560
rect 35403 15511 35445 15520
rect 35595 15560 35637 15569
rect 35595 15520 35596 15560
rect 35636 15520 35637 15560
rect 35595 15511 35637 15520
rect 35883 15560 35925 15569
rect 35883 15520 35884 15560
rect 35924 15520 35925 15560
rect 35883 15511 35925 15520
rect 35979 15560 36021 15569
rect 35979 15520 35980 15560
rect 36020 15520 36021 15560
rect 35979 15511 36021 15520
rect 36075 15560 36117 15569
rect 36075 15520 36076 15560
rect 36116 15520 36117 15560
rect 36363 15560 36405 15569
rect 36075 15511 36117 15520
rect 36259 15541 36317 15542
rect 36259 15501 36268 15541
rect 36308 15501 36317 15541
rect 36363 15520 36364 15560
rect 36404 15520 36405 15560
rect 36363 15511 36405 15520
rect 36555 15560 36597 15569
rect 36555 15520 36556 15560
rect 36596 15520 36597 15560
rect 36555 15511 36597 15520
rect 36739 15560 36797 15561
rect 36739 15520 36748 15560
rect 36788 15520 36797 15560
rect 36739 15519 36797 15520
rect 36843 15560 36885 15569
rect 36843 15520 36844 15560
rect 36884 15520 36885 15560
rect 36843 15511 36885 15520
rect 37515 15560 37557 15569
rect 37515 15520 37516 15560
rect 37556 15520 37557 15560
rect 37515 15511 37557 15520
rect 38091 15560 38133 15569
rect 38091 15520 38092 15560
rect 38132 15520 38133 15560
rect 38091 15511 38133 15520
rect 38179 15560 38237 15561
rect 38179 15520 38188 15560
rect 38228 15520 38237 15560
rect 38179 15519 38237 15520
rect 38659 15560 38717 15561
rect 38659 15520 38668 15560
rect 38708 15520 38717 15560
rect 38659 15519 38717 15520
rect 38859 15560 38901 15569
rect 38859 15520 38860 15560
rect 38900 15520 38901 15560
rect 38859 15511 38901 15520
rect 38947 15560 39005 15561
rect 38947 15520 38956 15560
rect 38996 15520 39005 15560
rect 38947 15519 39005 15520
rect 39523 15560 39581 15561
rect 39523 15520 39532 15560
rect 39572 15520 39581 15560
rect 39523 15519 39581 15520
rect 40395 15560 40437 15569
rect 40395 15520 40396 15560
rect 40436 15520 40437 15560
rect 40395 15511 40437 15520
rect 36259 15500 36317 15501
rect 31939 15490 31997 15491
rect 21571 15477 21629 15478
rect 7947 15436 7948 15476
rect 7988 15436 7989 15476
rect 7947 15427 7989 15436
rect 21963 15476 22005 15485
rect 21963 15436 21964 15476
rect 22004 15436 22005 15476
rect 21963 15427 22005 15436
rect 22827 15476 22869 15485
rect 22827 15436 22828 15476
rect 22868 15436 22869 15476
rect 22827 15427 22869 15436
rect 23019 15476 23061 15485
rect 23019 15436 23020 15476
rect 23060 15436 23061 15476
rect 23019 15427 23061 15436
rect 24843 15476 24885 15485
rect 24843 15436 24844 15476
rect 24884 15436 24885 15476
rect 24843 15427 24885 15436
rect 25035 15476 25077 15485
rect 25035 15436 25036 15476
rect 25076 15436 25077 15476
rect 25035 15427 25077 15436
rect 25899 15476 25941 15485
rect 25899 15436 25900 15476
rect 25940 15436 25941 15476
rect 25899 15427 25941 15436
rect 34627 15476 34685 15477
rect 34627 15436 34636 15476
rect 34676 15436 34685 15476
rect 34627 15435 34685 15436
rect 36939 15476 36981 15485
rect 36939 15436 36940 15476
rect 36980 15436 36981 15476
rect 36939 15427 36981 15436
rect 4587 15392 4629 15401
rect 4587 15352 4588 15392
rect 4628 15352 4629 15392
rect 4587 15343 4629 15352
rect 6795 15392 6837 15401
rect 6795 15352 6796 15392
rect 6836 15352 6837 15392
rect 6795 15343 6837 15352
rect 6891 15392 6933 15401
rect 6891 15352 6892 15392
rect 6932 15352 6933 15392
rect 6891 15343 6933 15352
rect 8803 15392 8861 15393
rect 8803 15352 8812 15392
rect 8852 15352 8861 15392
rect 8803 15351 8861 15352
rect 22923 15392 22965 15401
rect 22923 15352 22924 15392
rect 22964 15352 22965 15392
rect 22923 15343 22965 15352
rect 24171 15392 24213 15401
rect 24171 15352 24172 15392
rect 24212 15352 24213 15392
rect 24171 15343 24213 15352
rect 24939 15392 24981 15401
rect 24939 15352 24940 15392
rect 24980 15352 24981 15392
rect 24939 15343 24981 15352
rect 27627 15392 27669 15401
rect 27627 15352 27628 15392
rect 27668 15352 27669 15392
rect 27627 15343 27669 15352
rect 29835 15392 29877 15401
rect 29835 15352 29836 15392
rect 29876 15352 29877 15392
rect 29835 15343 29877 15352
rect 33387 15392 33429 15401
rect 33387 15352 33388 15392
rect 33428 15352 33429 15392
rect 33387 15343 33429 15352
rect 35595 15392 35637 15401
rect 35595 15352 35596 15392
rect 35636 15352 35637 15392
rect 35595 15343 35637 15352
rect 37035 15392 37077 15401
rect 37035 15352 37036 15392
rect 37076 15352 37077 15392
rect 37035 15343 37077 15352
rect 37515 15392 37557 15401
rect 37515 15352 37516 15392
rect 37556 15352 37557 15392
rect 37515 15343 37557 15352
rect 37707 15392 37749 15401
rect 37707 15352 37708 15392
rect 37748 15352 37749 15392
rect 37707 15343 37749 15352
rect 39147 15392 39189 15401
rect 39147 15352 39148 15392
rect 39188 15352 39189 15392
rect 39147 15343 39189 15352
rect 3339 15308 3381 15317
rect 3339 15268 3340 15308
rect 3380 15268 3381 15308
rect 3339 15259 3381 15268
rect 3811 15308 3869 15309
rect 3811 15268 3820 15308
rect 3860 15268 3869 15308
rect 3811 15267 3869 15268
rect 5443 15308 5501 15309
rect 5443 15268 5452 15308
rect 5492 15268 5501 15308
rect 5443 15267 5501 15268
rect 5635 15308 5693 15309
rect 5635 15268 5644 15308
rect 5684 15268 5693 15308
rect 5635 15267 5693 15268
rect 7179 15308 7221 15317
rect 7179 15268 7180 15308
rect 7220 15268 7221 15308
rect 7179 15259 7221 15268
rect 9003 15308 9045 15317
rect 9003 15268 9004 15308
rect 9044 15268 9045 15308
rect 9003 15259 9045 15268
rect 15619 15308 15677 15309
rect 15619 15268 15628 15308
rect 15668 15268 15677 15308
rect 15619 15267 15677 15268
rect 16971 15308 17013 15317
rect 16971 15268 16972 15308
rect 17012 15268 17013 15308
rect 16971 15259 17013 15268
rect 18891 15308 18933 15317
rect 18891 15268 18892 15308
rect 18932 15268 18933 15308
rect 18891 15259 18933 15268
rect 21195 15308 21237 15317
rect 21195 15268 21196 15308
rect 21236 15268 21237 15308
rect 21195 15259 21237 15268
rect 22251 15308 22293 15317
rect 22251 15268 22252 15308
rect 22292 15268 22293 15308
rect 22251 15259 22293 15268
rect 29059 15308 29117 15309
rect 29059 15268 29068 15308
rect 29108 15268 29117 15308
rect 29059 15267 29117 15268
rect 31563 15308 31605 15317
rect 31563 15268 31564 15308
rect 31604 15268 31605 15308
rect 31563 15259 31605 15268
rect 34539 15308 34581 15317
rect 34539 15268 34540 15308
rect 34580 15268 34581 15308
rect 34539 15259 34581 15268
rect 36555 15308 36597 15317
rect 36555 15268 36556 15308
rect 36596 15268 36597 15308
rect 36555 15259 36597 15268
rect 38379 15308 38421 15317
rect 38379 15268 38380 15308
rect 38420 15268 38421 15308
rect 38379 15259 38421 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 4675 14972 4733 14973
rect 4675 14932 4684 14972
rect 4724 14932 4733 14972
rect 4675 14931 4733 14932
rect 7075 14972 7133 14973
rect 7075 14932 7084 14972
rect 7124 14932 7133 14972
rect 7075 14931 7133 14932
rect 9099 14972 9141 14981
rect 9099 14932 9100 14972
rect 9140 14932 9141 14972
rect 9099 14923 9141 14932
rect 9283 14972 9341 14973
rect 9283 14932 9292 14972
rect 9332 14932 9341 14972
rect 9283 14931 9341 14932
rect 16011 14972 16053 14981
rect 16011 14932 16012 14972
rect 16052 14932 16053 14972
rect 16011 14923 16053 14932
rect 17547 14972 17589 14981
rect 17547 14932 17548 14972
rect 17588 14932 17589 14972
rect 17547 14923 17589 14932
rect 20139 14972 20181 14981
rect 20139 14932 20140 14972
rect 20180 14932 20181 14972
rect 20139 14923 20181 14932
rect 35691 14972 35733 14981
rect 35691 14932 35692 14972
rect 35732 14932 35733 14972
rect 35691 14923 35733 14932
rect 36075 14972 36117 14981
rect 36075 14932 36076 14972
rect 36116 14932 36117 14972
rect 36075 14923 36117 14932
rect 37131 14972 37173 14981
rect 37131 14932 37132 14972
rect 37172 14932 37173 14972
rect 37131 14923 37173 14932
rect 41547 14972 41589 14981
rect 41547 14932 41548 14972
rect 41588 14932 41589 14972
rect 41547 14923 41589 14932
rect 1515 14888 1557 14897
rect 1515 14848 1516 14888
rect 1556 14848 1557 14888
rect 1515 14839 1557 14848
rect 3435 14888 3477 14897
rect 3435 14848 3436 14888
rect 3476 14848 3477 14888
rect 3435 14839 3477 14848
rect 6595 14888 6653 14889
rect 6595 14848 6604 14888
rect 6644 14848 6653 14888
rect 6595 14847 6653 14848
rect 10155 14888 10197 14897
rect 10155 14848 10156 14888
rect 10196 14848 10197 14888
rect 10155 14839 10197 14848
rect 32331 14888 32373 14897
rect 32331 14848 32332 14888
rect 32372 14848 32373 14888
rect 32331 14839 32373 14848
rect 37603 14804 37661 14805
rect 37603 14764 37612 14804
rect 37652 14764 37661 14804
rect 37603 14763 37661 14764
rect 3723 14751 3765 14760
rect 2955 14720 2997 14729
rect 2955 14680 2956 14720
rect 2996 14680 2997 14720
rect 2955 14671 2997 14680
rect 3051 14720 3093 14729
rect 3051 14680 3052 14720
rect 3092 14680 3093 14720
rect 3051 14671 3093 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3627 14720 3669 14729
rect 3627 14680 3628 14720
rect 3668 14680 3669 14720
rect 3723 14711 3724 14751
rect 3764 14711 3765 14751
rect 3723 14702 3765 14711
rect 4203 14720 4245 14729
rect 3627 14671 3669 14680
rect 4203 14680 4204 14720
rect 4244 14680 4245 14720
rect 4203 14671 4245 14680
rect 4299 14720 4341 14729
rect 4299 14680 4300 14720
rect 4340 14680 4341 14720
rect 4299 14671 4341 14680
rect 4395 14720 4437 14729
rect 4395 14680 4396 14720
rect 4436 14680 4437 14720
rect 4395 14671 4437 14680
rect 4491 14720 4533 14729
rect 4491 14680 4492 14720
rect 4532 14680 4533 14720
rect 4491 14671 4533 14680
rect 5539 14720 5597 14721
rect 5539 14680 5548 14720
rect 5588 14680 5597 14720
rect 5539 14679 5597 14680
rect 6403 14720 6461 14721
rect 6403 14680 6412 14720
rect 6452 14680 6461 14720
rect 6403 14679 6461 14680
rect 6603 14720 6645 14729
rect 6603 14680 6604 14720
rect 6644 14680 6645 14720
rect 6603 14671 6645 14680
rect 6699 14720 6741 14729
rect 6699 14680 6700 14720
rect 6740 14680 6741 14720
rect 6699 14671 6741 14680
rect 6891 14720 6933 14729
rect 6891 14680 6892 14720
rect 6932 14680 6933 14720
rect 6891 14671 6933 14680
rect 7747 14720 7805 14721
rect 7747 14680 7756 14720
rect 7796 14680 7805 14720
rect 7747 14679 7805 14680
rect 7939 14720 7997 14721
rect 7939 14680 7948 14720
rect 7988 14680 7997 14720
rect 7939 14679 7997 14680
rect 8043 14720 8085 14729
rect 8043 14680 8044 14720
rect 8084 14680 8085 14720
rect 8043 14671 8085 14680
rect 8235 14720 8277 14729
rect 8235 14680 8236 14720
rect 8276 14680 8277 14720
rect 8235 14671 8277 14680
rect 8803 14720 8861 14721
rect 8803 14680 8812 14720
rect 8852 14680 8861 14720
rect 8803 14679 8861 14680
rect 8907 14720 8949 14729
rect 8907 14680 8908 14720
rect 8948 14680 8949 14720
rect 8907 14671 8949 14680
rect 9099 14720 9141 14729
rect 9099 14680 9100 14720
rect 9140 14680 9141 14720
rect 9099 14671 9141 14680
rect 9955 14720 10013 14721
rect 9955 14680 9964 14720
rect 10004 14680 10013 14720
rect 9955 14679 10013 14680
rect 11403 14720 11445 14729
rect 11403 14680 11404 14720
rect 11444 14680 11445 14720
rect 11403 14671 11445 14680
rect 13803 14720 13845 14729
rect 13803 14680 13804 14720
rect 13844 14680 13845 14720
rect 13803 14671 13845 14680
rect 13899 14720 13941 14729
rect 13899 14680 13900 14720
rect 13940 14680 13941 14720
rect 13899 14671 13941 14680
rect 13995 14720 14037 14729
rect 13995 14680 13996 14720
rect 14036 14680 14037 14720
rect 13995 14671 14037 14680
rect 14371 14720 14429 14721
rect 14371 14680 14380 14720
rect 14420 14680 14429 14720
rect 14371 14679 14429 14680
rect 14571 14720 14613 14729
rect 14571 14680 14572 14720
rect 14612 14680 14613 14720
rect 14571 14671 14613 14680
rect 15043 14720 15101 14721
rect 15043 14680 15052 14720
rect 15092 14680 15101 14720
rect 15043 14679 15101 14680
rect 15139 14720 15197 14721
rect 15139 14680 15148 14720
rect 15188 14680 15197 14720
rect 15139 14679 15197 14680
rect 15811 14720 15869 14721
rect 15811 14680 15820 14720
rect 15860 14680 15869 14720
rect 15811 14679 15869 14680
rect 15907 14720 15965 14721
rect 15907 14680 15916 14720
rect 15956 14680 15965 14720
rect 15907 14679 15965 14680
rect 17163 14720 17205 14729
rect 17163 14680 17164 14720
rect 17204 14680 17205 14720
rect 17163 14671 17205 14680
rect 17539 14720 17597 14721
rect 17539 14680 17548 14720
rect 17588 14680 17597 14720
rect 17539 14679 17597 14680
rect 17635 14720 17693 14721
rect 17635 14680 17644 14720
rect 17684 14680 17693 14720
rect 17635 14679 17693 14680
rect 17835 14720 17877 14729
rect 17835 14680 17836 14720
rect 17876 14680 17877 14720
rect 17835 14671 17877 14680
rect 17931 14720 17973 14729
rect 17931 14680 17932 14720
rect 17972 14680 17973 14720
rect 17931 14671 17973 14680
rect 18024 14720 18082 14721
rect 18024 14680 18033 14720
rect 18073 14680 18082 14720
rect 18024 14679 18082 14680
rect 18315 14720 18357 14729
rect 18315 14680 18316 14720
rect 18356 14680 18357 14720
rect 18315 14671 18357 14680
rect 18411 14720 18453 14729
rect 18411 14680 18412 14720
rect 18452 14680 18453 14720
rect 18411 14671 18453 14680
rect 18507 14720 18549 14729
rect 18507 14680 18508 14720
rect 18548 14680 18549 14720
rect 18507 14671 18549 14680
rect 18603 14720 18645 14729
rect 18603 14680 18604 14720
rect 18644 14680 18645 14720
rect 18603 14671 18645 14680
rect 19843 14720 19901 14721
rect 19843 14680 19852 14720
rect 19892 14680 19901 14720
rect 19843 14679 19901 14680
rect 19947 14720 19989 14729
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 20331 14720 20373 14729
rect 19947 14671 19989 14680
rect 20139 14678 20181 14687
rect 14475 14636 14517 14645
rect 20139 14638 20140 14678
rect 20180 14638 20181 14678
rect 20331 14680 20332 14720
rect 20372 14680 20373 14720
rect 20331 14671 20373 14680
rect 20619 14720 20661 14729
rect 20619 14680 20620 14720
rect 20660 14680 20661 14720
rect 20619 14671 20661 14680
rect 20803 14720 20861 14721
rect 20803 14680 20812 14720
rect 20852 14680 20861 14720
rect 20803 14679 20861 14680
rect 21675 14720 21717 14729
rect 21675 14680 21676 14720
rect 21716 14680 21717 14720
rect 21675 14671 21717 14680
rect 22051 14720 22109 14721
rect 22051 14680 22060 14720
rect 22100 14680 22109 14720
rect 22051 14679 22109 14680
rect 22923 14720 22965 14729
rect 22923 14680 22924 14720
rect 22964 14680 22965 14720
rect 22923 14671 22965 14680
rect 23299 14720 23357 14721
rect 23299 14680 23308 14720
rect 23348 14680 23357 14720
rect 23299 14679 23357 14680
rect 24259 14720 24317 14721
rect 24259 14680 24268 14720
rect 24308 14680 24317 14720
rect 24259 14679 24317 14680
rect 24747 14720 24789 14729
rect 24747 14680 24748 14720
rect 24788 14680 24789 14720
rect 24747 14671 24789 14680
rect 25603 14720 25661 14721
rect 25603 14680 25612 14720
rect 25652 14680 25661 14720
rect 25603 14679 25661 14680
rect 25987 14720 26045 14721
rect 25987 14680 25996 14720
rect 26036 14680 26045 14720
rect 25987 14679 26045 14680
rect 26379 14720 26421 14729
rect 26379 14680 26380 14720
rect 26420 14680 26421 14720
rect 26379 14671 26421 14680
rect 26571 14720 26613 14729
rect 26571 14680 26572 14720
rect 26612 14680 26613 14720
rect 26571 14671 26613 14680
rect 26859 14720 26901 14729
rect 26859 14680 26860 14720
rect 26900 14680 26901 14720
rect 26859 14671 26901 14680
rect 28107 14720 28149 14729
rect 28107 14680 28108 14720
rect 28148 14680 28149 14720
rect 28107 14671 28149 14680
rect 28299 14720 28341 14729
rect 28299 14680 28300 14720
rect 28340 14680 28341 14720
rect 28299 14671 28341 14680
rect 28483 14720 28541 14721
rect 28483 14680 28492 14720
rect 28532 14680 28541 14720
rect 28483 14679 28541 14680
rect 28587 14720 28629 14729
rect 28587 14680 28588 14720
rect 28628 14680 28629 14720
rect 28587 14671 28629 14680
rect 28779 14720 28821 14729
rect 28779 14680 28780 14720
rect 28820 14680 28821 14720
rect 28779 14671 28821 14680
rect 29059 14720 29117 14721
rect 29059 14680 29068 14720
rect 29108 14680 29117 14720
rect 29059 14679 29117 14680
rect 29355 14720 29397 14729
rect 29355 14680 29356 14720
rect 29396 14680 29397 14720
rect 29355 14671 29397 14680
rect 29547 14720 29589 14729
rect 29547 14680 29548 14720
rect 29588 14680 29589 14720
rect 29547 14671 29589 14680
rect 29635 14720 29693 14721
rect 29635 14680 29644 14720
rect 29684 14680 29693 14720
rect 29635 14679 29693 14680
rect 30115 14720 30173 14721
rect 30115 14680 30124 14720
rect 30164 14680 30173 14720
rect 30115 14679 30173 14680
rect 31371 14720 31413 14729
rect 31371 14680 31372 14720
rect 31412 14680 31413 14720
rect 31371 14671 31413 14680
rect 31467 14720 31509 14729
rect 31467 14680 31468 14720
rect 31508 14680 31509 14720
rect 31467 14671 31509 14680
rect 31563 14720 31605 14729
rect 31563 14680 31564 14720
rect 31604 14680 31605 14720
rect 31563 14671 31605 14680
rect 31659 14720 31701 14729
rect 31659 14680 31660 14720
rect 31700 14680 31701 14720
rect 31659 14671 31701 14680
rect 31843 14720 31901 14721
rect 31843 14680 31852 14720
rect 31892 14680 31901 14720
rect 32139 14720 32181 14729
rect 31843 14679 31901 14680
rect 31947 14706 31989 14715
rect 31947 14666 31948 14706
rect 31988 14666 31989 14706
rect 32139 14680 32140 14720
rect 32180 14680 32181 14720
rect 32139 14671 32181 14680
rect 32323 14720 32381 14721
rect 32323 14680 32332 14720
rect 32372 14680 32381 14720
rect 32323 14679 32381 14680
rect 32523 14720 32565 14729
rect 32523 14680 32524 14720
rect 32564 14680 32565 14720
rect 32523 14671 32565 14680
rect 32611 14720 32669 14721
rect 32611 14680 32620 14720
rect 32660 14680 32669 14720
rect 32611 14679 32669 14680
rect 33003 14720 33045 14729
rect 33003 14680 33004 14720
rect 33044 14680 33045 14720
rect 33003 14671 33045 14680
rect 33099 14720 33141 14729
rect 33099 14680 33100 14720
rect 33140 14680 33141 14720
rect 33099 14671 33141 14680
rect 33283 14720 33341 14721
rect 33283 14680 33292 14720
rect 33332 14680 33341 14720
rect 33283 14679 33341 14680
rect 34347 14720 34389 14729
rect 34347 14680 34348 14720
rect 34388 14680 34389 14720
rect 34347 14671 34389 14680
rect 34443 14720 34485 14729
rect 34443 14680 34444 14720
rect 34484 14680 34485 14720
rect 34443 14671 34485 14680
rect 35779 14720 35837 14721
rect 35779 14680 35788 14720
rect 35828 14680 35837 14720
rect 35779 14679 35837 14680
rect 36259 14720 36317 14721
rect 36259 14680 36268 14720
rect 36308 14680 36317 14720
rect 36259 14679 36317 14680
rect 36363 14720 36405 14729
rect 36363 14680 36364 14720
rect 36404 14680 36405 14720
rect 37323 14720 37365 14729
rect 36363 14671 36405 14680
rect 37131 14706 37173 14715
rect 31947 14657 31989 14666
rect 37131 14666 37132 14706
rect 37172 14666 37173 14706
rect 37323 14680 37324 14720
rect 37364 14680 37365 14720
rect 37323 14671 37365 14680
rect 37411 14720 37469 14721
rect 37411 14680 37420 14720
rect 37460 14680 37469 14720
rect 37411 14679 37469 14680
rect 37891 14720 37949 14721
rect 37891 14680 37900 14720
rect 37940 14680 37949 14720
rect 37891 14679 37949 14680
rect 37995 14720 38037 14729
rect 37995 14680 37996 14720
rect 38036 14680 38037 14720
rect 37995 14671 38037 14680
rect 38667 14720 38709 14729
rect 38667 14680 38668 14720
rect 38708 14680 38709 14720
rect 38667 14671 38709 14680
rect 38851 14720 38909 14721
rect 38851 14680 38860 14720
rect 38900 14680 38909 14720
rect 38851 14679 38909 14680
rect 39147 14720 39189 14729
rect 39147 14680 39148 14720
rect 39188 14680 39189 14720
rect 39147 14671 39189 14680
rect 39523 14720 39581 14721
rect 39523 14680 39532 14720
rect 39572 14680 39581 14720
rect 39523 14679 39581 14680
rect 40387 14720 40445 14721
rect 40387 14680 40396 14720
rect 40436 14680 40445 14720
rect 40387 14679 40445 14680
rect 37131 14657 37173 14666
rect 14475 14596 14476 14636
rect 14516 14596 14517 14636
rect 14475 14587 14517 14596
rect 16387 14636 16445 14637
rect 16387 14596 16396 14636
rect 16436 14596 16445 14636
rect 20139 14629 20181 14638
rect 25899 14636 25941 14645
rect 16387 14595 16445 14596
rect 25899 14596 25900 14636
rect 25940 14596 25941 14636
rect 25899 14587 25941 14596
rect 28683 14636 28725 14645
rect 28683 14596 28684 14636
rect 28724 14596 28725 14636
rect 28683 14587 28725 14596
rect 29451 14636 29493 14645
rect 29451 14596 29452 14636
rect 29492 14596 29493 14636
rect 29451 14587 29493 14596
rect 30307 14636 30365 14637
rect 30307 14596 30316 14636
rect 30356 14596 30365 14636
rect 30307 14595 30365 14596
rect 38763 14636 38805 14645
rect 38763 14596 38764 14636
rect 38804 14596 38805 14636
rect 38763 14587 38805 14596
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 1027 14552 1085 14553
rect 1027 14512 1036 14552
rect 1076 14512 1085 14552
rect 1027 14511 1085 14512
rect 3147 14552 3189 14561
rect 3147 14512 3148 14552
rect 3188 14512 3189 14552
rect 3147 14503 3189 14512
rect 3715 14552 3773 14553
rect 3715 14512 3724 14552
rect 3764 14512 3773 14552
rect 3715 14511 3773 14512
rect 4867 14552 4925 14553
rect 4867 14512 4876 14552
rect 4916 14512 4925 14552
rect 4867 14511 4925 14512
rect 5731 14552 5789 14553
rect 5731 14512 5740 14552
rect 5780 14512 5789 14552
rect 5731 14511 5789 14512
rect 8131 14552 8189 14553
rect 8131 14512 8140 14552
rect 8180 14512 8189 14552
rect 8131 14511 8189 14512
rect 11787 14552 11829 14561
rect 11787 14512 11788 14552
rect 11828 14512 11829 14552
rect 11787 14503 11829 14512
rect 13699 14552 13757 14553
rect 13699 14512 13708 14552
rect 13748 14512 13757 14552
rect 13699 14511 13757 14512
rect 15339 14552 15381 14561
rect 15339 14512 15340 14552
rect 15380 14512 15381 14552
rect 15339 14503 15381 14512
rect 20523 14552 20565 14561
rect 20523 14512 20524 14552
rect 20564 14512 20565 14552
rect 20523 14503 20565 14512
rect 25131 14552 25173 14561
rect 25131 14512 25132 14552
rect 25172 14512 25173 14552
rect 25131 14503 25173 14512
rect 26667 14552 26709 14561
rect 26667 14512 26668 14552
rect 26708 14512 26709 14552
rect 26667 14503 26709 14512
rect 28203 14552 28245 14561
rect 28203 14512 28204 14552
rect 28244 14512 28245 14552
rect 28203 14503 28245 14512
rect 28971 14552 29013 14561
rect 28971 14512 28972 14552
rect 29012 14512 29013 14552
rect 28971 14503 29013 14512
rect 30019 14552 30077 14553
rect 30019 14512 30028 14552
rect 30068 14512 30077 14552
rect 30019 14511 30077 14512
rect 32035 14552 32093 14553
rect 32035 14512 32044 14552
rect 32084 14512 32093 14552
rect 32035 14511 32093 14512
rect 32803 14552 32861 14553
rect 32803 14512 32812 14552
rect 32852 14512 32861 14552
rect 32803 14511 32861 14512
rect 33955 14552 34013 14553
rect 33955 14512 33964 14552
rect 34004 14512 34013 14552
rect 33955 14511 34013 14512
rect 34147 14552 34205 14553
rect 34147 14512 34156 14552
rect 34196 14512 34205 14552
rect 34147 14511 34205 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 4771 14216 4829 14217
rect 4771 14176 4780 14216
rect 4820 14176 4829 14216
rect 4771 14175 4829 14176
rect 8035 14216 8093 14217
rect 8035 14176 8044 14216
rect 8084 14176 8093 14216
rect 8035 14175 8093 14176
rect 8707 14216 8765 14217
rect 8707 14176 8716 14216
rect 8756 14176 8765 14216
rect 8707 14175 8765 14176
rect 15811 14216 15869 14217
rect 15811 14176 15820 14216
rect 15860 14176 15869 14216
rect 15811 14175 15869 14176
rect 19851 14216 19893 14225
rect 19851 14176 19852 14216
rect 19892 14176 19893 14216
rect 19851 14167 19893 14176
rect 25891 14216 25949 14217
rect 25891 14176 25900 14216
rect 25940 14176 25949 14216
rect 25891 14175 25949 14176
rect 27043 14216 27101 14217
rect 27043 14176 27052 14216
rect 27092 14176 27101 14216
rect 27043 14175 27101 14176
rect 27235 14216 27293 14217
rect 27235 14176 27244 14216
rect 27284 14176 27293 14216
rect 27235 14175 27293 14176
rect 28587 14216 28629 14225
rect 28587 14176 28588 14216
rect 28628 14176 28629 14216
rect 28587 14167 28629 14176
rect 29923 14216 29981 14217
rect 29923 14176 29932 14216
rect 29972 14176 29981 14216
rect 29923 14175 29981 14176
rect 33667 14216 33725 14217
rect 33667 14176 33676 14216
rect 33716 14176 33725 14216
rect 33667 14175 33725 14176
rect 35115 14216 35157 14225
rect 35115 14176 35116 14216
rect 35156 14176 35157 14216
rect 35115 14167 35157 14176
rect 38947 14216 39005 14217
rect 38947 14176 38956 14216
rect 38996 14176 39005 14216
rect 38947 14175 39005 14176
rect 5643 14132 5685 14141
rect 5643 14092 5644 14132
rect 5684 14092 5685 14132
rect 5643 14083 5685 14092
rect 9579 14132 9621 14141
rect 9579 14092 9580 14132
rect 9620 14092 9621 14132
rect 9579 14083 9621 14092
rect 13035 14132 13077 14141
rect 13035 14092 13036 14132
rect 13076 14092 13077 14132
rect 13035 14083 13077 14092
rect 17835 14132 17877 14141
rect 17835 14092 17836 14132
rect 17876 14092 17877 14132
rect 17835 14083 17877 14092
rect 20515 14132 20573 14133
rect 20515 14092 20524 14132
rect 20564 14092 20573 14132
rect 20515 14091 20573 14092
rect 21867 14132 21909 14141
rect 21867 14092 21868 14132
rect 21908 14092 21909 14132
rect 21867 14083 21909 14092
rect 29827 14132 29885 14133
rect 29827 14092 29836 14132
rect 29876 14092 29885 14132
rect 29827 14091 29885 14092
rect 1035 14048 1077 14057
rect 1035 14008 1036 14048
rect 1076 14008 1077 14048
rect 1035 13999 1077 14008
rect 1411 14048 1469 14049
rect 1411 14008 1420 14048
rect 1460 14008 1469 14048
rect 1411 14007 1469 14008
rect 2275 14048 2333 14049
rect 2275 14008 2284 14048
rect 2324 14008 2333 14048
rect 2275 14007 2333 14008
rect 3523 14048 3581 14049
rect 3523 14008 3532 14048
rect 3572 14008 3581 14048
rect 3523 14007 3581 14008
rect 4579 14048 4637 14049
rect 4579 14008 4588 14048
rect 4628 14008 4637 14048
rect 4579 14007 4637 14008
rect 5443 14048 5501 14049
rect 5443 14008 5452 14048
rect 5492 14008 5501 14048
rect 5443 14007 5501 14008
rect 6019 14048 6077 14049
rect 6019 14008 6028 14048
rect 6068 14008 6077 14048
rect 6019 14007 6077 14008
rect 6883 14048 6941 14049
rect 6883 14008 6892 14048
rect 6932 14008 6941 14048
rect 6883 14007 6941 14008
rect 9379 14048 9437 14049
rect 9379 14008 9388 14048
rect 9428 14008 9437 14048
rect 9379 14007 9437 14008
rect 9955 14048 10013 14049
rect 9955 14008 9964 14048
rect 10004 14008 10013 14048
rect 9955 14007 10013 14008
rect 10819 14048 10877 14049
rect 10819 14008 10828 14048
rect 10868 14008 10877 14048
rect 10819 14007 10877 14008
rect 12835 14048 12893 14049
rect 12835 14008 12844 14048
rect 12884 14008 12893 14048
rect 12835 14007 12893 14008
rect 13699 14048 13757 14049
rect 13699 14008 13708 14048
rect 13748 14008 13757 14048
rect 13699 14007 13757 14008
rect 14083 14048 14141 14049
rect 14083 14008 14092 14048
rect 14132 14008 14141 14048
rect 14083 14007 14141 14008
rect 14179 14048 14237 14049
rect 14179 14008 14188 14048
rect 14228 14008 14237 14048
rect 14179 14007 14237 14008
rect 14659 14048 14717 14049
rect 14659 14008 14668 14048
rect 14708 14008 14717 14048
rect 14659 14007 14717 14008
rect 14763 14048 14805 14057
rect 14763 14008 14764 14048
rect 14804 14008 14805 14048
rect 14763 13999 14805 14008
rect 14947 14048 15005 14049
rect 14947 14008 14956 14048
rect 14996 14008 15005 14048
rect 14947 14007 15005 14008
rect 15139 14048 15197 14049
rect 15139 14008 15148 14048
rect 15188 14008 15197 14048
rect 15139 14007 15197 14008
rect 15339 14048 15381 14057
rect 15339 14008 15340 14048
rect 15380 14008 15381 14048
rect 15339 13999 15381 14008
rect 15531 14048 15573 14057
rect 15531 14008 15532 14048
rect 15572 14008 15573 14048
rect 15531 13999 15573 14008
rect 15627 14048 15669 14057
rect 15627 14008 15628 14048
rect 15668 14008 15669 14048
rect 15627 13999 15669 14008
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 16875 14048 16917 14057
rect 16875 14008 16876 14048
rect 16916 14008 16917 14048
rect 16875 13999 16917 14008
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17355 14048 17397 14057
rect 17355 14008 17356 14048
rect 17396 14008 17397 14048
rect 17355 13999 17397 14008
rect 17451 14048 17493 14057
rect 17451 14008 17452 14048
rect 17492 14008 17493 14048
rect 17451 13999 17493 14008
rect 17547 14048 17589 14057
rect 17547 14008 17548 14048
rect 17588 14008 17589 14048
rect 17547 13999 17589 14008
rect 17739 14048 17781 14057
rect 17739 14008 17740 14048
rect 17780 14008 17781 14048
rect 17739 13999 17781 14008
rect 17923 14048 17981 14049
rect 17923 14008 17932 14048
rect 17972 14008 17981 14048
rect 17923 14007 17981 14008
rect 18795 14048 18837 14057
rect 18795 14008 18796 14048
rect 18836 14008 18837 14048
rect 18795 13999 18837 14008
rect 18891 14048 18933 14057
rect 18891 14008 18892 14048
rect 18932 14008 18933 14048
rect 18891 13999 18933 14008
rect 18987 14048 19029 14057
rect 18987 14008 18988 14048
rect 19028 14008 19029 14048
rect 18987 13999 19029 14008
rect 19083 14048 19125 14057
rect 19083 14008 19084 14048
rect 19124 14008 19125 14048
rect 19083 13999 19125 14008
rect 19467 14048 19509 14057
rect 19467 14008 19468 14048
rect 19508 14008 19509 14048
rect 19467 13999 19509 14008
rect 19555 14048 19613 14049
rect 19555 14008 19564 14048
rect 19604 14008 19613 14048
rect 19555 14007 19613 14008
rect 20035 14048 20093 14049
rect 20035 14008 20044 14048
rect 20084 14008 20093 14048
rect 20035 14007 20093 14008
rect 20419 14048 20477 14049
rect 20419 14008 20428 14048
rect 20468 14008 20477 14048
rect 20419 14007 20477 14008
rect 20995 14048 21053 14049
rect 20995 14008 21004 14048
rect 21044 14008 21053 14048
rect 20995 14007 21053 14008
rect 21099 14048 21141 14057
rect 21099 14008 21100 14048
rect 21140 14008 21141 14048
rect 21099 13999 21141 14008
rect 21291 14048 21333 14057
rect 21291 14008 21292 14048
rect 21332 14008 21333 14048
rect 21291 13999 21333 14008
rect 21579 14048 21621 14057
rect 21579 14008 21580 14048
rect 21620 14008 21621 14048
rect 21579 13999 21621 14008
rect 21675 14048 21717 14057
rect 21675 14008 21676 14048
rect 21716 14008 21717 14048
rect 21675 13999 21717 14008
rect 21771 14048 21813 14057
rect 21771 14008 21772 14048
rect 21812 14008 21813 14048
rect 21771 13999 21813 14008
rect 23011 14048 23069 14049
rect 23011 14008 23020 14048
rect 23060 14008 23069 14048
rect 23011 14007 23069 14008
rect 25411 14048 25469 14049
rect 25411 14008 25420 14048
rect 25460 14008 25469 14048
rect 25411 14007 25469 14008
rect 25515 14048 25557 14057
rect 25515 14008 25516 14048
rect 25556 14008 25557 14048
rect 25515 13999 25557 14008
rect 25707 14048 25749 14057
rect 25707 14008 25708 14048
rect 25748 14008 25749 14048
rect 25707 13999 25749 14008
rect 26091 14048 26133 14057
rect 26091 14008 26092 14048
rect 26132 14008 26133 14048
rect 26091 13999 26133 14008
rect 26187 14048 26229 14057
rect 26187 14008 26188 14048
rect 26228 14008 26229 14048
rect 26187 13999 26229 14008
rect 26763 14048 26805 14057
rect 26763 14008 26764 14048
rect 26804 14008 26805 14048
rect 26763 13999 26805 14008
rect 26859 14048 26901 14057
rect 26859 14008 26860 14048
rect 26900 14008 26901 14048
rect 26859 13999 26901 14008
rect 27435 14048 27477 14057
rect 27435 14008 27436 14048
rect 27476 14008 27477 14048
rect 27435 13999 27477 14008
rect 27531 14048 27573 14057
rect 27531 14008 27532 14048
rect 27572 14008 27573 14048
rect 27531 13999 27573 14008
rect 27627 14048 27669 14057
rect 27627 14008 27628 14048
rect 27668 14008 27669 14048
rect 27627 13999 27669 14008
rect 27723 14048 27765 14057
rect 27723 14008 27724 14048
rect 27764 14008 27765 14048
rect 27723 13999 27765 14008
rect 28203 14048 28245 14057
rect 28203 14008 28204 14048
rect 28244 14008 28245 14048
rect 28203 13999 28245 14008
rect 28291 14048 28349 14049
rect 28291 14008 28300 14048
rect 28340 14008 28349 14048
rect 28291 14007 28349 14008
rect 29059 14048 29117 14049
rect 29059 14008 29068 14048
rect 29108 14008 29117 14048
rect 29059 14007 29117 14008
rect 29155 14048 29213 14049
rect 29155 14008 29164 14048
rect 29204 14008 29213 14048
rect 29155 14007 29213 14008
rect 29643 14048 29685 14057
rect 29643 14008 29644 14048
rect 29684 14008 29685 14048
rect 29643 13999 29685 14008
rect 29739 14048 29781 14057
rect 29739 14008 29740 14048
rect 29780 14008 29781 14048
rect 29739 13999 29781 14008
rect 31947 14048 31989 14057
rect 31947 14008 31948 14048
rect 31988 14008 31989 14048
rect 31947 13999 31989 14008
rect 34339 14048 34397 14049
rect 34339 14008 34348 14048
rect 34388 14008 34397 14048
rect 34339 14007 34397 14008
rect 34627 14048 34685 14049
rect 34627 14008 34636 14048
rect 34676 14008 34685 14048
rect 34627 14007 34685 14008
rect 36835 14048 36893 14049
rect 36835 14008 36844 14048
rect 36884 14008 36893 14048
rect 36835 14007 36893 14008
rect 37795 14048 37853 14049
rect 37795 14008 37804 14048
rect 37844 14008 37853 14048
rect 37795 14007 37853 14008
rect 38755 14048 38813 14049
rect 38755 14008 38764 14048
rect 38804 14008 38813 14048
rect 38755 14007 38813 14008
rect 39147 14048 39189 14057
rect 39147 14008 39148 14048
rect 39188 14008 39189 14048
rect 39147 13999 39189 14008
rect 39243 14048 39285 14057
rect 39243 14008 39244 14048
rect 39284 14008 39285 14048
rect 39243 13999 39285 14008
rect 39819 14048 39861 14057
rect 39819 14008 39820 14048
rect 39860 14008 39861 14048
rect 39819 13999 39861 14008
rect 40483 14048 40541 14049
rect 40483 14008 40492 14048
rect 40532 14008 40541 14048
rect 40483 14007 40541 14008
rect 3907 13880 3965 13881
rect 3907 13840 3916 13880
rect 3956 13840 3965 13880
rect 3907 13839 3965 13840
rect 8235 13880 8277 13889
rect 8235 13840 8236 13880
rect 8276 13840 8277 13880
rect 8235 13831 8277 13840
rect 11971 13880 12029 13881
rect 11971 13840 11980 13880
rect 12020 13840 12029 13880
rect 11971 13839 12029 13840
rect 25707 13880 25749 13889
rect 25707 13840 25708 13880
rect 25748 13840 25749 13880
rect 25707 13831 25749 13840
rect 28971 13880 29013 13889
rect 28971 13840 28972 13880
rect 29012 13840 29013 13880
rect 28971 13831 29013 13840
rect 29731 13880 29789 13881
rect 29731 13840 29740 13880
rect 29780 13840 29789 13880
rect 29731 13839 29789 13840
rect 32139 13880 32181 13889
rect 32139 13840 32140 13880
rect 32180 13840 32181 13880
rect 32139 13831 32181 13840
rect 33483 13880 33525 13889
rect 33483 13840 33484 13880
rect 33524 13840 33525 13880
rect 33483 13831 33525 13840
rect 39627 13880 39669 13889
rect 39627 13840 39628 13880
rect 39668 13840 39669 13880
rect 39627 13831 39669 13840
rect 8707 13796 8765 13797
rect 8707 13756 8716 13796
rect 8756 13756 8765 13796
rect 8707 13755 8765 13756
rect 12163 13796 12221 13797
rect 12163 13756 12172 13796
rect 12212 13756 12221 13796
rect 12163 13755 12221 13756
rect 13995 13796 14037 13805
rect 13995 13756 13996 13796
rect 14036 13756 14037 13796
rect 13995 13747 14037 13756
rect 14763 13796 14805 13805
rect 14763 13756 14764 13796
rect 14804 13756 14805 13796
rect 14763 13747 14805 13756
rect 15243 13796 15285 13805
rect 15243 13756 15244 13796
rect 15284 13756 15285 13796
rect 15243 13747 15285 13756
rect 16299 13796 16341 13805
rect 16299 13756 16300 13796
rect 16340 13756 16341 13796
rect 16299 13747 16341 13756
rect 21291 13796 21333 13805
rect 21291 13756 21292 13796
rect 21332 13756 21333 13796
rect 21291 13747 21333 13756
rect 22539 13796 22581 13805
rect 22539 13756 22540 13796
rect 22580 13756 22581 13796
rect 22539 13747 22581 13756
rect 38083 13796 38141 13797
rect 38083 13756 38092 13796
rect 38132 13756 38141 13796
rect 38083 13755 38141 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 5635 13460 5693 13461
rect 5635 13420 5644 13460
rect 5684 13420 5693 13460
rect 5635 13419 5693 13420
rect 6507 13460 6549 13469
rect 6507 13420 6508 13460
rect 6548 13420 6549 13460
rect 6507 13411 6549 13420
rect 9579 13460 9621 13469
rect 9579 13420 9580 13460
rect 9620 13420 9621 13460
rect 9579 13411 9621 13420
rect 13323 13460 13365 13469
rect 13323 13420 13324 13460
rect 13364 13420 13365 13460
rect 13323 13411 13365 13420
rect 14763 13460 14805 13469
rect 14763 13420 14764 13460
rect 14804 13420 14805 13460
rect 14763 13411 14805 13420
rect 15243 13460 15285 13469
rect 15243 13420 15244 13460
rect 15284 13420 15285 13460
rect 15243 13411 15285 13420
rect 16299 13460 16341 13469
rect 16299 13420 16300 13460
rect 16340 13420 16341 13460
rect 16299 13411 16341 13420
rect 27723 13460 27765 13469
rect 27723 13420 27724 13460
rect 27764 13420 27765 13460
rect 27723 13411 27765 13420
rect 29259 13460 29301 13469
rect 29259 13420 29260 13460
rect 29300 13420 29301 13460
rect 29259 13411 29301 13420
rect 36171 13460 36213 13469
rect 36171 13420 36172 13460
rect 36212 13420 36213 13460
rect 36171 13411 36213 13420
rect 10059 13376 10101 13385
rect 10059 13336 10060 13376
rect 10100 13336 10101 13376
rect 10059 13327 10101 13336
rect 12267 13376 12309 13385
rect 12267 13336 12268 13376
rect 12308 13336 12309 13376
rect 12267 13327 12309 13336
rect 26667 13376 26709 13385
rect 26667 13336 26668 13376
rect 26708 13336 26709 13376
rect 26667 13327 26709 13336
rect 28203 13376 28245 13385
rect 28203 13336 28204 13376
rect 28244 13336 28245 13376
rect 28203 13327 28245 13336
rect 30219 13376 30261 13385
rect 30219 13336 30220 13376
rect 30260 13336 30261 13376
rect 30219 13327 30261 13336
rect 31555 13376 31613 13377
rect 31555 13336 31564 13376
rect 31604 13336 31613 13376
rect 31555 13335 31613 13336
rect 39339 13376 39381 13385
rect 39339 13336 39340 13376
rect 39380 13336 39381 13376
rect 39339 13327 39381 13336
rect 11203 13292 11261 13293
rect 11203 13252 11212 13292
rect 11252 13252 11261 13292
rect 11203 13251 11261 13252
rect 24843 13292 24885 13301
rect 24843 13252 24844 13292
rect 24884 13252 24885 13292
rect 24843 13243 24885 13252
rect 26571 13292 26613 13301
rect 26571 13252 26572 13292
rect 26612 13252 26613 13292
rect 26571 13243 26613 13252
rect 26763 13292 26805 13301
rect 26763 13252 26764 13292
rect 26804 13252 26805 13292
rect 26763 13243 26805 13252
rect 27915 13250 27957 13259
rect 21613 13223 21655 13232
rect 3243 13208 3285 13217
rect 3243 13168 3244 13208
rect 3284 13168 3285 13208
rect 3243 13159 3285 13168
rect 3619 13208 3677 13209
rect 3619 13168 3628 13208
rect 3668 13168 3677 13208
rect 3619 13167 3677 13168
rect 4483 13208 4541 13209
rect 4483 13168 4492 13208
rect 4532 13168 4541 13208
rect 4483 13167 4541 13168
rect 5827 13208 5885 13209
rect 5827 13168 5836 13208
rect 5876 13168 5885 13208
rect 5827 13167 5885 13168
rect 6787 13208 6845 13209
rect 6787 13168 6796 13208
rect 6836 13168 6845 13208
rect 6787 13167 6845 13168
rect 7179 13208 7221 13217
rect 7179 13168 7180 13208
rect 7220 13168 7221 13208
rect 7179 13159 7221 13168
rect 7555 13208 7613 13209
rect 7555 13168 7564 13208
rect 7604 13168 7613 13208
rect 7555 13167 7613 13168
rect 8419 13208 8477 13209
rect 8419 13168 8428 13208
rect 8468 13168 8477 13208
rect 8419 13167 8477 13168
rect 12459 13208 12501 13217
rect 12459 13168 12460 13208
rect 12500 13168 12501 13208
rect 12459 13159 12501 13168
rect 13027 13208 13085 13209
rect 13027 13168 13036 13208
rect 13076 13168 13085 13208
rect 13027 13167 13085 13168
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 13315 13208 13373 13209
rect 13315 13168 13324 13208
rect 13364 13168 13373 13208
rect 13315 13167 13373 13168
rect 13795 13208 13853 13209
rect 13795 13168 13804 13208
rect 13844 13168 13853 13208
rect 13795 13167 13853 13168
rect 13891 13208 13949 13209
rect 13891 13168 13900 13208
rect 13940 13168 13949 13208
rect 13891 13167 13949 13168
rect 14371 13208 14429 13209
rect 14371 13168 14380 13208
rect 14420 13168 14429 13208
rect 14371 13167 14429 13168
rect 14475 13208 14517 13217
rect 14475 13168 14476 13208
rect 14516 13168 14517 13208
rect 14475 13159 14517 13168
rect 14947 13208 15005 13209
rect 14947 13168 14956 13208
rect 14996 13168 15005 13208
rect 14947 13167 15005 13168
rect 15051 13208 15093 13217
rect 15051 13168 15052 13208
rect 15092 13168 15093 13208
rect 15051 13159 15093 13168
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15435 13208 15477 13217
rect 15435 13168 15436 13208
rect 15476 13168 15477 13208
rect 15435 13159 15477 13168
rect 15531 13208 15573 13217
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 15619 13208 15677 13209
rect 15619 13168 15628 13208
rect 15668 13168 15677 13208
rect 15619 13167 15677 13168
rect 16003 13208 16061 13209
rect 16003 13168 16012 13208
rect 16052 13168 16061 13208
rect 16003 13167 16061 13168
rect 16107 13208 16149 13217
rect 16107 13168 16108 13208
rect 16148 13168 16149 13208
rect 16107 13159 16149 13168
rect 16299 13208 16341 13217
rect 16299 13168 16300 13208
rect 16340 13168 16341 13208
rect 16299 13159 16341 13168
rect 16963 13208 17021 13209
rect 16963 13168 16972 13208
rect 17012 13168 17021 13208
rect 16963 13167 17021 13168
rect 17067 13208 17109 13217
rect 17067 13168 17068 13208
rect 17108 13168 17109 13208
rect 17067 13159 17109 13168
rect 17259 13208 17301 13217
rect 17259 13168 17260 13208
rect 17300 13168 17301 13208
rect 17259 13159 17301 13168
rect 17635 13208 17693 13209
rect 17635 13168 17644 13208
rect 17684 13168 17693 13208
rect 17635 13167 17693 13168
rect 17731 13208 17789 13209
rect 17731 13168 17740 13208
rect 17780 13168 17789 13208
rect 17731 13167 17789 13168
rect 17931 13208 17973 13217
rect 17931 13168 17932 13208
rect 17972 13168 17973 13208
rect 17931 13159 17973 13168
rect 18027 13208 18069 13217
rect 18027 13168 18028 13208
rect 18068 13168 18069 13208
rect 18027 13159 18069 13168
rect 18120 13208 18178 13209
rect 18120 13168 18129 13208
rect 18169 13168 18178 13208
rect 18120 13167 18178 13168
rect 19083 13208 19125 13217
rect 19083 13168 19084 13208
rect 19124 13168 19125 13208
rect 19083 13159 19125 13168
rect 19275 13208 19317 13217
rect 19275 13168 19276 13208
rect 19316 13168 19317 13208
rect 19275 13159 19317 13168
rect 19363 13208 19421 13209
rect 19363 13168 19372 13208
rect 19412 13168 19421 13208
rect 19363 13167 19421 13168
rect 19659 13208 19701 13217
rect 19659 13168 19660 13208
rect 19700 13168 19701 13208
rect 19659 13159 19701 13168
rect 19755 13208 19797 13217
rect 19755 13168 19756 13208
rect 19796 13168 19797 13208
rect 19755 13159 19797 13168
rect 19851 13208 19893 13217
rect 19851 13168 19852 13208
rect 19892 13168 19893 13208
rect 19851 13159 19893 13168
rect 20331 13208 20373 13217
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 20427 13208 20469 13217
rect 20427 13168 20428 13208
rect 20468 13168 20469 13208
rect 20427 13159 20469 13168
rect 21099 13208 21141 13217
rect 21099 13168 21100 13208
rect 21140 13168 21141 13208
rect 21099 13159 21141 13168
rect 21195 13208 21237 13217
rect 21195 13168 21196 13208
rect 21236 13168 21237 13208
rect 21195 13159 21237 13168
rect 21291 13208 21333 13217
rect 21291 13168 21292 13208
rect 21332 13168 21333 13208
rect 21613 13183 21614 13223
rect 21654 13183 21655 13223
rect 21613 13174 21655 13183
rect 21771 13208 21813 13217
rect 21291 13159 21333 13168
rect 21771 13168 21772 13208
rect 21812 13168 21813 13208
rect 21771 13159 21813 13168
rect 21867 13208 21909 13217
rect 21867 13168 21868 13208
rect 21908 13168 21909 13208
rect 21867 13159 21909 13168
rect 22051 13208 22109 13209
rect 22051 13168 22060 13208
rect 22100 13168 22109 13208
rect 22051 13167 22109 13168
rect 22147 13208 22205 13209
rect 22147 13168 22156 13208
rect 22196 13168 22205 13208
rect 22147 13167 22205 13168
rect 22443 13208 22485 13217
rect 22443 13168 22444 13208
rect 22484 13168 22485 13208
rect 22443 13159 22485 13168
rect 22819 13208 22877 13209
rect 22819 13168 22828 13208
rect 22868 13168 22877 13208
rect 22819 13167 22877 13168
rect 23683 13208 23741 13209
rect 23683 13168 23692 13208
rect 23732 13168 23741 13208
rect 23683 13167 23741 13168
rect 26083 13208 26141 13209
rect 26083 13168 26092 13208
rect 26132 13168 26141 13208
rect 26083 13167 26141 13168
rect 26859 13208 26901 13217
rect 26859 13168 26860 13208
rect 26900 13168 26901 13208
rect 26467 13166 26525 13167
rect 17163 13124 17205 13133
rect 17163 13084 17164 13124
rect 17204 13084 17205 13124
rect 17163 13075 17205 13084
rect 19179 13124 19221 13133
rect 26467 13126 26476 13166
rect 26516 13126 26525 13166
rect 26859 13159 26901 13168
rect 27051 13208 27093 13217
rect 27051 13168 27052 13208
rect 27092 13168 27093 13208
rect 27051 13159 27093 13168
rect 27147 13208 27189 13217
rect 27147 13168 27148 13208
rect 27188 13168 27189 13208
rect 27147 13159 27189 13168
rect 27243 13208 27285 13217
rect 27243 13168 27244 13208
rect 27284 13168 27285 13208
rect 27243 13159 27285 13168
rect 27339 13208 27381 13217
rect 27915 13210 27916 13250
rect 27956 13210 27957 13250
rect 27339 13168 27340 13208
rect 27380 13168 27381 13208
rect 27339 13159 27381 13168
rect 27715 13208 27773 13209
rect 27715 13168 27724 13208
rect 27764 13168 27773 13208
rect 27915 13201 27957 13210
rect 28003 13208 28061 13209
rect 27715 13167 27773 13168
rect 28003 13168 28012 13208
rect 28052 13168 28061 13208
rect 28395 13208 28437 13217
rect 28003 13167 28061 13168
rect 28203 13166 28245 13175
rect 26467 13125 26525 13126
rect 28203 13126 28204 13166
rect 28244 13126 28245 13166
rect 28395 13168 28396 13208
rect 28436 13168 28437 13208
rect 28395 13159 28437 13168
rect 28483 13208 28541 13209
rect 28483 13168 28492 13208
rect 28532 13168 28541 13208
rect 28483 13167 28541 13168
rect 28675 13208 28733 13209
rect 28675 13168 28684 13208
rect 28724 13168 28733 13208
rect 28675 13167 28733 13168
rect 28779 13208 28821 13217
rect 28779 13168 28780 13208
rect 28820 13168 28821 13208
rect 28779 13159 28821 13168
rect 28971 13208 29013 13217
rect 28971 13168 28972 13208
rect 29012 13168 29013 13208
rect 28971 13159 29013 13168
rect 29451 13208 29493 13217
rect 29451 13168 29452 13208
rect 29492 13168 29493 13208
rect 29451 13159 29493 13168
rect 29547 13208 29589 13217
rect 29547 13168 29548 13208
rect 29588 13168 29589 13208
rect 29547 13159 29589 13168
rect 29739 13208 29781 13217
rect 29739 13168 29740 13208
rect 29780 13168 29781 13208
rect 29739 13159 29781 13168
rect 29835 13208 29877 13217
rect 29835 13168 29836 13208
rect 29876 13168 29877 13208
rect 29835 13159 29877 13168
rect 30219 13208 30261 13217
rect 30219 13168 30220 13208
rect 30260 13168 30261 13208
rect 30219 13159 30261 13168
rect 30411 13208 30453 13217
rect 30411 13168 30412 13208
rect 30452 13168 30453 13208
rect 30411 13159 30453 13168
rect 30603 13208 30645 13217
rect 30603 13168 30604 13208
rect 30644 13168 30645 13208
rect 30603 13159 30645 13168
rect 30795 13208 30837 13217
rect 30795 13168 30796 13208
rect 30836 13168 30837 13208
rect 30795 13159 30837 13168
rect 31363 13208 31421 13209
rect 31363 13168 31372 13208
rect 31412 13168 31421 13208
rect 31363 13167 31421 13168
rect 31563 13208 31605 13217
rect 31563 13168 31564 13208
rect 31604 13168 31605 13208
rect 31563 13159 31605 13168
rect 31651 13208 31709 13209
rect 31651 13168 31660 13208
rect 31700 13168 31709 13208
rect 31651 13167 31709 13168
rect 32235 13208 32277 13217
rect 32235 13168 32236 13208
rect 32276 13168 32277 13208
rect 32235 13159 32277 13168
rect 32427 13208 32469 13217
rect 32427 13168 32428 13208
rect 32468 13168 32469 13208
rect 32427 13159 32469 13168
rect 32515 13208 32573 13209
rect 32515 13168 32524 13208
rect 32564 13168 32573 13208
rect 32515 13167 32573 13168
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 33003 13208 33045 13217
rect 33003 13168 33004 13208
rect 33044 13168 33045 13208
rect 33003 13159 33045 13168
rect 33099 13208 33141 13217
rect 33099 13168 33100 13208
rect 33140 13168 33141 13208
rect 33099 13159 33141 13168
rect 33291 13208 33333 13217
rect 33291 13168 33292 13208
rect 33332 13168 33333 13208
rect 33291 13159 33333 13168
rect 33483 13208 33525 13217
rect 33483 13168 33484 13208
rect 33524 13168 33525 13208
rect 33483 13159 33525 13168
rect 33571 13208 33629 13209
rect 33571 13168 33580 13208
rect 33620 13168 33629 13208
rect 33571 13167 33629 13168
rect 33771 13208 33813 13217
rect 33771 13168 33772 13208
rect 33812 13168 33813 13208
rect 33771 13159 33813 13168
rect 34147 13208 34205 13209
rect 34147 13168 34156 13208
rect 34196 13168 34205 13208
rect 34147 13167 34205 13168
rect 35011 13208 35069 13209
rect 35011 13168 35020 13208
rect 35060 13168 35069 13208
rect 35011 13167 35069 13168
rect 36939 13208 36981 13217
rect 36939 13168 36940 13208
rect 36980 13168 36981 13208
rect 36939 13159 36981 13168
rect 37315 13208 37373 13209
rect 37315 13168 37324 13208
rect 37364 13168 37373 13208
rect 37315 13167 37373 13168
rect 38179 13208 38237 13209
rect 38179 13168 38188 13208
rect 38228 13168 38237 13208
rect 38179 13167 38237 13168
rect 19179 13084 19180 13124
rect 19220 13084 19221 13124
rect 28203 13117 28245 13126
rect 28875 13124 28917 13133
rect 19179 13075 19221 13084
rect 28875 13084 28876 13124
rect 28916 13084 28917 13124
rect 20131 13082 20189 13083
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 12075 13040 12117 13049
rect 12075 13000 12076 13040
rect 12116 13000 12117 13040
rect 12075 12991 12117 13000
rect 14091 13040 14133 13049
rect 14091 13000 14092 13040
rect 14132 13000 14133 13040
rect 14091 12991 14133 13000
rect 14283 13036 14325 13045
rect 20131 13042 20140 13082
rect 20180 13042 20189 13082
rect 28875 13075 28917 13084
rect 29347 13124 29405 13125
rect 29347 13084 29356 13124
rect 29396 13084 29405 13124
rect 29347 13083 29405 13084
rect 32331 13124 32373 13133
rect 32331 13084 32332 13124
rect 32372 13084 32373 13124
rect 32331 13075 32373 13084
rect 33387 13124 33429 13133
rect 33387 13084 33388 13124
rect 33428 13084 33429 13124
rect 33387 13075 33429 13084
rect 20131 13041 20189 13042
rect 14283 12996 14284 13036
rect 14324 12996 14325 13036
rect 17827 13040 17885 13041
rect 17827 13000 17836 13040
rect 17876 13000 17885 13040
rect 17827 12999 17885 13000
rect 19555 13040 19613 13041
rect 19555 13000 19564 13040
rect 19604 13000 19613 13040
rect 19555 12999 19613 13000
rect 21379 13040 21437 13041
rect 21379 13000 21388 13040
rect 21428 13000 21437 13040
rect 21379 12999 21437 13000
rect 21667 13040 21725 13041
rect 21667 13000 21676 13040
rect 21716 13000 21725 13040
rect 21667 12999 21725 13000
rect 25411 13040 25469 13041
rect 25411 13000 25420 13040
rect 25460 13000 25469 13040
rect 25411 12999 25469 13000
rect 29251 13040 29309 13041
rect 29251 13000 29260 13040
rect 29300 13000 29309 13040
rect 29251 12999 29309 13000
rect 30019 13040 30077 13041
rect 30019 13000 30028 13040
rect 30068 13000 30077 13040
rect 30019 12999 30077 13000
rect 30699 13040 30741 13049
rect 30699 13000 30700 13040
rect 30740 13000 30741 13040
rect 14283 12987 14325 12996
rect 30699 12991 30741 13000
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 14947 12704 15005 12705
rect 14947 12664 14956 12704
rect 14996 12664 15005 12704
rect 14947 12663 15005 12664
rect 19363 12704 19421 12705
rect 19363 12664 19372 12704
rect 19412 12664 19421 12704
rect 19363 12663 19421 12664
rect 27051 12704 27093 12713
rect 27051 12664 27052 12704
rect 27092 12664 27093 12704
rect 27051 12655 27093 12664
rect 27235 12704 27293 12705
rect 27235 12664 27244 12704
rect 27284 12664 27293 12704
rect 27235 12663 27293 12664
rect 28675 12704 28733 12705
rect 28675 12664 28684 12704
rect 28724 12664 28733 12704
rect 28675 12663 28733 12664
rect 34723 12704 34781 12705
rect 34723 12664 34732 12704
rect 34772 12664 34781 12704
rect 34723 12663 34781 12664
rect 36931 12704 36989 12705
rect 36931 12664 36940 12704
rect 36980 12664 36989 12704
rect 36931 12663 36989 12664
rect 4299 12620 4341 12629
rect 4299 12580 4300 12620
rect 4340 12580 4341 12620
rect 4299 12571 4341 12580
rect 5355 12620 5397 12629
rect 5355 12580 5356 12620
rect 5396 12580 5397 12620
rect 5355 12571 5397 12580
rect 5835 12620 5877 12629
rect 5835 12580 5836 12620
rect 5876 12580 5877 12620
rect 5835 12571 5877 12580
rect 9675 12620 9717 12629
rect 9675 12580 9676 12620
rect 9716 12580 9717 12620
rect 9675 12571 9717 12580
rect 13803 12620 13845 12629
rect 13803 12580 13804 12620
rect 13844 12580 13845 12620
rect 13803 12571 13845 12580
rect 18603 12620 18645 12629
rect 18603 12580 18604 12620
rect 18644 12580 18645 12620
rect 18603 12571 18645 12580
rect 21195 12620 21237 12629
rect 21195 12580 21196 12620
rect 21236 12580 21237 12620
rect 21195 12571 21237 12580
rect 27819 12620 27861 12629
rect 27819 12580 27820 12620
rect 27860 12580 27861 12620
rect 35499 12620 35541 12629
rect 27819 12571 27861 12580
rect 29355 12578 29397 12587
rect 18507 12557 18549 12566
rect 3723 12536 3765 12545
rect 3723 12496 3724 12536
rect 3764 12496 3765 12536
rect 3723 12487 3765 12496
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 3915 12487 3957 12496
rect 4203 12536 4245 12545
rect 4203 12496 4204 12536
rect 4244 12496 4245 12536
rect 4203 12487 4245 12496
rect 4395 12536 4437 12545
rect 4395 12496 4396 12536
rect 4436 12496 4437 12536
rect 4395 12487 4437 12496
rect 4491 12536 4533 12545
rect 4491 12496 4492 12536
rect 4532 12496 4533 12536
rect 4491 12487 4533 12496
rect 5163 12536 5205 12545
rect 5163 12496 5164 12536
rect 5204 12496 5205 12536
rect 5163 12487 5205 12496
rect 5451 12536 5493 12545
rect 5451 12496 5452 12536
rect 5492 12496 5493 12536
rect 5451 12487 5493 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 5931 12536 5973 12545
rect 5931 12496 5932 12536
rect 5972 12496 5973 12536
rect 5931 12487 5973 12496
rect 6019 12536 6077 12537
rect 6019 12496 6028 12536
rect 6068 12496 6077 12536
rect 6019 12495 6077 12496
rect 7075 12536 7133 12537
rect 7075 12496 7084 12536
rect 7124 12496 7133 12536
rect 7075 12495 7133 12496
rect 8323 12536 8381 12537
rect 8323 12496 8332 12536
rect 8372 12496 8381 12536
rect 8323 12495 8381 12496
rect 8619 12536 8661 12545
rect 8619 12496 8620 12536
rect 8660 12496 8661 12536
rect 8619 12487 8661 12496
rect 9283 12536 9341 12537
rect 9283 12496 9292 12536
rect 9332 12496 9341 12536
rect 9283 12495 9341 12496
rect 9475 12536 9533 12537
rect 9475 12496 9484 12536
rect 9524 12496 9533 12536
rect 9475 12495 9533 12496
rect 9579 12536 9621 12545
rect 9579 12496 9580 12536
rect 9620 12496 9621 12536
rect 9579 12487 9621 12496
rect 9771 12536 9813 12545
rect 9771 12496 9772 12536
rect 9812 12496 9813 12536
rect 9771 12487 9813 12496
rect 10627 12536 10685 12537
rect 10627 12496 10636 12536
rect 10676 12496 10685 12536
rect 10627 12495 10685 12496
rect 12643 12536 12701 12537
rect 12643 12496 12652 12536
rect 12692 12496 12701 12536
rect 12643 12495 12701 12496
rect 13227 12536 13269 12545
rect 13227 12496 13228 12536
rect 13268 12496 13269 12536
rect 13227 12487 13269 12496
rect 13323 12536 13365 12545
rect 13323 12496 13324 12536
rect 13364 12496 13365 12536
rect 13323 12487 13365 12496
rect 13419 12536 13461 12545
rect 13419 12496 13420 12536
rect 13460 12496 13461 12536
rect 13419 12487 13461 12496
rect 13515 12536 13557 12545
rect 13515 12496 13516 12536
rect 13556 12496 13557 12536
rect 13515 12487 13557 12496
rect 13707 12536 13749 12545
rect 13707 12496 13708 12536
rect 13748 12496 13749 12536
rect 13707 12487 13749 12496
rect 13899 12536 13941 12545
rect 13899 12496 13900 12536
rect 13940 12496 13941 12536
rect 13899 12487 13941 12496
rect 13987 12536 14045 12537
rect 13987 12496 13996 12536
rect 14036 12496 14045 12536
rect 13987 12495 14045 12496
rect 14379 12536 14421 12545
rect 14379 12496 14380 12536
rect 14420 12496 14421 12536
rect 14379 12487 14421 12496
rect 14667 12536 14709 12545
rect 14667 12496 14668 12536
rect 14708 12496 14709 12536
rect 14667 12487 14709 12496
rect 14763 12536 14805 12545
rect 14763 12496 14764 12536
rect 14804 12496 14805 12536
rect 14763 12487 14805 12496
rect 14859 12536 14901 12545
rect 14859 12496 14860 12536
rect 14900 12496 14901 12536
rect 14859 12487 14901 12496
rect 15435 12536 15477 12545
rect 15435 12496 15436 12536
rect 15476 12496 15477 12536
rect 15435 12487 15477 12496
rect 15723 12536 15765 12545
rect 15723 12496 15724 12536
rect 15764 12496 15765 12536
rect 15523 12494 15581 12495
rect 3819 12452 3861 12461
rect 3819 12412 3820 12452
rect 3860 12412 3861 12452
rect 3819 12403 3861 12412
rect 11587 12452 11645 12453
rect 11587 12412 11596 12452
rect 11636 12412 11645 12452
rect 11587 12411 11645 12412
rect 15339 12452 15381 12461
rect 15523 12454 15532 12494
rect 15572 12454 15581 12494
rect 15723 12487 15765 12496
rect 15915 12536 15957 12545
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 15915 12487 15957 12496
rect 16003 12536 16061 12537
rect 16003 12496 16012 12536
rect 16052 12496 16061 12536
rect 16003 12495 16061 12496
rect 16203 12536 16245 12545
rect 16203 12496 16204 12536
rect 16244 12496 16245 12536
rect 16203 12487 16245 12496
rect 16395 12536 16437 12545
rect 16395 12496 16396 12536
rect 16436 12496 16437 12536
rect 16395 12487 16437 12496
rect 16579 12536 16637 12537
rect 16579 12496 16588 12536
rect 16628 12496 16637 12536
rect 16579 12495 16637 12496
rect 16683 12536 16725 12545
rect 16683 12496 16684 12536
rect 16724 12496 16725 12536
rect 16683 12487 16725 12496
rect 18315 12536 18357 12545
rect 18315 12496 18316 12536
rect 18356 12496 18357 12536
rect 18315 12487 18357 12496
rect 18411 12536 18453 12545
rect 18411 12496 18412 12536
rect 18452 12496 18453 12536
rect 18507 12517 18508 12557
rect 18548 12517 18549 12557
rect 18507 12508 18549 12517
rect 18795 12536 18837 12545
rect 18411 12487 18453 12496
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 18795 12487 18837 12496
rect 18987 12536 19029 12545
rect 18987 12496 18988 12536
rect 19028 12496 19029 12536
rect 18987 12487 19029 12496
rect 19075 12536 19133 12537
rect 19075 12496 19084 12536
rect 19124 12496 19133 12536
rect 19075 12495 19133 12496
rect 19358 12536 19416 12537
rect 19358 12496 19367 12536
rect 19407 12496 19416 12536
rect 19358 12495 19416 12496
rect 19467 12536 19509 12545
rect 19467 12496 19468 12536
rect 19508 12496 19509 12536
rect 19467 12487 19509 12496
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19747 12536 19805 12537
rect 19747 12496 19756 12536
rect 19796 12496 19805 12536
rect 19747 12495 19805 12496
rect 19843 12536 19901 12537
rect 19843 12496 19852 12536
rect 19892 12496 19901 12536
rect 19843 12495 19901 12496
rect 20043 12536 20085 12545
rect 20043 12496 20044 12536
rect 20084 12496 20085 12536
rect 20043 12487 20085 12496
rect 20139 12536 20181 12545
rect 20139 12496 20140 12536
rect 20180 12496 20181 12536
rect 20139 12487 20181 12496
rect 20235 12536 20277 12545
rect 20235 12496 20236 12536
rect 20276 12496 20277 12536
rect 20235 12487 20277 12496
rect 20331 12536 20373 12545
rect 20331 12496 20332 12536
rect 20372 12496 20373 12536
rect 20331 12487 20373 12496
rect 20619 12536 20661 12545
rect 20619 12496 20620 12536
rect 20660 12496 20661 12536
rect 20619 12487 20661 12496
rect 20715 12536 20757 12545
rect 20715 12496 20716 12536
rect 20756 12496 20757 12536
rect 20715 12487 20757 12496
rect 20811 12536 20853 12545
rect 20811 12496 20812 12536
rect 20852 12496 20853 12536
rect 20811 12487 20853 12496
rect 20907 12536 20949 12545
rect 20907 12496 20908 12536
rect 20948 12496 20949 12536
rect 20907 12487 20949 12496
rect 21099 12536 21141 12545
rect 21099 12496 21100 12536
rect 21140 12496 21141 12536
rect 21099 12487 21141 12496
rect 21291 12536 21333 12545
rect 21291 12496 21292 12536
rect 21332 12496 21333 12536
rect 21291 12487 21333 12496
rect 21379 12536 21437 12537
rect 21379 12496 21388 12536
rect 21428 12496 21437 12536
rect 21379 12495 21437 12496
rect 21571 12536 21629 12537
rect 21571 12496 21580 12536
rect 21620 12496 21629 12536
rect 21571 12495 21629 12496
rect 24739 12536 24797 12537
rect 24739 12496 24748 12536
rect 24788 12496 24797 12536
rect 24739 12495 24797 12496
rect 25611 12536 25653 12545
rect 25611 12496 25612 12536
rect 25652 12496 25653 12536
rect 25611 12487 25653 12496
rect 25987 12536 26045 12537
rect 25987 12496 25996 12536
rect 26036 12496 26045 12536
rect 25987 12495 26045 12496
rect 26379 12536 26421 12545
rect 26379 12496 26380 12536
rect 26420 12496 26421 12536
rect 26379 12487 26421 12496
rect 26667 12536 26709 12545
rect 26667 12496 26668 12536
rect 26708 12496 26709 12536
rect 26667 12487 26709 12496
rect 26859 12536 26901 12545
rect 26859 12496 26860 12536
rect 26900 12496 26901 12536
rect 26755 12494 26813 12495
rect 15523 12453 15581 12454
rect 15339 12412 15340 12452
rect 15380 12412 15381 12452
rect 15339 12403 15381 12412
rect 26091 12452 26133 12461
rect 26091 12412 26092 12452
rect 26132 12412 26133 12452
rect 26091 12403 26133 12412
rect 26283 12452 26325 12461
rect 26755 12454 26764 12494
rect 26804 12454 26813 12494
rect 26859 12487 26901 12496
rect 27435 12536 27477 12545
rect 27435 12496 27436 12536
rect 27476 12496 27477 12536
rect 27435 12487 27477 12496
rect 27531 12536 27573 12545
rect 27531 12496 27532 12536
rect 27572 12496 27573 12536
rect 27531 12487 27573 12496
rect 27723 12536 27765 12545
rect 27723 12496 27724 12536
rect 27764 12496 27765 12536
rect 27723 12487 27765 12496
rect 27907 12536 27965 12537
rect 27907 12496 27916 12536
rect 27956 12496 27965 12536
rect 27907 12495 27965 12496
rect 28387 12536 28445 12537
rect 28387 12496 28396 12536
rect 28436 12496 28445 12536
rect 28387 12495 28445 12496
rect 28875 12536 28917 12545
rect 28875 12496 28876 12536
rect 28916 12496 28917 12536
rect 28875 12487 28917 12496
rect 28971 12536 29013 12545
rect 28971 12496 28972 12536
rect 29012 12496 29013 12536
rect 28971 12487 29013 12496
rect 29163 12536 29205 12545
rect 29163 12496 29164 12536
rect 29204 12496 29205 12536
rect 29355 12538 29356 12578
rect 29396 12538 29397 12578
rect 35499 12580 35500 12620
rect 35540 12580 35541 12620
rect 35499 12571 35541 12580
rect 36259 12620 36317 12621
rect 36259 12580 36268 12620
rect 36308 12580 36317 12620
rect 36259 12579 36317 12580
rect 29355 12529 29397 12538
rect 29539 12536 29597 12537
rect 29163 12487 29205 12496
rect 29539 12496 29548 12536
rect 29588 12496 29597 12536
rect 29539 12495 29597 12496
rect 29931 12536 29973 12545
rect 29931 12496 29932 12536
rect 29972 12496 29973 12536
rect 29931 12487 29973 12496
rect 30027 12536 30069 12545
rect 30027 12496 30028 12536
rect 30068 12496 30069 12536
rect 30027 12487 30069 12496
rect 30123 12536 30165 12545
rect 30123 12496 30124 12536
rect 30164 12496 30165 12536
rect 30123 12487 30165 12496
rect 30219 12536 30261 12545
rect 30219 12496 30220 12536
rect 30260 12496 30261 12536
rect 30219 12487 30261 12496
rect 32035 12536 32093 12537
rect 32035 12496 32044 12536
rect 32084 12496 32093 12536
rect 32035 12495 32093 12496
rect 33283 12536 33341 12537
rect 33283 12496 33292 12536
rect 33332 12496 33341 12536
rect 33283 12495 33341 12496
rect 34443 12536 34485 12545
rect 34443 12496 34444 12536
rect 34484 12496 34485 12536
rect 34443 12487 34485 12496
rect 34539 12536 34581 12545
rect 34539 12496 34540 12536
rect 34580 12496 34581 12536
rect 34539 12487 34581 12496
rect 35395 12536 35453 12537
rect 35395 12496 35404 12536
rect 35444 12496 35453 12536
rect 35395 12495 35453 12496
rect 35683 12536 35741 12537
rect 35683 12496 35692 12536
rect 35732 12496 35741 12536
rect 35683 12495 35741 12496
rect 35787 12536 35829 12545
rect 35787 12496 35788 12536
rect 35828 12496 35829 12536
rect 35787 12487 35829 12496
rect 35979 12536 36021 12545
rect 35979 12496 35980 12536
rect 36020 12496 36021 12536
rect 35979 12487 36021 12496
rect 36355 12536 36413 12537
rect 36355 12496 36364 12536
rect 36404 12496 36413 12536
rect 36355 12495 36413 12496
rect 36739 12536 36797 12537
rect 36739 12496 36748 12536
rect 36788 12496 36797 12536
rect 36739 12495 36797 12496
rect 37603 12536 37661 12537
rect 37603 12496 37612 12536
rect 37652 12496 37661 12536
rect 37603 12495 37661 12496
rect 39043 12536 39101 12537
rect 39043 12496 39052 12536
rect 39092 12496 39101 12536
rect 39043 12495 39101 12496
rect 26755 12453 26813 12454
rect 26283 12412 26284 12452
rect 26324 12412 26325 12452
rect 26283 12403 26325 12412
rect 29259 12452 29301 12461
rect 29259 12412 29260 12452
rect 29300 12412 29301 12452
rect 29259 12403 29301 12412
rect 29451 12452 29493 12461
rect 29451 12412 29452 12452
rect 29492 12412 29493 12452
rect 29451 12403 29493 12412
rect 4683 12368 4725 12377
rect 4683 12328 4684 12368
rect 4724 12328 4725 12368
rect 4683 12319 4725 12328
rect 6219 12368 6261 12377
rect 6219 12328 6220 12368
rect 6260 12328 6261 12368
rect 6219 12319 6261 12328
rect 6603 12368 6645 12377
rect 6603 12328 6604 12368
rect 6644 12328 6645 12368
rect 6603 12319 6645 12328
rect 6987 12368 7029 12377
rect 6987 12328 6988 12368
rect 7028 12328 7029 12368
rect 6987 12319 7029 12328
rect 7467 12368 7509 12377
rect 7467 12328 7468 12368
rect 7508 12328 7509 12368
rect 7467 12319 7509 12328
rect 10827 12368 10869 12377
rect 10827 12328 10828 12368
rect 10868 12328 10869 12368
rect 10827 12319 10869 12328
rect 14187 12368 14229 12377
rect 14187 12328 14188 12368
rect 14228 12328 14229 12368
rect 14187 12319 14229 12328
rect 14379 12368 14421 12377
rect 14379 12328 14380 12368
rect 14420 12328 14421 12368
rect 14379 12319 14421 12328
rect 15147 12368 15189 12377
rect 15147 12328 15148 12368
rect 15188 12328 15189 12368
rect 15147 12319 15189 12328
rect 15243 12368 15285 12377
rect 15243 12328 15244 12368
rect 15284 12328 15285 12368
rect 15243 12319 15285 12328
rect 16203 12368 16245 12377
rect 16203 12328 16204 12368
rect 16244 12328 16245 12368
rect 16203 12319 16245 12328
rect 22923 12368 22965 12377
rect 22923 12328 22924 12368
rect 22964 12328 22965 12368
rect 22923 12319 22965 12328
rect 26187 12368 26229 12377
rect 26187 12328 26188 12368
rect 26228 12328 26229 12368
rect 26187 12319 26229 12328
rect 28491 12368 28533 12377
rect 28491 12328 28492 12368
rect 28532 12328 28533 12368
rect 28491 12319 28533 12328
rect 29731 12368 29789 12369
rect 29731 12328 29740 12368
rect 29780 12328 29789 12368
rect 29731 12327 29789 12328
rect 33579 12368 33621 12377
rect 33579 12328 33580 12368
rect 33620 12328 33621 12368
rect 33579 12319 33621 12328
rect 7651 12284 7709 12285
rect 7651 12244 7660 12284
rect 7700 12244 7709 12284
rect 7651 12243 7709 12244
rect 9955 12284 10013 12285
rect 9955 12244 9964 12284
rect 10004 12244 10013 12284
rect 9955 12243 10013 12244
rect 11787 12284 11829 12293
rect 11787 12244 11788 12284
rect 11828 12244 11829 12284
rect 11787 12235 11829 12244
rect 11971 12284 12029 12285
rect 11971 12244 11980 12284
rect 12020 12244 12029 12284
rect 11971 12243 12029 12244
rect 15723 12284 15765 12293
rect 15723 12244 15724 12284
rect 15764 12244 15765 12284
rect 15723 12235 15765 12244
rect 18795 12284 18837 12293
rect 18795 12244 18796 12284
rect 18836 12244 18837 12284
rect 18795 12235 18837 12244
rect 22243 12284 22301 12285
rect 22243 12244 22252 12284
rect 22292 12244 22301 12284
rect 22243 12243 22301 12244
rect 32331 12284 32373 12293
rect 32331 12244 32332 12284
rect 32372 12244 32373 12284
rect 32331 12235 32373 12244
rect 33771 12284 33813 12293
rect 33771 12244 33772 12284
rect 33812 12244 33813 12284
rect 33771 12235 33813 12244
rect 35979 12284 36021 12293
rect 35979 12244 35980 12284
rect 36020 12244 36021 12284
rect 35979 12235 36021 12244
rect 38379 12284 38421 12293
rect 38379 12244 38380 12284
rect 38420 12244 38421 12284
rect 38379 12235 38421 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 8419 11948 8477 11949
rect 8419 11908 8428 11948
rect 8468 11908 8477 11948
rect 8419 11907 8477 11908
rect 13707 11948 13749 11957
rect 13707 11908 13708 11948
rect 13748 11908 13749 11948
rect 13707 11899 13749 11908
rect 17835 11948 17877 11957
rect 17835 11908 17836 11948
rect 17876 11908 17877 11948
rect 17835 11899 17877 11908
rect 31083 11948 31125 11957
rect 31083 11908 31084 11948
rect 31124 11908 31125 11948
rect 31083 11899 31125 11908
rect 33195 11948 33237 11957
rect 33195 11908 33196 11948
rect 33236 11908 33237 11948
rect 33195 11899 33237 11908
rect 33963 11948 34005 11957
rect 33963 11908 33964 11948
rect 34004 11908 34005 11948
rect 33963 11899 34005 11908
rect 21195 11864 21237 11873
rect 21195 11824 21196 11864
rect 21236 11824 21237 11864
rect 21195 11815 21237 11824
rect 32715 11864 32757 11873
rect 32715 11824 32716 11864
rect 32756 11824 32757 11864
rect 32715 11815 32757 11824
rect 33483 11864 33525 11873
rect 33483 11824 33484 11864
rect 33524 11824 33525 11864
rect 33483 11815 33525 11824
rect 35019 11864 35061 11873
rect 35019 11824 35020 11864
rect 35060 11824 35061 11864
rect 33571 11822 33629 11823
rect 8811 11780 8853 11789
rect 33571 11782 33580 11822
rect 33620 11782 33629 11822
rect 35019 11815 35061 11824
rect 33571 11781 33629 11782
rect 8811 11740 8812 11780
rect 8852 11740 8853 11780
rect 8811 11731 8853 11740
rect 15523 11780 15581 11781
rect 15523 11740 15532 11780
rect 15572 11740 15581 11780
rect 15523 11739 15581 11740
rect 19267 11780 19325 11781
rect 19267 11740 19276 11780
rect 19316 11740 19325 11780
rect 19267 11739 19325 11740
rect 34923 11780 34965 11789
rect 34923 11740 34924 11780
rect 34964 11740 34965 11780
rect 34923 11731 34965 11740
rect 35115 11780 35157 11789
rect 35115 11740 35116 11780
rect 35156 11740 35157 11780
rect 35115 11731 35157 11740
rect 18376 11711 18418 11720
rect 6027 11696 6069 11705
rect 6027 11656 6028 11696
rect 6068 11656 6069 11696
rect 6027 11647 6069 11656
rect 6403 11696 6461 11697
rect 6403 11656 6412 11696
rect 6452 11656 6461 11696
rect 6403 11655 6461 11656
rect 7267 11696 7325 11697
rect 7267 11656 7276 11696
rect 7316 11656 7325 11696
rect 7267 11655 7325 11656
rect 9579 11696 9621 11705
rect 9579 11656 9580 11696
rect 9620 11656 9621 11696
rect 9579 11647 9621 11656
rect 10059 11696 10101 11705
rect 10059 11656 10060 11696
rect 10100 11656 10101 11696
rect 10059 11647 10101 11656
rect 10435 11696 10493 11697
rect 10435 11656 10444 11696
rect 10484 11656 10493 11696
rect 10435 11655 10493 11656
rect 11299 11696 11357 11697
rect 11299 11656 11308 11696
rect 11348 11656 11357 11696
rect 11299 11655 11357 11656
rect 12835 11696 12893 11697
rect 12835 11656 12844 11696
rect 12884 11656 12893 11696
rect 12835 11655 12893 11656
rect 13707 11696 13749 11705
rect 13707 11656 13708 11696
rect 13748 11656 13749 11696
rect 13707 11647 13749 11656
rect 13899 11696 13941 11705
rect 13899 11656 13900 11696
rect 13940 11656 13941 11696
rect 13899 11647 13941 11656
rect 13987 11696 14045 11697
rect 13987 11656 13996 11696
rect 14036 11656 14045 11696
rect 13987 11655 14045 11656
rect 14475 11696 14517 11705
rect 14475 11656 14476 11696
rect 14516 11656 14517 11696
rect 14475 11647 14517 11656
rect 14571 11696 14613 11705
rect 14571 11656 14572 11696
rect 14612 11656 14613 11696
rect 14571 11647 14613 11656
rect 14667 11696 14709 11705
rect 14667 11656 14668 11696
rect 14708 11656 14709 11696
rect 14667 11647 14709 11656
rect 14763 11696 14805 11705
rect 14763 11656 14764 11696
rect 14804 11656 14805 11696
rect 14763 11647 14805 11656
rect 15235 11696 15293 11697
rect 15235 11656 15244 11696
rect 15284 11656 15293 11696
rect 15235 11655 15293 11656
rect 15331 11696 15389 11697
rect 15331 11656 15340 11696
rect 15380 11656 15389 11696
rect 15331 11655 15389 11656
rect 15723 11696 15765 11705
rect 15723 11656 15724 11696
rect 15764 11656 15765 11696
rect 15723 11647 15765 11656
rect 15907 11696 15965 11697
rect 15907 11656 15916 11696
rect 15956 11656 15965 11696
rect 15907 11655 15965 11656
rect 16299 11696 16341 11705
rect 16299 11656 16300 11696
rect 16340 11656 16341 11696
rect 16299 11647 16341 11656
rect 16395 11696 16437 11705
rect 16395 11656 16396 11696
rect 16436 11656 16437 11696
rect 16395 11647 16437 11656
rect 16587 11696 16629 11705
rect 16587 11656 16588 11696
rect 16628 11656 16629 11696
rect 16587 11647 16629 11656
rect 16683 11696 16725 11705
rect 18075 11700 18117 11709
rect 16683 11656 16684 11696
rect 16724 11656 16725 11696
rect 16683 11647 16725 11656
rect 17827 11696 17885 11697
rect 17827 11656 17836 11696
rect 17876 11656 17885 11696
rect 17827 11655 17885 11656
rect 17923 11696 17981 11697
rect 17923 11656 17932 11696
rect 17972 11656 17981 11696
rect 17923 11655 17981 11656
rect 18075 11660 18076 11700
rect 18116 11660 18117 11700
rect 18075 11651 18117 11660
rect 18219 11696 18261 11705
rect 18219 11656 18220 11696
rect 18260 11656 18261 11696
rect 18376 11671 18377 11711
rect 18417 11671 18418 11711
rect 20200 11711 20242 11720
rect 18376 11662 18418 11671
rect 19651 11696 19709 11697
rect 18219 11647 18261 11656
rect 19651 11656 19660 11696
rect 19700 11656 19709 11696
rect 19651 11655 19709 11656
rect 19747 11696 19805 11697
rect 19747 11656 19756 11696
rect 19796 11656 19805 11696
rect 19747 11655 19805 11656
rect 19947 11696 19989 11705
rect 19947 11656 19948 11696
rect 19988 11656 19989 11696
rect 19947 11647 19989 11656
rect 20043 11696 20085 11705
rect 20043 11656 20044 11696
rect 20084 11656 20085 11696
rect 20200 11671 20201 11711
rect 20241 11671 20242 11711
rect 20200 11662 20242 11671
rect 21771 11696 21813 11705
rect 20043 11647 20085 11656
rect 21771 11656 21772 11696
rect 21812 11656 21813 11696
rect 21771 11647 21813 11656
rect 22147 11696 22205 11697
rect 22147 11656 22156 11696
rect 22196 11656 22205 11696
rect 22147 11655 22205 11656
rect 23011 11696 23069 11697
rect 23011 11656 23020 11696
rect 23060 11656 23069 11696
rect 23011 11655 23069 11656
rect 24355 11696 24413 11697
rect 24355 11656 24364 11696
rect 24404 11656 24413 11696
rect 25899 11696 25941 11705
rect 24355 11655 24413 11656
rect 25792 11685 25850 11686
rect 25792 11645 25801 11685
rect 25841 11645 25850 11685
rect 25899 11656 25900 11696
rect 25940 11656 25941 11696
rect 25899 11647 25941 11656
rect 26091 11696 26133 11705
rect 26091 11656 26092 11696
rect 26132 11656 26133 11696
rect 26091 11647 26133 11656
rect 26187 11696 26229 11705
rect 26187 11656 26188 11696
rect 26228 11656 26229 11696
rect 26187 11647 26229 11656
rect 26283 11696 26325 11705
rect 26283 11656 26284 11696
rect 26324 11656 26325 11696
rect 26283 11647 26325 11656
rect 26379 11696 26421 11705
rect 26379 11656 26380 11696
rect 26420 11656 26421 11696
rect 26379 11647 26421 11656
rect 26571 11696 26613 11705
rect 26571 11656 26572 11696
rect 26612 11656 26613 11696
rect 26571 11647 26613 11656
rect 26667 11696 26709 11705
rect 26667 11656 26668 11696
rect 26708 11656 26709 11696
rect 26667 11647 26709 11656
rect 26763 11696 26805 11705
rect 26763 11656 26764 11696
rect 26804 11656 26805 11696
rect 26763 11647 26805 11656
rect 26859 11696 26901 11705
rect 26859 11656 26860 11696
rect 26900 11656 26901 11696
rect 26859 11647 26901 11656
rect 27051 11696 27093 11705
rect 27051 11656 27052 11696
rect 27092 11656 27093 11696
rect 27051 11647 27093 11656
rect 27147 11696 27189 11705
rect 27147 11656 27148 11696
rect 27188 11656 27189 11696
rect 27147 11647 27189 11656
rect 27243 11696 27285 11705
rect 27243 11656 27244 11696
rect 27284 11656 27285 11696
rect 27243 11647 27285 11656
rect 27339 11696 27381 11705
rect 27339 11656 27340 11696
rect 27380 11656 27381 11696
rect 27339 11647 27381 11656
rect 28971 11696 29013 11705
rect 28971 11656 28972 11696
rect 29012 11656 29013 11696
rect 28971 11647 29013 11656
rect 29067 11696 29109 11705
rect 29067 11656 29068 11696
rect 29108 11656 29109 11696
rect 29067 11647 29109 11656
rect 29163 11696 29205 11705
rect 29163 11656 29164 11696
rect 29204 11656 29205 11696
rect 29163 11647 29205 11656
rect 29259 11696 29301 11705
rect 29259 11656 29260 11696
rect 29300 11656 29301 11696
rect 29259 11647 29301 11656
rect 29643 11696 29685 11705
rect 29643 11656 29644 11696
rect 29684 11656 29685 11696
rect 29643 11647 29685 11656
rect 29739 11696 29781 11705
rect 29739 11656 29740 11696
rect 29780 11656 29781 11696
rect 29739 11647 29781 11656
rect 30123 11696 30165 11705
rect 30123 11656 30124 11696
rect 30164 11656 30165 11696
rect 30123 11647 30165 11656
rect 30219 11696 30261 11705
rect 30219 11656 30220 11696
rect 30260 11656 30261 11696
rect 30219 11647 30261 11656
rect 30403 11696 30461 11697
rect 30403 11656 30412 11696
rect 30452 11656 30461 11696
rect 30403 11655 30461 11656
rect 31363 11696 31421 11697
rect 31363 11656 31372 11696
rect 31412 11656 31421 11696
rect 31363 11655 31421 11656
rect 32323 11696 32381 11697
rect 32323 11656 32332 11696
rect 32372 11656 32381 11696
rect 32323 11655 32381 11656
rect 32523 11696 32565 11705
rect 32523 11656 32524 11696
rect 32564 11656 32565 11696
rect 32523 11647 32565 11656
rect 32715 11696 32757 11705
rect 32715 11656 32716 11696
rect 32756 11656 32757 11696
rect 32715 11647 32757 11656
rect 32907 11696 32949 11705
rect 32907 11656 32908 11696
rect 32948 11656 32949 11696
rect 32907 11647 32949 11656
rect 33195 11696 33237 11705
rect 33195 11656 33196 11696
rect 33236 11656 33237 11696
rect 33195 11647 33237 11656
rect 33675 11696 33717 11705
rect 33675 11656 33676 11696
rect 33716 11656 33717 11696
rect 33675 11647 33717 11656
rect 33763 11696 33821 11697
rect 33763 11656 33772 11696
rect 33812 11656 33821 11696
rect 33763 11655 33821 11656
rect 33963 11696 34005 11705
rect 33963 11656 33964 11696
rect 34004 11656 34005 11696
rect 33963 11647 34005 11656
rect 34251 11696 34293 11705
rect 34251 11656 34252 11696
rect 34292 11656 34293 11696
rect 34251 11647 34293 11656
rect 34819 11696 34877 11697
rect 34819 11656 34828 11696
rect 34868 11656 34877 11696
rect 36067 11696 36125 11697
rect 34819 11655 34877 11656
rect 35211 11654 35253 11663
rect 36067 11656 36076 11696
rect 36116 11656 36125 11696
rect 36067 11655 36125 11656
rect 36259 11696 36317 11697
rect 36259 11656 36268 11696
rect 36308 11656 36317 11696
rect 36259 11655 36317 11656
rect 36939 11696 36981 11705
rect 36939 11656 36940 11696
rect 36980 11656 36981 11696
rect 25792 11644 25850 11645
rect 15819 11612 15861 11621
rect 15819 11572 15820 11612
rect 15860 11572 15861 11612
rect 35211 11614 35212 11654
rect 35252 11614 35253 11654
rect 36939 11647 36981 11656
rect 37131 11696 37173 11705
rect 37131 11656 37132 11696
rect 37172 11656 37173 11696
rect 37131 11647 37173 11656
rect 37507 11696 37565 11697
rect 37507 11656 37516 11696
rect 37556 11656 37565 11696
rect 37507 11655 37565 11656
rect 38371 11696 38429 11697
rect 38371 11656 38380 11696
rect 38420 11656 38429 11696
rect 38371 11655 38429 11656
rect 39531 11696 39573 11705
rect 39531 11656 39532 11696
rect 39572 11656 39573 11696
rect 39531 11647 39573 11656
rect 35211 11605 35253 11614
rect 15819 11563 15861 11572
rect 643 11528 701 11529
rect 643 11488 652 11528
rect 692 11488 701 11528
rect 643 11487 701 11488
rect 12451 11528 12509 11529
rect 12451 11488 12460 11528
rect 12500 11488 12509 11528
rect 12451 11487 12509 11488
rect 13507 11528 13565 11529
rect 13507 11488 13516 11528
rect 13556 11488 13565 11528
rect 13507 11487 13565 11488
rect 16099 11528 16157 11529
rect 16099 11488 16108 11528
rect 16148 11488 16157 11528
rect 16099 11487 16157 11488
rect 16867 11528 16925 11529
rect 16867 11488 16876 11528
rect 16916 11488 16925 11528
rect 16867 11487 16925 11488
rect 19843 11528 19901 11529
rect 19843 11488 19852 11528
rect 19892 11488 19901 11528
rect 19843 11487 19901 11488
rect 24163 11528 24221 11529
rect 24163 11488 24172 11528
rect 24212 11488 24221 11528
rect 24163 11487 24221 11488
rect 25027 11528 25085 11529
rect 25027 11488 25036 11528
rect 25076 11488 25085 11528
rect 25027 11487 25085 11488
rect 29443 11528 29501 11529
rect 29443 11488 29452 11528
rect 29492 11488 29501 11528
rect 29443 11487 29501 11488
rect 29923 11528 29981 11529
rect 29923 11488 29932 11528
rect 29972 11488 29981 11528
rect 29923 11487 29981 11488
rect 32235 11528 32277 11537
rect 32235 11488 32236 11528
rect 32276 11488 32277 11528
rect 32235 11479 32277 11488
rect 33675 11528 33717 11537
rect 33675 11488 33676 11528
rect 33716 11488 33717 11528
rect 33675 11479 33717 11488
rect 35395 11528 35453 11529
rect 35395 11488 35404 11528
rect 35444 11488 35453 11528
rect 35395 11487 35453 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 16299 11196 16341 11205
rect 643 11192 701 11193
rect 643 11152 652 11192
rect 692 11152 701 11192
rect 643 11151 701 11152
rect 16299 11156 16300 11196
rect 16340 11156 16341 11196
rect 16299 11147 16341 11156
rect 17251 11192 17309 11193
rect 17251 11152 17260 11192
rect 17300 11152 17309 11192
rect 17251 11151 17309 11152
rect 25707 11192 25749 11201
rect 25707 11152 25708 11192
rect 25748 11152 25749 11192
rect 25707 11143 25749 11152
rect 25987 11192 26045 11193
rect 25987 11152 25996 11192
rect 26036 11152 26045 11192
rect 25987 11151 26045 11152
rect 28779 11192 28821 11201
rect 28779 11152 28780 11192
rect 28820 11152 28821 11192
rect 28779 11143 28821 11152
rect 29347 11192 29405 11193
rect 29347 11152 29356 11192
rect 29396 11152 29405 11192
rect 29347 11151 29405 11152
rect 30019 11192 30077 11193
rect 30019 11152 30028 11192
rect 30068 11152 30077 11192
rect 30019 11151 30077 11152
rect 31459 11192 31517 11193
rect 31459 11152 31468 11192
rect 31508 11152 31517 11192
rect 31459 11151 31517 11152
rect 34443 11192 34485 11201
rect 34443 11152 34444 11192
rect 34484 11152 34485 11192
rect 34443 11143 34485 11152
rect 9675 11108 9717 11117
rect 9675 11068 9676 11108
rect 9716 11068 9717 11108
rect 9675 11059 9717 11068
rect 27339 11108 27381 11117
rect 27339 11068 27340 11108
rect 27380 11068 27381 11108
rect 27339 11059 27381 11068
rect 26851 11045 26909 11046
rect 8419 11024 8477 11025
rect 8419 10984 8428 11024
rect 8468 10984 8477 11024
rect 8419 10983 8477 10984
rect 9283 11024 9341 11025
rect 9283 10984 9292 11024
rect 9332 10984 9341 11024
rect 9283 10983 9341 10984
rect 10051 11024 10109 11025
rect 10051 10984 10060 11024
rect 10100 10984 10109 11024
rect 10051 10983 10109 10984
rect 10155 11024 10197 11033
rect 10155 10984 10156 11024
rect 10196 10984 10197 11024
rect 10155 10975 10197 10984
rect 10347 11024 10389 11033
rect 10347 10984 10348 11024
rect 10388 10984 10389 11024
rect 10347 10975 10389 10984
rect 10531 11024 10589 11025
rect 10531 10984 10540 11024
rect 10580 10984 10589 11024
rect 10531 10983 10589 10984
rect 11403 11024 11445 11033
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11403 10975 11445 10984
rect 11499 11024 11541 11033
rect 11499 10984 11500 11024
rect 11540 10984 11541 11024
rect 11499 10975 11541 10984
rect 11595 11024 11637 11033
rect 11595 10984 11596 11024
rect 11636 10984 11637 11024
rect 11595 10975 11637 10984
rect 11691 11024 11733 11033
rect 11691 10984 11692 11024
rect 11732 10984 11733 11024
rect 11691 10975 11733 10984
rect 12451 11024 12509 11025
rect 12451 10984 12460 11024
rect 12500 10984 12509 11024
rect 12451 10983 12509 10984
rect 12643 11024 12701 11025
rect 12643 10984 12652 11024
rect 12692 10984 12701 11024
rect 12643 10983 12701 10984
rect 13891 11024 13949 11025
rect 13891 10984 13900 11024
rect 13940 10984 13949 11024
rect 13891 10983 13949 10984
rect 14859 11024 14901 11033
rect 14859 10984 14860 11024
rect 14900 10984 14901 11024
rect 14859 10975 14901 10984
rect 14947 11024 15005 11025
rect 14947 10984 14956 11024
rect 14996 10984 15005 11024
rect 14947 10983 15005 10984
rect 16195 11024 16253 11025
rect 16195 10984 16204 11024
rect 16244 10984 16253 11024
rect 16195 10983 16253 10984
rect 16958 11024 17016 11025
rect 16958 10984 16967 11024
rect 17007 10984 17016 11024
rect 16958 10983 17016 10984
rect 17067 11024 17109 11033
rect 17067 10984 17068 11024
rect 17108 10984 17109 11024
rect 16099 10982 16157 10983
rect 16099 10942 16108 10982
rect 16148 10942 16157 10982
rect 17067 10975 17109 10984
rect 17163 11024 17205 11033
rect 17163 10984 17164 11024
rect 17204 10984 17205 11024
rect 17163 10975 17205 10984
rect 17347 11024 17405 11025
rect 17347 10984 17356 11024
rect 17396 10984 17405 11024
rect 17347 10983 17405 10984
rect 17443 11024 17501 11025
rect 17443 10984 17452 11024
rect 17492 10984 17501 11024
rect 17443 10983 17501 10984
rect 17635 11024 17693 11025
rect 17635 10984 17644 11024
rect 17684 10984 17693 11024
rect 17635 10983 17693 10984
rect 18507 11024 18549 11033
rect 18507 10984 18508 11024
rect 18548 10984 18549 11024
rect 18507 10975 18549 10984
rect 18883 11024 18941 11025
rect 18883 10984 18892 11024
rect 18932 10984 18941 11024
rect 18883 10983 18941 10984
rect 18979 11024 19037 11025
rect 18979 10984 18988 11024
rect 19028 10984 19037 11024
rect 18979 10983 19037 10984
rect 19179 11024 19221 11033
rect 19179 10984 19180 11024
rect 19220 10984 19221 11024
rect 19179 10975 19221 10984
rect 19275 11024 19317 11033
rect 19275 10984 19276 11024
rect 19316 10984 19317 11024
rect 19275 10975 19317 10984
rect 19368 11024 19426 11025
rect 19368 10984 19377 11024
rect 19417 10984 19426 11024
rect 19368 10983 19426 10984
rect 19843 11024 19901 11025
rect 19843 10984 19852 11024
rect 19892 10984 19901 11024
rect 19843 10983 19901 10984
rect 20803 11024 20861 11025
rect 20803 10984 20812 11024
rect 20852 10984 20861 11024
rect 20803 10983 20861 10984
rect 21667 11024 21725 11025
rect 21667 10984 21676 11024
rect 21716 10984 21725 11024
rect 21667 10983 21725 10984
rect 21867 11024 21909 11033
rect 21867 10984 21868 11024
rect 21908 10984 21909 11024
rect 21867 10975 21909 10984
rect 22059 11024 22101 11033
rect 22059 10984 22060 11024
rect 22100 10984 22101 11024
rect 22059 10975 22101 10984
rect 22147 11024 22205 11025
rect 22147 10984 22156 11024
rect 22196 10984 22205 11024
rect 22147 10983 22205 10984
rect 23683 11024 23741 11025
rect 23683 10984 23692 11024
rect 23732 10984 23741 11024
rect 23683 10983 23741 10984
rect 23787 11024 23829 11033
rect 23787 10984 23788 11024
rect 23828 10984 23829 11024
rect 23787 10975 23829 10984
rect 24163 11024 24221 11025
rect 24163 10984 24172 11024
rect 24212 10984 24221 11024
rect 24163 10983 24221 10984
rect 25035 11024 25077 11033
rect 25035 10984 25036 11024
rect 25076 10984 25077 11024
rect 25035 10975 25077 10984
rect 25795 11024 25853 11025
rect 25795 10984 25804 11024
rect 25844 10984 25853 11024
rect 25795 10983 25853 10984
rect 26091 11024 26133 11033
rect 26091 10984 26092 11024
rect 26132 10984 26133 11024
rect 26091 10975 26133 10984
rect 26187 11024 26229 11033
rect 26187 10984 26188 11024
rect 26228 10984 26229 11024
rect 26187 10975 26229 10984
rect 26283 11024 26325 11033
rect 26283 10984 26284 11024
rect 26324 10984 26325 11024
rect 26283 10975 26325 10984
rect 26475 11024 26517 11033
rect 26475 10984 26476 11024
rect 26516 10984 26517 11024
rect 26475 10975 26517 10984
rect 26667 11024 26709 11033
rect 26667 10984 26668 11024
rect 26708 10984 26709 11024
rect 26851 11005 26860 11045
rect 26900 11005 26909 11045
rect 26851 11004 26909 11005
rect 27051 11024 27093 11033
rect 26667 10975 26709 10984
rect 27051 10984 27052 11024
rect 27092 10984 27093 11024
rect 27051 10975 27093 10984
rect 27243 11024 27285 11033
rect 27243 10984 27244 11024
rect 27284 10984 27285 11024
rect 27243 10975 27285 10984
rect 27435 11024 27477 11033
rect 27435 10984 27436 11024
rect 27476 10984 27477 11024
rect 27435 10975 27477 10984
rect 28683 11024 28725 11033
rect 28683 10984 28684 11024
rect 28724 10984 28725 11024
rect 28683 10975 28725 10984
rect 28875 11024 28917 11033
rect 28875 10984 28876 11024
rect 28916 10984 28917 11024
rect 28875 10975 28917 10984
rect 29067 11024 29109 11033
rect 29067 10984 29068 11024
rect 29108 10984 29109 11024
rect 29067 10975 29109 10984
rect 29163 11024 29205 11033
rect 29163 10984 29164 11024
rect 29204 10984 29205 11024
rect 29163 10975 29205 10984
rect 29547 11024 29589 11033
rect 29547 10984 29548 11024
rect 29588 10984 29589 11024
rect 29251 10982 29309 10983
rect 16099 10941 16157 10942
rect 29251 10942 29260 10982
rect 29300 10942 29309 10982
rect 29547 10975 29589 10984
rect 29739 11024 29781 11033
rect 29739 10984 29740 11024
rect 29780 10984 29781 11024
rect 29635 10982 29693 10983
rect 29251 10941 29309 10942
rect 29635 10942 29644 10982
rect 29684 10942 29693 10982
rect 29739 10975 29781 10984
rect 29835 11024 29877 11033
rect 29835 10984 29836 11024
rect 29876 10984 29877 11024
rect 29835 10975 29877 10984
rect 30219 11024 30261 11033
rect 30219 10984 30220 11024
rect 30260 10984 30261 11024
rect 30219 10975 30261 10984
rect 30315 11024 30357 11033
rect 30315 10984 30316 11024
rect 30356 10984 30357 11024
rect 30315 10975 30357 10984
rect 30507 11024 30549 11033
rect 30507 10984 30508 11024
rect 30548 10984 30549 11024
rect 30507 10975 30549 10984
rect 30691 11024 30749 11025
rect 30691 10984 30700 11024
rect 30740 10984 30749 11024
rect 30691 10983 30749 10984
rect 31171 11024 31229 11025
rect 31171 10984 31180 11024
rect 31220 10984 31229 11024
rect 31171 10983 31229 10984
rect 31267 11024 31325 11025
rect 31267 10984 31276 11024
rect 31316 10984 31325 11024
rect 31267 10983 31325 10984
rect 31467 11024 31509 11033
rect 31467 10984 31468 11024
rect 31508 10984 31509 11024
rect 31467 10975 31509 10984
rect 31563 11024 31605 11033
rect 31563 10984 31564 11024
rect 31604 10984 31605 11024
rect 31563 10975 31605 10984
rect 31656 11024 31714 11025
rect 31656 10984 31665 11024
rect 31705 10984 31714 11024
rect 31656 10983 31714 10984
rect 32419 11024 32477 11025
rect 32419 10984 32428 11024
rect 32468 10984 32477 11024
rect 32419 10983 32477 10984
rect 32707 11024 32765 11025
rect 32707 10984 32716 11024
rect 32756 10984 32765 11024
rect 32707 10983 32765 10984
rect 33099 11024 33141 11033
rect 33099 10984 33100 11024
rect 33140 10984 33141 11024
rect 33099 10975 33141 10984
rect 34339 11024 34397 11025
rect 34339 10984 34348 11024
rect 34388 10984 34397 11024
rect 34339 10983 34397 10984
rect 34731 11024 34773 11033
rect 34731 10984 34732 11024
rect 34772 10984 34773 11024
rect 34731 10975 34773 10984
rect 34827 11024 34869 11033
rect 34827 10984 34828 11024
rect 34868 10984 34869 11024
rect 34827 10975 34869 10984
rect 34923 11024 34965 11033
rect 34923 10984 34924 11024
rect 34964 10984 34965 11024
rect 34923 10975 34965 10984
rect 35019 11024 35061 11033
rect 35019 10984 35020 11024
rect 35060 10984 35061 11024
rect 35019 10975 35061 10984
rect 35403 11024 35445 11033
rect 35403 10984 35404 11024
rect 35444 10984 35445 11024
rect 35403 10975 35445 10984
rect 35779 11024 35837 11025
rect 35779 10984 35788 11024
rect 35828 10984 35837 11024
rect 35779 10983 35837 10984
rect 36643 11024 36701 11025
rect 36643 10984 36652 11024
rect 36692 10984 36701 11024
rect 36643 10983 36701 10984
rect 37803 11024 37845 11033
rect 37803 10984 37804 11024
rect 37844 10984 37845 11024
rect 37803 10975 37845 10984
rect 38091 11024 38133 11033
rect 38091 10984 38092 11024
rect 38132 10984 38133 11024
rect 38091 10975 38133 10984
rect 38755 11024 38813 11025
rect 38755 10984 38764 11024
rect 38804 10984 38813 11024
rect 38755 10983 38813 10984
rect 29635 10941 29693 10942
rect 15235 10940 15293 10941
rect 15235 10900 15244 10940
rect 15284 10900 15293 10940
rect 15235 10899 15293 10900
rect 15619 10940 15677 10941
rect 15619 10900 15628 10940
rect 15668 10900 15677 10940
rect 15619 10899 15677 10900
rect 23299 10940 23357 10941
rect 23299 10900 23308 10940
rect 23348 10900 23357 10940
rect 23299 10899 23357 10900
rect 30603 10940 30645 10949
rect 30603 10900 30604 10940
rect 30644 10900 30645 10940
rect 30603 10891 30645 10900
rect 32811 10940 32853 10949
rect 32811 10900 32812 10940
rect 32852 10900 32853 10940
rect 32811 10891 32853 10900
rect 33003 10940 33045 10949
rect 33003 10900 33004 10940
rect 33044 10900 33045 10940
rect 33003 10891 33045 10900
rect 10347 10856 10389 10865
rect 10347 10816 10348 10856
rect 10388 10816 10389 10856
rect 10347 10807 10389 10816
rect 11883 10856 11925 10865
rect 11883 10816 11884 10856
rect 11924 10816 11925 10856
rect 11883 10807 11925 10816
rect 13227 10856 13269 10865
rect 13227 10816 13228 10856
rect 13268 10816 13269 10856
rect 13227 10807 13269 10816
rect 13611 10856 13653 10865
rect 13611 10816 13612 10856
rect 13652 10816 13653 10856
rect 13611 10807 13653 10816
rect 18315 10856 18357 10865
rect 18315 10816 18316 10856
rect 18356 10816 18357 10856
rect 18315 10807 18357 10816
rect 22347 10856 22389 10865
rect 22347 10816 22348 10856
rect 22388 10816 22389 10856
rect 22347 10807 22389 10816
rect 26475 10856 26517 10865
rect 26475 10816 26476 10856
rect 26516 10816 26517 10856
rect 26475 10807 26517 10816
rect 32523 10856 32565 10865
rect 32523 10816 32524 10856
rect 32564 10816 32565 10856
rect 32523 10807 32565 10816
rect 32907 10856 32949 10865
rect 32907 10816 32908 10856
rect 32948 10816 32949 10856
rect 32907 10807 32949 10816
rect 7267 10772 7325 10773
rect 7267 10732 7276 10772
rect 7316 10732 7325 10772
rect 7267 10731 7325 10732
rect 11203 10772 11261 10773
rect 11203 10732 11212 10772
rect 11252 10732 11261 10772
rect 11203 10731 11261 10732
rect 15435 10772 15477 10781
rect 15435 10732 15436 10772
rect 15476 10732 15477 10772
rect 15435 10723 15477 10732
rect 15819 10772 15861 10781
rect 15819 10732 15820 10772
rect 15860 10732 15861 10772
rect 15819 10723 15861 10732
rect 18891 10772 18933 10781
rect 18891 10732 18892 10772
rect 18932 10732 18933 10772
rect 18891 10723 18933 10732
rect 20139 10772 20181 10781
rect 20139 10732 20140 10772
rect 20180 10732 20181 10772
rect 20139 10723 20181 10732
rect 20995 10772 21053 10773
rect 20995 10732 21004 10772
rect 21044 10732 21053 10772
rect 20995 10731 21053 10732
rect 21867 10772 21909 10781
rect 21867 10732 21868 10772
rect 21908 10732 21909 10772
rect 21867 10723 21909 10732
rect 23499 10772 23541 10781
rect 23499 10732 23500 10772
rect 23540 10732 23541 10772
rect 23499 10723 23541 10732
rect 24459 10772 24501 10781
rect 24459 10732 24460 10772
rect 24500 10732 24501 10772
rect 24459 10723 24501 10732
rect 26955 10772 26997 10781
rect 26955 10732 26956 10772
rect 26996 10732 26997 10772
rect 26955 10723 26997 10732
rect 35203 10772 35261 10773
rect 35203 10732 35212 10772
rect 35252 10732 35261 10772
rect 35203 10731 35261 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 13515 10436 13557 10445
rect 13515 10396 13516 10436
rect 13556 10396 13557 10436
rect 13515 10387 13557 10396
rect 26667 10436 26709 10445
rect 26667 10396 26668 10436
rect 26708 10396 26709 10436
rect 26667 10387 26709 10396
rect 29355 10436 29397 10445
rect 29355 10396 29356 10436
rect 29396 10396 29397 10436
rect 29355 10387 29397 10396
rect 30987 10436 31029 10445
rect 30987 10396 30988 10436
rect 31028 10396 31029 10436
rect 30987 10387 31029 10396
rect 31275 10436 31317 10445
rect 31275 10396 31276 10436
rect 31316 10396 31317 10436
rect 31275 10387 31317 10396
rect 32715 10436 32757 10445
rect 32715 10396 32716 10436
rect 32756 10396 32757 10436
rect 32715 10387 32757 10396
rect 34627 10436 34685 10437
rect 34627 10396 34636 10436
rect 34676 10396 34685 10436
rect 34627 10395 34685 10396
rect 35019 10436 35061 10445
rect 35019 10396 35020 10436
rect 35060 10396 35061 10436
rect 35019 10387 35061 10396
rect 35307 10436 35349 10445
rect 35307 10396 35308 10436
rect 35348 10396 35349 10436
rect 35307 10387 35349 10396
rect 6027 10352 6069 10361
rect 6027 10312 6028 10352
rect 6068 10312 6069 10352
rect 6027 10303 6069 10312
rect 6795 10352 6837 10361
rect 6795 10312 6796 10352
rect 6836 10312 6837 10352
rect 6795 10303 6837 10312
rect 9003 10352 9045 10361
rect 9003 10312 9004 10352
rect 9044 10312 9045 10352
rect 9003 10303 9045 10312
rect 9955 10352 10013 10353
rect 9955 10312 9964 10352
rect 10004 10312 10013 10352
rect 9955 10311 10013 10312
rect 23107 10352 23165 10353
rect 23107 10312 23116 10352
rect 23156 10312 23165 10352
rect 23107 10311 23165 10312
rect 29155 10352 29213 10353
rect 29155 10312 29164 10352
rect 29204 10312 29213 10352
rect 29155 10311 29213 10312
rect 20331 10268 20373 10277
rect 20331 10228 20332 10268
rect 20372 10228 20373 10268
rect 20331 10219 20373 10228
rect 25123 10268 25181 10269
rect 25123 10228 25132 10268
rect 25172 10228 25181 10268
rect 25123 10227 25181 10228
rect 30994 10197 31036 10206
rect 7651 10184 7709 10185
rect 7651 10144 7660 10184
rect 7700 10144 7709 10184
rect 7651 10143 7709 10144
rect 7843 10184 7901 10185
rect 7843 10144 7852 10184
rect 7892 10144 7901 10184
rect 7843 10143 7901 10144
rect 9667 10184 9725 10185
rect 9667 10144 9676 10184
rect 9716 10144 9725 10184
rect 9667 10143 9725 10144
rect 11107 10184 11165 10185
rect 11107 10144 11116 10184
rect 11156 10144 11165 10184
rect 11107 10143 11165 10144
rect 11971 10184 12029 10185
rect 11971 10144 11980 10184
rect 12020 10144 12029 10184
rect 11971 10143 12029 10144
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12547 10184 12605 10185
rect 12547 10144 12556 10184
rect 12596 10144 12605 10184
rect 12547 10143 12605 10144
rect 13227 10184 13269 10193
rect 13227 10144 13228 10184
rect 13268 10144 13269 10184
rect 13227 10135 13269 10144
rect 13411 10184 13469 10185
rect 13411 10144 13420 10184
rect 13460 10144 13469 10184
rect 13411 10143 13469 10144
rect 14659 10184 14717 10185
rect 14659 10144 14668 10184
rect 14708 10144 14717 10184
rect 14659 10143 14717 10144
rect 15619 10184 15677 10185
rect 15619 10144 15628 10184
rect 15668 10144 15677 10184
rect 15619 10143 15677 10144
rect 16099 10184 16157 10185
rect 16099 10144 16108 10184
rect 16148 10144 16157 10184
rect 16099 10143 16157 10144
rect 16203 10184 16245 10193
rect 16203 10144 16204 10184
rect 16244 10144 16245 10184
rect 16203 10135 16245 10144
rect 16387 10184 16445 10185
rect 16387 10144 16396 10184
rect 16436 10144 16445 10184
rect 16387 10143 16445 10144
rect 16587 10184 16629 10193
rect 16587 10144 16588 10184
rect 16628 10144 16629 10184
rect 16587 10135 16629 10144
rect 16779 10184 16821 10193
rect 16779 10144 16780 10184
rect 16820 10144 16821 10184
rect 16779 10135 16821 10144
rect 16867 10184 16925 10185
rect 16867 10144 16876 10184
rect 16916 10144 16925 10184
rect 16867 10143 16925 10144
rect 17059 10184 17117 10185
rect 17059 10144 17068 10184
rect 17108 10144 17117 10184
rect 17059 10143 17117 10144
rect 18307 10184 18365 10185
rect 18307 10144 18316 10184
rect 18356 10144 18365 10184
rect 18307 10143 18365 10144
rect 19171 10184 19229 10185
rect 19171 10144 19180 10184
rect 19220 10144 19229 10184
rect 19171 10143 19229 10144
rect 20715 10184 20757 10193
rect 20715 10144 20716 10184
rect 20756 10144 20757 10184
rect 20715 10135 20757 10144
rect 21091 10184 21149 10185
rect 21091 10144 21100 10184
rect 21140 10144 21149 10184
rect 21091 10143 21149 10144
rect 21955 10184 22013 10185
rect 21955 10144 21964 10184
rect 22004 10144 22013 10184
rect 21955 10143 22013 10144
rect 23299 10184 23357 10185
rect 23299 10144 23308 10184
rect 23348 10144 23357 10184
rect 23299 10143 23357 10144
rect 24363 10184 24405 10193
rect 24363 10144 24364 10184
rect 24404 10144 24405 10184
rect 24363 10135 24405 10144
rect 24459 10184 24501 10193
rect 24459 10144 24460 10184
rect 24500 10144 24501 10184
rect 24459 10135 24501 10144
rect 24651 10184 24693 10193
rect 24651 10144 24652 10184
rect 24692 10144 24693 10184
rect 24651 10135 24693 10144
rect 24747 10184 24789 10193
rect 24747 10144 24748 10184
rect 24788 10144 24789 10184
rect 24747 10135 24789 10144
rect 24939 10184 24981 10193
rect 24939 10144 24940 10184
rect 24980 10144 24981 10184
rect 24939 10135 24981 10144
rect 26187 10184 26229 10193
rect 26187 10144 26188 10184
rect 26228 10144 26229 10184
rect 26187 10135 26229 10144
rect 26283 10184 26325 10193
rect 26283 10144 26284 10184
rect 26324 10144 26325 10184
rect 26283 10135 26325 10144
rect 26379 10184 26421 10193
rect 26379 10144 26380 10184
rect 26420 10144 26421 10184
rect 26379 10135 26421 10144
rect 26475 10184 26517 10193
rect 26475 10144 26476 10184
rect 26516 10144 26517 10184
rect 26475 10135 26517 10144
rect 26659 10184 26717 10185
rect 26659 10144 26668 10184
rect 26708 10144 26717 10184
rect 26659 10143 26717 10144
rect 26755 10184 26813 10185
rect 26755 10144 26764 10184
rect 26804 10144 26813 10184
rect 26755 10143 26813 10144
rect 26955 10184 26997 10193
rect 26955 10144 26956 10184
rect 26996 10144 26997 10184
rect 26955 10135 26997 10144
rect 27051 10184 27093 10193
rect 27051 10144 27052 10184
rect 27092 10144 27093 10184
rect 27051 10135 27093 10144
rect 27144 10184 27202 10185
rect 27144 10144 27153 10184
rect 27193 10144 27202 10184
rect 27144 10143 27202 10144
rect 28875 10184 28917 10193
rect 28875 10144 28876 10184
rect 28916 10144 28917 10184
rect 28875 10135 28917 10144
rect 29067 10184 29109 10193
rect 29067 10144 29068 10184
rect 29108 10144 29109 10184
rect 29067 10135 29109 10144
rect 29163 10184 29205 10193
rect 29163 10144 29164 10184
rect 29204 10144 29205 10184
rect 29163 10135 29205 10144
rect 29347 10184 29405 10185
rect 29347 10144 29356 10184
rect 29396 10144 29405 10184
rect 29347 10143 29405 10144
rect 29443 10184 29501 10185
rect 29443 10144 29452 10184
rect 29492 10144 29501 10184
rect 29443 10143 29501 10144
rect 29643 10184 29685 10193
rect 29643 10144 29644 10184
rect 29684 10144 29685 10184
rect 29832 10184 29890 10185
rect 29643 10135 29685 10144
rect 29739 10142 29781 10151
rect 29832 10144 29841 10184
rect 29881 10144 29890 10184
rect 29832 10143 29890 10144
rect 30123 10184 30165 10193
rect 30123 10144 30124 10184
rect 30164 10144 30165 10184
rect 6987 10100 7029 10109
rect 6987 10060 6988 10100
rect 7028 10060 7029 10100
rect 6987 10051 7029 10060
rect 16683 10100 16725 10109
rect 16683 10060 16684 10100
rect 16724 10060 16725 10100
rect 16683 10051 16725 10060
rect 17739 10100 17781 10109
rect 17739 10060 17740 10100
rect 17780 10060 17781 10100
rect 17739 10051 17781 10060
rect 17931 10100 17973 10109
rect 17931 10060 17932 10100
rect 17972 10060 17973 10100
rect 17931 10051 17973 10060
rect 23979 10100 24021 10109
rect 23979 10060 23980 10100
rect 24020 10060 24021 10100
rect 23979 10051 24021 10060
rect 24843 10100 24885 10109
rect 24843 10060 24844 10100
rect 24884 10060 24885 10100
rect 29739 10102 29740 10142
rect 29780 10102 29781 10142
rect 30123 10135 30165 10144
rect 30411 10184 30453 10193
rect 30411 10144 30412 10184
rect 30452 10144 30453 10184
rect 30411 10135 30453 10144
rect 30795 10184 30837 10193
rect 30795 10144 30796 10184
rect 30836 10144 30837 10184
rect 30994 10157 30995 10197
rect 31035 10157 31036 10197
rect 30994 10148 31036 10157
rect 31179 10184 31221 10193
rect 30795 10135 30837 10144
rect 31179 10144 31180 10184
rect 31220 10144 31221 10184
rect 31179 10135 31221 10144
rect 31363 10184 31421 10185
rect 31363 10144 31372 10184
rect 31412 10144 31421 10184
rect 31363 10143 31421 10144
rect 32139 10184 32181 10193
rect 32139 10144 32140 10184
rect 32180 10144 32181 10184
rect 32139 10135 32181 10144
rect 32235 10184 32277 10193
rect 32235 10144 32236 10184
rect 32276 10144 32277 10184
rect 32235 10135 32277 10144
rect 32331 10184 32373 10193
rect 32331 10144 32332 10184
rect 32372 10144 32373 10184
rect 32331 10135 32373 10144
rect 32427 10184 32469 10193
rect 32427 10144 32428 10184
rect 32468 10144 32469 10184
rect 32427 10135 32469 10144
rect 32619 10184 32661 10193
rect 32619 10144 32620 10184
rect 32660 10144 32661 10184
rect 32619 10135 32661 10144
rect 32803 10184 32861 10185
rect 32803 10144 32812 10184
rect 32852 10144 32861 10184
rect 32803 10143 32861 10144
rect 33091 10184 33149 10185
rect 33091 10144 33100 10184
rect 33140 10144 33149 10184
rect 33091 10143 33149 10144
rect 34435 10184 34493 10185
rect 34435 10144 34444 10184
rect 34484 10144 34493 10184
rect 34435 10143 34493 10144
rect 34819 10184 34877 10185
rect 34819 10144 34828 10184
rect 34868 10144 34877 10184
rect 34819 10143 34877 10144
rect 35019 10184 35061 10193
rect 35019 10144 35020 10184
rect 35060 10144 35061 10184
rect 35019 10135 35061 10144
rect 35107 10184 35165 10185
rect 35107 10144 35116 10184
rect 35156 10144 35165 10184
rect 35107 10143 35165 10144
rect 35299 10184 35357 10185
rect 35299 10144 35308 10184
rect 35348 10144 35357 10184
rect 35299 10143 35357 10144
rect 35499 10184 35541 10193
rect 35499 10144 35500 10184
rect 35540 10144 35541 10184
rect 35499 10135 35541 10144
rect 35587 10184 35645 10185
rect 35587 10144 35596 10184
rect 35636 10144 35645 10184
rect 35587 10143 35645 10144
rect 35779 10184 35837 10185
rect 35779 10144 35788 10184
rect 35828 10144 35837 10184
rect 35779 10143 35837 10144
rect 36067 10184 36125 10185
rect 36067 10144 36076 10184
rect 36116 10144 36125 10184
rect 36067 10143 36125 10144
rect 36547 10184 36605 10185
rect 36547 10144 36556 10184
rect 36596 10144 36605 10184
rect 36547 10143 36605 10144
rect 37227 10184 37269 10193
rect 37227 10144 37228 10184
rect 37268 10144 37269 10184
rect 37227 10135 37269 10144
rect 37419 10184 37461 10193
rect 37419 10144 37420 10184
rect 37460 10144 37461 10184
rect 37419 10135 37461 10144
rect 37795 10184 37853 10185
rect 37795 10144 37804 10184
rect 37844 10144 37853 10184
rect 37795 10143 37853 10144
rect 38659 10184 38717 10185
rect 38659 10144 38668 10184
rect 38708 10144 38717 10184
rect 38659 10143 38717 10144
rect 39819 10184 39861 10193
rect 39819 10144 39820 10184
rect 39860 10144 39861 10184
rect 39819 10135 39861 10144
rect 29739 10093 29781 10102
rect 30315 10100 30357 10109
rect 24843 10051 24885 10060
rect 30315 10060 30316 10100
rect 30356 10060 30357 10100
rect 30315 10051 30357 10060
rect 33003 10100 33045 10109
rect 33003 10060 33004 10100
rect 33044 10060 33045 10100
rect 33003 10051 33045 10060
rect 36259 10100 36317 10101
rect 36259 10060 36268 10100
rect 36308 10060 36317 10100
rect 36259 10059 36317 10060
rect 643 10016 701 10017
rect 643 9976 652 10016
rect 692 9976 701 10016
rect 643 9975 701 9976
rect 8515 10016 8573 10017
rect 8515 9976 8524 10016
rect 8564 9976 8573 10016
rect 8515 9975 8573 9976
rect 16395 10016 16437 10025
rect 16395 9976 16396 10016
rect 16436 9976 16437 10016
rect 16395 9967 16437 9976
rect 24163 10016 24221 10017
rect 24163 9976 24172 10016
rect 24212 9976 24221 10016
rect 24163 9975 24221 9976
rect 25323 10016 25365 10025
rect 25323 9976 25324 10016
rect 25364 9976 25365 10016
rect 25323 9967 25365 9976
rect 34339 10016 34397 10017
rect 34339 9976 34348 10016
rect 34388 9976 34397 10016
rect 34339 9975 34397 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 643 9680 701 9681
rect 643 9640 652 9680
rect 692 9640 701 9680
rect 643 9639 701 9640
rect 9475 9680 9533 9681
rect 9475 9640 9484 9680
rect 9524 9640 9533 9680
rect 9475 9639 9533 9640
rect 10051 9680 10109 9681
rect 10051 9640 10060 9680
rect 10100 9640 10109 9680
rect 10051 9639 10109 9640
rect 11011 9680 11069 9681
rect 11011 9640 11020 9680
rect 11060 9640 11069 9680
rect 11011 9639 11069 9640
rect 11491 9680 11549 9681
rect 11491 9640 11500 9680
rect 11540 9640 11549 9680
rect 11491 9639 11549 9640
rect 13315 9680 13373 9681
rect 13315 9640 13324 9680
rect 13364 9640 13373 9680
rect 13315 9639 13373 9640
rect 27331 9680 27389 9681
rect 27331 9640 27340 9680
rect 27380 9640 27389 9680
rect 27331 9639 27389 9640
rect 27819 9680 27861 9689
rect 27819 9640 27820 9680
rect 27860 9640 27861 9680
rect 27819 9631 27861 9640
rect 28195 9680 28253 9681
rect 28195 9640 28204 9680
rect 28244 9640 28253 9680
rect 28195 9639 28253 9640
rect 29539 9680 29597 9681
rect 29539 9640 29548 9680
rect 29588 9640 29597 9680
rect 29539 9639 29597 9640
rect 30603 9680 30645 9689
rect 30603 9640 30604 9680
rect 30644 9640 30645 9680
rect 30603 9631 30645 9640
rect 32131 9680 32189 9681
rect 32131 9640 32140 9680
rect 32180 9640 32189 9680
rect 32131 9639 32189 9640
rect 33187 9680 33245 9681
rect 33187 9640 33196 9680
rect 33236 9640 33245 9680
rect 33187 9639 33245 9640
rect 35203 9680 35261 9681
rect 35203 9640 35212 9680
rect 35252 9640 35261 9680
rect 35203 9639 35261 9640
rect 35587 9680 35645 9681
rect 35587 9640 35596 9680
rect 35636 9640 35645 9680
rect 35587 9639 35645 9640
rect 35875 9680 35933 9681
rect 35875 9640 35884 9680
rect 35924 9640 35933 9680
rect 35875 9639 35933 9640
rect 38179 9680 38237 9681
rect 38179 9640 38188 9680
rect 38228 9640 38237 9680
rect 38179 9639 38237 9640
rect 5547 9596 5589 9605
rect 5547 9556 5548 9596
rect 5588 9556 5589 9596
rect 5547 9547 5589 9556
rect 13803 9596 13845 9605
rect 13803 9556 13804 9596
rect 13844 9556 13845 9596
rect 13803 9547 13845 9556
rect 24843 9596 24885 9605
rect 24843 9556 24844 9596
rect 24884 9556 24885 9596
rect 24843 9547 24885 9556
rect 15723 9533 15765 9542
rect 5923 9512 5981 9513
rect 5923 9472 5932 9512
rect 5972 9472 5981 9512
rect 5923 9471 5981 9472
rect 6787 9512 6845 9513
rect 6787 9472 6796 9512
rect 6836 9472 6845 9512
rect 6787 9471 6845 9472
rect 8139 9512 8181 9521
rect 8139 9472 8140 9512
rect 8180 9472 8181 9512
rect 8139 9463 8181 9472
rect 8227 9512 8285 9513
rect 8227 9472 8236 9512
rect 8276 9472 8285 9512
rect 8227 9471 8285 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 9091 9512 9149 9513
rect 9091 9472 9100 9512
rect 9140 9472 9149 9512
rect 9091 9471 9149 9472
rect 9283 9512 9341 9513
rect 9283 9472 9292 9512
rect 9332 9472 9341 9512
rect 9283 9471 9341 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9859 9512 9917 9513
rect 9859 9472 9868 9512
rect 9908 9472 9917 9512
rect 9859 9471 9917 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10155 9512 10197 9521
rect 10155 9472 10156 9512
rect 10196 9472 10197 9512
rect 10155 9463 10197 9472
rect 10339 9512 10397 9513
rect 10339 9472 10348 9512
rect 10388 9472 10397 9512
rect 10339 9471 10397 9472
rect 10443 9512 10485 9521
rect 10443 9472 10444 9512
rect 10484 9472 10485 9512
rect 10443 9463 10485 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11211 9512 11253 9521
rect 11211 9472 11212 9512
rect 11252 9472 11253 9512
rect 11211 9463 11253 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11595 9512 11637 9521
rect 11595 9472 11596 9512
rect 11636 9472 11637 9512
rect 11595 9463 11637 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 11787 9512 11829 9521
rect 11787 9472 11788 9512
rect 11828 9472 11829 9512
rect 11787 9463 11829 9472
rect 12643 9512 12701 9513
rect 12643 9472 12652 9512
rect 12692 9472 12701 9512
rect 12643 9471 12701 9472
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13123 9512 13181 9513
rect 13123 9472 13132 9512
rect 13172 9472 13181 9512
rect 13123 9471 13181 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13515 9512 13557 9521
rect 13515 9472 13516 9512
rect 13556 9472 13557 9512
rect 13515 9463 13557 9472
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13899 9512 13941 9521
rect 13899 9472 13900 9512
rect 13940 9472 13941 9512
rect 13899 9463 13941 9472
rect 13995 9512 14037 9521
rect 13995 9472 13996 9512
rect 14036 9472 14037 9512
rect 13995 9463 14037 9472
rect 14091 9512 14133 9521
rect 14091 9472 14092 9512
rect 14132 9472 14133 9512
rect 14091 9463 14133 9472
rect 14275 9512 14333 9513
rect 14275 9472 14284 9512
rect 14324 9472 14333 9512
rect 14275 9471 14333 9472
rect 14379 9512 14421 9521
rect 14379 9472 14380 9512
rect 14420 9472 14421 9512
rect 14379 9463 14421 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 14859 9512 14901 9521
rect 14859 9472 14860 9512
rect 14900 9472 14901 9512
rect 14859 9463 14901 9472
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15243 9512 15285 9521
rect 15243 9472 15244 9512
rect 15284 9472 15285 9512
rect 15243 9463 15285 9472
rect 15339 9512 15381 9521
rect 15339 9472 15340 9512
rect 15380 9472 15381 9512
rect 15339 9463 15381 9472
rect 15435 9512 15477 9521
rect 15435 9472 15436 9512
rect 15476 9472 15477 9512
rect 15435 9463 15477 9472
rect 15531 9512 15573 9521
rect 15531 9472 15532 9512
rect 15572 9472 15573 9512
rect 15723 9493 15724 9533
rect 15764 9493 15765 9533
rect 15723 9484 15765 9493
rect 15819 9512 15861 9521
rect 15531 9463 15573 9472
rect 15819 9472 15820 9512
rect 15860 9472 15861 9512
rect 15819 9463 15861 9472
rect 15915 9512 15957 9521
rect 15915 9472 15916 9512
rect 15956 9472 15957 9512
rect 15915 9463 15957 9472
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 16195 9512 16253 9513
rect 16195 9472 16204 9512
rect 16244 9472 16253 9512
rect 16195 9471 16253 9472
rect 16299 9512 16341 9521
rect 16299 9472 16300 9512
rect 16340 9472 16341 9512
rect 16299 9463 16341 9472
rect 16483 9512 16541 9513
rect 16483 9472 16492 9512
rect 16532 9472 16541 9512
rect 16483 9471 16541 9472
rect 16971 9512 17013 9521
rect 16971 9472 16972 9512
rect 17012 9472 17013 9512
rect 16971 9463 17013 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17251 9512 17309 9513
rect 17251 9472 17260 9512
rect 17300 9472 17309 9512
rect 17251 9471 17309 9472
rect 17539 9512 17597 9513
rect 17539 9472 17548 9512
rect 17588 9472 17597 9512
rect 17539 9471 17597 9472
rect 21099 9512 21141 9521
rect 21099 9472 21100 9512
rect 21140 9472 21141 9512
rect 21099 9463 21141 9472
rect 21475 9512 21533 9513
rect 21475 9472 21484 9512
rect 21524 9472 21533 9512
rect 21475 9471 21533 9472
rect 21667 9512 21725 9513
rect 21667 9472 21676 9512
rect 21716 9472 21725 9512
rect 21667 9471 21725 9472
rect 22435 9512 22493 9513
rect 22435 9472 22444 9512
rect 22484 9472 22493 9512
rect 22435 9471 22493 9472
rect 23683 9512 23741 9513
rect 23683 9472 23692 9512
rect 23732 9472 23741 9512
rect 23683 9471 23741 9472
rect 24075 9512 24117 9521
rect 24075 9472 24076 9512
rect 24116 9472 24117 9512
rect 24075 9463 24117 9472
rect 24171 9512 24213 9521
rect 24171 9472 24172 9512
rect 24212 9472 24213 9512
rect 24171 9463 24213 9472
rect 24267 9512 24309 9521
rect 24267 9472 24268 9512
rect 24308 9472 24309 9512
rect 24267 9463 24309 9472
rect 24363 9512 24405 9521
rect 24363 9472 24364 9512
rect 24404 9472 24405 9512
rect 24363 9463 24405 9472
rect 24555 9512 24597 9521
rect 24555 9472 24556 9512
rect 24596 9472 24597 9512
rect 24555 9463 24597 9472
rect 24651 9512 24693 9521
rect 24651 9472 24652 9512
rect 24692 9472 24693 9512
rect 24651 9463 24693 9472
rect 24747 9512 24789 9521
rect 24747 9472 24748 9512
rect 24788 9472 24789 9512
rect 24747 9463 24789 9472
rect 25219 9512 25277 9513
rect 25219 9472 25228 9512
rect 25268 9472 25277 9512
rect 25219 9471 25277 9472
rect 27243 9512 27285 9521
rect 27243 9472 27244 9512
rect 27284 9472 27285 9512
rect 27243 9463 27285 9472
rect 27435 9512 27477 9521
rect 27435 9472 27436 9512
rect 27476 9472 27477 9512
rect 27435 9463 27477 9472
rect 27523 9512 27581 9513
rect 27523 9472 27532 9512
rect 27572 9472 27581 9512
rect 27523 9471 27581 9472
rect 27907 9512 27965 9513
rect 27907 9472 27916 9512
rect 27956 9472 27965 9512
rect 27907 9471 27965 9472
rect 28299 9512 28341 9521
rect 28299 9472 28300 9512
rect 28340 9472 28341 9512
rect 28299 9463 28341 9472
rect 28395 9512 28437 9521
rect 28395 9472 28396 9512
rect 28436 9472 28437 9512
rect 28395 9463 28437 9472
rect 28491 9512 28533 9521
rect 28491 9472 28492 9512
rect 28532 9472 28533 9512
rect 28491 9463 28533 9472
rect 28683 9512 28725 9521
rect 28683 9472 28684 9512
rect 28724 9472 28725 9512
rect 28683 9463 28725 9472
rect 28779 9512 28821 9521
rect 28779 9472 28780 9512
rect 28820 9472 28821 9512
rect 28779 9463 28821 9472
rect 28875 9512 28917 9521
rect 28875 9472 28876 9512
rect 28916 9472 28917 9512
rect 28875 9463 28917 9472
rect 28971 9512 29013 9521
rect 28971 9472 28972 9512
rect 29012 9472 29013 9512
rect 28971 9463 29013 9472
rect 29246 9512 29304 9513
rect 29246 9472 29255 9512
rect 29295 9472 29304 9512
rect 29246 9471 29304 9472
rect 29355 9512 29397 9521
rect 29355 9472 29356 9512
rect 29396 9472 29397 9512
rect 29355 9463 29397 9472
rect 29451 9512 29493 9521
rect 29451 9472 29452 9512
rect 29492 9472 29493 9512
rect 29451 9463 29493 9472
rect 29635 9512 29693 9513
rect 29635 9472 29644 9512
rect 29684 9472 29693 9512
rect 29635 9471 29693 9472
rect 29731 9512 29789 9513
rect 29731 9472 29740 9512
rect 29780 9472 29789 9512
rect 29731 9471 29789 9472
rect 29923 9512 29981 9513
rect 29923 9472 29932 9512
rect 29972 9472 29981 9512
rect 29923 9471 29981 9472
rect 30315 9512 30357 9521
rect 30315 9472 30316 9512
rect 30356 9472 30357 9512
rect 30315 9463 30357 9472
rect 30507 9512 30549 9521
rect 30507 9472 30508 9512
rect 30548 9472 30549 9512
rect 30507 9463 30549 9472
rect 30699 9512 30741 9521
rect 30699 9472 30700 9512
rect 30740 9472 30741 9512
rect 30699 9463 30741 9472
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 31947 9512 31989 9521
rect 31947 9472 31948 9512
rect 31988 9472 31989 9512
rect 31947 9463 31989 9472
rect 32043 9512 32085 9521
rect 32043 9472 32044 9512
rect 32084 9472 32085 9512
rect 32043 9463 32085 9472
rect 32611 9512 32669 9513
rect 32611 9472 32620 9512
rect 32660 9472 32669 9512
rect 32611 9471 32669 9472
rect 32907 9512 32949 9521
rect 32907 9472 32908 9512
rect 32948 9472 32949 9512
rect 32907 9463 32949 9472
rect 33003 9512 33045 9521
rect 33003 9472 33004 9512
rect 33044 9472 33045 9512
rect 33003 9463 33045 9472
rect 33099 9512 33141 9521
rect 33099 9472 33100 9512
rect 33140 9472 33141 9512
rect 33099 9463 33141 9472
rect 34243 9512 34301 9513
rect 34243 9472 34252 9512
rect 34292 9472 34301 9512
rect 34243 9471 34301 9472
rect 34435 9512 34493 9513
rect 34435 9472 34444 9512
rect 34484 9472 34493 9512
rect 34435 9471 34493 9472
rect 34635 9512 34677 9521
rect 34635 9472 34636 9512
rect 34676 9472 34677 9512
rect 34635 9463 34677 9472
rect 34723 9512 34781 9513
rect 34723 9472 34732 9512
rect 34772 9472 34781 9512
rect 34723 9471 34781 9472
rect 34923 9512 34965 9521
rect 34923 9472 34924 9512
rect 34964 9472 34965 9512
rect 34923 9463 34965 9472
rect 35115 9512 35157 9521
rect 35115 9472 35116 9512
rect 35156 9472 35157 9512
rect 35115 9463 35157 9472
rect 35211 9512 35253 9521
rect 35211 9472 35212 9512
rect 35252 9472 35253 9512
rect 35211 9463 35253 9472
rect 35683 9512 35741 9513
rect 35683 9472 35692 9512
rect 35732 9472 35741 9512
rect 35683 9471 35741 9472
rect 36259 9512 36317 9513
rect 36259 9472 36268 9512
rect 36308 9472 36317 9512
rect 36259 9471 36317 9472
rect 37323 9512 37365 9521
rect 37323 9472 37324 9512
rect 37364 9472 37365 9512
rect 37323 9463 37365 9472
rect 37987 9512 38045 9513
rect 37987 9472 37996 9512
rect 38036 9472 38045 9512
rect 37987 9471 38045 9472
rect 38851 9512 38909 9513
rect 38851 9472 38860 9512
rect 38900 9472 38909 9512
rect 38851 9471 38909 9472
rect 7947 9428 7989 9437
rect 7947 9388 7948 9428
rect 7988 9388 7989 9428
rect 7947 9379 7989 9388
rect 22827 9428 22869 9437
rect 22827 9388 22828 9428
rect 22868 9388 22869 9428
rect 22827 9379 22869 9388
rect 30027 9428 30069 9437
rect 30027 9388 30028 9428
rect 30068 9388 30069 9428
rect 30027 9379 30069 9388
rect 30219 9428 30261 9437
rect 30219 9388 30220 9428
rect 30260 9388 30261 9428
rect 30219 9379 30261 9388
rect 3915 9344 3957 9353
rect 3915 9304 3916 9344
rect 3956 9304 3957 9344
rect 3915 9295 3957 9304
rect 12843 9344 12885 9353
rect 12843 9304 12844 9344
rect 12884 9304 12885 9344
rect 12843 9295 12885 9304
rect 16491 9344 16533 9353
rect 16491 9304 16492 9344
rect 16532 9304 16533 9344
rect 16491 9295 16533 9304
rect 18699 9344 18741 9353
rect 18699 9304 18700 9344
rect 18740 9304 18741 9344
rect 18699 9295 18741 9304
rect 20907 9344 20949 9353
rect 20907 9304 20908 9344
rect 20948 9304 20949 9344
rect 20907 9295 20949 9304
rect 23403 9344 23445 9353
rect 23403 9304 23404 9344
rect 23444 9304 23445 9344
rect 23403 9295 23445 9304
rect 30123 9344 30165 9353
rect 30123 9304 30124 9344
rect 30164 9304 30165 9344
rect 30123 9295 30165 9304
rect 11971 9260 12029 9261
rect 11971 9220 11980 9260
rect 12020 9220 12029 9260
rect 11971 9219 12029 9220
rect 14571 9260 14613 9269
rect 14571 9220 14572 9260
rect 14612 9220 14613 9260
rect 14571 9211 14613 9220
rect 16971 9260 17013 9269
rect 16971 9220 16972 9260
rect 17012 9220 17013 9260
rect 16971 9211 17013 9220
rect 18219 9260 18261 9269
rect 18219 9220 18220 9260
rect 18260 9220 18261 9260
rect 18219 9211 18261 9220
rect 22539 9260 22581 9269
rect 22539 9220 22540 9260
rect 22580 9220 22581 9260
rect 22539 9211 22581 9220
rect 25323 9260 25365 9269
rect 25323 9220 25324 9260
rect 25364 9220 25365 9260
rect 25323 9211 25365 9220
rect 32715 9260 32757 9269
rect 32715 9220 32716 9260
rect 32756 9220 32757 9260
rect 32715 9211 32757 9220
rect 34155 9260 34197 9269
rect 34155 9220 34156 9260
rect 34196 9220 34197 9260
rect 34155 9211 34197 9220
rect 34443 9260 34485 9269
rect 34443 9220 34444 9260
rect 34484 9220 34485 9260
rect 34443 9211 34485 9220
rect 35875 9260 35933 9261
rect 35875 9220 35884 9260
rect 35924 9220 35933 9260
rect 35875 9219 35933 9220
rect 36931 9260 36989 9261
rect 36931 9220 36940 9260
rect 36980 9220 36989 9260
rect 36931 9219 36989 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 16299 8924 16341 8933
rect 16299 8884 16300 8924
rect 16340 8884 16341 8924
rect 16299 8875 16341 8884
rect 24171 8924 24213 8933
rect 24171 8884 24172 8924
rect 24212 8884 24213 8924
rect 31467 8924 31509 8933
rect 24171 8875 24213 8884
rect 24843 8882 24885 8891
rect 6123 8840 6165 8849
rect 6123 8800 6124 8840
rect 6164 8800 6165 8840
rect 6123 8791 6165 8800
rect 18027 8840 18069 8849
rect 18027 8800 18028 8840
rect 18068 8800 18069 8840
rect 18027 8791 18069 8800
rect 19755 8840 19797 8849
rect 19755 8800 19756 8840
rect 19796 8800 19797 8840
rect 24843 8842 24844 8882
rect 24884 8842 24885 8882
rect 31467 8884 31468 8924
rect 31508 8884 31509 8924
rect 31467 8875 31509 8884
rect 32139 8924 32181 8933
rect 32139 8884 32140 8924
rect 32180 8884 32181 8924
rect 32139 8875 32181 8884
rect 39051 8924 39093 8933
rect 39051 8884 39052 8924
rect 39092 8884 39093 8924
rect 39051 8875 39093 8884
rect 24843 8833 24885 8842
rect 26379 8840 26421 8849
rect 19755 8791 19797 8800
rect 26379 8800 26380 8840
rect 26420 8800 26421 8840
rect 26379 8791 26421 8800
rect 27139 8840 27197 8841
rect 27139 8800 27148 8840
rect 27188 8800 27197 8840
rect 27139 8799 27197 8800
rect 30027 8840 30069 8849
rect 30027 8800 30028 8840
rect 30068 8800 30069 8840
rect 30027 8791 30069 8800
rect 32523 8840 32565 8849
rect 32523 8800 32524 8840
rect 32564 8800 32565 8840
rect 32523 8791 32565 8800
rect 35595 8840 35637 8849
rect 35595 8800 35596 8840
rect 35636 8800 35637 8840
rect 35595 8791 35637 8800
rect 13419 8756 13461 8765
rect 13419 8716 13420 8756
rect 13460 8716 13461 8756
rect 13419 8707 13461 8716
rect 24747 8756 24789 8765
rect 24747 8716 24748 8756
rect 24788 8716 24789 8756
rect 24747 8707 24789 8716
rect 24939 8756 24981 8765
rect 24939 8716 24940 8756
rect 24980 8716 24981 8756
rect 24939 8707 24981 8716
rect 32427 8756 32469 8765
rect 32427 8716 32428 8756
rect 32468 8716 32469 8756
rect 25699 8714 25757 8715
rect 3435 8672 3477 8681
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 3811 8672 3869 8673
rect 3811 8632 3820 8672
rect 3860 8632 3869 8672
rect 3811 8631 3869 8632
rect 4675 8672 4733 8673
rect 4675 8632 4684 8672
rect 4724 8632 4733 8672
rect 4675 8631 4733 8632
rect 5923 8672 5981 8673
rect 5923 8632 5932 8672
rect 5972 8632 5981 8672
rect 5923 8631 5981 8632
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 6315 8672 6357 8681
rect 6315 8632 6316 8672
rect 6356 8632 6357 8672
rect 6315 8623 6357 8632
rect 7075 8672 7133 8673
rect 7075 8632 7084 8672
rect 7124 8632 7133 8672
rect 7075 8631 7133 8632
rect 7939 8672 7997 8673
rect 7939 8632 7948 8672
rect 7988 8632 7997 8672
rect 7939 8631 7997 8632
rect 9475 8672 9533 8673
rect 9475 8632 9484 8672
rect 9524 8632 9533 8672
rect 9475 8631 9533 8632
rect 10339 8672 10397 8673
rect 10339 8632 10348 8672
rect 10388 8632 10397 8672
rect 10339 8631 10397 8632
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10635 8672 10677 8681
rect 10635 8632 10636 8672
rect 10676 8632 10677 8672
rect 10635 8623 10677 8632
rect 11019 8672 11061 8681
rect 11019 8632 11020 8672
rect 11060 8632 11061 8672
rect 11019 8623 11061 8632
rect 11395 8672 11453 8673
rect 11395 8632 11404 8672
rect 11444 8632 11453 8672
rect 11395 8631 11453 8632
rect 12259 8672 12317 8673
rect 12259 8632 12268 8672
rect 12308 8632 12317 8672
rect 12259 8631 12317 8632
rect 14275 8672 14333 8673
rect 14275 8632 14284 8672
rect 14324 8632 14333 8672
rect 14275 8631 14333 8632
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14859 8672 14901 8681
rect 14859 8632 14860 8672
rect 14900 8632 14901 8672
rect 14859 8623 14901 8632
rect 14955 8672 14997 8681
rect 14955 8632 14956 8672
rect 14996 8632 14997 8672
rect 14955 8623 14997 8632
rect 15811 8672 15869 8673
rect 15811 8632 15820 8672
rect 15860 8632 15869 8672
rect 15811 8631 15869 8632
rect 16003 8672 16061 8673
rect 16003 8632 16012 8672
rect 16052 8632 16061 8672
rect 16003 8631 16061 8632
rect 16107 8672 16149 8681
rect 16107 8632 16108 8672
rect 16148 8632 16149 8672
rect 16107 8623 16149 8632
rect 16291 8672 16349 8673
rect 16291 8632 16300 8672
rect 16340 8632 16349 8672
rect 16291 8631 16349 8632
rect 16683 8672 16725 8681
rect 16683 8632 16684 8672
rect 16724 8632 16725 8672
rect 16683 8623 16725 8632
rect 16779 8672 16821 8681
rect 16779 8632 16780 8672
rect 16820 8632 16821 8672
rect 16779 8623 16821 8632
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 16875 8623 16917 8632
rect 16971 8672 17013 8681
rect 16971 8632 16972 8672
rect 17012 8632 17013 8672
rect 16971 8623 17013 8632
rect 17155 8672 17213 8673
rect 17155 8632 17164 8672
rect 17204 8632 17213 8672
rect 17155 8631 17213 8632
rect 21003 8672 21045 8681
rect 21003 8632 21004 8672
rect 21044 8632 21045 8672
rect 21003 8623 21045 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22347 8672 22389 8681
rect 22347 8632 22348 8672
rect 22388 8632 22389 8672
rect 22347 8623 22389 8632
rect 23115 8672 23157 8681
rect 23115 8632 23116 8672
rect 23156 8632 23157 8672
rect 23115 8623 23157 8632
rect 23211 8672 23253 8681
rect 23211 8632 23212 8672
rect 23252 8632 23253 8672
rect 23211 8623 23253 8632
rect 23403 8672 23445 8681
rect 23403 8632 23404 8672
rect 23444 8632 23445 8672
rect 23403 8623 23445 8632
rect 23499 8672 23541 8681
rect 23499 8632 23500 8672
rect 23540 8632 23541 8672
rect 23499 8623 23541 8632
rect 23875 8672 23933 8673
rect 23875 8632 23884 8672
rect 23924 8632 23933 8672
rect 23875 8631 23933 8632
rect 23979 8672 24021 8681
rect 23979 8632 23980 8672
rect 24020 8632 24021 8672
rect 23979 8623 24021 8632
rect 24171 8672 24213 8681
rect 24171 8632 24172 8672
rect 24212 8632 24213 8672
rect 24171 8623 24213 8632
rect 24651 8672 24693 8681
rect 24651 8632 24652 8672
rect 24692 8632 24693 8672
rect 24651 8623 24693 8632
rect 25027 8672 25085 8673
rect 25027 8632 25036 8672
rect 25076 8632 25085 8672
rect 25027 8631 25085 8632
rect 25315 8672 25373 8673
rect 25315 8632 25324 8672
rect 25364 8632 25373 8672
rect 25315 8631 25373 8632
rect 25611 8672 25653 8681
rect 25699 8674 25708 8714
rect 25748 8674 25757 8714
rect 32427 8707 32469 8716
rect 32619 8756 32661 8765
rect 32619 8716 32620 8756
rect 32660 8716 32661 8756
rect 32619 8707 32661 8716
rect 34155 8756 34197 8765
rect 34155 8716 34156 8756
rect 34196 8716 34197 8756
rect 34155 8707 34197 8716
rect 34731 8697 34773 8706
rect 25699 8673 25757 8674
rect 25611 8632 25612 8672
rect 25652 8632 25653 8672
rect 25611 8623 25653 8632
rect 25803 8672 25845 8681
rect 25803 8632 25804 8672
rect 25844 8632 25845 8672
rect 25803 8623 25845 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 26379 8672 26421 8681
rect 26379 8632 26380 8672
rect 26420 8632 26421 8672
rect 26379 8623 26421 8632
rect 26571 8672 26613 8681
rect 26571 8632 26572 8672
rect 26612 8632 26613 8672
rect 26571 8623 26613 8632
rect 26763 8672 26805 8681
rect 26763 8632 26764 8672
rect 26804 8632 26805 8672
rect 26763 8623 26805 8632
rect 26859 8672 26901 8681
rect 26859 8632 26860 8672
rect 26900 8632 26901 8672
rect 26859 8623 26901 8632
rect 27051 8672 27093 8681
rect 27051 8632 27052 8672
rect 27092 8632 27093 8672
rect 27051 8623 27093 8632
rect 27147 8672 27189 8681
rect 27147 8632 27148 8672
rect 27188 8632 27189 8672
rect 27147 8623 27189 8632
rect 27339 8672 27381 8681
rect 27339 8632 27340 8672
rect 27380 8632 27381 8672
rect 27339 8623 27381 8632
rect 28771 8672 28829 8673
rect 28771 8632 28780 8672
rect 28820 8632 28829 8672
rect 28771 8631 28829 8632
rect 29067 8672 29109 8681
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 29739 8672 29781 8681
rect 29739 8632 29740 8672
rect 29780 8632 29781 8672
rect 29739 8623 29781 8632
rect 29835 8672 29877 8681
rect 29835 8632 29836 8672
rect 29876 8632 29877 8672
rect 29835 8623 29877 8632
rect 30115 8672 30173 8673
rect 30115 8632 30124 8672
rect 30164 8632 30173 8672
rect 30115 8631 30173 8632
rect 31075 8672 31133 8673
rect 31075 8632 31084 8672
rect 31124 8632 31133 8672
rect 31075 8631 31133 8632
rect 31363 8672 31421 8673
rect 31363 8632 31372 8672
rect 31412 8632 31421 8672
rect 31363 8631 31421 8632
rect 31467 8672 31509 8681
rect 31467 8632 31468 8672
rect 31508 8632 31509 8672
rect 31467 8623 31509 8632
rect 31651 8672 31709 8673
rect 31651 8632 31660 8672
rect 31700 8632 31709 8672
rect 31651 8631 31709 8632
rect 31843 8672 31901 8673
rect 31843 8632 31852 8672
rect 31892 8632 31901 8672
rect 31843 8631 31901 8632
rect 31947 8672 31989 8681
rect 31947 8632 31948 8672
rect 31988 8632 31989 8672
rect 31947 8623 31989 8632
rect 32139 8672 32181 8681
rect 32139 8632 32140 8672
rect 32180 8632 32181 8672
rect 32139 8623 32181 8632
rect 32331 8672 32373 8681
rect 32331 8632 32332 8672
rect 32372 8632 32373 8672
rect 32331 8623 32373 8632
rect 32707 8672 32765 8673
rect 32707 8632 32716 8672
rect 32756 8632 32765 8672
rect 32707 8631 32765 8632
rect 32907 8672 32949 8681
rect 32907 8632 32908 8672
rect 32948 8632 32949 8672
rect 32907 8623 32949 8632
rect 33003 8672 33045 8681
rect 33003 8632 33004 8672
rect 33044 8632 33045 8672
rect 33003 8623 33045 8632
rect 33475 8672 33533 8673
rect 33475 8632 33484 8672
rect 33524 8632 33533 8672
rect 33963 8672 34005 8681
rect 33475 8631 33533 8632
rect 33667 8669 33725 8670
rect 33667 8629 33676 8669
rect 33716 8629 33725 8669
rect 33667 8628 33725 8629
rect 33963 8632 33964 8672
rect 34004 8632 34005 8672
rect 33963 8623 34005 8632
rect 34251 8672 34293 8681
rect 34251 8632 34252 8672
rect 34292 8632 34293 8672
rect 34251 8623 34293 8632
rect 34443 8672 34485 8681
rect 34443 8632 34444 8672
rect 34484 8632 34485 8672
rect 34443 8623 34485 8632
rect 34635 8672 34677 8681
rect 34635 8632 34636 8672
rect 34676 8632 34677 8672
rect 34731 8657 34732 8697
rect 34772 8657 34773 8697
rect 34731 8648 34773 8657
rect 35299 8672 35357 8673
rect 34635 8623 34677 8632
rect 35299 8632 35308 8672
rect 35348 8632 35357 8672
rect 35299 8631 35357 8632
rect 35403 8672 35445 8681
rect 35403 8632 35404 8672
rect 35444 8632 35445 8672
rect 35403 8623 35445 8632
rect 35595 8672 35637 8681
rect 35595 8632 35596 8672
rect 35636 8632 35637 8672
rect 35595 8623 35637 8632
rect 35779 8672 35837 8673
rect 35779 8632 35788 8672
rect 35828 8632 35837 8672
rect 35779 8631 35837 8632
rect 36459 8672 36501 8681
rect 36459 8632 36460 8672
rect 36500 8632 36501 8672
rect 36459 8623 36501 8632
rect 36651 8672 36693 8681
rect 36651 8632 36652 8672
rect 36692 8632 36693 8672
rect 36651 8623 36693 8632
rect 37027 8672 37085 8673
rect 37027 8632 37036 8672
rect 37076 8632 37085 8672
rect 37027 8631 37085 8632
rect 37891 8672 37949 8673
rect 37891 8632 37900 8672
rect 37940 8632 37949 8672
rect 37891 8631 37949 8632
rect 6699 8588 6741 8597
rect 6699 8548 6700 8588
rect 6740 8548 6741 8588
rect 6699 8539 6741 8548
rect 643 8504 701 8505
rect 643 8464 652 8504
rect 692 8464 701 8504
rect 643 8463 701 8464
rect 9091 8504 9149 8505
rect 9091 8464 9100 8504
rect 9140 8464 9149 8504
rect 9091 8463 9149 8464
rect 10147 8504 10205 8505
rect 10147 8464 10156 8504
rect 10196 8464 10205 8504
rect 10147 8463 10205 8464
rect 10531 8504 10589 8505
rect 10531 8464 10540 8504
rect 10580 8464 10589 8504
rect 10531 8463 10589 8464
rect 13603 8504 13661 8505
rect 13603 8464 13612 8504
rect 13652 8464 13661 8504
rect 13603 8463 13661 8464
rect 14659 8504 14717 8505
rect 14659 8464 14668 8504
rect 14708 8464 14717 8504
rect 14659 8463 14717 8464
rect 15139 8504 15197 8505
rect 15139 8464 15148 8504
rect 15188 8464 15197 8504
rect 15139 8463 15197 8464
rect 17827 8504 17885 8505
rect 17827 8464 17836 8504
rect 17876 8464 17885 8504
rect 17827 8463 17885 8464
rect 20619 8504 20661 8513
rect 20619 8464 20620 8504
rect 20660 8464 20661 8504
rect 20619 8455 20661 8464
rect 22251 8504 22293 8513
rect 22251 8464 22252 8504
rect 22292 8464 22293 8504
rect 22251 8455 22293 8464
rect 22915 8504 22973 8505
rect 22915 8464 22924 8504
rect 22964 8464 22973 8504
rect 22915 8463 22973 8464
rect 23683 8504 23741 8505
rect 23683 8464 23692 8504
rect 23732 8464 23741 8504
rect 23683 8463 23741 8464
rect 25227 8504 25269 8513
rect 25227 8464 25228 8504
rect 25268 8464 25269 8504
rect 25227 8455 25269 8464
rect 25891 8504 25949 8505
rect 25891 8464 25900 8504
rect 25940 8464 25949 8504
rect 25891 8463 25949 8464
rect 26667 8504 26709 8513
rect 26667 8464 26668 8504
rect 26708 8464 26709 8504
rect 26667 8455 26709 8464
rect 28875 8504 28917 8513
rect 28875 8464 28876 8504
rect 28916 8464 28917 8504
rect 28875 8455 28917 8464
rect 29347 8504 29405 8505
rect 29347 8464 29356 8504
rect 29396 8464 29405 8504
rect 29347 8463 29405 8464
rect 29539 8504 29597 8505
rect 29539 8464 29548 8504
rect 29588 8464 29597 8504
rect 29539 8463 29597 8464
rect 31179 8504 31221 8513
rect 31179 8464 31180 8504
rect 31220 8464 31221 8504
rect 31179 8455 31221 8464
rect 33187 8504 33245 8505
rect 33187 8464 33196 8504
rect 33236 8464 33245 8504
rect 33187 8463 33245 8464
rect 34723 8462 34781 8463
rect 34723 8422 34732 8462
rect 34772 8422 34781 8462
rect 34723 8421 34781 8422
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 643 8168 701 8169
rect 643 8128 652 8168
rect 692 8128 701 8168
rect 643 8127 701 8128
rect 5635 8168 5693 8169
rect 5635 8128 5644 8168
rect 5684 8128 5693 8168
rect 5635 8127 5693 8128
rect 8227 8168 8285 8169
rect 8227 8128 8236 8168
rect 8276 8128 8285 8168
rect 8227 8127 8285 8128
rect 9283 8168 9341 8169
rect 9283 8128 9292 8168
rect 9332 8128 9341 8168
rect 9283 8127 9341 8128
rect 13035 8168 13077 8177
rect 13035 8128 13036 8168
rect 13076 8128 13077 8168
rect 13035 8119 13077 8128
rect 13611 8168 13653 8177
rect 13611 8128 13612 8168
rect 13652 8128 13653 8168
rect 13611 8119 13653 8128
rect 14467 8168 14525 8169
rect 14467 8128 14476 8168
rect 14516 8128 14525 8168
rect 14467 8127 14525 8128
rect 17347 8168 17405 8169
rect 17347 8128 17356 8168
rect 17396 8128 17405 8168
rect 17347 8127 17405 8128
rect 20899 8168 20957 8169
rect 20899 8128 20908 8168
rect 20948 8128 20957 8168
rect 20899 8127 20957 8128
rect 22819 8168 22877 8169
rect 22819 8128 22828 8168
rect 22868 8128 22877 8168
rect 22819 8127 22877 8128
rect 23403 8168 23445 8177
rect 23403 8128 23404 8168
rect 23444 8128 23445 8168
rect 23403 8119 23445 8128
rect 26571 8168 26613 8177
rect 26571 8128 26572 8168
rect 26612 8128 26613 8168
rect 26571 8119 26613 8128
rect 26955 8168 26997 8177
rect 26955 8128 26956 8168
rect 26996 8128 26997 8168
rect 26955 8119 26997 8128
rect 28387 8168 28445 8169
rect 28387 8128 28396 8168
rect 28436 8128 28445 8168
rect 28387 8127 28445 8128
rect 30211 8168 30269 8169
rect 30211 8128 30220 8168
rect 30260 8128 30269 8168
rect 30211 8127 30269 8128
rect 30787 8168 30845 8169
rect 30787 8128 30796 8168
rect 30836 8128 30845 8168
rect 30787 8127 30845 8128
rect 32131 8168 32189 8169
rect 32131 8128 32140 8168
rect 32180 8128 32189 8168
rect 32131 8127 32189 8128
rect 32715 8168 32757 8177
rect 32715 8128 32716 8168
rect 32756 8128 32757 8168
rect 32715 8119 32757 8128
rect 34627 8168 34685 8169
rect 34627 8128 34636 8168
rect 34676 8128 34685 8168
rect 34627 8127 34685 8128
rect 35683 8168 35741 8169
rect 35683 8128 35692 8168
rect 35732 8128 35741 8168
rect 35683 8127 35741 8128
rect 14955 8084 14997 8093
rect 14955 8044 14956 8084
rect 14996 8044 14997 8084
rect 14955 8035 14997 8044
rect 17547 8084 17589 8093
rect 17547 8044 17548 8084
rect 17588 8044 17589 8084
rect 17547 8035 17589 8044
rect 28875 8084 28917 8093
rect 28875 8044 28876 8084
rect 28916 8044 28917 8084
rect 28875 8035 28917 8044
rect 31851 8084 31893 8093
rect 31851 8044 31852 8084
rect 31892 8044 31893 8084
rect 31851 8035 31893 8044
rect 4483 8000 4541 8001
rect 4483 7960 4492 8000
rect 4532 7960 4541 8000
rect 4483 7959 4541 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4875 8000 4917 8009
rect 4875 7960 4876 8000
rect 4916 7960 4917 8000
rect 4875 7951 4917 7960
rect 4963 8000 5021 8001
rect 4963 7960 4972 8000
rect 5012 7960 5021 8000
rect 4963 7959 5021 7960
rect 5163 8000 5205 8009
rect 5163 7960 5164 8000
rect 5204 7960 5205 8000
rect 5163 7951 5205 7960
rect 5259 8000 5301 8009
rect 5259 7960 5260 8000
rect 5300 7960 5301 8000
rect 5259 7951 5301 7960
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5451 8000 5493 8009
rect 5451 7960 5452 8000
rect 5492 7960 5493 8000
rect 5451 7951 5493 7960
rect 5739 8000 5781 8009
rect 5739 7960 5740 8000
rect 5780 7960 5781 8000
rect 5739 7951 5781 7960
rect 5835 8000 5877 8009
rect 5835 7960 5836 8000
rect 5876 7960 5877 8000
rect 5835 7951 5877 7960
rect 5931 8000 5973 8009
rect 5931 7960 5932 8000
rect 5972 7960 5973 8000
rect 5931 7951 5973 7960
rect 7459 8000 7517 8001
rect 7459 7960 7468 8000
rect 7508 7960 7517 8000
rect 7459 7959 7517 7960
rect 7563 8000 7605 8009
rect 7563 7960 7564 8000
rect 7604 7960 7605 8000
rect 7563 7951 7605 7960
rect 7755 8000 7797 8009
rect 7755 7960 7756 8000
rect 7796 7960 7797 8000
rect 7755 7951 7797 7960
rect 8043 8000 8085 8009
rect 8043 7960 8044 8000
rect 8084 7960 8085 8000
rect 8043 7951 8085 7960
rect 8899 8000 8957 8001
rect 8899 7960 8908 8000
rect 8948 7960 8957 8000
rect 8899 7959 8957 7960
rect 9091 8000 9149 8001
rect 9091 7960 9100 8000
rect 9140 7960 9149 8000
rect 9091 7959 9149 7960
rect 9187 8000 9245 8001
rect 9187 7960 9196 8000
rect 9236 7960 9245 8000
rect 9187 7959 9245 7960
rect 9387 8000 9429 8009
rect 9387 7960 9388 8000
rect 9428 7960 9429 8000
rect 9387 7951 9429 7960
rect 9483 8000 9525 8009
rect 9483 7960 9484 8000
rect 9524 7960 9525 8000
rect 9483 7951 9525 7960
rect 9630 8000 9688 8001
rect 9630 7960 9639 8000
rect 9679 7960 9688 8000
rect 9630 7959 9688 7960
rect 9955 8000 10013 8001
rect 9955 7960 9964 8000
rect 10004 7960 10013 8000
rect 9955 7959 10013 7960
rect 10147 8000 10205 8001
rect 10147 7960 10156 8000
rect 10196 7960 10205 8000
rect 10147 7959 10205 7960
rect 11779 8000 11837 8001
rect 11779 7960 11788 8000
rect 11828 7960 11837 8000
rect 11779 7959 11837 7960
rect 12651 8000 12693 8009
rect 12651 7960 12652 8000
rect 12692 7960 12693 8000
rect 12651 7951 12693 7960
rect 13123 8000 13181 8001
rect 13123 7960 13132 8000
rect 13172 7960 13181 8000
rect 13123 7959 13181 7960
rect 13995 8000 14037 8009
rect 13995 7960 13996 8000
rect 14036 7960 14037 8000
rect 13995 7951 14037 7960
rect 14091 8000 14133 8009
rect 14091 7960 14092 8000
rect 14132 7960 14133 8000
rect 14091 7951 14133 7960
rect 14187 8000 14229 8009
rect 14187 7960 14188 8000
rect 14228 7960 14229 8000
rect 14187 7951 14229 7960
rect 14283 8000 14325 8009
rect 14283 7960 14284 8000
rect 14324 7960 14325 8000
rect 14283 7951 14325 7960
rect 14571 8000 14613 8009
rect 14571 7960 14572 8000
rect 14612 7960 14613 8000
rect 14571 7951 14613 7960
rect 14667 8000 14709 8009
rect 14667 7960 14668 8000
rect 14708 7960 14709 8000
rect 14667 7951 14709 7960
rect 14763 8000 14805 8009
rect 14763 7960 14764 8000
rect 14804 7960 14805 8000
rect 14763 7951 14805 7960
rect 15331 8000 15389 8001
rect 15331 7960 15340 8000
rect 15380 7960 15389 8000
rect 15331 7959 15389 7960
rect 16195 8000 16253 8001
rect 16195 7960 16204 8000
rect 16244 7960 16253 8000
rect 16195 7959 16253 7960
rect 17923 8000 17981 8001
rect 17923 7960 17932 8000
rect 17972 7960 17981 8000
rect 17923 7959 17981 7960
rect 18787 8000 18845 8001
rect 18787 7960 18796 8000
rect 18836 7960 18845 8000
rect 18787 7959 18845 7960
rect 20227 8000 20285 8001
rect 20227 7960 20236 8000
rect 20276 7960 20285 8000
rect 20227 7959 20285 7960
rect 21195 8000 21237 8009
rect 21195 7960 21196 8000
rect 21236 7960 21237 8000
rect 21195 7951 21237 7960
rect 21483 8000 21525 8009
rect 21483 7960 21484 8000
rect 21524 7960 21525 8000
rect 21483 7951 21525 7960
rect 21667 8000 21725 8001
rect 21667 7960 21676 8000
rect 21716 7960 21725 8000
rect 21667 7959 21725 7960
rect 22539 8000 22581 8009
rect 22539 7960 22540 8000
rect 22580 7960 22581 8000
rect 22539 7951 22581 7960
rect 22635 8000 22677 8009
rect 22635 7960 22636 8000
rect 22676 7960 22677 8000
rect 22635 7951 22677 7960
rect 23211 8000 23253 8009
rect 23211 7960 23212 8000
rect 23252 7960 23253 8000
rect 23211 7951 23253 7960
rect 23499 8000 23541 8009
rect 24075 8000 24117 8009
rect 23499 7960 23500 8000
rect 23540 7960 23541 8000
rect 23499 7951 23541 7960
rect 23787 7991 23829 8000
rect 23787 7951 23788 7991
rect 23828 7951 23829 7991
rect 24075 7960 24076 8000
rect 24116 7960 24117 8000
rect 24075 7951 24117 7960
rect 24747 8000 24789 8009
rect 24747 7960 24748 8000
rect 24788 7960 24789 8000
rect 24747 7951 24789 7960
rect 25035 8000 25077 8009
rect 25035 7960 25036 8000
rect 25076 7960 25077 8000
rect 25035 7951 25077 7960
rect 25219 8000 25277 8001
rect 25219 7960 25228 8000
rect 25268 7960 25277 8000
rect 25219 7959 25277 7960
rect 25315 8000 25373 8001
rect 25315 7960 25324 8000
rect 25364 7960 25373 8000
rect 25315 7959 25373 7960
rect 25515 8000 25557 8009
rect 25515 7960 25516 8000
rect 25556 7960 25557 8000
rect 25515 7951 25557 7960
rect 25611 8000 25653 8009
rect 25611 7960 25612 8000
rect 25652 7960 25653 8000
rect 25611 7951 25653 7960
rect 25758 8000 25816 8001
rect 25758 7960 25767 8000
rect 25807 7960 25816 8000
rect 25758 7959 25816 7960
rect 26379 8000 26421 8009
rect 26379 7960 26380 8000
rect 26420 7960 26421 8000
rect 26379 7951 26421 7960
rect 26667 8000 26709 8009
rect 26667 7960 26668 8000
rect 26708 7960 26709 8000
rect 26667 7951 26709 7960
rect 27139 8000 27197 8001
rect 27139 7960 27148 8000
rect 27188 7960 27197 8000
rect 27139 7959 27197 7960
rect 27427 8000 27485 8001
rect 27427 7960 27436 8000
rect 27476 7960 27485 8000
rect 27427 7959 27485 7960
rect 28107 8000 28149 8009
rect 28107 7960 28108 8000
rect 28148 7960 28149 8000
rect 28107 7951 28149 7960
rect 28203 8000 28245 8009
rect 28203 7960 28204 8000
rect 28244 7960 28245 8000
rect 28203 7951 28245 7960
rect 28299 8000 28341 8009
rect 28299 7960 28300 8000
rect 28340 7960 28341 8000
rect 28299 7951 28341 7960
rect 28587 8000 28629 8009
rect 28587 7960 28588 8000
rect 28628 7960 28629 8000
rect 28587 7951 28629 7960
rect 28683 8000 28725 8009
rect 28683 7960 28684 8000
rect 28724 7960 28725 8000
rect 28683 7951 28725 7960
rect 28779 8000 28821 8009
rect 28779 7960 28780 8000
rect 28820 7960 28821 8000
rect 28779 7951 28821 7960
rect 29059 8000 29117 8001
rect 29059 7960 29068 8000
rect 29108 7960 29117 8000
rect 29059 7959 29117 7960
rect 29451 8000 29493 8009
rect 29451 7960 29452 8000
rect 29492 7960 29493 8000
rect 29451 7951 29493 7960
rect 29731 8000 29789 8001
rect 29731 7960 29740 8000
rect 29780 7960 29789 8000
rect 29731 7959 29789 7960
rect 29827 8000 29885 8001
rect 29827 7960 29836 8000
rect 29876 7960 29885 8000
rect 29827 7959 29885 7960
rect 30027 8000 30069 8009
rect 30027 7960 30028 8000
rect 30068 7960 30069 8000
rect 30027 7951 30069 7960
rect 30123 8000 30165 8009
rect 30123 7960 30124 8000
rect 30164 7960 30165 8000
rect 30507 8000 30549 8009
rect 30123 7951 30165 7960
rect 30280 7985 30322 7994
rect 23787 7942 23829 7951
rect 30280 7945 30281 7985
rect 30321 7945 30322 7985
rect 30507 7960 30508 8000
rect 30548 7960 30549 8000
rect 30507 7951 30549 7960
rect 30603 8000 30645 8009
rect 30603 7960 30604 8000
rect 30644 7960 30645 8000
rect 30603 7951 30645 7960
rect 30699 8000 30741 8009
rect 30699 7960 30700 8000
rect 30740 7960 30741 8000
rect 30699 7951 30741 7960
rect 31083 8000 31125 8009
rect 31083 7960 31084 8000
rect 31124 7960 31125 8000
rect 31083 7951 31125 7960
rect 31459 8000 31517 8001
rect 31459 7960 31468 8000
rect 31508 7960 31517 8000
rect 31459 7959 31517 7960
rect 31755 8000 31797 8009
rect 31755 7960 31756 8000
rect 31796 7960 31797 8000
rect 31755 7951 31797 7960
rect 31939 8000 31997 8001
rect 31939 7960 31948 8000
rect 31988 7960 31997 8000
rect 31939 7959 31997 7960
rect 32331 8000 32373 8009
rect 32331 7960 32332 8000
rect 32372 7960 32373 8000
rect 32331 7951 32373 7960
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 32619 8000 32661 8009
rect 32619 7960 32620 8000
rect 32660 7960 32661 8000
rect 32619 7951 32661 7960
rect 32907 8000 32949 8009
rect 32907 7960 32908 8000
rect 32948 7960 32949 8000
rect 32907 7951 32949 7960
rect 33283 8000 33341 8001
rect 33283 7960 33292 8000
rect 33332 7960 33341 8000
rect 33283 7959 33341 7960
rect 33475 8000 33533 8001
rect 33475 7960 33484 8000
rect 33524 7960 33533 8000
rect 33475 7959 33533 7960
rect 33579 8000 33621 8009
rect 33579 7960 33580 8000
rect 33620 7960 33621 8000
rect 33579 7951 33621 7960
rect 33771 8000 33813 8009
rect 33771 7960 33772 8000
rect 33812 7960 33813 8000
rect 33771 7951 33813 7960
rect 33955 8000 34013 8001
rect 33955 7960 33964 8000
rect 34004 7960 34013 8000
rect 33955 7959 34013 7960
rect 34819 8000 34877 8001
rect 34819 7960 34828 8000
rect 34868 7960 34877 8000
rect 34819 7959 34877 7960
rect 36355 8000 36413 8001
rect 36355 7960 36364 8000
rect 36404 7960 36413 8000
rect 36355 7959 36413 7960
rect 36555 8000 36597 8009
rect 36555 7960 36556 8000
rect 36596 7960 36597 8000
rect 36555 7951 36597 7960
rect 36931 8000 36989 8001
rect 36931 7960 36940 8000
rect 36980 7960 36989 8000
rect 36931 7959 36989 7960
rect 37795 8000 37853 8001
rect 37795 7960 37804 8000
rect 37844 7960 37853 8000
rect 37795 7959 37853 7960
rect 6115 7941 6173 7942
rect 6115 7901 6124 7941
rect 6164 7901 6173 7941
rect 30280 7936 30322 7945
rect 6115 7900 6173 7901
rect 13795 7916 13853 7917
rect 13795 7876 13804 7916
rect 13844 7876 13853 7916
rect 13795 7875 13853 7876
rect 19947 7916 19989 7925
rect 19947 7876 19948 7916
rect 19988 7876 19989 7916
rect 19947 7867 19989 7876
rect 24939 7916 24981 7925
rect 24939 7876 24940 7916
rect 24980 7876 24981 7916
rect 24939 7867 24981 7876
rect 29163 7916 29205 7925
rect 29163 7876 29164 7916
rect 29204 7876 29205 7916
rect 29163 7867 29205 7876
rect 29355 7916 29397 7925
rect 29355 7876 29356 7916
rect 29396 7876 29397 7916
rect 29355 7867 29397 7876
rect 31179 7916 31221 7925
rect 31179 7876 31180 7916
rect 31220 7876 31221 7916
rect 31179 7867 31221 7876
rect 31371 7916 31413 7925
rect 31371 7876 31372 7916
rect 31412 7876 31413 7916
rect 31371 7867 31413 7876
rect 2859 7832 2901 7841
rect 2859 7792 2860 7832
rect 2900 7792 2901 7832
rect 2859 7783 2901 7792
rect 4683 7832 4725 7841
rect 4683 7792 4684 7832
rect 4724 7792 4725 7832
rect 4683 7783 4725 7792
rect 9867 7832 9909 7841
rect 9867 7792 9868 7832
rect 9908 7792 9909 7832
rect 9867 7783 9909 7792
rect 11403 7832 11445 7841
rect 11403 7792 11404 7832
rect 11444 7792 11445 7832
rect 11403 7783 11445 7792
rect 29259 7832 29301 7841
rect 29259 7792 29260 7832
rect 29300 7792 29301 7832
rect 29259 7783 29301 7792
rect 31275 7832 31317 7841
rect 31275 7792 31276 7832
rect 31316 7792 31317 7832
rect 31275 7783 31317 7792
rect 33771 7832 33813 7841
rect 33771 7792 33772 7832
rect 33812 7792 33813 7832
rect 33771 7783 33813 7792
rect 3811 7748 3869 7749
rect 3811 7708 3820 7748
rect 3860 7708 3869 7748
rect 3811 7707 3869 7708
rect 6787 7748 6845 7749
rect 6787 7708 6796 7748
rect 6836 7708 6845 7748
rect 6787 7707 6845 7708
rect 7755 7748 7797 7757
rect 7755 7708 7756 7748
rect 7796 7708 7797 7748
rect 7755 7699 7797 7708
rect 10251 7748 10293 7757
rect 10251 7708 10252 7748
rect 10292 7708 10293 7748
rect 10251 7699 10293 7708
rect 21483 7748 21525 7757
rect 21483 7708 21484 7748
rect 21524 7708 21525 7748
rect 21483 7699 21525 7708
rect 22339 7748 22397 7749
rect 22339 7708 22348 7748
rect 22388 7708 22397 7748
rect 22339 7707 22397 7708
rect 24075 7748 24117 7757
rect 24075 7708 24076 7748
rect 24116 7708 24117 7748
rect 24075 7699 24117 7708
rect 25227 7748 25269 7757
rect 25227 7708 25228 7748
rect 25268 7708 25269 7748
rect 25227 7699 25269 7708
rect 33195 7748 33237 7757
rect 33195 7708 33196 7748
rect 33236 7708 33237 7748
rect 33195 7699 33237 7708
rect 35491 7748 35549 7749
rect 35491 7708 35500 7748
rect 35540 7708 35549 7748
rect 35491 7707 35549 7708
rect 38955 7748 38997 7757
rect 38955 7708 38956 7748
rect 38996 7708 38997 7748
rect 38955 7699 38997 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 4779 7412 4821 7421
rect 4779 7372 4780 7412
rect 4820 7372 4821 7412
rect 4779 7363 4821 7372
rect 5827 7412 5885 7413
rect 5827 7372 5836 7412
rect 5876 7372 5885 7412
rect 5827 7371 5885 7372
rect 6987 7412 7029 7421
rect 6987 7372 6988 7412
rect 7028 7372 7029 7412
rect 6987 7363 7029 7372
rect 8139 7412 8181 7421
rect 8139 7372 8140 7412
rect 8180 7372 8181 7412
rect 8139 7363 8181 7372
rect 13035 7412 13077 7421
rect 13035 7372 13036 7412
rect 13076 7372 13077 7412
rect 13035 7363 13077 7372
rect 22059 7412 22101 7421
rect 22059 7372 22060 7412
rect 22100 7372 22101 7412
rect 22059 7363 22101 7372
rect 24171 7412 24213 7421
rect 24171 7372 24172 7412
rect 24212 7372 24213 7412
rect 24171 7363 24213 7372
rect 26667 7412 26709 7421
rect 26667 7372 26668 7412
rect 26708 7372 26709 7412
rect 26667 7363 26709 7372
rect 31179 7412 31221 7421
rect 31179 7372 31180 7412
rect 31220 7372 31221 7412
rect 31179 7363 31221 7372
rect 31563 7412 31605 7421
rect 31563 7372 31564 7412
rect 31604 7372 31605 7412
rect 31563 7363 31605 7372
rect 33771 7412 33813 7421
rect 33771 7372 33772 7412
rect 33812 7372 33813 7412
rect 33771 7363 33813 7372
rect 36547 7412 36605 7413
rect 36547 7372 36556 7412
rect 36596 7372 36605 7412
rect 36547 7371 36605 7372
rect 37411 7412 37469 7413
rect 37411 7372 37420 7412
rect 37460 7372 37469 7412
rect 37411 7371 37469 7372
rect 10059 7328 10101 7337
rect 10059 7288 10060 7328
rect 10100 7288 10101 7328
rect 10059 7279 10101 7288
rect 14475 7328 14517 7337
rect 14475 7288 14476 7328
rect 14516 7288 14517 7328
rect 14475 7279 14517 7288
rect 15435 7328 15477 7337
rect 15435 7288 15436 7328
rect 15476 7288 15477 7328
rect 15435 7279 15477 7288
rect 16491 7328 16533 7337
rect 16491 7288 16492 7328
rect 16532 7288 16533 7328
rect 16491 7279 16533 7288
rect 29259 7328 29301 7337
rect 29259 7288 29260 7328
rect 29300 7288 29301 7328
rect 29259 7279 29301 7288
rect 10723 7244 10781 7245
rect 10723 7204 10732 7244
rect 10772 7204 10781 7244
rect 10723 7203 10781 7204
rect 14379 7244 14421 7253
rect 14379 7204 14380 7244
rect 14420 7204 14421 7244
rect 14379 7195 14421 7204
rect 29643 7244 29685 7253
rect 29643 7204 29644 7244
rect 29684 7204 29685 7244
rect 29643 7195 29685 7204
rect 23464 7175 23506 7184
rect 2379 7160 2421 7169
rect 2379 7120 2380 7160
rect 2420 7120 2421 7160
rect 2379 7111 2421 7120
rect 2755 7160 2813 7161
rect 2755 7120 2764 7160
rect 2804 7120 2813 7160
rect 2755 7119 2813 7120
rect 3619 7160 3677 7161
rect 3619 7120 3628 7160
rect 3668 7120 3677 7160
rect 3619 7119 3677 7120
rect 5155 7160 5213 7161
rect 5155 7120 5164 7160
rect 5204 7120 5213 7160
rect 5155 7119 5213 7120
rect 6211 7160 6269 7161
rect 6211 7120 6220 7160
rect 6260 7120 6269 7160
rect 6211 7119 6269 7120
rect 6499 7160 6557 7161
rect 6499 7120 6508 7160
rect 6548 7120 6557 7160
rect 6499 7119 6557 7120
rect 7459 7160 7517 7161
rect 7459 7120 7468 7160
rect 7508 7120 7517 7160
rect 7459 7119 7517 7120
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 8139 7160 8181 7169
rect 8139 7120 8140 7160
rect 8180 7120 8181 7160
rect 8139 7111 8181 7120
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 8427 7160 8469 7169
rect 8427 7120 8428 7160
rect 8468 7120 8469 7160
rect 8427 7111 8469 7120
rect 8803 7160 8861 7161
rect 8803 7120 8812 7160
rect 8852 7120 8861 7160
rect 8803 7119 8861 7120
rect 8899 7160 8957 7161
rect 8899 7120 8908 7160
rect 8948 7120 8957 7160
rect 8899 7119 8957 7120
rect 9099 7160 9141 7169
rect 9099 7120 9100 7160
rect 9140 7120 9141 7160
rect 9099 7111 9141 7120
rect 9195 7160 9237 7169
rect 9195 7120 9196 7160
rect 9236 7120 9237 7160
rect 9195 7111 9237 7120
rect 9288 7160 9346 7161
rect 9288 7120 9297 7160
rect 9337 7120 9346 7160
rect 9288 7119 9346 7120
rect 9667 7160 9725 7161
rect 9667 7120 9676 7160
rect 9716 7120 9725 7160
rect 9667 7119 9725 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 10251 7160 10293 7169
rect 10251 7120 10252 7160
rect 10292 7120 10293 7160
rect 10251 7111 10293 7120
rect 10347 7160 10389 7169
rect 10347 7120 10348 7160
rect 10388 7120 10389 7160
rect 10347 7111 10389 7120
rect 11307 7160 11349 7169
rect 11307 7120 11308 7160
rect 11348 7120 11349 7160
rect 11307 7111 11349 7120
rect 11403 7160 11445 7169
rect 11403 7120 11404 7160
rect 11444 7120 11445 7160
rect 11403 7111 11445 7120
rect 11787 7160 11829 7169
rect 11787 7120 11788 7160
rect 11828 7120 11829 7160
rect 11787 7111 11829 7120
rect 11883 7160 11925 7169
rect 11883 7120 11884 7160
rect 11924 7120 11925 7160
rect 11883 7111 11925 7120
rect 12355 7160 12413 7161
rect 12355 7120 12364 7160
rect 12404 7120 12413 7160
rect 12355 7119 12413 7120
rect 13603 7160 13661 7161
rect 13603 7120 13612 7160
rect 13652 7120 13661 7160
rect 13603 7119 13661 7120
rect 14179 7160 14237 7161
rect 14179 7120 14188 7160
rect 14228 7120 14237 7160
rect 14179 7119 14237 7120
rect 14283 7160 14325 7169
rect 14283 7120 14284 7160
rect 14324 7120 14325 7160
rect 14283 7111 14325 7120
rect 14763 7160 14805 7169
rect 14763 7120 14764 7160
rect 14804 7120 14805 7160
rect 14763 7111 14805 7120
rect 15051 7160 15093 7169
rect 15051 7120 15052 7160
rect 15092 7120 15093 7160
rect 15051 7111 15093 7120
rect 15619 7160 15677 7161
rect 15619 7120 15628 7160
rect 15668 7120 15677 7160
rect 15619 7119 15677 7120
rect 17539 7160 17597 7161
rect 17539 7120 17548 7160
rect 17588 7120 17597 7160
rect 17539 7119 17597 7120
rect 17827 7160 17885 7161
rect 17827 7120 17836 7160
rect 17876 7120 17885 7160
rect 17827 7119 17885 7120
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 19363 7160 19421 7161
rect 19363 7120 19372 7160
rect 19412 7120 19421 7160
rect 19363 7119 19421 7120
rect 20227 7160 20285 7161
rect 20227 7120 20236 7160
rect 20276 7120 20285 7160
rect 20227 7119 20285 7120
rect 22443 7160 22485 7169
rect 22443 7120 22444 7160
rect 22484 7120 22485 7160
rect 22443 7111 22485 7120
rect 22915 7160 22973 7161
rect 22915 7120 22924 7160
rect 22964 7120 22973 7160
rect 22915 7119 22973 7120
rect 23011 7160 23069 7161
rect 23011 7120 23020 7160
rect 23060 7120 23069 7160
rect 23011 7119 23069 7120
rect 23211 7160 23253 7169
rect 23211 7120 23212 7160
rect 23252 7120 23253 7160
rect 23211 7111 23253 7120
rect 23307 7160 23349 7169
rect 23307 7120 23308 7160
rect 23348 7120 23349 7160
rect 23464 7135 23465 7175
rect 23505 7135 23506 7175
rect 24712 7175 24754 7184
rect 23464 7126 23506 7135
rect 23691 7160 23733 7169
rect 23307 7111 23349 7120
rect 23691 7120 23692 7160
rect 23732 7120 23733 7160
rect 23691 7111 23733 7120
rect 23787 7160 23829 7169
rect 23787 7120 23788 7160
rect 23828 7120 23829 7160
rect 23787 7111 23829 7120
rect 24163 7160 24221 7161
rect 24163 7120 24172 7160
rect 24212 7120 24221 7160
rect 24163 7119 24221 7120
rect 24259 7160 24317 7161
rect 24259 7120 24268 7160
rect 24308 7120 24317 7160
rect 24259 7119 24317 7120
rect 24459 7160 24501 7169
rect 24459 7120 24460 7160
rect 24500 7120 24501 7160
rect 24459 7111 24501 7120
rect 24555 7160 24597 7169
rect 24555 7120 24556 7160
rect 24596 7120 24597 7160
rect 24712 7135 24713 7175
rect 24753 7135 24754 7175
rect 24712 7126 24754 7135
rect 25227 7160 25269 7169
rect 24555 7111 24597 7120
rect 25227 7120 25228 7160
rect 25268 7120 25269 7160
rect 25227 7111 25269 7120
rect 25419 7160 25461 7169
rect 25419 7120 25420 7160
rect 25460 7120 25461 7160
rect 25419 7111 25461 7120
rect 25515 7160 25557 7169
rect 25515 7120 25516 7160
rect 25556 7120 25557 7160
rect 25515 7111 25557 7120
rect 25899 7160 25941 7169
rect 25899 7120 25900 7160
rect 25940 7120 25941 7160
rect 25899 7111 25941 7120
rect 25995 7160 26037 7169
rect 25995 7120 25996 7160
rect 26036 7120 26037 7160
rect 25995 7111 26037 7120
rect 26187 7160 26229 7169
rect 26187 7120 26188 7160
rect 26228 7120 26229 7160
rect 26187 7111 26229 7120
rect 26283 7160 26325 7169
rect 26283 7120 26284 7160
rect 26324 7120 26325 7160
rect 26283 7111 26325 7120
rect 26379 7160 26421 7169
rect 26379 7120 26380 7160
rect 26420 7120 26421 7160
rect 26379 7111 26421 7120
rect 26659 7160 26717 7161
rect 26659 7120 26668 7160
rect 26708 7120 26717 7160
rect 26659 7119 26717 7120
rect 26755 7160 26813 7161
rect 26755 7120 26764 7160
rect 26804 7120 26813 7160
rect 26755 7119 26813 7120
rect 26955 7160 26997 7169
rect 26955 7120 26956 7160
rect 26996 7120 26997 7160
rect 26955 7111 26997 7120
rect 27051 7160 27093 7169
rect 27051 7120 27052 7160
rect 27092 7120 27093 7160
rect 27051 7111 27093 7120
rect 27198 7160 27256 7161
rect 27198 7120 27207 7160
rect 27247 7120 27256 7160
rect 27198 7119 27256 7120
rect 28011 7160 28053 7169
rect 28011 7120 28012 7160
rect 28052 7120 28053 7160
rect 28011 7111 28053 7120
rect 28107 7160 28149 7169
rect 28107 7120 28108 7160
rect 28148 7120 28149 7160
rect 28107 7111 28149 7120
rect 28203 7160 28245 7169
rect 28203 7120 28204 7160
rect 28244 7120 28245 7160
rect 28203 7111 28245 7120
rect 28683 7160 28725 7169
rect 28683 7120 28684 7160
rect 28724 7120 28725 7160
rect 28683 7111 28725 7120
rect 28779 7160 28821 7169
rect 28779 7120 28780 7160
rect 28820 7120 28821 7160
rect 28779 7111 28821 7120
rect 28971 7160 29013 7169
rect 28971 7120 28972 7160
rect 29012 7120 29013 7160
rect 28971 7111 29013 7120
rect 29259 7160 29301 7169
rect 29259 7120 29260 7160
rect 29300 7120 29301 7160
rect 29259 7111 29301 7120
rect 29451 7160 29493 7169
rect 29451 7120 29452 7160
rect 29492 7120 29493 7160
rect 29451 7111 29493 7120
rect 29739 7160 29781 7169
rect 29739 7120 29740 7160
rect 29780 7120 29781 7160
rect 29739 7111 29781 7120
rect 30123 7160 30165 7169
rect 30123 7120 30124 7160
rect 30164 7120 30165 7160
rect 30123 7111 30165 7120
rect 30219 7160 30261 7169
rect 30219 7120 30220 7160
rect 30260 7120 30261 7160
rect 30219 7111 30261 7120
rect 31267 7160 31325 7161
rect 31267 7120 31276 7160
rect 31316 7120 31325 7160
rect 31267 7119 31325 7120
rect 31651 7160 31709 7161
rect 31651 7120 31660 7160
rect 31700 7120 31709 7160
rect 31651 7119 31709 7120
rect 32515 7160 32573 7161
rect 32515 7120 32524 7160
rect 32564 7120 32573 7160
rect 32515 7119 32573 7120
rect 34915 7160 34973 7161
rect 34915 7120 34924 7160
rect 34964 7120 34973 7160
rect 34915 7119 34973 7120
rect 35779 7160 35837 7161
rect 35779 7120 35788 7160
rect 35828 7120 35837 7160
rect 35779 7119 35837 7120
rect 36171 7160 36213 7169
rect 36171 7120 36172 7160
rect 36212 7120 36213 7160
rect 36171 7111 36213 7120
rect 37219 7160 37277 7161
rect 37219 7120 37228 7160
rect 37268 7120 37277 7160
rect 37219 7119 37277 7120
rect 38083 7160 38141 7161
rect 38083 7120 38092 7160
rect 38132 7120 38141 7160
rect 38083 7119 38141 7120
rect 643 6992 701 6993
rect 643 6952 652 6992
rect 692 6952 701 6992
rect 643 6951 701 6952
rect 5827 6992 5885 6993
rect 5827 6952 5836 6992
rect 5876 6952 5885 6992
rect 5827 6951 5885 6952
rect 6019 6992 6077 6993
rect 6019 6952 6028 6992
rect 6068 6952 6077 6992
rect 6019 6951 6077 6952
rect 6307 6992 6365 6993
rect 6307 6952 6316 6992
rect 6356 6952 6365 6992
rect 6307 6951 6365 6952
rect 8043 6992 8085 7001
rect 8043 6952 8044 6992
rect 8084 6952 8085 6992
rect 8043 6943 8085 6952
rect 8611 6992 8669 6993
rect 8611 6952 8620 6992
rect 8660 6952 8669 6992
rect 8611 6951 8669 6952
rect 9283 6992 9341 6993
rect 9283 6952 9292 6992
rect 9332 6952 9341 6992
rect 9283 6951 9341 6952
rect 9579 6988 9621 6997
rect 9579 6948 9580 6988
rect 9620 6948 9621 6988
rect 10531 6992 10589 6993
rect 10531 6952 10540 6992
rect 10580 6952 10589 6992
rect 10531 6951 10589 6952
rect 11587 6992 11645 6993
rect 11587 6952 11596 6992
rect 11636 6952 11645 6992
rect 11587 6951 11645 6952
rect 12067 6992 12125 6993
rect 12067 6952 12076 6992
rect 12116 6952 12125 6992
rect 12067 6951 12125 6952
rect 13507 6992 13565 6993
rect 13507 6952 13516 6992
rect 13556 6952 13565 6992
rect 13507 6951 13565 6952
rect 13795 6992 13853 6993
rect 13795 6952 13804 6992
rect 13844 6952 13853 6992
rect 13795 6951 13853 6952
rect 14283 6992 14325 7001
rect 14283 6952 14284 6992
rect 14324 6952 14325 6992
rect 9579 6939 9621 6948
rect 14283 6943 14325 6952
rect 14955 6992 14997 7001
rect 14955 6952 14956 6992
rect 14996 6952 14997 6992
rect 14955 6943 14997 6952
rect 16291 6992 16349 6993
rect 16291 6952 16300 6992
rect 16340 6952 16349 6992
rect 16291 6951 16349 6952
rect 16867 6992 16925 6993
rect 16867 6952 16876 6992
rect 16916 6952 16925 6992
rect 16867 6951 16925 6952
rect 17739 6992 17781 7001
rect 17739 6952 17740 6992
rect 17780 6952 17781 6992
rect 17739 6943 17781 6952
rect 21379 6992 21437 6993
rect 21379 6952 21388 6992
rect 21428 6952 21437 6992
rect 21379 6951 21437 6952
rect 23395 6992 23453 6993
rect 23395 6952 23404 6992
rect 23444 6952 23453 6992
rect 23395 6951 23453 6952
rect 23971 6992 24029 6993
rect 23971 6952 23980 6992
rect 24020 6952 24029 6992
rect 23971 6951 24029 6952
rect 25699 6992 25757 6993
rect 25699 6952 25708 6992
rect 25748 6952 25757 6992
rect 25699 6951 25757 6952
rect 26467 6992 26525 6993
rect 26467 6952 26476 6992
rect 26516 6952 26525 6992
rect 26467 6951 26525 6952
rect 28291 6992 28349 6993
rect 28291 6952 28300 6992
rect 28340 6952 28349 6992
rect 28291 6951 28349 6952
rect 28483 6992 28541 6993
rect 28483 6952 28492 6992
rect 28532 6952 28541 6992
rect 28483 6951 28541 6952
rect 29923 6992 29981 6993
rect 29923 6952 29932 6992
rect 29972 6952 29981 6992
rect 29923 6951 29981 6952
rect 31843 6992 31901 6993
rect 31843 6952 31852 6992
rect 31892 6952 31901 6992
rect 31843 6951 31901 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 15051 6714 15093 6723
rect 15051 6674 15052 6714
rect 15092 6674 15093 6714
rect 15051 6665 15093 6674
rect 8427 6656 8469 6665
rect 8427 6616 8428 6656
rect 8468 6616 8469 6656
rect 8427 6607 8469 6616
rect 8707 6656 8765 6657
rect 8707 6616 8716 6656
rect 8756 6616 8765 6656
rect 8707 6615 8765 6616
rect 10051 6656 10109 6657
rect 10051 6616 10060 6656
rect 10100 6616 10109 6656
rect 10051 6615 10109 6616
rect 12355 6656 12413 6657
rect 12355 6616 12364 6656
rect 12404 6616 12413 6656
rect 12355 6615 12413 6616
rect 13123 6656 13181 6657
rect 13123 6616 13132 6656
rect 13172 6616 13181 6656
rect 13123 6615 13181 6616
rect 13227 6656 13269 6665
rect 13227 6616 13228 6656
rect 13268 6616 13269 6656
rect 13227 6607 13269 6616
rect 14179 6656 14237 6657
rect 14179 6616 14188 6656
rect 14228 6616 14237 6656
rect 14179 6615 14237 6616
rect 15331 6656 15389 6657
rect 15331 6616 15340 6656
rect 15380 6616 15389 6656
rect 15331 6615 15389 6616
rect 22155 6656 22197 6665
rect 22155 6616 22156 6656
rect 22196 6616 22197 6656
rect 22155 6607 22197 6616
rect 23107 6656 23165 6657
rect 23107 6616 23116 6656
rect 23156 6616 23165 6656
rect 23107 6615 23165 6616
rect 23499 6656 23541 6665
rect 23499 6616 23500 6656
rect 23540 6616 23541 6656
rect 23499 6607 23541 6616
rect 23883 6656 23925 6665
rect 23883 6616 23884 6656
rect 23924 6616 23925 6656
rect 23883 6607 23925 6616
rect 24451 6656 24509 6657
rect 24451 6616 24460 6656
rect 24500 6616 24509 6656
rect 24451 6615 24509 6616
rect 25987 6656 26045 6657
rect 25987 6616 25996 6656
rect 26036 6616 26045 6656
rect 25987 6615 26045 6616
rect 26563 6656 26621 6657
rect 26563 6616 26572 6656
rect 26612 6616 26621 6656
rect 26563 6615 26621 6616
rect 27139 6656 27197 6657
rect 27139 6616 27148 6656
rect 27188 6616 27197 6656
rect 27139 6615 27197 6616
rect 28299 6656 28341 6665
rect 28299 6616 28300 6656
rect 28340 6616 28341 6656
rect 28299 6607 28341 6616
rect 35299 6656 35357 6657
rect 35299 6616 35308 6656
rect 35348 6616 35357 6656
rect 35299 6615 35357 6616
rect 9955 6572 10013 6573
rect 9955 6532 9964 6572
rect 10004 6532 10013 6572
rect 9955 6531 10013 6532
rect 13027 6572 13085 6573
rect 13027 6532 13036 6572
rect 13076 6532 13085 6572
rect 13027 6531 13085 6532
rect 15723 6572 15765 6581
rect 15723 6532 15724 6572
rect 15764 6532 15765 6572
rect 15723 6523 15765 6532
rect 21859 6572 21917 6573
rect 21859 6532 21868 6572
rect 21908 6532 21917 6572
rect 21859 6531 21917 6532
rect 25891 6572 25949 6573
rect 25891 6532 25900 6572
rect 25940 6532 25949 6572
rect 25891 6531 25949 6532
rect 26467 6572 26525 6573
rect 26467 6532 26476 6572
rect 26516 6532 26525 6572
rect 26467 6531 26525 6532
rect 29923 6572 29981 6573
rect 29923 6532 29932 6572
rect 29972 6532 29981 6572
rect 29923 6531 29981 6532
rect 3723 6488 3765 6497
rect 3723 6448 3724 6488
rect 3764 6448 3765 6488
rect 3723 6439 3765 6448
rect 4099 6488 4157 6489
rect 4099 6448 4108 6488
rect 4148 6448 4157 6488
rect 4099 6447 4157 6448
rect 4963 6488 5021 6489
rect 4963 6448 4972 6488
rect 5012 6448 5021 6488
rect 4963 6447 5021 6448
rect 6211 6488 6269 6489
rect 6211 6448 6220 6488
rect 6260 6448 6269 6488
rect 7467 6488 7509 6497
rect 6211 6447 6269 6448
rect 6403 6475 6461 6476
rect 6403 6435 6412 6475
rect 6452 6435 6461 6475
rect 7467 6448 7468 6488
rect 7508 6448 7509 6488
rect 7467 6439 7509 6448
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 7659 6488 7701 6497
rect 7659 6448 7660 6488
rect 7700 6448 7701 6488
rect 7659 6439 7701 6448
rect 7755 6488 7797 6497
rect 7755 6448 7756 6488
rect 7796 6448 7797 6488
rect 7755 6439 7797 6448
rect 8235 6488 8277 6497
rect 8235 6448 8236 6488
rect 8276 6448 8277 6488
rect 8235 6439 8277 6448
rect 8523 6488 8565 6497
rect 8523 6448 8524 6488
rect 8564 6448 8565 6488
rect 8523 6439 8565 6448
rect 8907 6488 8949 6497
rect 8907 6448 8908 6488
rect 8948 6448 8949 6488
rect 8907 6439 8949 6448
rect 9003 6488 9045 6497
rect 9003 6448 9004 6488
rect 9044 6448 9045 6488
rect 9003 6439 9045 6448
rect 9187 6488 9245 6489
rect 9187 6448 9196 6488
rect 9236 6448 9245 6488
rect 9187 6447 9245 6448
rect 9291 6488 9333 6497
rect 9291 6448 9292 6488
rect 9332 6448 9333 6488
rect 9291 6439 9333 6448
rect 9771 6488 9813 6497
rect 9771 6448 9772 6488
rect 9812 6448 9813 6488
rect 9771 6439 9813 6448
rect 9867 6488 9909 6497
rect 9867 6448 9868 6488
rect 9908 6448 9909 6488
rect 9867 6439 9909 6448
rect 10339 6488 10397 6489
rect 10339 6448 10348 6488
rect 10388 6448 10397 6488
rect 10339 6447 10397 6448
rect 10539 6488 10581 6497
rect 10539 6448 10540 6488
rect 10580 6448 10581 6488
rect 10539 6439 10581 6448
rect 10627 6488 10685 6489
rect 10627 6448 10636 6488
rect 10676 6448 10685 6488
rect 10627 6447 10685 6448
rect 10915 6488 10973 6489
rect 10915 6448 10924 6488
rect 10964 6448 10973 6488
rect 10915 6447 10973 6448
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12651 6488 12693 6497
rect 12651 6448 12652 6488
rect 12692 6448 12693 6488
rect 12651 6439 12693 6448
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12843 6439 12885 6448
rect 12939 6488 12981 6497
rect 12939 6448 12940 6488
rect 12980 6448 12981 6488
rect 12939 6439 12981 6448
rect 13699 6488 13757 6489
rect 13699 6448 13708 6488
rect 13748 6448 13757 6488
rect 13699 6447 13757 6448
rect 13795 6488 13853 6489
rect 13795 6448 13804 6488
rect 13844 6448 13853 6488
rect 13795 6447 13853 6448
rect 13995 6488 14037 6497
rect 13995 6448 13996 6488
rect 14036 6448 14037 6488
rect 13995 6439 14037 6448
rect 14091 6488 14133 6497
rect 14091 6448 14092 6488
rect 14132 6448 14133 6488
rect 14091 6439 14133 6448
rect 14184 6488 14242 6489
rect 14184 6448 14193 6488
rect 14233 6448 14242 6488
rect 14184 6447 14242 6448
rect 14859 6488 14901 6497
rect 14859 6448 14860 6488
rect 14900 6448 14901 6488
rect 14859 6439 14901 6448
rect 14947 6488 15005 6489
rect 14947 6448 14956 6488
rect 14996 6448 15005 6488
rect 14947 6447 15005 6448
rect 15243 6488 15285 6497
rect 15243 6448 15244 6488
rect 15284 6448 15285 6488
rect 15243 6439 15285 6448
rect 15435 6488 15477 6497
rect 15435 6448 15436 6488
rect 15476 6448 15477 6488
rect 15435 6439 15477 6448
rect 15523 6488 15581 6489
rect 15523 6448 15532 6488
rect 15572 6448 15581 6488
rect 15523 6447 15581 6448
rect 16099 6488 16157 6489
rect 16099 6448 16108 6488
rect 16148 6448 16157 6488
rect 16099 6447 16157 6448
rect 16963 6488 17021 6489
rect 16963 6448 16972 6488
rect 17012 6448 17021 6488
rect 16963 6447 17021 6448
rect 19555 6488 19613 6489
rect 19555 6448 19564 6488
rect 19604 6448 19613 6488
rect 19555 6447 19613 6448
rect 20995 6488 21053 6489
rect 20995 6448 21004 6488
rect 21044 6448 21053 6488
rect 20995 6447 21053 6448
rect 22243 6488 22301 6489
rect 22243 6448 22252 6488
rect 22292 6448 22301 6488
rect 22243 6447 22301 6448
rect 22435 6488 22493 6489
rect 22435 6448 22444 6488
rect 22484 6448 22493 6488
rect 22435 6447 22493 6448
rect 23691 6488 23733 6497
rect 23691 6448 23692 6488
rect 23732 6448 23733 6488
rect 23691 6439 23733 6448
rect 23979 6488 24021 6497
rect 23979 6448 23980 6488
rect 24020 6448 24021 6488
rect 23979 6439 24021 6448
rect 24171 6488 24213 6497
rect 24171 6448 24172 6488
rect 24212 6448 24213 6488
rect 24171 6439 24213 6448
rect 24267 6488 24309 6497
rect 24267 6448 24268 6488
rect 24308 6448 24309 6488
rect 24267 6439 24309 6448
rect 24643 6488 24701 6489
rect 24643 6448 24652 6488
rect 24692 6448 24701 6488
rect 24643 6447 24701 6448
rect 24747 6488 24789 6497
rect 24747 6448 24748 6488
rect 24788 6448 24789 6488
rect 24747 6439 24789 6448
rect 24939 6488 24981 6497
rect 24939 6448 24940 6488
rect 24980 6448 24981 6488
rect 24939 6439 24981 6448
rect 25123 6488 25181 6489
rect 25123 6448 25132 6488
rect 25172 6448 25181 6488
rect 25123 6447 25181 6448
rect 25515 6488 25557 6497
rect 25515 6448 25516 6488
rect 25556 6448 25557 6488
rect 25515 6439 25557 6448
rect 25707 6488 25749 6497
rect 25707 6448 25708 6488
rect 25748 6448 25749 6488
rect 25707 6439 25749 6448
rect 25803 6488 25845 6497
rect 25803 6448 25804 6488
rect 25844 6448 25845 6488
rect 25803 6439 25845 6448
rect 26283 6488 26325 6497
rect 26283 6448 26284 6488
rect 26324 6448 26325 6488
rect 26283 6439 26325 6448
rect 26379 6488 26421 6497
rect 26379 6448 26380 6488
rect 26420 6448 26421 6488
rect 26379 6439 26421 6448
rect 26859 6488 26901 6497
rect 26859 6448 26860 6488
rect 26900 6448 26901 6488
rect 26859 6439 26901 6448
rect 26955 6488 26997 6497
rect 26955 6448 26956 6488
rect 26996 6448 26997 6488
rect 26955 6439 26997 6448
rect 28387 6488 28445 6489
rect 28387 6448 28396 6488
rect 28436 6448 28445 6488
rect 28387 6447 28445 6448
rect 28587 6488 28629 6497
rect 28587 6448 28588 6488
rect 28628 6448 28629 6488
rect 28587 6439 28629 6448
rect 28779 6488 28821 6497
rect 28779 6448 28780 6488
rect 28820 6448 28821 6488
rect 28779 6439 28821 6448
rect 28963 6488 29021 6489
rect 28963 6448 28972 6488
rect 29012 6448 29021 6488
rect 28963 6447 29021 6448
rect 29067 6488 29109 6497
rect 29067 6448 29068 6488
rect 29108 6448 29109 6488
rect 29067 6439 29109 6448
rect 29259 6488 29301 6497
rect 29259 6448 29260 6488
rect 29300 6448 29301 6488
rect 29259 6439 29301 6448
rect 29443 6488 29501 6489
rect 29443 6448 29452 6488
rect 29492 6448 29501 6488
rect 29443 6447 29501 6448
rect 29731 6488 29789 6489
rect 29731 6448 29740 6488
rect 29780 6448 29789 6488
rect 29731 6447 29789 6448
rect 30211 6488 30269 6489
rect 30211 6448 30220 6488
rect 30260 6448 30269 6488
rect 30211 6447 30269 6448
rect 30891 6488 30933 6497
rect 30891 6448 30892 6488
rect 30932 6448 30933 6488
rect 30891 6439 30933 6448
rect 31083 6488 31125 6497
rect 31083 6448 31084 6488
rect 31124 6448 31125 6488
rect 31083 6439 31125 6448
rect 31459 6488 31517 6489
rect 31459 6448 31468 6488
rect 31508 6448 31517 6488
rect 31459 6447 31517 6448
rect 32323 6488 32381 6489
rect 32323 6448 32332 6488
rect 32372 6448 32381 6488
rect 32323 6447 32381 6448
rect 33483 6488 33525 6497
rect 33483 6448 33484 6488
rect 33524 6448 33525 6488
rect 33483 6439 33525 6448
rect 34435 6488 34493 6489
rect 34435 6448 34444 6488
rect 34484 6448 34493 6488
rect 34435 6447 34493 6448
rect 34627 6488 34685 6489
rect 34627 6448 34636 6488
rect 34676 6448 34685 6488
rect 34627 6447 34685 6448
rect 35499 6488 35541 6497
rect 35499 6448 35500 6488
rect 35540 6448 35541 6488
rect 35499 6439 35541 6448
rect 35875 6488 35933 6489
rect 35875 6448 35884 6488
rect 35924 6448 35933 6488
rect 35875 6447 35933 6448
rect 36739 6488 36797 6489
rect 36739 6448 36748 6488
rect 36788 6448 36797 6488
rect 36739 6447 36797 6448
rect 37899 6488 37941 6497
rect 37899 6448 37900 6488
rect 37940 6448 37941 6488
rect 37899 6439 37941 6448
rect 6403 6434 6461 6435
rect 9387 6404 9429 6413
rect 9387 6364 9388 6404
rect 9428 6364 9429 6404
rect 9387 6355 9429 6364
rect 18787 6404 18845 6405
rect 18787 6364 18796 6404
rect 18836 6364 18845 6404
rect 18787 6363 18845 6364
rect 23299 6404 23357 6405
rect 23299 6364 23308 6404
rect 23348 6364 23357 6404
rect 23299 6363 23357 6364
rect 25227 6404 25269 6413
rect 25227 6364 25228 6404
rect 25268 6364 25269 6404
rect 25227 6355 25269 6364
rect 25419 6404 25461 6413
rect 25419 6364 25420 6404
rect 25460 6364 25461 6404
rect 25419 6355 25461 6364
rect 7075 6320 7133 6321
rect 7075 6280 7084 6320
rect 7124 6280 7133 6320
rect 7075 6279 7133 6280
rect 9483 6320 9525 6329
rect 9483 6280 9484 6320
rect 9524 6280 9525 6320
rect 9483 6271 9525 6280
rect 11211 6320 11253 6329
rect 11211 6280 11212 6320
rect 11252 6280 11253 6320
rect 11211 6271 11253 6280
rect 14571 6320 14613 6329
rect 14571 6280 14572 6320
rect 14612 6280 14613 6320
rect 14571 6271 14613 6280
rect 18115 6320 18173 6321
rect 18115 6280 18124 6320
rect 18164 6280 18173 6320
rect 18115 6279 18173 6280
rect 18411 6320 18453 6329
rect 18411 6280 18412 6320
rect 18452 6280 18453 6320
rect 18411 6271 18453 6280
rect 24939 6320 24981 6329
rect 24939 6280 24940 6320
rect 24980 6280 24981 6320
rect 24939 6271 24981 6280
rect 25323 6320 25365 6329
rect 25323 6280 25324 6320
rect 25364 6280 25365 6320
rect 25323 6271 25365 6280
rect 26571 6320 26613 6329
rect 26571 6280 26572 6320
rect 26612 6280 26613 6320
rect 26571 6271 26613 6280
rect 7267 6236 7325 6237
rect 7267 6196 7276 6236
rect 7316 6196 7325 6236
rect 7267 6195 7325 6196
rect 9579 6236 9621 6245
rect 9579 6196 9580 6236
rect 9620 6196 9621 6236
rect 9579 6187 9621 6196
rect 10059 6236 10101 6245
rect 10059 6196 10060 6236
rect 10100 6196 10101 6236
rect 10059 6187 10101 6196
rect 10539 6236 10581 6245
rect 10539 6196 10540 6236
rect 10580 6196 10581 6236
rect 10539 6187 10581 6196
rect 20235 6236 20277 6245
rect 20235 6196 20236 6236
rect 20276 6196 20277 6236
rect 20235 6187 20277 6196
rect 25995 6236 26037 6245
rect 25995 6196 25996 6236
rect 26036 6196 26037 6236
rect 25995 6187 26037 6196
rect 28779 6236 28821 6245
rect 28779 6196 28780 6236
rect 28820 6196 28821 6236
rect 28779 6187 28821 6196
rect 29259 6236 29301 6245
rect 29259 6196 29260 6236
rect 29300 6196 29301 6236
rect 29259 6187 29301 6196
rect 33763 6236 33821 6237
rect 33763 6196 33772 6236
rect 33812 6196 33821 6236
rect 33763 6195 33821 6196
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 4867 5900 4925 5901
rect 4867 5860 4876 5900
rect 4916 5860 4925 5900
rect 4867 5859 4925 5860
rect 8235 5900 8277 5909
rect 8235 5860 8236 5900
rect 8276 5860 8277 5900
rect 8235 5851 8277 5860
rect 11211 5900 11253 5909
rect 11211 5860 11212 5900
rect 11252 5860 11253 5900
rect 11211 5851 11253 5860
rect 23307 5900 23349 5909
rect 23307 5860 23308 5900
rect 23348 5860 23349 5900
rect 23307 5851 23349 5860
rect 28299 5900 28341 5909
rect 28299 5860 28300 5900
rect 28340 5860 28341 5900
rect 28299 5851 28341 5860
rect 29347 5900 29405 5901
rect 29347 5860 29356 5900
rect 29396 5860 29405 5900
rect 29347 5859 29405 5860
rect 31075 5900 31133 5901
rect 31075 5860 31084 5900
rect 31124 5860 31133 5900
rect 31075 5859 31133 5860
rect 34251 5900 34293 5909
rect 34251 5860 34252 5900
rect 34292 5860 34293 5900
rect 34251 5851 34293 5860
rect 4203 5816 4245 5825
rect 4203 5776 4204 5816
rect 4244 5776 4245 5816
rect 4203 5767 4245 5776
rect 4675 5816 4733 5817
rect 4675 5776 4684 5816
rect 4724 5776 4733 5816
rect 4675 5775 4733 5776
rect 10723 5816 10781 5817
rect 10723 5776 10732 5816
rect 10772 5776 10781 5816
rect 10723 5775 10781 5776
rect 11499 5816 11541 5825
rect 11499 5776 11500 5816
rect 11540 5776 11541 5816
rect 11499 5767 11541 5776
rect 11595 5816 11637 5825
rect 11595 5776 11596 5816
rect 11636 5776 11637 5816
rect 11595 5767 11637 5776
rect 17451 5816 17493 5825
rect 17451 5776 17452 5816
rect 17492 5776 17493 5816
rect 17451 5767 17493 5776
rect 24931 5816 24989 5817
rect 24931 5776 24940 5816
rect 24980 5776 24989 5816
rect 24931 5775 24989 5776
rect 35115 5816 35157 5825
rect 35115 5776 35116 5816
rect 35156 5776 35157 5816
rect 35115 5767 35157 5776
rect 11691 5732 11733 5741
rect 11691 5692 11692 5732
rect 11732 5692 11733 5732
rect 11691 5683 11733 5692
rect 13707 5732 13749 5741
rect 13707 5692 13708 5732
rect 13748 5692 13749 5732
rect 11875 5690 11933 5691
rect 4395 5648 4437 5657
rect 4395 5608 4396 5648
rect 4436 5608 4437 5648
rect 4395 5599 4437 5608
rect 4587 5648 4629 5657
rect 4587 5608 4588 5648
rect 4628 5608 4629 5648
rect 4587 5599 4629 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 5539 5648 5597 5649
rect 5539 5608 5548 5648
rect 5588 5608 5597 5648
rect 5539 5607 5597 5608
rect 5827 5648 5885 5649
rect 5827 5608 5836 5648
rect 5876 5608 5885 5648
rect 5827 5607 5885 5608
rect 6123 5648 6165 5657
rect 6123 5608 6124 5648
rect 6164 5608 6165 5648
rect 6123 5599 6165 5608
rect 6787 5648 6845 5649
rect 6787 5608 6796 5648
rect 6836 5608 6845 5648
rect 6787 5607 6845 5608
rect 7171 5648 7229 5649
rect 7171 5608 7180 5648
rect 7220 5608 7229 5648
rect 7171 5607 7229 5608
rect 7267 5648 7325 5649
rect 7267 5608 7276 5648
rect 7316 5608 7325 5648
rect 7267 5607 7325 5608
rect 7755 5648 7797 5657
rect 7755 5608 7756 5648
rect 7796 5608 7797 5648
rect 7755 5599 7797 5608
rect 7851 5648 7893 5657
rect 7851 5608 7852 5648
rect 7892 5608 7893 5648
rect 7851 5599 7893 5608
rect 7947 5648 7989 5657
rect 7947 5608 7948 5648
rect 7988 5608 7989 5648
rect 7947 5599 7989 5608
rect 8235 5648 8277 5657
rect 8235 5608 8236 5648
rect 8276 5608 8277 5648
rect 8235 5599 8277 5608
rect 8427 5648 8469 5657
rect 8427 5608 8428 5648
rect 8468 5608 8469 5648
rect 8427 5599 8469 5608
rect 8515 5648 8573 5649
rect 8515 5608 8524 5648
rect 8564 5608 8573 5648
rect 8515 5607 8573 5608
rect 9379 5648 9437 5649
rect 9379 5608 9388 5648
rect 9428 5608 9437 5648
rect 9379 5607 9437 5608
rect 10339 5648 10397 5649
rect 10339 5608 10348 5648
rect 10388 5608 10397 5648
rect 10339 5607 10397 5608
rect 10539 5648 10581 5657
rect 10539 5608 10540 5648
rect 10580 5608 10581 5648
rect 10539 5599 10581 5608
rect 10731 5648 10773 5657
rect 10731 5608 10732 5648
rect 10772 5608 10773 5648
rect 10731 5599 10773 5608
rect 10827 5648 10869 5657
rect 10827 5608 10828 5648
rect 10868 5608 10869 5648
rect 10827 5599 10869 5608
rect 11115 5648 11157 5657
rect 11115 5608 11116 5648
rect 11156 5608 11157 5648
rect 11115 5599 11157 5608
rect 11299 5648 11357 5649
rect 11299 5608 11308 5648
rect 11348 5608 11357 5648
rect 11299 5607 11357 5608
rect 11787 5648 11829 5657
rect 11875 5650 11884 5690
rect 11924 5650 11933 5690
rect 13707 5683 13749 5692
rect 14091 5732 14133 5741
rect 14091 5692 14092 5732
rect 14132 5692 14133 5732
rect 14091 5683 14133 5692
rect 23787 5732 23829 5741
rect 23787 5692 23788 5732
rect 23828 5692 23829 5732
rect 23787 5683 23829 5692
rect 35019 5732 35061 5741
rect 35019 5692 35020 5732
rect 35060 5692 35061 5732
rect 35019 5683 35061 5692
rect 35211 5732 35253 5741
rect 35211 5692 35212 5732
rect 35252 5692 35253 5732
rect 35211 5683 35253 5692
rect 15716 5665 15774 5666
rect 11875 5649 11933 5650
rect 11787 5608 11788 5648
rect 11828 5608 11829 5648
rect 11787 5599 11829 5608
rect 12171 5648 12213 5657
rect 12171 5608 12172 5648
rect 12212 5608 12213 5648
rect 12171 5599 12213 5608
rect 12267 5648 12309 5657
rect 12267 5608 12268 5648
rect 12308 5608 12309 5648
rect 12267 5599 12309 5608
rect 13411 5648 13469 5649
rect 13411 5608 13420 5648
rect 13460 5608 13469 5648
rect 13411 5607 13469 5608
rect 13611 5648 13653 5657
rect 13611 5608 13612 5648
rect 13652 5608 13653 5648
rect 13611 5599 13653 5608
rect 13803 5648 13845 5657
rect 13803 5608 13804 5648
rect 13844 5608 13845 5648
rect 13803 5599 13845 5608
rect 13995 5648 14037 5657
rect 13995 5608 13996 5648
rect 14036 5608 14037 5648
rect 13995 5599 14037 5608
rect 14187 5648 14229 5657
rect 14187 5608 14188 5648
rect 14228 5608 14229 5648
rect 14187 5599 14229 5608
rect 14371 5648 14429 5649
rect 14371 5608 14380 5648
rect 14420 5608 14429 5648
rect 14371 5607 14429 5608
rect 15051 5648 15093 5657
rect 15051 5608 15052 5648
rect 15092 5608 15093 5648
rect 15051 5599 15093 5608
rect 15427 5648 15485 5649
rect 15427 5608 15436 5648
rect 15476 5608 15485 5648
rect 15716 5625 15725 5665
rect 15765 5625 15774 5665
rect 15716 5624 15774 5625
rect 16011 5648 16053 5657
rect 15427 5607 15485 5608
rect 16011 5608 16012 5648
rect 16052 5608 16053 5648
rect 16011 5599 16053 5608
rect 16291 5648 16349 5649
rect 16291 5608 16300 5648
rect 16340 5608 16349 5648
rect 16291 5607 16349 5608
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 17931 5599 17973 5608
rect 18307 5648 18365 5649
rect 18307 5608 18316 5648
rect 18356 5608 18365 5648
rect 18307 5607 18365 5608
rect 19171 5648 19229 5649
rect 19171 5608 19180 5648
rect 19220 5608 19229 5648
rect 19171 5607 19229 5608
rect 20331 5648 20373 5657
rect 20331 5608 20332 5648
rect 20372 5608 20373 5648
rect 20331 5599 20373 5608
rect 20907 5648 20949 5657
rect 20907 5608 20908 5648
rect 20948 5608 20949 5648
rect 20907 5599 20949 5608
rect 21283 5648 21341 5649
rect 21283 5608 21292 5648
rect 21332 5608 21341 5648
rect 21283 5607 21341 5608
rect 22147 5648 22205 5649
rect 22147 5608 22156 5648
rect 22196 5608 22205 5648
rect 22147 5607 22205 5608
rect 23395 5648 23453 5649
rect 23395 5608 23404 5648
rect 23444 5608 23453 5648
rect 23395 5607 23453 5608
rect 23691 5648 23733 5657
rect 23691 5608 23692 5648
rect 23732 5608 23733 5648
rect 23691 5599 23733 5608
rect 23979 5648 24021 5657
rect 23979 5608 23980 5648
rect 24020 5608 24021 5648
rect 23979 5599 24021 5608
rect 24259 5648 24317 5649
rect 24259 5608 24268 5648
rect 24308 5608 24317 5648
rect 24259 5607 24317 5608
rect 25323 5648 25365 5657
rect 25323 5608 25324 5648
rect 25364 5608 25365 5648
rect 25323 5599 25365 5608
rect 25419 5648 25461 5657
rect 25419 5608 25420 5648
rect 25460 5608 25461 5648
rect 25419 5599 25461 5608
rect 25603 5648 25661 5649
rect 25603 5608 25612 5648
rect 25652 5608 25661 5648
rect 27243 5648 27285 5657
rect 25603 5607 25661 5608
rect 27134 5643 27192 5644
rect 27134 5603 27143 5643
rect 27183 5603 27192 5643
rect 27134 5602 27192 5603
rect 27243 5608 27244 5648
rect 27284 5608 27285 5648
rect 27243 5599 27285 5608
rect 27811 5648 27869 5649
rect 27811 5608 27820 5648
rect 27860 5608 27869 5648
rect 27811 5607 27869 5608
rect 27915 5648 27957 5657
rect 27915 5608 27916 5648
rect 27956 5608 27957 5648
rect 27915 5599 27957 5608
rect 28107 5648 28149 5657
rect 28107 5608 28108 5648
rect 28148 5608 28149 5648
rect 28107 5599 28149 5608
rect 28299 5648 28341 5657
rect 28299 5608 28300 5648
rect 28340 5608 28341 5648
rect 28299 5599 28341 5608
rect 28483 5648 28541 5649
rect 28483 5608 28492 5648
rect 28532 5608 28541 5648
rect 28483 5607 28541 5608
rect 30019 5648 30077 5649
rect 30019 5608 30028 5648
rect 30068 5608 30077 5648
rect 30019 5607 30077 5608
rect 30883 5648 30941 5649
rect 30883 5608 30892 5648
rect 30932 5608 30941 5648
rect 30883 5607 30941 5608
rect 31747 5648 31805 5649
rect 31747 5608 31756 5648
rect 31796 5608 31805 5648
rect 31747 5607 31805 5608
rect 33483 5648 33525 5657
rect 33483 5608 33484 5648
rect 33524 5608 33525 5648
rect 33483 5599 33525 5608
rect 33771 5648 33813 5657
rect 33771 5608 33772 5648
rect 33812 5608 33813 5648
rect 33771 5599 33813 5608
rect 33955 5648 34013 5649
rect 33955 5608 33964 5648
rect 34004 5608 34013 5648
rect 33955 5607 34013 5608
rect 34059 5648 34101 5657
rect 34059 5608 34060 5648
rect 34100 5608 34101 5648
rect 34059 5599 34101 5608
rect 34251 5648 34293 5657
rect 34251 5608 34252 5648
rect 34292 5608 34293 5648
rect 34251 5599 34293 5608
rect 34435 5648 34493 5649
rect 34435 5608 34444 5648
rect 34484 5608 34493 5648
rect 34435 5607 34493 5608
rect 34635 5648 34677 5657
rect 34635 5608 34636 5648
rect 34676 5608 34677 5648
rect 34635 5599 34677 5608
rect 34723 5648 34781 5649
rect 34723 5608 34732 5648
rect 34772 5608 34781 5648
rect 34723 5607 34781 5608
rect 34923 5648 34965 5657
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 35299 5648 35357 5649
rect 35299 5608 35308 5648
rect 35348 5608 35357 5648
rect 35299 5607 35357 5608
rect 12747 5564 12789 5573
rect 12747 5524 12748 5564
rect 12788 5524 12789 5564
rect 12747 5515 12789 5524
rect 27043 5564 27101 5565
rect 27043 5524 27052 5564
rect 27092 5524 27101 5564
rect 27043 5523 27101 5524
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 5739 5480 5781 5489
rect 5739 5440 5740 5480
rect 5780 5440 5781 5480
rect 5739 5431 5781 5440
rect 6987 5480 7029 5489
rect 6987 5440 6988 5480
rect 7028 5440 7029 5480
rect 6987 5431 7029 5440
rect 8035 5480 8093 5481
rect 8035 5440 8044 5480
rect 8084 5440 8093 5480
rect 8035 5439 8093 5440
rect 8707 5480 8765 5481
rect 8707 5440 8716 5480
rect 8756 5440 8765 5480
rect 8707 5439 8765 5440
rect 9667 5480 9725 5481
rect 9667 5440 9676 5480
rect 9716 5440 9725 5480
rect 9667 5439 9725 5440
rect 12451 5480 12509 5481
rect 12451 5440 12460 5480
rect 12500 5440 12509 5480
rect 12451 5439 12509 5440
rect 15339 5480 15381 5489
rect 15339 5440 15340 5480
rect 15380 5440 15381 5480
rect 15339 5431 15381 5440
rect 15819 5480 15861 5489
rect 15819 5440 15820 5480
rect 15860 5440 15861 5480
rect 15819 5431 15861 5440
rect 16203 5480 16245 5489
rect 16203 5440 16204 5480
rect 16244 5440 16245 5480
rect 16203 5431 16245 5440
rect 25123 5480 25181 5481
rect 25123 5440 25132 5480
rect 25172 5440 25181 5480
rect 25123 5439 25181 5440
rect 26275 5480 26333 5481
rect 26275 5440 26284 5480
rect 26324 5440 26333 5480
rect 26275 5439 26333 5440
rect 26859 5480 26901 5489
rect 26859 5440 26860 5480
rect 26900 5440 26901 5480
rect 26859 5431 26901 5440
rect 26947 5480 27005 5481
rect 26947 5440 26956 5480
rect 26996 5440 27005 5480
rect 26947 5439 27005 5440
rect 29155 5480 29213 5481
rect 29155 5440 29164 5480
rect 29204 5440 29213 5480
rect 29155 5439 29213 5440
rect 30211 5480 30269 5481
rect 30211 5440 30220 5480
rect 30260 5440 30269 5480
rect 30211 5439 30269 5440
rect 33675 5480 33717 5489
rect 33675 5440 33676 5480
rect 33716 5440 33717 5480
rect 33675 5431 33717 5440
rect 34443 5480 34485 5489
rect 34443 5440 34444 5480
rect 34484 5440 34485 5480
rect 34443 5431 34485 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 22155 5202 22197 5211
rect 22155 5162 22156 5202
rect 22196 5162 22197 5202
rect 22155 5153 22197 5162
rect 643 5144 701 5145
rect 643 5104 652 5144
rect 692 5104 701 5144
rect 643 5103 701 5104
rect 11971 5144 12029 5145
rect 11971 5104 11980 5144
rect 12020 5104 12029 5144
rect 11971 5103 12029 5104
rect 12075 5144 12117 5153
rect 12075 5104 12076 5144
rect 12116 5104 12117 5144
rect 12075 5095 12117 5104
rect 14755 5144 14813 5145
rect 14755 5104 14764 5144
rect 14804 5104 14813 5144
rect 14755 5103 14813 5104
rect 14859 5144 14901 5153
rect 14859 5104 14860 5144
rect 14900 5104 14901 5144
rect 14859 5095 14901 5104
rect 20611 5144 20669 5145
rect 20611 5104 20620 5144
rect 20660 5104 20669 5144
rect 20611 5103 20669 5104
rect 26667 5144 26709 5153
rect 26667 5104 26668 5144
rect 26708 5104 26709 5144
rect 26667 5095 26709 5104
rect 27331 5144 27389 5145
rect 27331 5104 27340 5144
rect 27380 5104 27389 5144
rect 27331 5103 27389 5104
rect 28395 5144 28437 5153
rect 28395 5104 28396 5144
rect 28436 5104 28437 5144
rect 28395 5095 28437 5104
rect 5931 5060 5973 5069
rect 5931 5020 5932 5060
rect 5972 5020 5973 5060
rect 5931 5011 5973 5020
rect 11875 5060 11933 5061
rect 11875 5020 11884 5060
rect 11924 5020 11933 5060
rect 11875 5019 11933 5020
rect 13803 5060 13845 5069
rect 13803 5020 13804 5060
rect 13844 5020 13845 5060
rect 13803 5011 13845 5020
rect 14659 5060 14717 5061
rect 14659 5020 14668 5060
rect 14708 5020 14717 5060
rect 14659 5019 14717 5020
rect 17739 5060 17781 5069
rect 17739 5020 17740 5060
rect 17780 5020 17781 5060
rect 17739 5011 17781 5020
rect 20811 5060 20853 5069
rect 20811 5020 20812 5060
rect 20852 5020 20853 5060
rect 20811 5011 20853 5020
rect 27427 5060 27485 5061
rect 27427 5020 27436 5060
rect 27476 5020 27485 5060
rect 27427 5019 27485 5020
rect 4203 4976 4245 4985
rect 4203 4936 4204 4976
rect 4244 4936 4245 4976
rect 4203 4927 4245 4936
rect 4395 4976 4437 4985
rect 4395 4936 4396 4976
rect 4436 4936 4437 4976
rect 4395 4927 4437 4936
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 5347 4976 5405 4977
rect 5347 4936 5356 4976
rect 5396 4936 5405 4976
rect 5347 4935 5405 4936
rect 5731 4976 5789 4977
rect 5731 4936 5740 4976
rect 5780 4936 5789 4976
rect 5731 4935 5789 4936
rect 5835 4976 5877 4985
rect 5835 4936 5836 4976
rect 5876 4936 5877 4976
rect 5835 4927 5877 4936
rect 6027 4976 6069 4985
rect 6027 4936 6028 4976
rect 6068 4936 6069 4976
rect 6027 4927 6069 4936
rect 6219 4976 6261 4985
rect 6219 4936 6220 4976
rect 6260 4936 6261 4976
rect 6219 4927 6261 4936
rect 6883 4976 6941 4977
rect 6883 4936 6892 4976
rect 6932 4936 6941 4976
rect 6883 4935 6941 4936
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7371 4976 7413 4985
rect 7371 4936 7372 4976
rect 7412 4936 7413 4976
rect 7371 4927 7413 4936
rect 7467 4976 7509 4985
rect 7467 4936 7468 4976
rect 7508 4936 7509 4976
rect 7467 4927 7509 4936
rect 7843 4976 7901 4977
rect 7843 4936 7852 4976
rect 7892 4936 7901 4976
rect 7843 4935 7901 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 9091 4976 9149 4977
rect 9091 4936 9100 4976
rect 9140 4936 9149 4976
rect 9091 4935 9149 4936
rect 9955 4976 10013 4977
rect 9955 4936 9964 4976
rect 10004 4936 10013 4976
rect 9955 4935 10013 4936
rect 11115 4976 11157 4985
rect 11115 4936 11116 4976
rect 11156 4936 11157 4976
rect 11115 4927 11157 4936
rect 11691 4976 11733 4985
rect 11691 4936 11692 4976
rect 11732 4936 11733 4976
rect 11691 4927 11733 4936
rect 11787 4976 11829 4985
rect 11787 4936 11788 4976
rect 11828 4936 11829 4976
rect 11787 4927 11829 4936
rect 12931 4976 12989 4977
rect 12931 4936 12940 4976
rect 12980 4936 12989 4976
rect 12931 4935 12989 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 13411 4976 13469 4977
rect 13411 4936 13420 4976
rect 13460 4936 13469 4976
rect 13411 4935 13469 4936
rect 13707 4976 13749 4985
rect 13707 4936 13708 4976
rect 13748 4936 13749 4976
rect 13707 4927 13749 4936
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 14091 4976 14133 4985
rect 14091 4936 14092 4976
rect 14132 4936 14133 4976
rect 14091 4927 14133 4936
rect 14275 4976 14333 4977
rect 14275 4936 14284 4976
rect 14324 4936 14333 4976
rect 14275 4935 14333 4936
rect 14475 4976 14517 4985
rect 14475 4936 14476 4976
rect 14516 4936 14517 4976
rect 14475 4927 14517 4936
rect 14571 4976 14613 4985
rect 14571 4936 14572 4976
rect 14612 4936 14613 4976
rect 14571 4927 14613 4936
rect 15139 4976 15197 4977
rect 15139 4936 15148 4976
rect 15188 4936 15197 4976
rect 15139 4935 15197 4936
rect 16011 4976 16053 4985
rect 16011 4936 16012 4976
rect 16052 4936 16053 4976
rect 16011 4927 16053 4936
rect 16099 4976 16157 4977
rect 16099 4936 16108 4976
rect 16148 4936 16157 4976
rect 16099 4935 16157 4936
rect 16291 4976 16349 4977
rect 16291 4936 16300 4976
rect 16340 4936 16349 4976
rect 16291 4935 16349 4936
rect 16395 4976 16437 4985
rect 16395 4936 16396 4976
rect 16436 4936 16437 4976
rect 16395 4927 16437 4936
rect 16587 4976 16629 4985
rect 16587 4936 16588 4976
rect 16628 4936 16629 4976
rect 16587 4927 16629 4936
rect 16771 4976 16829 4977
rect 16771 4936 16780 4976
rect 16820 4936 16829 4976
rect 16771 4935 16829 4936
rect 18403 4976 18461 4977
rect 18403 4936 18412 4976
rect 18452 4936 18461 4976
rect 18403 4935 18461 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 19939 4976 19997 4977
rect 19939 4936 19948 4976
rect 19988 4936 19997 4976
rect 19939 4935 19997 4936
rect 21475 4976 21533 4977
rect 21475 4936 21484 4976
rect 21524 4936 21533 4976
rect 21475 4935 21533 4936
rect 21963 4976 22005 4985
rect 21963 4936 21964 4976
rect 22004 4936 22005 4976
rect 21963 4927 22005 4936
rect 22051 4976 22109 4977
rect 22051 4936 22060 4976
rect 22100 4936 22109 4976
rect 22051 4935 22109 4936
rect 22339 4976 22397 4977
rect 22339 4936 22348 4976
rect 22388 4936 22397 4976
rect 22339 4935 22397 4936
rect 23019 4976 23061 4985
rect 23019 4936 23020 4976
rect 23060 4936 23061 4976
rect 23019 4927 23061 4936
rect 23307 4976 23349 4985
rect 23307 4936 23308 4976
rect 23348 4936 23349 4976
rect 23307 4927 23349 4936
rect 24451 4976 24509 4977
rect 24451 4936 24460 4976
rect 24500 4936 24509 4976
rect 24451 4935 24509 4936
rect 25315 4976 25373 4977
rect 25315 4936 25324 4976
rect 25364 4936 25373 4976
rect 25315 4935 25373 4936
rect 25707 4976 25749 4985
rect 25707 4936 25708 4976
rect 25748 4936 25749 4976
rect 25707 4927 25749 4936
rect 25987 4976 26045 4977
rect 25987 4936 25996 4976
rect 26036 4936 26045 4976
rect 25987 4935 26045 4936
rect 26091 4976 26133 4985
rect 26091 4936 26092 4976
rect 26132 4936 26133 4976
rect 26091 4927 26133 4936
rect 26467 4976 26525 4977
rect 26467 4936 26476 4976
rect 26516 4936 26525 4976
rect 26467 4935 26525 4936
rect 26755 4976 26813 4977
rect 26755 4936 26764 4976
rect 26804 4936 26813 4976
rect 26755 4935 26813 4936
rect 26947 4976 27005 4977
rect 26947 4936 26956 4976
rect 26996 4936 27005 4976
rect 26947 4935 27005 4936
rect 27531 4976 27573 4985
rect 27531 4936 27532 4976
rect 27572 4936 27573 4976
rect 27531 4927 27573 4936
rect 27627 4976 27669 4985
rect 27627 4936 27628 4976
rect 27668 4936 27669 4976
rect 27627 4927 27669 4936
rect 27907 4976 27965 4977
rect 27907 4936 27916 4976
rect 27956 4936 27965 4976
rect 27907 4935 27965 4936
rect 28011 4976 28053 4985
rect 28011 4936 28012 4976
rect 28052 4936 28053 4976
rect 28011 4927 28053 4936
rect 28203 4976 28245 4985
rect 28203 4936 28204 4976
rect 28244 4936 28245 4976
rect 28203 4927 28245 4936
rect 28579 4976 28637 4977
rect 28579 4936 28588 4976
rect 28628 4936 28637 4976
rect 28579 4935 28637 4936
rect 28675 4976 28733 4977
rect 28675 4936 28684 4976
rect 28724 4936 28733 4976
rect 28675 4935 28733 4936
rect 29163 4976 29205 4985
rect 29163 4936 29164 4976
rect 29204 4936 29205 4976
rect 29163 4927 29205 4936
rect 29539 4976 29597 4977
rect 29539 4936 29548 4976
rect 29588 4936 29597 4976
rect 29539 4935 29597 4936
rect 30403 4976 30461 4977
rect 30403 4936 30412 4976
rect 30452 4936 30461 4976
rect 30403 4935 30461 4936
rect 31563 4976 31605 4985
rect 31563 4936 31564 4976
rect 31604 4936 31605 4976
rect 31563 4927 31605 4936
rect 3819 4808 3861 4817
rect 3819 4768 3820 4808
rect 3860 4768 3861 4808
rect 3819 4759 3861 4768
rect 4483 4808 4541 4809
rect 4483 4768 4492 4808
rect 4532 4768 4541 4808
rect 4483 4767 4541 4768
rect 15811 4808 15869 4809
rect 15811 4768 15820 4808
rect 15860 4768 15869 4808
rect 15811 4767 15869 4768
rect 16587 4808 16629 4817
rect 16587 4768 16588 4808
rect 16628 4768 16629 4808
rect 16587 4759 16629 4768
rect 27339 4808 27381 4817
rect 27339 4768 27340 4808
rect 27380 4768 27381 4808
rect 27339 4759 27381 4768
rect 4675 4724 4733 4725
rect 4675 4684 4684 4724
rect 4724 4684 4733 4724
rect 4675 4683 4733 4684
rect 7651 4724 7709 4725
rect 7651 4684 7660 4724
rect 7700 4684 7709 4724
rect 7651 4683 7709 4684
rect 8515 4724 8573 4725
rect 8515 4684 8524 4724
rect 8564 4684 8573 4724
rect 8515 4683 8573 4684
rect 12259 4724 12317 4725
rect 12259 4684 12268 4724
rect 12308 4684 12317 4724
rect 12259 4683 12317 4684
rect 13131 4724 13173 4733
rect 13131 4684 13132 4724
rect 13172 4684 13173 4724
rect 13131 4675 13173 4684
rect 14187 4724 14229 4733
rect 14187 4684 14188 4724
rect 14228 4684 14229 4724
rect 14187 4675 14229 4684
rect 17443 4724 17501 4725
rect 17443 4684 17452 4724
rect 17492 4684 17501 4724
rect 17443 4683 17501 4684
rect 18891 4724 18933 4733
rect 18891 4684 18892 4724
rect 18932 4684 18933 4724
rect 18891 4675 18933 4684
rect 21675 4724 21717 4733
rect 21675 4684 21676 4724
rect 21716 4684 21717 4724
rect 21675 4675 21717 4684
rect 28203 4724 28245 4733
rect 28203 4684 28204 4724
rect 28244 4684 28245 4724
rect 28203 4675 28245 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 7563 4388 7605 4397
rect 7563 4348 7564 4388
rect 7604 4348 7605 4388
rect 7563 4339 7605 4348
rect 11211 4388 11253 4397
rect 11211 4348 11212 4388
rect 11252 4348 11253 4388
rect 11211 4339 11253 4348
rect 19363 4388 19421 4389
rect 19363 4348 19372 4388
rect 19412 4348 19421 4388
rect 19363 4347 19421 4348
rect 23307 4388 23349 4397
rect 23307 4348 23308 4388
rect 23348 4348 23349 4388
rect 23307 4339 23349 4348
rect 25227 4388 25269 4397
rect 25227 4348 25228 4388
rect 25268 4348 25269 4388
rect 25227 4339 25269 4348
rect 25515 4388 25557 4397
rect 25515 4348 25516 4388
rect 25556 4348 25557 4388
rect 25515 4339 25557 4348
rect 8139 4304 8181 4313
rect 8139 4264 8140 4304
rect 8180 4264 8181 4304
rect 8139 4255 8181 4264
rect 9195 4304 9237 4313
rect 9195 4264 9196 4304
rect 9236 4264 9237 4304
rect 9195 4255 9237 4264
rect 11019 4304 11061 4313
rect 11019 4264 11020 4304
rect 11060 4264 11061 4304
rect 11019 4255 11061 4264
rect 11403 4304 11445 4313
rect 11403 4264 11404 4304
rect 11444 4264 11445 4304
rect 11403 4255 11445 4264
rect 14563 4304 14621 4305
rect 14563 4264 14572 4304
rect 14612 4264 14621 4304
rect 14563 4263 14621 4264
rect 29059 4304 29117 4305
rect 29059 4264 29068 4304
rect 29108 4264 29117 4304
rect 29059 4263 29117 4264
rect 3339 4136 3381 4145
rect 3339 4096 3340 4136
rect 3380 4096 3381 4136
rect 3339 4087 3381 4096
rect 3715 4136 3773 4137
rect 3715 4096 3724 4136
rect 3764 4096 3773 4136
rect 3715 4095 3773 4096
rect 4579 4136 4637 4137
rect 4579 4096 4588 4136
rect 4628 4096 4637 4136
rect 4579 4095 4637 4096
rect 5827 4136 5885 4137
rect 5827 4096 5836 4136
rect 5876 4096 5885 4136
rect 5827 4095 5885 4096
rect 6211 4136 6269 4137
rect 6211 4096 6220 4136
rect 6260 4096 6269 4136
rect 6211 4095 6269 4096
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 7371 4136 7413 4145
rect 7371 4096 7372 4136
rect 7412 4096 7413 4136
rect 7371 4087 7413 4096
rect 7843 4136 7901 4137
rect 7843 4096 7852 4136
rect 7892 4096 7901 4136
rect 7843 4095 7901 4096
rect 9379 4136 9437 4137
rect 9379 4096 9388 4136
rect 9428 4096 9437 4136
rect 9379 4095 9437 4096
rect 9483 4136 9525 4145
rect 9483 4096 9484 4136
rect 9524 4096 9525 4136
rect 9483 4087 9525 4096
rect 9667 4136 9725 4137
rect 9667 4096 9676 4136
rect 9716 4096 9725 4136
rect 9667 4095 9725 4096
rect 10435 4136 10493 4137
rect 10435 4096 10444 4136
rect 10484 4096 10493 4136
rect 10435 4095 10493 4096
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 11403 4136 11445 4145
rect 11403 4096 11404 4136
rect 11444 4096 11445 4136
rect 11403 4087 11445 4096
rect 11691 4136 11733 4145
rect 11691 4096 11692 4136
rect 11732 4096 11733 4136
rect 11691 4087 11733 4096
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 12171 4136 12213 4145
rect 12171 4096 12172 4136
rect 12212 4096 12213 4136
rect 12171 4087 12213 4096
rect 12547 4136 12605 4137
rect 12547 4096 12556 4136
rect 12596 4096 12605 4136
rect 12547 4095 12605 4096
rect 13411 4136 13469 4137
rect 13411 4096 13420 4136
rect 13460 4096 13469 4136
rect 13411 4095 13469 4096
rect 14763 4136 14805 4145
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 14859 4136 14901 4145
rect 14859 4096 14860 4136
rect 14900 4096 14901 4136
rect 14859 4087 14901 4096
rect 14955 4136 14997 4145
rect 14955 4096 14956 4136
rect 14996 4096 14997 4136
rect 14955 4087 14997 4096
rect 15051 4136 15093 4145
rect 15051 4096 15052 4136
rect 15092 4096 15093 4136
rect 15051 4087 15093 4096
rect 15235 4136 15293 4137
rect 15235 4096 15244 4136
rect 15284 4096 15293 4136
rect 15235 4095 15293 4096
rect 16099 4136 16157 4137
rect 16099 4096 16108 4136
rect 16148 4096 16157 4136
rect 16099 4095 16157 4096
rect 17347 4136 17405 4137
rect 17347 4096 17356 4136
rect 17396 4096 17405 4136
rect 17347 4095 17405 4096
rect 18211 4136 18269 4137
rect 18211 4096 18220 4136
rect 18260 4096 18269 4136
rect 18211 4095 18269 4096
rect 19747 4136 19805 4137
rect 19747 4096 19756 4136
rect 19796 4096 19805 4136
rect 19747 4095 19805 4096
rect 20043 4136 20085 4145
rect 20043 4096 20044 4136
rect 20084 4096 20085 4136
rect 20043 4087 20085 4096
rect 20707 4136 20765 4137
rect 20707 4096 20716 4136
rect 20756 4096 20765 4136
rect 20707 4095 20765 4096
rect 20907 4136 20949 4145
rect 20907 4096 20908 4136
rect 20948 4096 20949 4136
rect 20907 4087 20949 4096
rect 21283 4136 21341 4137
rect 21283 4096 21292 4136
rect 21332 4096 21341 4136
rect 21283 4095 21341 4096
rect 22147 4136 22205 4137
rect 22147 4096 22156 4136
rect 22196 4096 22205 4136
rect 22147 4095 22205 4096
rect 23587 4136 23645 4137
rect 23587 4096 23596 4136
rect 23636 4096 23645 4136
rect 23587 4095 23645 4096
rect 23691 4136 23733 4145
rect 23691 4096 23692 4136
rect 23732 4096 23733 4136
rect 23691 4087 23733 4096
rect 23875 4136 23933 4137
rect 23875 4096 23884 4136
rect 23924 4096 23933 4136
rect 23875 4095 23933 4096
rect 25123 4136 25181 4137
rect 25123 4096 25132 4136
rect 25172 4096 25181 4136
rect 25123 4095 25181 4096
rect 25707 4136 25749 4145
rect 25707 4096 25708 4136
rect 25748 4096 25749 4136
rect 25707 4087 25749 4096
rect 25803 4136 25845 4145
rect 25803 4096 25804 4136
rect 25844 4096 25845 4136
rect 25803 4087 25845 4096
rect 25995 4136 26037 4145
rect 25995 4096 25996 4136
rect 26036 4096 26037 4136
rect 25995 4087 26037 4096
rect 26187 4136 26229 4145
rect 26187 4096 26188 4136
rect 26228 4096 26229 4136
rect 26187 4087 26229 4096
rect 26467 4136 26525 4137
rect 26467 4096 26476 4136
rect 26516 4096 26525 4136
rect 26467 4095 26525 4096
rect 26659 4136 26717 4137
rect 26659 4096 26668 4136
rect 26708 4096 26717 4136
rect 26659 4095 26717 4096
rect 26947 4136 27005 4137
rect 26947 4096 26956 4136
rect 26996 4096 27005 4136
rect 26947 4095 27005 4096
rect 28195 4136 28253 4137
rect 28195 4096 28204 4136
rect 28244 4096 28253 4136
rect 28195 4095 28253 4096
rect 28387 4136 28445 4137
rect 28387 4096 28396 4136
rect 28436 4096 28445 4136
rect 28387 4095 28445 4096
rect 29251 4136 29309 4137
rect 29251 4096 29260 4136
rect 29300 4096 29309 4136
rect 29251 4095 29309 4096
rect 29931 4136 29973 4145
rect 29931 4096 29932 4136
rect 29972 4096 29973 4136
rect 29931 4087 29973 4096
rect 30123 4136 30165 4145
rect 30123 4096 30124 4136
rect 30164 4096 30165 4136
rect 30123 4087 30165 4096
rect 30499 4136 30557 4137
rect 30499 4096 30508 4136
rect 30548 4096 30557 4136
rect 30499 4095 30557 4096
rect 31363 4136 31421 4137
rect 31363 4096 31372 4136
rect 31412 4096 31421 4136
rect 31363 4095 31421 4096
rect 32611 4136 32669 4137
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32611 4095 32669 4096
rect 10539 4052 10581 4061
rect 10539 4012 10540 4052
rect 10580 4012 10581 4052
rect 10539 4003 10581 4012
rect 16971 4052 17013 4061
rect 16971 4012 16972 4052
rect 17012 4012 17013 4052
rect 16971 4003 17013 4012
rect 25603 4052 25661 4053
rect 25603 4012 25612 4052
rect 25652 4012 25661 4052
rect 25603 4011 25661 4012
rect 26091 4052 26133 4061
rect 26091 4012 26092 4052
rect 26132 4012 26133 4052
rect 26091 4003 26133 4012
rect 643 3968 701 3969
rect 643 3928 652 3968
rect 692 3928 701 3968
rect 643 3927 701 3928
rect 6883 3968 6941 3969
rect 6883 3928 6892 3968
rect 6932 3928 6941 3968
rect 6883 3927 6941 3928
rect 7267 3968 7325 3969
rect 7267 3928 7276 3968
rect 7316 3928 7325 3968
rect 7267 3927 7325 3928
rect 9675 3968 9717 3977
rect 9675 3928 9676 3968
rect 9716 3928 9717 3968
rect 9675 3919 9717 3928
rect 11211 3968 11253 3977
rect 11211 3928 11212 3968
rect 11252 3928 11253 3968
rect 11211 3919 11253 3928
rect 15907 3968 15965 3969
rect 15907 3928 15916 3968
rect 15956 3928 15965 3968
rect 15907 3927 15965 3928
rect 16771 3968 16829 3969
rect 16771 3928 16780 3968
rect 16820 3928 16829 3968
rect 16771 3927 16829 3928
rect 19555 3968 19613 3969
rect 19555 3928 19564 3968
rect 19604 3928 19613 3968
rect 19555 3927 19613 3928
rect 19843 3968 19901 3969
rect 19843 3928 19852 3968
rect 19892 3928 19901 3968
rect 19843 3927 19901 3928
rect 23883 3968 23925 3977
rect 23883 3928 23884 3968
rect 23924 3928 23925 3968
rect 23883 3919 23925 3928
rect 25507 3968 25565 3969
rect 25507 3928 25516 3968
rect 25556 3928 25565 3968
rect 25507 3927 25565 3928
rect 26763 3968 26805 3977
rect 26763 3928 26764 3968
rect 26804 3928 26805 3968
rect 26763 3919 26805 3928
rect 27523 3968 27581 3969
rect 27523 3928 27532 3968
rect 27572 3928 27581 3968
rect 27523 3927 27581 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 25611 3690 25653 3699
rect 25611 3650 25612 3690
rect 25652 3650 25653 3690
rect 25611 3641 25653 3650
rect 643 3632 701 3633
rect 643 3592 652 3632
rect 692 3592 701 3632
rect 643 3591 701 3592
rect 8035 3632 8093 3633
rect 8035 3592 8044 3632
rect 8084 3592 8093 3632
rect 8035 3591 8093 3592
rect 9379 3632 9437 3633
rect 9379 3592 9388 3632
rect 9428 3592 9437 3632
rect 9379 3591 9437 3592
rect 11395 3632 11453 3633
rect 11395 3592 11404 3632
rect 11444 3592 11453 3632
rect 11395 3591 11453 3592
rect 12355 3632 12413 3633
rect 12355 3592 12364 3632
rect 12404 3592 12413 3632
rect 12355 3591 12413 3592
rect 14467 3632 14525 3633
rect 14467 3592 14476 3632
rect 14516 3592 14525 3632
rect 14467 3591 14525 3592
rect 15043 3632 15101 3633
rect 15043 3592 15052 3632
rect 15092 3592 15101 3632
rect 15043 3591 15101 3592
rect 16291 3632 16349 3633
rect 16291 3592 16300 3632
rect 16340 3592 16349 3632
rect 16291 3591 16349 3592
rect 26571 3632 26613 3641
rect 26571 3592 26572 3632
rect 26612 3592 26613 3632
rect 26571 3583 26613 3592
rect 27339 3632 27381 3641
rect 27339 3592 27340 3632
rect 27380 3592 27381 3632
rect 27339 3583 27381 3592
rect 27619 3632 27677 3633
rect 27619 3592 27628 3632
rect 27668 3592 27677 3632
rect 27619 3591 27677 3592
rect 16779 3548 16821 3557
rect 16779 3508 16780 3548
rect 16820 3508 16821 3548
rect 16779 3499 16821 3508
rect 24931 3548 24989 3549
rect 24931 3508 24940 3548
rect 24980 3508 24989 3548
rect 24931 3507 24989 3508
rect 11008 3485 11066 3486
rect 5451 3464 5493 3473
rect 5451 3424 5452 3464
rect 5492 3424 5493 3464
rect 5451 3415 5493 3424
rect 5827 3464 5885 3465
rect 5827 3424 5836 3464
rect 5876 3424 5885 3464
rect 5827 3423 5885 3424
rect 6691 3464 6749 3465
rect 6691 3424 6700 3464
rect 6740 3424 6749 3464
rect 6691 3423 6749 3424
rect 8707 3464 8765 3465
rect 8707 3424 8716 3464
rect 8756 3424 8765 3464
rect 8707 3423 8765 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 9483 3464 9525 3473
rect 9483 3424 9484 3464
rect 9524 3424 9525 3464
rect 9483 3415 9525 3424
rect 10531 3464 10589 3465
rect 10531 3424 10540 3464
rect 10580 3424 10589 3464
rect 11008 3445 11017 3485
rect 11057 3445 11066 3485
rect 11008 3444 11066 3445
rect 11211 3464 11253 3473
rect 10531 3423 10589 3424
rect 11211 3424 11212 3464
rect 11252 3424 11253 3464
rect 11211 3415 11253 3424
rect 12067 3464 12125 3465
rect 12067 3424 12076 3464
rect 12116 3424 12125 3464
rect 12067 3423 12125 3424
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 12459 3464 12501 3473
rect 12459 3424 12460 3464
rect 12500 3424 12501 3464
rect 12459 3415 12501 3424
rect 12547 3464 12605 3465
rect 12547 3424 12556 3464
rect 12596 3424 12605 3464
rect 12547 3423 12605 3424
rect 14563 3464 14621 3465
rect 14563 3424 14572 3464
rect 14612 3424 14621 3464
rect 14563 3423 14621 3424
rect 14955 3464 14997 3473
rect 14955 3424 14956 3464
rect 14996 3424 14997 3464
rect 14955 3415 14997 3424
rect 15147 3464 15189 3473
rect 15147 3424 15148 3464
rect 15188 3424 15189 3464
rect 15147 3415 15189 3424
rect 15235 3464 15293 3465
rect 15235 3424 15244 3464
rect 15284 3424 15293 3464
rect 15235 3423 15293 3424
rect 15427 3464 15485 3465
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 16203 3464 16245 3473
rect 16203 3424 16204 3464
rect 16244 3424 16245 3464
rect 16203 3415 16245 3424
rect 16395 3464 16437 3473
rect 16395 3424 16396 3464
rect 16436 3424 16437 3464
rect 16395 3415 16437 3424
rect 16483 3464 16541 3465
rect 16483 3424 16492 3464
rect 16532 3424 16541 3464
rect 16483 3423 16541 3424
rect 17155 3464 17213 3465
rect 17155 3424 17164 3464
rect 17204 3424 17213 3464
rect 17155 3423 17213 3424
rect 18019 3464 18077 3465
rect 18019 3424 18028 3464
rect 18068 3424 18077 3464
rect 18019 3423 18077 3424
rect 19747 3464 19805 3465
rect 19747 3424 19756 3464
rect 19796 3424 19805 3464
rect 19747 3423 19805 3424
rect 20427 3464 20469 3473
rect 20427 3424 20428 3464
rect 20468 3424 20469 3464
rect 20427 3415 20469 3424
rect 20619 3464 20661 3473
rect 20619 3424 20620 3464
rect 20660 3424 20661 3464
rect 20619 3415 20661 3424
rect 20995 3464 21053 3465
rect 20995 3424 21004 3464
rect 21044 3424 21053 3464
rect 20995 3423 21053 3424
rect 21859 3464 21917 3465
rect 21859 3424 21868 3464
rect 21908 3424 21917 3464
rect 21859 3423 21917 3424
rect 23019 3464 23061 3473
rect 23019 3424 23020 3464
rect 23060 3424 23061 3464
rect 23019 3415 23061 3424
rect 23299 3464 23357 3465
rect 23299 3424 23308 3464
rect 23348 3424 23357 3464
rect 23299 3423 23357 3424
rect 25123 3464 25181 3465
rect 25123 3424 25132 3464
rect 25172 3424 25181 3464
rect 25123 3423 25181 3424
rect 25411 3464 25469 3465
rect 25411 3424 25420 3464
rect 25460 3424 25469 3464
rect 25411 3423 25469 3424
rect 25803 3464 25845 3473
rect 25803 3424 25804 3464
rect 25844 3424 25845 3464
rect 25699 3422 25757 3423
rect 7851 3380 7893 3389
rect 7851 3340 7852 3380
rect 7892 3340 7893 3380
rect 7851 3331 7893 3340
rect 15531 3380 15573 3389
rect 15531 3340 15532 3380
rect 15572 3340 15573 3380
rect 15531 3331 15573 3340
rect 15723 3380 15765 3389
rect 25699 3382 25708 3422
rect 25748 3382 25757 3422
rect 25803 3415 25845 3424
rect 26475 3464 26517 3473
rect 26475 3424 26476 3464
rect 26516 3424 26517 3464
rect 26475 3415 26517 3424
rect 26667 3464 26709 3473
rect 26667 3424 26668 3464
rect 26708 3424 26709 3464
rect 26667 3415 26709 3424
rect 26851 3464 26909 3465
rect 26851 3424 26860 3464
rect 26900 3424 26909 3464
rect 26851 3423 26909 3424
rect 27235 3464 27293 3465
rect 27235 3424 27244 3464
rect 27284 3424 27293 3464
rect 27235 3423 27293 3424
rect 28291 3464 28349 3465
rect 28291 3424 28300 3464
rect 28340 3424 28349 3464
rect 28291 3423 28349 3424
rect 28491 3464 28533 3473
rect 28491 3424 28492 3464
rect 28532 3424 28533 3464
rect 28491 3415 28533 3424
rect 29155 3464 29213 3465
rect 29155 3424 29164 3464
rect 29204 3424 29213 3464
rect 29155 3423 29213 3424
rect 29355 3464 29397 3473
rect 29355 3424 29356 3464
rect 29396 3424 29397 3464
rect 29355 3415 29397 3424
rect 29731 3464 29789 3465
rect 29731 3424 29740 3464
rect 29780 3424 29789 3464
rect 29731 3423 29789 3424
rect 30595 3464 30653 3465
rect 30595 3424 30604 3464
rect 30644 3424 30653 3464
rect 30595 3423 30653 3424
rect 31843 3464 31901 3465
rect 31843 3424 31852 3464
rect 31892 3424 31901 3464
rect 31843 3423 31901 3424
rect 25699 3381 25757 3382
rect 15723 3340 15724 3380
rect 15764 3340 15765 3380
rect 15723 3331 15765 3340
rect 12747 3296 12789 3305
rect 12747 3256 12748 3296
rect 12788 3256 12789 3296
rect 12747 3247 12789 3256
rect 13323 3296 13365 3305
rect 13323 3256 13324 3296
rect 13364 3256 13365 3296
rect 13323 3247 13365 3256
rect 15627 3296 15669 3305
rect 15627 3256 15628 3296
rect 15668 3256 15669 3296
rect 15627 3247 15669 3256
rect 9675 3212 9717 3221
rect 9675 3172 9676 3212
rect 9716 3172 9717 3212
rect 9675 3163 9717 3172
rect 9859 3212 9917 3213
rect 9859 3172 9868 3212
rect 9908 3172 9917 3212
rect 9859 3171 9917 3172
rect 11115 3212 11157 3221
rect 11115 3172 11116 3212
rect 11156 3172 11157 3212
rect 11115 3163 11157 3172
rect 14755 3212 14813 3213
rect 14755 3172 14764 3212
rect 14804 3172 14813 3212
rect 14755 3171 14813 3172
rect 19171 3212 19229 3213
rect 19171 3172 19180 3212
rect 19220 3172 19229 3212
rect 19171 3171 19229 3172
rect 23971 3212 24029 3213
rect 23971 3172 23980 3212
rect 24020 3172 24029 3212
rect 23971 3171 24029 3172
rect 26091 3212 26133 3221
rect 26091 3172 26092 3212
rect 26132 3172 26133 3212
rect 26091 3163 26133 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 6699 2876 6741 2885
rect 6699 2836 6700 2876
rect 6740 2836 6741 2876
rect 6699 2827 6741 2836
rect 9387 2876 9429 2885
rect 9387 2836 9388 2876
rect 9428 2836 9429 2876
rect 9387 2827 9429 2836
rect 11979 2876 12021 2885
rect 11979 2836 11980 2876
rect 12020 2836 12021 2876
rect 11979 2827 12021 2836
rect 15235 2876 15293 2877
rect 15235 2836 15244 2876
rect 15284 2836 15293 2876
rect 15235 2835 15293 2836
rect 16875 2876 16917 2885
rect 16875 2836 16876 2876
rect 16916 2836 16917 2876
rect 16875 2827 16917 2836
rect 21379 2876 21437 2877
rect 21379 2836 21388 2876
rect 21428 2836 21437 2876
rect 21379 2835 21437 2836
rect 26371 2876 26429 2877
rect 26371 2836 26380 2876
rect 26420 2836 26429 2876
rect 26371 2835 26429 2836
rect 26563 2876 26621 2877
rect 26563 2836 26572 2876
rect 26612 2836 26621 2876
rect 26563 2835 26621 2836
rect 29835 2876 29877 2885
rect 29835 2836 29836 2876
rect 29876 2836 29877 2876
rect 29835 2827 29877 2836
rect 30211 2876 30269 2877
rect 30211 2836 30220 2876
rect 30260 2836 30269 2876
rect 30211 2835 30269 2836
rect 6891 2792 6933 2801
rect 6891 2752 6892 2792
rect 6932 2752 6933 2792
rect 6891 2743 6933 2752
rect 9195 2792 9237 2801
rect 9195 2752 9196 2792
rect 9236 2752 9237 2792
rect 9195 2743 9237 2752
rect 17259 2792 17301 2801
rect 17259 2752 17260 2792
rect 17300 2752 17301 2792
rect 17259 2743 17301 2752
rect 25515 2792 25557 2801
rect 25515 2752 25516 2792
rect 25556 2752 25557 2792
rect 25515 2743 25557 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 6123 2708 6165 2717
rect 6123 2668 6124 2708
rect 6164 2668 6165 2708
rect 6123 2659 6165 2668
rect 8523 2708 8565 2717
rect 8523 2668 8524 2708
rect 8564 2668 8565 2708
rect 8523 2659 8565 2668
rect 19939 2708 19997 2709
rect 19939 2668 19948 2708
rect 19988 2668 19997 2708
rect 19939 2667 19997 2668
rect 21963 2708 22005 2717
rect 21963 2668 21964 2708
rect 22004 2668 22005 2708
rect 21963 2659 22005 2668
rect 24555 2708 24597 2717
rect 24555 2668 24556 2708
rect 24596 2668 24597 2708
rect 24555 2659 24597 2668
rect 6027 2624 6069 2633
rect 6027 2584 6028 2624
rect 6068 2584 6069 2624
rect 6027 2575 6069 2584
rect 6219 2624 6261 2633
rect 6219 2584 6220 2624
rect 6260 2584 6261 2624
rect 6219 2575 6261 2584
rect 6403 2624 6461 2625
rect 6403 2584 6412 2624
rect 6452 2584 6461 2624
rect 6403 2583 6461 2584
rect 6507 2624 6549 2633
rect 6507 2584 6508 2624
rect 6548 2584 6549 2624
rect 6507 2575 6549 2584
rect 6699 2624 6741 2633
rect 6699 2584 6700 2624
rect 6740 2584 6741 2624
rect 6699 2575 6741 2584
rect 8043 2624 8085 2633
rect 8043 2584 8044 2624
rect 8084 2584 8085 2624
rect 8043 2575 8085 2584
rect 8139 2624 8181 2633
rect 8139 2584 8140 2624
rect 8180 2584 8181 2624
rect 8139 2575 8181 2584
rect 8227 2624 8285 2625
rect 8227 2584 8236 2624
rect 8276 2584 8285 2624
rect 8227 2583 8285 2584
rect 8427 2624 8469 2633
rect 8427 2584 8428 2624
rect 8468 2584 8469 2624
rect 8427 2575 8469 2584
rect 8619 2624 8661 2633
rect 8619 2584 8620 2624
rect 8660 2584 8661 2624
rect 8619 2575 8661 2584
rect 9195 2624 9237 2633
rect 9195 2584 9196 2624
rect 9236 2584 9237 2624
rect 9195 2575 9237 2584
rect 9579 2624 9621 2633
rect 9579 2584 9580 2624
rect 9620 2584 9621 2624
rect 9579 2575 9621 2584
rect 9955 2624 10013 2625
rect 9955 2584 9964 2624
rect 10004 2584 10013 2624
rect 9955 2583 10013 2584
rect 10819 2624 10877 2625
rect 10819 2584 10828 2624
rect 10868 2584 10877 2624
rect 10819 2583 10877 2584
rect 12067 2624 12125 2625
rect 12067 2584 12076 2624
rect 12116 2584 12125 2624
rect 12067 2583 12125 2584
rect 12843 2624 12885 2633
rect 12843 2584 12844 2624
rect 12884 2584 12885 2624
rect 12843 2575 12885 2584
rect 13219 2624 13277 2625
rect 13219 2584 13228 2624
rect 13268 2584 13277 2624
rect 13219 2583 13277 2584
rect 14083 2624 14141 2625
rect 14083 2584 14092 2624
rect 14132 2584 14141 2624
rect 14083 2583 14141 2584
rect 15715 2624 15773 2625
rect 15715 2584 15724 2624
rect 15764 2584 15773 2624
rect 15715 2583 15773 2584
rect 15907 2624 15965 2625
rect 15907 2584 15916 2624
rect 15956 2584 15965 2624
rect 15907 2583 15965 2584
rect 16099 2624 16157 2625
rect 16099 2584 16108 2624
rect 16148 2584 16157 2624
rect 16099 2583 16157 2584
rect 16299 2624 16341 2633
rect 16299 2584 16300 2624
rect 16340 2584 16341 2624
rect 16299 2575 16341 2584
rect 16483 2624 16541 2625
rect 16483 2584 16492 2624
rect 16532 2584 16541 2624
rect 16483 2583 16541 2584
rect 16683 2624 16725 2633
rect 16683 2584 16684 2624
rect 16724 2584 16725 2624
rect 16683 2575 16725 2584
rect 16963 2624 17021 2625
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 16963 2583 17021 2584
rect 18691 2624 18749 2625
rect 18691 2584 18700 2624
rect 18740 2584 18749 2624
rect 18691 2583 18749 2584
rect 20227 2624 20285 2625
rect 20227 2584 20236 2624
rect 20276 2584 20285 2624
rect 20227 2583 20285 2584
rect 20331 2624 20373 2633
rect 20331 2584 20332 2624
rect 20372 2584 20373 2624
rect 20331 2575 20373 2584
rect 20707 2624 20765 2625
rect 20707 2584 20716 2624
rect 20756 2584 20765 2624
rect 20707 2583 20765 2584
rect 23107 2624 23165 2625
rect 23107 2584 23116 2624
rect 23156 2584 23165 2624
rect 23107 2583 23165 2584
rect 23971 2624 24029 2625
rect 23971 2584 23980 2624
rect 24020 2584 24029 2624
rect 23971 2583 24029 2584
rect 24363 2624 24405 2633
rect 24363 2584 24364 2624
rect 24404 2584 24405 2624
rect 24363 2575 24405 2584
rect 25219 2624 25277 2625
rect 25219 2584 25228 2624
rect 25268 2584 25277 2624
rect 25219 2583 25277 2584
rect 25411 2624 25469 2625
rect 25411 2584 25420 2624
rect 25460 2584 25469 2624
rect 25411 2583 25469 2584
rect 25699 2624 25757 2625
rect 25699 2584 25708 2624
rect 25748 2584 25757 2624
rect 25699 2583 25757 2584
rect 27235 2624 27293 2625
rect 27235 2584 27244 2624
rect 27284 2584 27293 2624
rect 27235 2583 27293 2584
rect 27435 2624 27477 2633
rect 27435 2584 27436 2624
rect 27476 2584 27477 2624
rect 27435 2575 27477 2584
rect 27811 2624 27869 2625
rect 27811 2584 27820 2624
rect 27860 2584 27869 2624
rect 27811 2583 27869 2584
rect 28675 2624 28733 2625
rect 28675 2584 28684 2624
rect 28724 2584 28733 2624
rect 28675 2583 28733 2584
rect 30883 2624 30941 2625
rect 30883 2584 30892 2624
rect 30932 2584 30941 2624
rect 30883 2583 30941 2584
rect 16203 2540 16245 2549
rect 16203 2500 16204 2540
rect 16244 2500 16245 2540
rect 16203 2491 16245 2500
rect 16587 2540 16629 2549
rect 16587 2500 16588 2540
rect 16628 2500 16629 2540
rect 16587 2491 16629 2500
rect 18027 2540 18069 2549
rect 18027 2500 18028 2540
rect 18068 2500 18069 2540
rect 18027 2491 18069 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 26371 2456 26429 2457
rect 26371 2416 26380 2456
rect 26420 2416 26429 2456
rect 26371 2415 26429 2416
rect 26563 2456 26621 2457
rect 26563 2416 26572 2456
rect 26612 2416 26621 2456
rect 26563 2415 26621 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 20811 2120 20853 2129
rect 20811 2080 20812 2120
rect 20852 2080 20853 2120
rect 20811 2071 20853 2080
rect 22059 2120 22101 2129
rect 22059 2080 22060 2120
rect 22100 2080 22101 2120
rect 22059 2071 22101 2080
rect 29355 2120 29397 2129
rect 29355 2080 29356 2120
rect 29396 2080 29397 2120
rect 29355 2071 29397 2080
rect 15051 2036 15093 2045
rect 15051 1996 15052 2036
rect 15092 1996 15093 2036
rect 15051 1987 15093 1996
rect 9667 1952 9725 1953
rect 9667 1912 9676 1952
rect 9716 1912 9725 1952
rect 9667 1911 9725 1912
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 9963 1952 10005 1961
rect 9963 1912 9964 1952
rect 10004 1912 10005 1952
rect 9963 1903 10005 1912
rect 10731 1952 10773 1961
rect 10731 1912 10732 1952
rect 10772 1912 10773 1952
rect 10731 1903 10773 1912
rect 11107 1952 11165 1953
rect 11107 1912 11116 1952
rect 11156 1912 11165 1952
rect 11107 1911 11165 1912
rect 11971 1952 12029 1953
rect 11971 1912 11980 1952
rect 12020 1912 12029 1952
rect 11971 1911 12029 1912
rect 13131 1952 13173 1961
rect 13131 1912 13132 1952
rect 13172 1912 13173 1952
rect 13131 1903 13173 1912
rect 15427 1952 15485 1953
rect 15427 1912 15436 1952
rect 15476 1912 15485 1952
rect 15427 1911 15485 1912
rect 16291 1952 16349 1953
rect 16291 1912 16300 1952
rect 16340 1912 16349 1952
rect 16291 1911 16349 1912
rect 20995 1952 21053 1953
rect 20995 1912 21004 1952
rect 21044 1912 21053 1952
rect 20995 1911 21053 1912
rect 21283 1952 21341 1953
rect 21283 1912 21292 1952
rect 21332 1912 21341 1952
rect 21283 1911 21341 1912
rect 22531 1952 22589 1953
rect 22531 1912 22540 1952
rect 22580 1912 22589 1952
rect 22531 1911 22589 1912
rect 23595 1952 23637 1961
rect 23595 1912 23596 1952
rect 23636 1912 23637 1952
rect 23595 1903 23637 1912
rect 23971 1952 24029 1953
rect 23971 1912 23980 1952
rect 24020 1912 24029 1952
rect 23971 1911 24029 1912
rect 24835 1952 24893 1953
rect 24835 1912 24844 1952
rect 24884 1912 24893 1952
rect 24835 1911 24893 1912
rect 25995 1952 26037 1961
rect 25995 1912 25996 1952
rect 26036 1912 26037 1952
rect 25995 1903 26037 1912
rect 26283 1952 26325 1961
rect 26283 1912 26284 1952
rect 26324 1912 26325 1952
rect 26283 1903 26325 1912
rect 26659 1952 26717 1953
rect 26659 1912 26668 1952
rect 26708 1912 26717 1952
rect 26659 1911 26717 1912
rect 27523 1952 27581 1953
rect 27523 1912 27532 1952
rect 27572 1912 27581 1952
rect 27523 1911 27581 1912
rect 28771 1952 28829 1953
rect 28771 1912 28780 1952
rect 28820 1912 28829 1952
rect 28771 1911 28829 1912
rect 29443 1952 29501 1953
rect 29443 1912 29452 1952
rect 29492 1912 29501 1952
rect 29443 1911 29501 1912
rect 9963 1784 10005 1793
rect 9963 1744 9964 1784
rect 10004 1744 10005 1784
rect 9963 1735 10005 1744
rect 10155 1784 10197 1793
rect 10155 1744 10156 1784
rect 10196 1744 10197 1784
rect 10155 1735 10197 1744
rect 17443 1700 17501 1701
rect 17443 1660 17452 1700
rect 17492 1660 17501 1700
rect 17443 1659 17501 1660
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 26275 1364 26333 1365
rect 26275 1324 26284 1364
rect 26324 1324 26333 1364
rect 26275 1323 26333 1324
rect 10155 1280 10197 1289
rect 10155 1240 10156 1280
rect 10196 1240 10197 1280
rect 10155 1231 10197 1240
rect 11203 1280 11261 1281
rect 11203 1240 11212 1280
rect 11252 1240 11261 1280
rect 11203 1239 11261 1240
rect 15531 1280 15573 1289
rect 15531 1240 15532 1280
rect 15572 1240 15573 1280
rect 15531 1231 15573 1240
rect 24355 1280 24413 1281
rect 24355 1240 24364 1280
rect 24404 1240 24413 1280
rect 24355 1239 24413 1240
rect 25219 1196 25277 1197
rect 25219 1156 25228 1196
rect 25268 1156 25277 1196
rect 25219 1155 25277 1156
rect 10243 1112 10301 1113
rect 10243 1072 10252 1112
rect 10292 1072 10301 1112
rect 10243 1071 10301 1072
rect 11875 1112 11933 1113
rect 11875 1072 11884 1112
rect 11924 1072 11933 1112
rect 11875 1071 11933 1072
rect 23299 1112 23357 1113
rect 23299 1072 23308 1112
rect 23348 1072 23357 1112
rect 23299 1071 23357 1072
rect 23979 1112 24021 1121
rect 23979 1072 23980 1112
rect 24020 1072 24021 1112
rect 23979 1063 24021 1072
rect 25027 1112 25085 1113
rect 25027 1072 25036 1112
rect 25076 1072 25085 1112
rect 25027 1071 25085 1072
rect 25507 1112 25565 1113
rect 25507 1072 25516 1112
rect 25556 1072 25565 1112
rect 25507 1071 25565 1072
rect 25611 1112 25653 1121
rect 25611 1072 25612 1112
rect 25652 1072 25653 1112
rect 25611 1063 25653 1072
rect 26083 1112 26141 1113
rect 26083 1072 26092 1112
rect 26132 1072 26141 1112
rect 26083 1071 26141 1072
rect 26467 1112 26525 1113
rect 26467 1072 26476 1112
rect 26516 1072 26525 1112
rect 26467 1071 26525 1072
rect 26667 1112 26709 1121
rect 26667 1072 26668 1112
rect 26708 1072 26709 1112
rect 26667 1063 26709 1072
rect 26755 1112 26813 1113
rect 26755 1072 26764 1112
rect 26804 1072 26813 1112
rect 26755 1071 26813 1072
rect 25987 944 26045 945
rect 25987 904 25996 944
rect 26036 904 26045 944
rect 25987 903 26045 904
rect 26475 944 26517 953
rect 26475 904 26476 944
rect 26516 904 26517 944
rect 26475 895 26517 904
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 27820 37528 27860 37568
rect 27628 37360 27668 37400
rect 30988 37360 31028 37400
rect 31756 37360 31796 37400
rect 32428 37360 32468 37400
rect 27532 37192 27572 37232
rect 30892 37192 30932 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 31660 36856 31700 36896
rect 33292 36772 33332 36812
rect 12556 36688 12596 36728
rect 12652 36688 12692 36728
rect 12844 36688 12884 36728
rect 13708 36688 13748 36728
rect 16108 36688 16148 36728
rect 25612 36688 25652 36728
rect 25708 36688 25748 36728
rect 25900 36688 25940 36728
rect 26092 36688 26132 36728
rect 26188 36688 26228 36728
rect 26284 36688 26324 36728
rect 26380 36688 26420 36728
rect 27724 36688 27764 36728
rect 28012 36688 28052 36728
rect 28684 36688 28724 36728
rect 28972 36688 29012 36728
rect 30508 36688 30548 36728
rect 30796 36688 30836 36728
rect 32332 36688 32372 36728
rect 32620 36688 32660 36728
rect 36076 36688 36116 36728
rect 40012 36688 40052 36728
rect 41068 36688 41108 36728
rect 9964 36520 10004 36560
rect 12844 36520 12884 36560
rect 13900 36520 13940 36560
rect 16300 36520 16340 36560
rect 24940 36520 24980 36560
rect 25900 36520 25940 36560
rect 29644 36520 29684 36560
rect 33484 36520 33524 36560
rect 36460 36520 36500 36560
rect 39148 36520 39188 36560
rect 13036 36436 13076 36476
rect 15436 36436 15476 36476
rect 27052 36436 27092 36476
rect 29068 36436 29108 36476
rect 29836 36436 29876 36476
rect 31468 36436 31508 36476
rect 35404 36436 35444 36476
rect 39340 36436 39380 36476
rect 40396 36436 40436 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 12556 36100 12596 36140
rect 29452 36100 29492 36140
rect 32044 36100 32084 36140
rect 32236 36100 32276 36140
rect 35596 36100 35636 36140
rect 19756 36016 19796 36056
rect 23884 36016 23924 36056
rect 9868 35848 9908 35888
rect 10732 35848 10772 35888
rect 12460 35848 12500 35888
rect 12748 35848 12788 35888
rect 13132 35848 13172 35888
rect 13996 35848 14036 35888
rect 15340 35848 15380 35888
rect 15724 35848 15764 35888
rect 16588 35848 16628 35888
rect 19564 35848 19604 35888
rect 21772 35848 21812 35888
rect 24460 35848 24500 35888
rect 24844 35848 24884 35888
rect 25708 35848 25748 35888
rect 27436 35848 27476 35888
rect 28300 35848 28340 35888
rect 29644 35848 29684 35888
rect 30028 35848 30068 35888
rect 30892 35848 30932 35888
rect 32236 35848 32276 35888
rect 32428 35848 32468 35888
rect 32524 35848 32564 35888
rect 32716 35848 32756 35888
rect 33100 35848 33140 35888
rect 33964 35848 34004 35888
rect 35212 35848 35252 35888
rect 36748 35848 36788 35888
rect 37612 35848 37652 35888
rect 37996 35848 38036 35888
rect 38188 35848 38228 35888
rect 38860 35848 38900 35888
rect 39052 35848 39092 35888
rect 39436 35848 39476 35888
rect 40300 35848 40340 35888
rect 9484 35764 9524 35804
rect 27052 35764 27092 35804
rect 11884 35680 11924 35720
rect 15148 35680 15188 35720
rect 17740 35680 17780 35720
rect 18892 35680 18932 35720
rect 21100 35680 21140 35720
rect 26860 35680 26900 35720
rect 32044 35680 32084 35720
rect 41452 35680 41492 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 9004 35344 9044 35384
rect 12268 35344 12308 35384
rect 27244 35344 27284 35384
rect 37612 35344 37652 35384
rect 38476 35344 38516 35384
rect 5932 35260 5972 35300
rect 13996 35260 14036 35300
rect 18796 35260 18836 35300
rect 23404 35260 23444 35300
rect 26380 35260 26420 35300
rect 29740 35260 29780 35300
rect 31372 35260 31412 35300
rect 33196 35260 33236 35300
rect 34636 35260 34676 35300
rect 36076 35260 36116 35300
rect 39052 35260 39092 35300
rect 39436 35260 39476 35300
rect 5356 35176 5396 35216
rect 5452 35176 5492 35216
rect 5644 35176 5684 35216
rect 5836 35176 5876 35216
rect 6028 35176 6068 35216
rect 6124 35176 6164 35216
rect 6988 35176 7028 35216
rect 8332 35176 8372 35216
rect 8812 35176 8852 35216
rect 8908 35176 8948 35216
rect 9100 35176 9140 35216
rect 9292 35176 9332 35216
rect 9676 35176 9716 35216
rect 10540 35176 10580 35216
rect 12940 35176 12980 35216
rect 13804 35176 13844 35216
rect 14092 35176 14132 35216
rect 14284 35176 14324 35216
rect 14380 35176 14420 35216
rect 14476 35176 14516 35216
rect 14572 35176 14612 35216
rect 15436 35176 15476 35216
rect 16300 35176 16340 35216
rect 16492 35176 16532 35216
rect 16684 35176 16724 35216
rect 16780 35176 16820 35216
rect 16972 35176 17012 35216
rect 17068 35176 17108 35216
rect 17164 35176 17204 35216
rect 17260 35176 17300 35216
rect 18316 35176 18356 35216
rect 19180 35176 19220 35216
rect 20044 35176 20084 35216
rect 22252 35176 22292 35216
rect 23788 35176 23828 35216
rect 24652 35176 24692 35216
rect 25996 35176 26036 35216
rect 26092 35176 26132 35216
rect 26284 35176 26324 35216
rect 26476 35176 26516 35216
rect 26572 35176 26612 35216
rect 26764 35176 26804 35216
rect 26860 35176 26900 35216
rect 27052 35176 27092 35216
rect 27916 35176 27956 35216
rect 29548 35176 29588 35216
rect 29644 35176 29684 35216
rect 29836 35176 29876 35216
rect 30412 35176 30452 35216
rect 30508 35176 30548 35216
rect 30604 35176 30644 35216
rect 30700 35176 30740 35216
rect 30988 35176 31028 35216
rect 31276 35176 31316 35216
rect 31948 35176 31988 35216
rect 32908 35176 32948 35216
rect 33100 35176 33140 35216
rect 34252 35176 34292 35216
rect 34732 35176 34772 35216
rect 35308 35176 35348 35216
rect 35404 35176 35444 35216
rect 35596 35176 35636 35216
rect 35788 35176 35828 35216
rect 35884 35176 35924 35216
rect 35980 35176 36020 35216
rect 36940 35176 36980 35216
rect 38092 35176 38132 35216
rect 38380 35176 38420 35216
rect 38572 35176 38612 35216
rect 38668 35176 38708 35216
rect 39148 35176 39188 35216
rect 39340 35176 39380 35216
rect 39532 35176 39572 35216
rect 39628 35176 39668 35216
rect 40108 35176 40148 35216
rect 40300 35176 40340 35216
rect 40876 35176 40916 35216
rect 41260 35176 41300 35216
rect 42124 35176 42164 35216
rect 44428 35176 44468 35216
rect 11692 35092 11732 35132
rect 25804 35092 25844 35132
rect 28492 35092 28532 35132
rect 37228 35092 37268 35132
rect 4492 35008 4532 35048
rect 7180 35008 7220 35048
rect 12076 35008 12116 35048
rect 17452 35008 17492 35048
rect 22444 35008 22484 35048
rect 27052 35008 27092 35048
rect 28300 35008 28340 35048
rect 28876 35008 28916 35048
rect 29260 35008 29300 35048
rect 30220 35008 30260 35048
rect 35116 35008 35156 35048
rect 40684 35008 40724 35048
rect 5644 34924 5684 34964
rect 6316 34924 6356 34964
rect 7660 34924 7700 34964
rect 12268 34924 12308 34964
rect 13132 34924 13172 34964
rect 14764 34924 14804 34964
rect 15628 34924 15668 34964
rect 16492 34924 16532 34964
rect 18412 34924 18452 34964
rect 21196 34924 21236 34964
rect 21580 34924 21620 34964
rect 31660 34924 31700 34964
rect 32236 34924 32276 34964
rect 33868 34924 33908 34964
rect 35596 34924 35636 34964
rect 36268 34924 36308 34964
rect 40204 34924 40244 34964
rect 43276 34924 43316 34964
rect 43756 34924 43796 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 6028 34588 6068 34628
rect 9388 34588 9428 34628
rect 10924 34588 10964 34628
rect 18316 34588 18356 34628
rect 24076 34588 24116 34628
rect 32524 34588 32564 34628
rect 41452 34588 41492 34628
rect 2572 34504 2612 34544
rect 10444 34504 10484 34544
rect 14188 34504 14228 34544
rect 28588 34504 28628 34544
rect 42604 34504 42644 34544
rect 43660 34504 43700 34544
rect 18124 34420 18164 34460
rect 42124 34420 42164 34460
rect 3628 34336 3668 34376
rect 4012 34336 4052 34376
rect 4876 34336 4916 34376
rect 6220 34336 6260 34376
rect 6604 34336 6644 34376
rect 7468 34336 7508 34376
rect 8812 34336 8852 34376
rect 8908 34336 8948 34376
rect 9100 34336 9140 34376
rect 9196 34336 9236 34376
rect 9388 34336 9428 34376
rect 9580 34336 9620 34376
rect 10252 34336 10292 34376
rect 10828 34336 10868 34376
rect 11212 34336 11252 34376
rect 11500 34336 11540 34376
rect 11596 34336 11636 34376
rect 11692 34336 11732 34376
rect 11884 34336 11924 34376
rect 11980 34336 12020 34376
rect 12076 34336 12116 34376
rect 12172 34336 12212 34376
rect 12364 34336 12404 34376
rect 12460 34336 12500 34376
rect 12556 34336 12596 34376
rect 12940 34336 12980 34376
rect 13036 34336 13076 34376
rect 13132 34336 13172 34376
rect 13228 34336 13268 34376
rect 13516 34336 13556 34376
rect 13804 34336 13844 34376
rect 14380 34336 14420 34376
rect 14476 34336 14516 34376
rect 14668 34336 14708 34376
rect 14764 34336 14804 34376
rect 14956 34336 14996 34376
rect 15148 34336 15188 34376
rect 15340 34336 15380 34376
rect 15436 34336 15476 34376
rect 16108 34336 16148 34376
rect 16972 34336 17012 34376
rect 19372 34378 19412 34418
rect 18988 34311 19028 34351
rect 19276 34336 19316 34376
rect 19468 34336 19508 34376
rect 21388 34336 21428 34376
rect 21772 34336 21812 34376
rect 22636 34336 22676 34376
rect 24172 34336 24212 34376
rect 24364 34336 24404 34376
rect 25036 34336 25076 34376
rect 25420 34336 25460 34376
rect 25516 34336 25556 34376
rect 25612 34336 25652 34376
rect 25708 34336 25748 34376
rect 25900 34336 25940 34376
rect 26860 34336 26900 34376
rect 27340 34336 27380 34376
rect 27436 34336 27476 34376
rect 27532 34336 27572 34376
rect 27628 34336 27668 34376
rect 27916 34336 27956 34376
rect 28204 34336 28244 34376
rect 28300 34336 28340 34376
rect 28780 34336 28820 34376
rect 29836 34336 29876 34376
rect 29932 34336 29972 34376
rect 30028 34336 30068 34376
rect 30124 34336 30164 34376
rect 31276 34336 31316 34376
rect 31660 34336 31700 34376
rect 31756 34336 31796 34376
rect 31948 34336 31988 34376
rect 32236 34336 32276 34376
rect 33196 34336 33236 34376
rect 33388 34336 33428 34376
rect 33772 34336 33812 34376
rect 34636 34336 34676 34376
rect 35980 34336 36020 34376
rect 36364 34336 36404 34376
rect 37228 34336 37268 34376
rect 38860 34336 38900 34376
rect 38956 34336 38996 34376
rect 39052 34336 39092 34376
rect 39148 34336 39188 34376
rect 39340 34336 39380 34376
rect 39436 34336 39476 34376
rect 39532 34336 39572 34376
rect 39628 34336 39668 34376
rect 39820 34336 39860 34376
rect 40012 34336 40052 34376
rect 40108 34336 40148 34376
rect 40396 34336 40436 34376
rect 40492 34336 40532 34376
rect 40588 34336 40628 34376
rect 40780 34336 40820 34376
rect 41644 34336 41684 34376
rect 41836 34336 41876 34376
rect 41932 34336 41972 34376
rect 42220 34336 42260 34376
rect 42796 34336 42836 34376
rect 42892 34336 42932 34376
rect 42988 34336 43028 34376
rect 44524 34336 44564 34376
rect 13900 34252 13940 34292
rect 14860 34252 14900 34292
rect 15724 34252 15764 34292
rect 39916 34252 39956 34292
rect 8620 34168 8660 34208
rect 11116 34168 11156 34208
rect 11404 34168 11444 34208
rect 12652 34168 12692 34208
rect 15244 34168 15284 34208
rect 19180 34168 19220 34208
rect 23788 34168 23828 34208
rect 29452 34168 29492 34208
rect 30796 34168 30836 34208
rect 31852 34168 31892 34208
rect 35788 34168 35828 34208
rect 38380 34168 38420 34208
rect 40300 34168 40340 34208
rect 41740 34168 41780 34208
rect 43084 34168 43124 34208
rect 43852 34168 43892 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 4588 33832 4628 33872
rect 6316 33832 6356 33872
rect 9484 33832 9524 33872
rect 11788 33832 11828 33872
rect 18796 33832 18836 33872
rect 21772 33832 21812 33872
rect 33868 33832 33908 33872
rect 36364 33832 36404 33872
rect 45964 33832 46004 33872
rect 4876 33748 4916 33788
rect 6988 33748 7028 33788
rect 9004 33748 9044 33788
rect 17644 33748 17684 33788
rect 25996 33748 26036 33788
rect 30412 33748 30452 33788
rect 32428 33748 32468 33788
rect 42124 33748 42164 33788
rect 1996 33664 2036 33704
rect 2380 33664 2420 33704
rect 3244 33664 3284 33704
rect 4684 33664 4724 33704
rect 4972 33664 5012 33704
rect 5068 33664 5108 33704
rect 5164 33664 5204 33704
rect 5356 33664 5396 33704
rect 6028 33664 6068 33704
rect 6412 33664 6452 33704
rect 6508 33664 6548 33704
rect 6604 33664 6644 33704
rect 7852 33664 7892 33704
rect 8620 33664 8660 33704
rect 8908 33664 8948 33704
rect 10444 33664 10484 33704
rect 10636 33664 10676 33704
rect 11596 33664 11636 33704
rect 12940 33664 12980 33704
rect 13804 33664 13844 33704
rect 14188 33664 14228 33704
rect 14380 33664 14420 33704
rect 15052 33664 15092 33704
rect 15916 33664 15956 33704
rect 17740 33664 17780 33704
rect 18028 33664 18068 33704
rect 18604 33664 18644 33704
rect 18700 33664 18740 33704
rect 18892 33664 18932 33704
rect 19276 33664 19316 33704
rect 20332 33664 20372 33704
rect 20908 33664 20948 33704
rect 21100 33664 21140 33704
rect 21196 33664 21236 33704
rect 21292 33664 21332 33704
rect 21388 33664 21428 33704
rect 21580 33664 21620 33704
rect 21676 33664 21716 33704
rect 21868 33664 21908 33704
rect 24172 33664 24212 33704
rect 25612 33664 25652 33704
rect 25900 33664 25940 33704
rect 26764 33664 26804 33704
rect 27628 33664 27668 33704
rect 29164 33664 29204 33704
rect 30028 33664 30068 33704
rect 30604 33664 30644 33704
rect 32140 33664 32180 33704
rect 33196 33664 33236 33704
rect 33676 33664 33716 33704
rect 33772 33664 33812 33704
rect 33964 33664 34004 33704
rect 34156 33664 34196 33704
rect 34252 33664 34292 33704
rect 34348 33664 34388 33704
rect 34444 33664 34484 33704
rect 36460 33664 36500 33704
rect 36556 33664 36596 33704
rect 36652 33664 36692 33704
rect 36844 33664 36884 33704
rect 37996 33664 38036 33704
rect 38092 33664 38132 33704
rect 38284 33664 38324 33704
rect 38476 33664 38516 33704
rect 38572 33664 38612 33704
rect 38764 33664 38804 33704
rect 38860 33664 38900 33704
rect 38956 33664 38996 33704
rect 39052 33664 39092 33704
rect 39244 33664 39284 33704
rect 40108 33664 40148 33704
rect 40780 33664 40820 33704
rect 41164 33664 41204 33704
rect 42892 33664 42932 33704
rect 43372 33664 43412 33704
rect 43564 33664 43604 33704
rect 43948 33664 43988 33704
rect 44812 33664 44852 33704
rect 4396 33580 4436 33620
rect 9676 33580 9716 33620
rect 20044 33580 20084 33620
rect 20812 33580 20852 33620
rect 25036 33580 25076 33620
rect 28012 33580 28052 33620
rect 37516 33580 37556 33620
rect 24364 33496 24404 33536
rect 27436 33496 27476 33536
rect 34636 33496 34676 33536
rect 39916 33496 39956 33536
rect 9292 33412 9332 33452
rect 10924 33412 10964 33452
rect 11788 33412 11828 33452
rect 15244 33412 15284 33452
rect 17356 33412 17396 33452
rect 19468 33412 19508 33452
rect 20428 33412 20468 33452
rect 23500 33412 23540 33452
rect 26284 33412 26324 33452
rect 31276 33412 31316 33452
rect 31468 33412 31508 33452
rect 38284 33412 38324 33452
rect 41836 33412 41876 33452
rect 43276 33412 43316 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4492 33076 4532 33116
rect 12940 33076 12980 33116
rect 13804 33076 13844 33116
rect 20332 33076 20372 33116
rect 30220 33076 30260 33116
rect 44140 33076 44180 33116
rect 1708 32992 1748 33032
rect 2380 32992 2420 33032
rect 5164 32992 5204 33032
rect 7084 32992 7124 33032
rect 21388 32992 21428 33032
rect 28684 32992 28724 33032
rect 34636 32992 34676 33032
rect 36940 32992 36980 33032
rect 41068 32992 41108 33032
rect 44812 32992 44852 33032
rect 47884 32992 47924 33032
rect 3052 32908 3092 32948
rect 11980 32908 12020 32948
rect 17260 32908 17300 32948
rect 18604 32908 18644 32948
rect 18700 32908 18740 32948
rect 25708 32908 25748 32948
rect 40300 32908 40340 32948
rect 2092 32824 2132 32864
rect 2188 32824 2228 32864
rect 2380 32824 2420 32864
rect 2572 32824 2612 32864
rect 2668 32824 2708 32864
rect 2764 32824 2804 32864
rect 2860 32824 2900 32864
rect 3724 32824 3764 32864
rect 4012 32824 4052 32864
rect 4108 32824 4148 32864
rect 4204 32824 4244 32864
rect 4300 32824 4340 32864
rect 4492 32824 4532 32864
rect 4684 32824 4724 32864
rect 4780 32824 4820 32864
rect 6028 32824 6068 32864
rect 6412 32824 6452 32864
rect 6508 32824 6548 32864
rect 6604 32824 6644 32864
rect 6796 32824 6836 32864
rect 6892 32824 6932 32864
rect 7084 32824 7124 32864
rect 7276 32824 7316 32864
rect 8140 32824 8180 32864
rect 9004 32824 9044 32864
rect 9964 32824 10004 32864
rect 10252 32824 10292 32864
rect 10444 32824 10484 32864
rect 11116 32824 11156 32864
rect 13228 32824 13268 32864
rect 13516 32824 13556 32864
rect 13612 32824 13652 32864
rect 13804 32824 13844 32864
rect 14668 32824 14708 32864
rect 14860 32824 14900 32864
rect 15244 32824 15284 32864
rect 16108 32824 16148 32864
rect 17644 32833 17684 32873
rect 18124 32824 18164 32864
rect 19084 32824 19124 32864
rect 19180 32824 19220 32864
rect 19468 32824 19508 32864
rect 19660 32824 19700 32864
rect 19756 32824 19796 32864
rect 20044 32824 20084 32864
rect 23308 32824 23348 32864
rect 23692 32824 23732 32864
rect 24556 32824 24596 32864
rect 25996 32824 26036 32864
rect 26092 32824 26132 32864
rect 26188 32824 26228 32864
rect 26380 32824 26420 32864
rect 27052 32824 27092 32864
rect 27244 32824 27284 32864
rect 27532 32824 27572 32864
rect 27628 32824 27668 32864
rect 27724 32824 27764 32864
rect 28012 32824 28052 32864
rect 29068 32824 29108 32864
rect 29164 32824 29204 32864
rect 29356 32824 29396 32864
rect 30508 32824 30548 32864
rect 30892 32824 30932 32864
rect 31084 32824 31124 32864
rect 31468 32824 31508 32864
rect 32332 32824 32372 32864
rect 34444 32824 34484 32864
rect 36076 32824 36116 32864
rect 37324 32824 37364 32864
rect 37612 32824 37652 32864
rect 37900 32824 37940 32864
rect 38284 32824 38324 32864
rect 39148 32824 39188 32864
rect 40492 32824 40532 32864
rect 40684 32824 40724 32864
rect 41260 32824 41300 32864
rect 41356 32824 41396 32864
rect 41452 32824 41492 32864
rect 41548 32824 41588 32864
rect 41740 32824 41780 32864
rect 42124 32824 42164 32864
rect 42988 32824 43028 32864
rect 45676 32824 45716 32864
rect 47692 32824 47732 32864
rect 5356 32740 5396 32780
rect 8812 32740 8852 32780
rect 17452 32740 17492 32780
rect 20908 32740 20948 32780
rect 37228 32740 37268 32780
rect 40588 32740 40628 32780
rect 6316 32656 6356 32696
rect 7948 32656 7988 32696
rect 13996 32656 14036 32696
rect 19564 32656 19604 32696
rect 25900 32656 25940 32696
rect 27340 32656 27380 32696
rect 27820 32656 27860 32696
rect 29260 32656 29300 32696
rect 30796 32656 30836 32696
rect 33484 32656 33524 32696
rect 33772 32656 33812 32696
rect 36748 32656 36788 32696
rect 45004 32656 45044 32696
rect 47020 32656 47060 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 4108 32320 4148 32360
rect 7372 32320 7412 32360
rect 7564 32320 7604 32360
rect 7948 32320 7988 32360
rect 14284 32320 14324 32360
rect 14956 32320 14996 32360
rect 15148 32320 15188 32360
rect 18220 32320 18260 32360
rect 19084 32320 19124 32360
rect 20140 32320 20180 32360
rect 23596 32320 23636 32360
rect 27244 32320 27284 32360
rect 28492 32320 28532 32360
rect 31852 32320 31892 32360
rect 36076 32320 36116 32360
rect 37708 32320 37748 32360
rect 40204 32320 40244 32360
rect 42124 32320 42164 32360
rect 43948 32320 43988 32360
rect 47116 32320 47156 32360
rect 1324 32236 1364 32276
rect 4972 32236 5012 32276
rect 8428 32236 8468 32276
rect 22540 32236 22580 32276
rect 33676 32236 33716 32276
rect 44716 32236 44756 32276
rect 1708 32152 1748 32192
rect 2572 32152 2612 32192
rect 4780 32177 4820 32217
rect 5356 32152 5396 32192
rect 6220 32152 6260 32192
rect 7660 32152 7700 32192
rect 8044 32152 8084 32192
rect 8140 32152 8180 32192
rect 8236 32152 8276 32192
rect 8812 32152 8852 32192
rect 9676 32152 9716 32192
rect 11020 32152 11060 32192
rect 11884 32152 11924 32192
rect 12268 32152 12308 32192
rect 13132 32152 13172 32192
rect 14860 32152 14900 32192
rect 15340 32152 15380 32192
rect 3724 32068 3764 32108
rect 15244 32110 15284 32150
rect 15436 32152 15476 32192
rect 15628 32152 15668 32192
rect 15724 32152 15764 32192
rect 15820 32152 15860 32192
rect 15916 32152 15956 32192
rect 16108 32152 16148 32192
rect 16780 32152 16820 32192
rect 17644 32152 17684 32192
rect 17932 32152 17972 32192
rect 18028 32152 18068 32192
rect 18124 32152 18164 32192
rect 18412 32152 18452 32192
rect 19276 32152 19316 32192
rect 19948 32152 19988 32192
rect 21292 32152 21332 32192
rect 22156 32152 22196 32192
rect 23500 32152 23540 32192
rect 23692 32152 23732 32192
rect 23788 32152 23828 32192
rect 24844 32152 24884 32192
rect 25228 32152 25268 32192
rect 26092 32152 26132 32192
rect 27532 32152 27572 32192
rect 27820 32152 27860 32192
rect 27916 32152 27956 32192
rect 28396 32152 28436 32192
rect 29356 32152 29396 32192
rect 30508 32152 30548 32192
rect 30892 32152 30932 32192
rect 31180 32152 31220 32192
rect 31276 32152 31316 32192
rect 31948 32152 31988 32192
rect 32044 32152 32084 32192
rect 32140 32152 32180 32192
rect 32332 32152 32372 32192
rect 32428 32152 32468 32192
rect 32524 32152 32564 32192
rect 32620 32152 32660 32192
rect 33484 32152 33524 32192
rect 34060 32152 34100 32192
rect 34924 32152 34964 32192
rect 36652 32152 36692 32192
rect 37612 32152 37652 32192
rect 37996 32152 38036 32192
rect 38188 32152 38228 32192
rect 39244 32152 39284 32192
rect 40108 32152 40148 32192
rect 40492 32152 40532 32192
rect 41452 32152 41492 32192
rect 41932 32152 41972 32192
rect 42028 32152 42068 32192
rect 42220 32152 42260 32192
rect 42412 32152 42452 32192
rect 42508 32152 42548 32192
rect 42700 32152 42740 32192
rect 42892 32152 42932 32192
rect 42988 32152 43028 32192
rect 43084 32152 43124 32192
rect 43180 32152 43220 32192
rect 43468 32152 43508 32192
rect 45100 32152 45140 32192
rect 45964 32152 46004 32192
rect 48076 32152 48116 32192
rect 48268 32152 48308 32192
rect 48364 32152 48404 32192
rect 48460 32152 48500 32192
rect 48556 32152 48596 32192
rect 49804 32152 49844 32192
rect 10828 32068 10868 32108
rect 14668 31984 14708 32024
rect 38380 31984 38420 32024
rect 39052 31984 39092 32024
rect 4108 31900 4148 31940
rect 7372 31900 7412 31940
rect 11692 31900 11732 31940
rect 16972 31900 17012 31940
rect 28204 31900 28244 31940
rect 28684 31900 28724 31940
rect 30028 31900 30068 31940
rect 31564 31900 31604 31940
rect 32812 31900 32852 31940
rect 36556 31900 36596 31940
rect 39916 31900 39956 31940
rect 42700 31900 42740 31940
rect 47116 31900 47156 31940
rect 47404 31900 47444 31940
rect 49132 31900 49172 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 11500 31564 11540 31604
rect 12268 31564 12308 31604
rect 42028 31564 42068 31604
rect 49708 31564 49748 31604
rect 1900 31480 1940 31520
rect 3436 31480 3476 31520
rect 5548 31480 5588 31520
rect 6700 31480 6740 31520
rect 7372 31480 7412 31520
rect 7660 31480 7700 31520
rect 7852 31480 7892 31520
rect 8332 31480 8372 31520
rect 9964 31480 10004 31520
rect 10444 31480 10484 31520
rect 11692 31480 11732 31520
rect 14092 31480 14132 31520
rect 16780 31480 16820 31520
rect 19372 31480 19412 31520
rect 19756 31480 19796 31520
rect 20812 31480 20852 31520
rect 23020 31480 23060 31520
rect 24076 31480 24116 31520
rect 24556 31480 24596 31520
rect 28780 31480 28820 31520
rect 33100 31480 33140 31520
rect 34540 31480 34580 31520
rect 45100 31480 45140 31520
rect 46444 31480 46484 31520
rect 10828 31396 10868 31436
rect 13324 31396 13364 31436
rect 3532 31312 3572 31352
rect 3820 31312 3860 31352
rect 4012 31312 4052 31352
rect 4108 31312 4148 31352
rect 4204 31312 4244 31352
rect 4300 31312 4340 31352
rect 4492 31312 4532 31352
rect 4684 31312 4724 31352
rect 4780 31312 4820 31352
rect 4972 31312 5012 31352
rect 5068 31312 5108 31352
rect 5260 31312 5300 31352
rect 5356 31312 5396 31352
rect 5548 31312 5588 31352
rect 6124 31312 6164 31352
rect 6988 31312 7028 31352
rect 7564 31312 7604 31352
rect 7948 31312 7988 31352
rect 8524 31312 8564 31352
rect 8620 31312 8660 31352
rect 8812 31312 8852 31352
rect 9676 31312 9716 31352
rect 10060 31312 10100 31352
rect 11884 31312 11924 31352
rect 12268 31312 12308 31352
rect 12460 31312 12500 31352
rect 12556 31312 12596 31352
rect 12748 31312 12788 31352
rect 12844 31312 12884 31352
rect 12940 31312 12980 31352
rect 13036 31312 13076 31352
rect 13228 31312 13268 31352
rect 13612 31312 13652 31352
rect 13804 31312 13844 31352
rect 14380 31312 14420 31352
rect 14476 31312 14516 31352
rect 14764 31312 14804 31352
rect 15244 31312 15284 31352
rect 15916 31312 15956 31352
rect 16204 31312 16244 31352
rect 16492 31312 16532 31352
rect 16588 31312 16628 31352
rect 16780 31312 16820 31352
rect 16972 31312 17012 31352
rect 17356 31312 17396 31352
rect 18220 31312 18260 31352
rect 20620 31312 20660 31352
rect 20812 31312 20852 31352
rect 21004 31312 21044 31352
rect 21100 31312 21140 31352
rect 21292 31312 21332 31352
rect 24172 31312 24212 31352
rect 25420 31312 25460 31352
rect 25900 31312 25940 31352
rect 26092 31312 26132 31352
rect 26188 31312 26228 31352
rect 26380 31312 26420 31352
rect 27052 31312 27092 31352
rect 27340 31312 27380 31352
rect 27436 31312 27476 31352
rect 27532 31312 27572 31352
rect 27628 31312 27668 31352
rect 27820 31312 27860 31352
rect 27916 31312 27956 31352
rect 28108 31312 28148 31352
rect 28300 31312 28340 31352
rect 28972 31312 29012 31352
rect 29356 31312 29396 31352
rect 30220 31312 30260 31352
rect 31564 31312 31604 31352
rect 32524 31312 32564 31352
rect 33292 31312 33332 31352
rect 33388 31312 33428 31352
rect 33580 31312 33620 31352
rect 33868 31312 33908 31352
rect 33964 31312 34004 31352
rect 34060 31312 34100 31352
rect 34252 31312 34292 31352
rect 34348 31312 34388 31352
rect 34540 31312 34580 31352
rect 35020 31312 35060 31352
rect 35404 31312 35444 31352
rect 36268 31312 36308 31352
rect 38284 31312 38324 31352
rect 39724 31312 39764 31352
rect 40588 31312 40628 31352
rect 41932 31312 41972 31352
rect 42892 31312 42932 31352
rect 43084 31312 43124 31352
rect 44620 31312 44660 31352
rect 44812 31312 44852 31352
rect 44908 31312 44948 31352
rect 45100 31312 45140 31352
rect 45292 31312 45332 31352
rect 45580 31312 45620 31352
rect 45676 31312 45716 31352
rect 45772 31312 45812 31352
rect 45868 31312 45908 31352
rect 46252 31312 46292 31352
rect 47308 31312 47348 31352
rect 47692 31312 47732 31352
rect 48556 31312 48596 31352
rect 8716 31228 8756 31268
rect 13900 31228 13940 31268
rect 25996 31228 26036 31268
rect 28012 31228 28052 31268
rect 28396 31228 28436 31268
rect 33484 31228 33524 31268
rect 39340 31228 39380 31268
rect 45388 31228 45428 31268
rect 3724 31144 3764 31184
rect 4588 31144 4628 31184
rect 9004 31144 9044 31184
rect 13516 31144 13556 31184
rect 16108 31144 16148 31184
rect 19948 31144 19988 31184
rect 21388 31144 21428 31184
rect 24748 31144 24788 31184
rect 31372 31144 31412 31184
rect 32236 31144 32276 31184
rect 32428 31144 32468 31184
rect 33772 31144 33812 31184
rect 37420 31144 37460 31184
rect 38668 31144 38708 31184
rect 41740 31144 41780 31184
rect 42220 31144 42260 31184
rect 43756 31144 43796 31184
rect 43948 31144 43988 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 4012 30808 4052 30848
rect 4876 30808 4916 30848
rect 12940 30808 12980 30848
rect 25036 30808 25076 30848
rect 31084 30808 31124 30848
rect 31276 30808 31316 30848
rect 31564 30808 31604 30848
rect 38668 30808 38708 30848
rect 40972 30808 41012 30848
rect 44620 30808 44660 30848
rect 47212 30808 47252 30848
rect 8620 30724 8660 30764
rect 27724 30724 27764 30764
rect 42220 30724 42260 30764
rect 1324 30640 1364 30680
rect 1708 30640 1748 30680
rect 2572 30640 2612 30680
rect 4684 30640 4724 30680
rect 5548 30640 5588 30680
rect 6604 30640 6644 30680
rect 6892 30640 6932 30680
rect 6988 30640 7028 30680
rect 7372 30640 7412 30680
rect 7948 30640 7988 30680
rect 8428 30626 8468 30666
rect 9676 30640 9716 30680
rect 10924 30640 10964 30680
rect 11020 30640 11060 30680
rect 11116 30640 11156 30680
rect 11212 30640 11252 30680
rect 12076 30640 12116 30680
rect 12268 30640 12308 30680
rect 13132 30640 13172 30680
rect 13324 30640 13364 30680
rect 13516 30640 13556 30680
rect 13612 30640 13652 30680
rect 13804 30640 13844 30680
rect 13996 30640 14036 30680
rect 14956 30640 14996 30680
rect 15916 30640 15956 30680
rect 19660 30640 19700 30680
rect 19948 30640 19988 30680
rect 20332 30640 20372 30680
rect 21196 30640 21236 30680
rect 22636 30640 22676 30680
rect 23020 30640 23060 30680
rect 23884 30640 23924 30680
rect 25516 30640 25556 30680
rect 25612 30640 25652 30680
rect 25708 30640 25748 30680
rect 25804 30640 25844 30680
rect 25996 30640 26036 30680
rect 26956 30640 26996 30680
rect 27340 30640 27380 30680
rect 27628 30640 27668 30680
rect 28396 30640 28436 30680
rect 28492 30640 28532 30680
rect 28588 30640 28628 30680
rect 28684 30640 28724 30680
rect 29740 30640 29780 30680
rect 30604 30640 30644 30680
rect 30796 30640 30836 30680
rect 30892 30640 30932 30680
rect 30988 30640 31028 30680
rect 31372 30640 31412 30680
rect 31660 30640 31700 30680
rect 32428 30640 32468 30680
rect 34252 30640 34292 30680
rect 35116 30640 35156 30680
rect 35308 30640 35348 30680
rect 35404 30640 35444 30680
rect 35500 30640 35540 30680
rect 35596 30640 35636 30680
rect 36652 30640 36692 30680
rect 37036 30640 37076 30680
rect 37228 30640 37268 30680
rect 38092 30640 38132 30680
rect 38188 30640 38228 30680
rect 38380 30640 38420 30680
rect 38572 30640 38612 30680
rect 38764 30640 38804 30680
rect 38860 30640 38900 30680
rect 39052 30640 39092 30680
rect 39148 30640 39188 30680
rect 39244 30640 39284 30680
rect 39340 30640 39380 30680
rect 39532 30640 39572 30680
rect 40492 30640 40532 30680
rect 41644 30640 41684 30680
rect 41740 30640 41780 30680
rect 41836 30640 41876 30680
rect 41932 30640 41972 30680
rect 42604 30640 42644 30680
rect 43468 30640 43508 30680
rect 44812 30640 44852 30680
rect 45004 30640 45044 30680
rect 45100 30640 45140 30680
rect 46540 30640 46580 30680
rect 46828 30640 46868 30680
rect 47020 30640 47060 30680
rect 47116 30640 47156 30680
rect 47308 30640 47348 30680
rect 47692 30640 47732 30680
rect 47788 30640 47828 30680
rect 47884 30640 47924 30680
rect 47980 30640 48020 30680
rect 48268 30640 48308 30680
rect 48460 30640 48500 30680
rect 48556 30640 48596 30680
rect 48940 30640 48980 30680
rect 3724 30556 3764 30596
rect 7468 30556 7508 30596
rect 16300 30556 16340 30596
rect 31948 30556 31988 30596
rect 35980 30556 36020 30596
rect 9868 30472 9908 30512
rect 13804 30472 13844 30512
rect 17452 30472 17492 30512
rect 45292 30472 45332 30512
rect 48268 30472 48308 30512
rect 49996 30472 50036 30512
rect 50188 30472 50228 30512
rect 4012 30388 4052 30428
rect 5932 30388 5972 30428
rect 9004 30388 9044 30428
rect 11404 30388 11444 30428
rect 13228 30388 13268 30428
rect 14668 30388 14708 30428
rect 16108 30388 16148 30428
rect 18988 30388 19028 30428
rect 22348 30388 22388 30428
rect 28012 30388 28052 30428
rect 29068 30388 29108 30428
rect 29932 30388 29972 30428
rect 32716 30388 32756 30428
rect 33580 30388 33620 30428
rect 34444 30388 34484 30428
rect 37132 30388 37172 30428
rect 38380 30388 38420 30428
rect 40204 30388 40244 30428
rect 44812 30388 44852 30428
rect 46444 30388 46484 30428
rect 46732 30388 46772 30428
rect 49612 30388 49652 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 8044 30052 8084 30092
rect 11596 30052 11636 30092
rect 23308 30052 23348 30092
rect 24172 30052 24212 30092
rect 31276 30052 31316 30092
rect 35596 30052 35636 30092
rect 36268 30052 36308 30092
rect 1036 29968 1076 30008
rect 12844 29968 12884 30008
rect 13804 29968 13844 30008
rect 19468 29968 19508 30008
rect 22348 29968 22388 30008
rect 26956 29968 26996 30008
rect 38764 29968 38804 30008
rect 42316 29968 42356 30008
rect 46924 29968 46964 30008
rect 3628 29884 3668 29924
rect 5068 29884 5108 29924
rect 11308 29884 11348 29924
rect 17356 29884 17396 29924
rect 42124 29884 42164 29924
rect 1228 29800 1268 29840
rect 1612 29800 1652 29840
rect 2476 29800 2516 29840
rect 4108 29800 4148 29840
rect 4204 29800 4244 29840
rect 4300 29800 4340 29840
rect 4588 29800 4628 29840
rect 4684 29800 4724 29840
rect 5164 29800 5204 29840
rect 5644 29800 5684 29840
rect 6124 29814 6164 29854
rect 6508 29800 6548 29840
rect 7564 29800 7604 29840
rect 7660 29800 7700 29840
rect 7756 29800 7796 29840
rect 7852 29800 7892 29840
rect 8716 29800 8756 29840
rect 8908 29800 8948 29840
rect 9292 29800 9332 29840
rect 10156 29800 10196 29840
rect 11596 29800 11636 29840
rect 11788 29800 11828 29840
rect 11884 29800 11924 29840
rect 12172 29800 12212 29840
rect 12460 29800 12500 29840
rect 12556 29800 12596 29840
rect 13132 29800 13172 29840
rect 13420 29800 13460 29840
rect 13516 29800 13556 29840
rect 13996 29800 14036 29840
rect 14188 29800 14228 29840
rect 14476 29800 14516 29840
rect 14572 29800 14612 29840
rect 14668 29800 14708 29840
rect 14764 29800 14804 29840
rect 14956 29800 14996 29840
rect 15340 29800 15380 29840
rect 16204 29800 16244 29840
rect 18604 29800 18644 29840
rect 18700 29800 18740 29840
rect 18796 29800 18836 29840
rect 18892 29800 18932 29840
rect 19180 29800 19220 29840
rect 20140 29800 20180 29840
rect 20428 29800 20468 29840
rect 21964 29800 22004 29840
rect 23020 29800 23060 29840
rect 25324 29800 25364 29840
rect 26188 29800 26228 29840
rect 27340 29800 27380 29840
rect 27628 29800 27668 29840
rect 28588 29800 28628 29840
rect 28876 29800 28916 29840
rect 29260 29800 29300 29840
rect 30124 29800 30164 29840
rect 31468 29800 31508 29840
rect 31660 29800 31700 29840
rect 31756 29800 31796 29840
rect 31948 29800 31988 29840
rect 32908 29800 32948 29840
rect 33196 29800 33236 29840
rect 33580 29800 33620 29840
rect 34444 29800 34484 29840
rect 35980 29800 36020 29840
rect 36076 29800 36116 29840
rect 36268 29800 36308 29840
rect 37132 29800 37172 29840
rect 37420 29800 37460 29840
rect 37516 29800 37556 29840
rect 37612 29800 37652 29840
rect 38284 29800 38324 29840
rect 38380 29800 38420 29840
rect 38476 29800 38516 29840
rect 38572 29800 38612 29840
rect 39052 29800 39092 29840
rect 39148 29800 39188 29840
rect 39436 29800 39476 29840
rect 39724 29800 39764 29840
rect 40108 29800 40148 29840
rect 40972 29800 41012 29840
rect 42988 29800 43028 29840
rect 43180 29800 43220 29840
rect 43276 29800 43316 29840
rect 43372 29800 43412 29840
rect 43660 29800 43700 29840
rect 44908 29800 44948 29840
rect 45772 29800 45812 29840
rect 47788 29800 47828 29840
rect 48556 29800 48596 29840
rect 49420 29800 49460 29840
rect 14092 29716 14132 29756
rect 26572 29716 26612 29756
rect 27244 29716 27284 29756
rect 27916 29716 27956 29756
rect 44332 29716 44372 29756
rect 44524 29716 44564 29756
rect 48172 29716 48212 29756
rect 4012 29632 4052 29672
rect 6316 29632 6356 29672
rect 7180 29632 7220 29672
rect 21100 29632 21140 29672
rect 21292 29632 21332 29672
rect 23500 29632 23540 29672
rect 31564 29632 31604 29672
rect 36460 29632 36500 29672
rect 37708 29632 37748 29672
rect 43468 29632 43508 29672
rect 47116 29632 47156 29672
rect 50572 29632 50612 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 5548 29296 5588 29336
rect 6028 29296 6068 29336
rect 13324 29296 13364 29336
rect 20524 29296 20564 29336
rect 33196 29296 33236 29336
rect 33580 29296 33620 29336
rect 41260 29296 41300 29336
rect 42508 29296 42548 29336
rect 45100 29296 45140 29336
rect 47596 29296 47636 29336
rect 49228 29296 49268 29336
rect 2764 29170 2804 29210
rect 3244 29212 3284 29252
rect 5260 29212 5300 29252
rect 8428 29212 8468 29252
rect 10924 29212 10964 29252
rect 14380 29212 14420 29252
rect 22924 29212 22964 29252
rect 2956 29128 2996 29168
rect 3052 29128 3092 29168
rect 3340 29128 3380 29168
rect 3436 29128 3476 29168
rect 3532 29128 3572 29168
rect 3724 29128 3764 29168
rect 4684 29128 4724 29168
rect 5068 29128 5108 29168
rect 5164 29128 5204 29168
rect 5356 29128 5396 29168
rect 5644 29128 5684 29168
rect 5740 29128 5780 29168
rect 5836 29128 5876 29168
rect 7180 29128 7220 29168
rect 8044 29128 8084 29168
rect 8716 29128 8756 29168
rect 9100 29128 9140 29168
rect 9964 29128 10004 29168
rect 11308 29128 11348 29168
rect 12172 29128 12212 29168
rect 13996 29128 14036 29168
rect 14284 29128 14324 29168
rect 16108 29128 16148 29168
rect 17740 29128 17780 29168
rect 18604 29128 18644 29168
rect 18988 29128 19028 29168
rect 19180 29128 19220 29168
rect 19852 29128 19892 29168
rect 20044 29128 20084 29168
rect 20236 29128 20276 29168
rect 20332 29128 20372 29168
rect 21676 29128 21716 29168
rect 22540 29128 22580 29168
rect 26284 29128 26324 29168
rect 26380 29128 26420 29168
rect 26476 29128 26516 29168
rect 26572 29128 26612 29168
rect 26764 29128 26804 29168
rect 26956 29128 26996 29168
rect 27052 29128 27092 29168
rect 27244 29128 27284 29168
rect 27916 29170 27956 29210
rect 35980 29212 36020 29252
rect 51628 29212 51668 29252
rect 27436 29128 27476 29168
rect 27532 29128 27572 29168
rect 28108 29128 28148 29168
rect 28204 29128 28244 29168
rect 28396 29128 28436 29168
rect 28492 29128 28532 29168
rect 29068 29128 29108 29168
rect 29260 29128 29300 29168
rect 29356 29128 29396 29168
rect 29836 29128 29876 29168
rect 29932 29128 29972 29168
rect 30124 29128 30164 29168
rect 30220 29128 30260 29168
rect 30412 29128 30452 29168
rect 30604 29128 30644 29168
rect 30700 29128 30740 29168
rect 30796 29128 30836 29168
rect 30892 29128 30932 29168
rect 31084 29128 31124 29168
rect 31948 29128 31988 29168
rect 32620 29128 32660 29168
rect 33292 29128 33332 29168
rect 33484 29128 33524 29168
rect 33676 29128 33716 29168
rect 33772 29128 33812 29168
rect 33964 29128 34004 29168
rect 34828 29128 34868 29168
rect 36364 29128 36404 29168
rect 37228 29128 37268 29168
rect 39820 29128 39860 29168
rect 41644 29128 41684 29168
rect 41836 29128 41876 29168
rect 42892 29128 42932 29168
rect 43276 29128 43316 29168
rect 44140 29128 44180 29168
rect 44620 29128 44660 29168
rect 45868 29128 45908 29168
rect 47116 29128 47156 29168
rect 49036 29128 49076 29168
rect 50380 29128 50420 29168
rect 51244 29128 51284 29168
rect 8620 29044 8660 29084
rect 15436 29044 15476 29084
rect 31756 29044 31796 29084
rect 35788 29044 35828 29084
rect 38956 29044 38996 29084
rect 41452 29044 41492 29084
rect 41740 29044 41780 29084
rect 1804 28960 1844 29000
rect 2764 28960 2804 29000
rect 15244 28960 15284 29000
rect 16588 28960 16628 29000
rect 20044 28960 20084 29000
rect 25420 28960 25460 29000
rect 27244 28960 27284 29000
rect 27916 28960 27956 29000
rect 29068 28960 29108 29000
rect 33004 28960 33044 29000
rect 35404 28960 35444 29000
rect 35596 28960 35636 29000
rect 40876 28960 40916 29000
rect 9292 28876 9332 28916
rect 14668 28876 14708 28916
rect 20524 28876 20564 28916
rect 26764 28876 26804 28916
rect 30412 28876 30452 28916
rect 38380 28876 38420 28916
rect 45772 28876 45812 28916
rect 47788 28876 47828 28916
rect 48364 28876 48404 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 3724 28540 3764 28580
rect 20044 28540 20084 28580
rect 27532 28540 27572 28580
rect 31084 28540 31124 28580
rect 34252 28540 34292 28580
rect 39052 28540 39092 28580
rect 39340 28540 39380 28580
rect 47308 28540 47348 28580
rect 6412 28456 6452 28496
rect 8908 28456 8948 28496
rect 11404 28456 11444 28496
rect 16300 28456 16340 28496
rect 19276 28456 19316 28496
rect 22348 28456 22388 28496
rect 35308 28456 35348 28496
rect 36460 28456 36500 28496
rect 42220 28456 42260 28496
rect 47500 28456 47540 28496
rect 50860 28456 50900 28496
rect 51244 28456 51284 28496
rect 41068 28372 41108 28412
rect 45100 28372 45140 28412
rect 1708 28288 1748 28328
rect 2572 28288 2612 28328
rect 4012 28288 4052 28328
rect 4204 28288 4244 28328
rect 4300 28288 4340 28328
rect 5164 28288 5204 28328
rect 5356 28288 5396 28328
rect 6604 28288 6644 28328
rect 6700 28288 6740 28328
rect 6796 28288 6836 28328
rect 6892 28288 6932 28328
rect 7084 28288 7124 28328
rect 7276 28288 7316 28328
rect 7372 28288 7412 28328
rect 8236 28288 8276 28328
rect 8716 28288 8756 28328
rect 10156 28288 10196 28328
rect 11884 28288 11924 28328
rect 12076 28288 12116 28328
rect 12268 28288 12308 28328
rect 12460 28288 12500 28328
rect 12652 28288 12692 28328
rect 12748 28288 12788 28328
rect 12940 28288 12980 28328
rect 13132 28288 13172 28328
rect 13804 28288 13844 28328
rect 14092 28288 14132 28328
rect 17932 28288 17972 28328
rect 18700 28288 18740 28328
rect 18796 28288 18836 28328
rect 18892 28288 18932 28328
rect 18988 28288 19028 28328
rect 19372 28288 19412 28328
rect 19564 28288 19604 28328
rect 19660 28288 19700 28328
rect 19756 28288 19796 28328
rect 19852 28288 19892 28328
rect 20044 28288 20084 28328
rect 20236 28288 20276 28328
rect 20332 28288 20372 28328
rect 20524 28288 20564 28328
rect 20620 28288 20660 28328
rect 20716 28288 20756 28328
rect 21100 28288 21140 28328
rect 23404 28288 23444 28328
rect 24364 28288 24404 28328
rect 25324 28288 25364 28328
rect 25996 28288 26036 28328
rect 26476 28288 26516 28328
rect 26572 28288 26612 28328
rect 26668 28288 26708 28328
rect 27724 28288 27764 28328
rect 28492 28288 28532 28328
rect 28588 28288 28628 28328
rect 28780 28288 28820 28328
rect 28876 28288 28916 28328
rect 29068 28288 29108 28328
rect 30604 28288 30644 28328
rect 30700 28288 30740 28328
rect 30796 28288 30836 28328
rect 30892 28288 30932 28328
rect 32236 28288 32276 28328
rect 33100 28288 33140 28328
rect 33484 28288 33524 28328
rect 34348 28288 34388 28328
rect 35692 28288 35732 28328
rect 35980 28288 36020 28328
rect 37132 28288 37172 28328
rect 37228 28288 37268 28328
rect 37324 28288 37364 28328
rect 37420 28288 37460 28328
rect 38860 28288 38900 28328
rect 39148 28288 39188 28328
rect 39436 28288 39476 28328
rect 40012 28293 40052 28333
rect 40492 28288 40532 28328
rect 40972 28288 41012 28328
rect 41452 28288 41492 28328
rect 41548 28288 41588 28328
rect 41932 28288 41972 28328
rect 43180 28288 43220 28328
rect 43372 28288 43412 28328
rect 43468 28288 43508 28328
rect 43564 28288 43604 28328
rect 43660 28288 43700 28328
rect 44044 28302 44084 28342
rect 44524 28288 44564 28328
rect 45004 28288 45044 28328
rect 45484 28288 45524 28328
rect 45580 28288 45620 28328
rect 46444 28288 46484 28328
rect 46540 28288 46580 28328
rect 46828 28288 46868 28328
rect 47020 28288 47060 28328
rect 47116 28288 47156 28328
rect 47308 28288 47348 28328
rect 48172 28288 48212 28328
rect 48364 28288 48404 28328
rect 48460 28288 48500 28328
rect 48748 28288 48788 28328
rect 48844 28288 48884 28328
rect 48940 28288 48980 28328
rect 49132 28288 49172 28328
rect 50668 28288 50708 28328
rect 1324 28204 1364 28244
rect 4108 28204 4148 28244
rect 7180 28204 7220 28244
rect 11980 28204 12020 28244
rect 12364 28204 12404 28244
rect 17068 28204 17108 28244
rect 21004 28204 21044 28244
rect 28972 28204 29012 28244
rect 35596 28204 35636 28244
rect 49996 28204 50036 28244
rect 4492 28120 4532 28160
rect 6028 28120 6068 28160
rect 7564 28120 7604 28160
rect 10060 28120 10100 28160
rect 12844 28120 12884 28160
rect 14572 28120 14612 28160
rect 20812 28120 20852 28160
rect 22732 28120 22772 28160
rect 26092 28120 26132 28160
rect 26380 28120 26420 28160
rect 28300 28120 28340 28160
rect 38188 28120 38228 28160
rect 39820 28120 39860 28160
rect 43084 28120 43124 28160
rect 43852 28120 43892 28160
rect 46732 28120 46772 28160
rect 48652 28120 48692 28160
rect 49804 28120 49844 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 4684 27784 4724 27824
rect 12172 27784 12212 27824
rect 42892 27784 42932 27824
rect 2668 27700 2708 27740
rect 7468 27700 7508 27740
rect 19852 27700 19892 27740
rect 29740 27700 29780 27740
rect 36364 27700 36404 27740
rect 44428 27700 44468 27740
rect 51628 27700 51668 27740
rect 2764 27616 2804 27656
rect 3052 27616 3092 27656
rect 3340 27616 3380 27656
rect 3532 27616 3572 27656
rect 3628 27616 3668 27656
rect 3820 27616 3860 27656
rect 4204 27616 4244 27656
rect 5932 27616 5972 27656
rect 6988 27616 7028 27656
rect 7372 27616 7412 27656
rect 7660 27616 7700 27656
rect 7756 27616 7796 27656
rect 7852 27616 7892 27656
rect 7948 27616 7988 27656
rect 8140 27616 8180 27656
rect 8812 27616 8852 27656
rect 9004 27616 9044 27656
rect 9388 27616 9428 27656
rect 10252 27616 10292 27656
rect 11692 27616 11732 27656
rect 12652 27616 12692 27656
rect 13132 27616 13172 27656
rect 13324 27616 13364 27656
rect 13420 27616 13460 27656
rect 13612 27616 13652 27656
rect 13708 27616 13748 27656
rect 13900 27616 13940 27656
rect 13996 27587 14036 27627
rect 14151 27616 14191 27656
rect 14764 27616 14804 27656
rect 14860 27616 14900 27656
rect 15052 27616 15092 27656
rect 15148 27616 15188 27656
rect 15305 27601 15345 27641
rect 16012 27616 16052 27656
rect 16204 27616 16244 27656
rect 16300 27616 16340 27656
rect 17452 27616 17492 27656
rect 18412 27616 18452 27656
rect 19948 27616 19988 27656
rect 20236 27616 20276 27656
rect 20524 27616 20564 27656
rect 20716 27616 20756 27656
rect 20812 27616 20852 27656
rect 21004 27616 21044 27656
rect 21196 27616 21236 27656
rect 21292 27616 21332 27656
rect 21484 27616 21524 27656
rect 21580 27616 21620 27656
rect 21868 27616 21908 27656
rect 22252 27616 22292 27656
rect 23116 27616 23156 27656
rect 24652 27616 24692 27656
rect 24748 27581 24788 27621
rect 24844 27616 24884 27656
rect 26284 27616 26324 27656
rect 26764 27616 26804 27656
rect 27724 27616 27764 27656
rect 28012 27616 28052 27656
rect 28108 27616 28148 27656
rect 28492 27616 28532 27656
rect 29068 27616 29108 27656
rect 29548 27611 29588 27651
rect 30508 27616 30548 27656
rect 30700 27616 30740 27656
rect 30796 27616 30836 27656
rect 30988 27616 31028 27656
rect 31180 27616 31220 27656
rect 31276 27616 31316 27656
rect 31468 27616 31508 27656
rect 31564 27616 31604 27656
rect 31660 27616 31700 27656
rect 31756 27616 31796 27656
rect 31948 27616 31988 27656
rect 32151 27629 32191 27669
rect 33292 27616 33332 27656
rect 34156 27616 34196 27656
rect 34252 27616 34292 27656
rect 34348 27616 34388 27656
rect 34444 27616 34484 27656
rect 35212 27616 35252 27656
rect 36076 27616 36116 27656
rect 36268 27616 36308 27656
rect 36460 27616 36500 27656
rect 37804 27616 37844 27656
rect 38188 27616 38228 27656
rect 38284 27616 38324 27656
rect 38380 27616 38420 27656
rect 38476 27616 38516 27656
rect 38956 27616 38996 27656
rect 39916 27616 39956 27656
rect 40108 27616 40148 27656
rect 42988 27616 43028 27656
rect 43180 27597 43220 27637
rect 43276 27616 43316 27656
rect 43468 27616 43508 27656
rect 43660 27616 43700 27656
rect 43756 27616 43796 27656
rect 43852 27616 43892 27656
rect 43948 27616 43988 27656
rect 44332 27616 44372 27656
rect 44524 27616 44564 27656
rect 45100 27616 45140 27656
rect 45196 27616 45236 27656
rect 45292 27616 45332 27656
rect 45388 27616 45428 27656
rect 45964 27616 46004 27656
rect 46156 27616 46196 27656
rect 46252 27616 46292 27656
rect 46924 27616 46964 27656
rect 47212 27616 47252 27656
rect 47500 27616 47540 27656
rect 47596 27616 47636 27656
rect 47692 27616 47732 27656
rect 47788 27616 47828 27656
rect 48172 27616 48212 27656
rect 48268 27616 48308 27656
rect 48364 27616 48404 27656
rect 48460 27616 48500 27656
rect 48652 27616 48692 27656
rect 48748 27616 48788 27656
rect 48940 27616 48980 27656
rect 50380 27616 50420 27656
rect 51244 27616 51284 27656
rect 5644 27532 5684 27572
rect 19180 27532 19220 27572
rect 24268 27532 24308 27572
rect 25516 27532 25556 27572
rect 28588 27532 28628 27572
rect 49228 27532 49268 27572
rect 1708 27448 1748 27488
rect 3244 27448 3284 27488
rect 19564 27448 19604 27488
rect 21004 27448 21044 27488
rect 26092 27448 26132 27488
rect 32044 27448 32084 27488
rect 33100 27448 33140 27488
rect 36940 27448 36980 27488
rect 42220 27448 42260 27488
rect 46444 27448 46484 27488
rect 2956 27364 2996 27404
rect 3820 27364 3860 27404
rect 5452 27364 5492 27404
rect 5836 27364 5876 27404
rect 6796 27364 6836 27404
rect 11404 27364 11444 27404
rect 13132 27364 13172 27404
rect 13612 27364 13652 27404
rect 14764 27364 14804 27404
rect 16012 27364 16052 27404
rect 19372 27364 19412 27404
rect 20524 27364 20564 27404
rect 25132 27364 25172 27404
rect 30508 27364 30548 27404
rect 30988 27364 31028 27404
rect 33964 27364 34004 27404
rect 37708 27364 37748 27404
rect 39628 27364 39668 27404
rect 43468 27364 43508 27404
rect 45964 27364 46004 27404
rect 47020 27364 47060 27404
rect 47308 27364 47348 27404
rect 48940 27364 48980 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 3628 27028 3668 27068
rect 4684 27028 4724 27068
rect 7852 27028 7892 27068
rect 9196 27028 9236 27068
rect 11980 27028 12020 27068
rect 13516 27028 13556 27068
rect 14380 27028 14420 27068
rect 15052 27028 15092 27068
rect 21292 27028 21332 27068
rect 27916 27028 27956 27068
rect 31372 27028 31412 27068
rect 31852 27028 31892 27068
rect 32812 27028 32852 27068
rect 38764 27028 38804 27068
rect 39628 27028 39668 27068
rect 47980 27028 48020 27068
rect 48172 27028 48212 27068
rect 49324 27028 49364 27068
rect 10060 26944 10100 26984
rect 18028 26944 18068 26984
rect 19276 26944 19316 26984
rect 22348 26944 22388 26984
rect 24940 26944 24980 26984
rect 26188 26944 26228 26984
rect 44140 26860 44180 26900
rect 1228 26776 1268 26816
rect 1612 26776 1652 26816
rect 2476 26776 2516 26816
rect 4492 26776 4532 26816
rect 5836 26776 5876 26816
rect 6700 26776 6740 26816
rect 7084 26776 7124 26816
rect 8428 26776 8468 26816
rect 9868 26776 9908 26816
rect 10540 26776 10580 26816
rect 10732 26776 10772 26816
rect 10828 26776 10868 26816
rect 11020 26776 11060 26816
rect 11308 26776 11348 26816
rect 11596 26776 11636 26816
rect 12172 26776 12212 26816
rect 12268 26776 12308 26816
rect 12364 26776 12404 26816
rect 12460 26776 12500 26816
rect 13708 26776 13748 26816
rect 14092 26776 14132 26816
rect 14188 26776 14228 26816
rect 14380 26776 14420 26816
rect 14572 26776 14612 26816
rect 14668 26776 14708 26816
rect 14860 26776 14900 26816
rect 15052 26776 15092 26816
rect 15244 26776 15284 26816
rect 15340 26776 15380 26816
rect 16780 26776 16820 26816
rect 16972 26776 17012 26816
rect 17164 26776 17204 26816
rect 17356 26776 17396 26816
rect 17548 26776 17588 26816
rect 17644 26776 17684 26816
rect 17740 26776 17780 26816
rect 18700 26776 18740 26816
rect 19660 26776 19700 26816
rect 19948 26776 19988 26816
rect 20428 26776 20468 26816
rect 21964 26776 22004 26816
rect 24268 26776 24308 26816
rect 24460 26776 24500 26816
rect 24748 26776 24788 26816
rect 27340 26776 27380 26816
rect 28780 26776 28820 26816
rect 28972 26776 29012 26816
rect 29068 26776 29108 26816
rect 29452 26776 29492 26816
rect 29548 26776 29588 26816
rect 29644 26776 29684 26816
rect 30316 26776 30356 26816
rect 30412 26811 30452 26851
rect 30508 26776 30548 26816
rect 30892 26776 30932 26816
rect 31084 26776 31124 26816
rect 31180 26776 31220 26816
rect 31372 26776 31412 26816
rect 31564 26776 31604 26816
rect 31660 26776 31700 26816
rect 32140 26776 32180 26816
rect 32236 26776 32276 26816
rect 32524 26776 32564 26816
rect 33964 26776 34004 26816
rect 34828 26776 34868 26816
rect 35500 26776 35540 26816
rect 35596 26776 35636 26816
rect 35692 26776 35732 26816
rect 35884 26776 35924 26816
rect 36076 26776 36116 26816
rect 36172 26776 36212 26816
rect 36748 26776 36788 26816
rect 37612 26776 37652 26816
rect 38956 26776 38996 26816
rect 40300 26776 40340 26816
rect 41740 26776 41780 26816
rect 42124 26776 42164 26816
rect 42988 26776 43028 26816
rect 45004 26776 45044 26816
rect 45580 26776 45620 26816
rect 45964 26776 46004 26816
rect 46828 26776 46868 26816
rect 48844 26776 48884 26816
rect 49036 26776 49076 26816
rect 49132 26776 49172 26816
rect 49324 26776 49364 26816
rect 49612 26776 49652 26816
rect 49996 26776 50036 26816
rect 50860 26776 50900 26816
rect 11692 26692 11732 26732
rect 16876 26692 16916 26732
rect 17260 26692 17300 26732
rect 19564 26692 19604 26732
rect 24364 26692 24404 26732
rect 35212 26692 35252 26732
rect 36364 26692 36404 26732
rect 3820 26608 3860 26648
rect 8044 26608 8084 26648
rect 10444 26608 10484 26648
rect 10924 26608 10964 26648
rect 14764 26608 14804 26648
rect 17836 26608 17876 26648
rect 21100 26608 21140 26648
rect 28876 26608 28916 26648
rect 30028 26608 30068 26648
rect 30988 26608 31028 26648
rect 35404 26608 35444 26648
rect 35980 26608 36020 26648
rect 40684 26608 40724 26648
rect 44332 26608 44372 26648
rect 52012 26608 52052 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3628 26272 3668 26312
rect 3820 26272 3860 26312
rect 9196 26272 9236 26312
rect 20620 26272 20660 26312
rect 29644 26272 29684 26312
rect 31756 26272 31796 26312
rect 43564 26272 43604 26312
rect 45676 26272 45716 26312
rect 49804 26272 49844 26312
rect 1228 26188 1268 26228
rect 4396 26188 4436 26228
rect 7852 26188 7892 26228
rect 15148 26188 15188 26228
rect 17164 26188 17204 26228
rect 39148 26188 39188 26228
rect 44236 26188 44276 26228
rect 1612 26104 1652 26144
rect 2476 26104 2516 26144
rect 4012 26125 4052 26165
rect 4108 26104 4148 26144
rect 3916 26062 3956 26102
rect 4300 26104 4340 26144
rect 4492 26104 4532 26144
rect 4588 26104 4628 26144
rect 4972 26104 5012 26144
rect 5068 26104 5108 26144
rect 5260 26104 5300 26144
rect 6988 26104 7028 26144
rect 7468 26104 7508 26144
rect 7756 26104 7796 26144
rect 9100 26104 9140 26144
rect 9292 26104 9332 26144
rect 9388 26104 9428 26144
rect 10732 26104 10772 26144
rect 10924 26104 10964 26144
rect 11116 26104 11156 26144
rect 11308 26104 11348 26144
rect 12268 26104 12308 26144
rect 12556 26104 12596 26144
rect 12652 26104 12692 26144
rect 12844 26104 12884 26144
rect 13132 26104 13172 26144
rect 13358 26097 13398 26137
rect 13516 26104 13556 26144
rect 13612 26104 13652 26144
rect 13804 26104 13844 26144
rect 13900 26104 13940 26144
rect 14284 26104 14324 26144
rect 14380 26104 14420 26144
rect 14572 26104 14612 26144
rect 14668 26104 14708 26144
rect 14769 26104 14809 26144
rect 15052 26104 15092 26144
rect 15244 26104 15284 26144
rect 15436 26104 15476 26144
rect 15628 26104 15668 26144
rect 15916 26104 15956 26144
rect 16012 26104 16052 26144
rect 16108 26104 16148 26144
rect 16204 26104 16244 26144
rect 16396 26104 16436 26144
rect 16588 26104 16628 26144
rect 16684 26104 16724 26144
rect 17260 26104 17300 26144
rect 17548 26104 17588 26144
rect 18124 26104 18164 26144
rect 18220 26104 18260 26144
rect 18412 26104 18452 26144
rect 18700 26104 18740 26144
rect 18796 26104 18836 26144
rect 18892 26104 18932 26144
rect 18988 26104 19028 26144
rect 19180 26104 19220 26144
rect 19276 26104 19316 26144
rect 19468 26104 19508 26144
rect 9676 26020 9716 26060
rect 19372 26062 19412 26102
rect 19660 26104 19700 26144
rect 20524 26104 20564 26144
rect 20908 26104 20948 26144
rect 22060 26104 22100 26144
rect 22924 26104 22964 26144
rect 23308 26104 23348 26144
rect 23692 26104 23732 26144
rect 23788 26104 23828 26144
rect 23884 26104 23924 26144
rect 23980 26104 24020 26144
rect 25132 26104 25172 26144
rect 25804 26104 25844 26144
rect 25900 26099 25940 26139
rect 25996 26104 26036 26144
rect 26956 26104 26996 26144
rect 27532 26104 27572 26144
rect 27628 26099 27668 26139
rect 27724 26104 27764 26144
rect 28396 26104 28436 26144
rect 29356 26104 29396 26144
rect 29548 26104 29588 26144
rect 29740 26104 29780 26144
rect 29836 26104 29876 26144
rect 30892 26104 30932 26144
rect 30988 26069 31028 26109
rect 31084 26104 31124 26144
rect 32140 26104 32180 26144
rect 33676 26104 33716 26144
rect 33868 26119 33908 26159
rect 33964 26104 34004 26144
rect 34156 26104 34196 26144
rect 35980 26104 36020 26144
rect 39340 26099 39380 26139
rect 39820 26104 39860 26144
rect 40300 26104 40340 26144
rect 40396 26104 40436 26144
rect 40780 26104 40820 26144
rect 40876 26104 40916 26144
rect 42220 26104 42260 26144
rect 42316 26104 42356 26144
rect 42412 26104 42452 26144
rect 42508 26104 42548 26144
rect 42796 26104 42836 26144
rect 42892 26104 42932 26144
rect 43084 26104 43124 26144
rect 43180 26104 43220 26144
rect 43372 26104 43412 26144
rect 43660 26104 43700 26144
rect 43756 26104 43796 26144
rect 43852 26104 43892 26144
rect 44332 26104 44372 26144
rect 44428 26104 44468 26144
rect 44524 26104 44564 26144
rect 44716 26104 44756 26144
rect 44908 26104 44948 26144
rect 46060 26104 46100 26144
rect 46156 26104 46196 26144
rect 46348 26104 46388 26144
rect 47212 26104 47252 26144
rect 47404 26104 47444 26144
rect 47500 26104 47540 26144
rect 47596 26104 47636 26144
rect 47692 26104 47732 26144
rect 47884 26104 47924 26144
rect 48076 26104 48116 26144
rect 48172 26104 48212 26144
rect 48940 26104 48980 26144
rect 49900 26104 49940 26144
rect 50764 26104 50804 26144
rect 50956 26104 50996 26144
rect 51628 26104 51668 26144
rect 11020 26020 11060 26060
rect 24268 26020 24308 26060
rect 45868 26020 45908 26060
rect 1036 25936 1076 25976
rect 5260 25936 5300 25976
rect 5644 25936 5684 25976
rect 6412 25936 6452 25976
rect 8908 25936 8948 25976
rect 12844 25936 12884 25976
rect 16876 25936 16916 25976
rect 18412 25936 18452 25976
rect 29068 25936 29108 25976
rect 34156 25936 34196 25976
rect 36844 25936 36884 25976
rect 44812 25936 44852 25976
rect 45292 25936 45332 25976
rect 48748 25936 48788 25976
rect 8140 25852 8180 25892
rect 10060 25852 10100 25892
rect 13036 25852 13076 25892
rect 13900 25852 13940 25892
rect 14284 25852 14324 25892
rect 15436 25852 15476 25892
rect 16396 25852 16436 25892
rect 20332 25852 20372 25892
rect 25516 25852 25556 25892
rect 26284 25852 26324 25892
rect 27244 25852 27284 25892
rect 30604 25852 30644 25892
rect 33580 25852 33620 25892
rect 36652 25852 36692 25892
rect 43372 25852 43412 25892
rect 46348 25852 46388 25892
rect 46540 25852 46580 25892
rect 47884 25852 47924 25892
rect 49612 25852 49652 25892
rect 50092 25852 50132 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 11500 25516 11540 25556
rect 13132 25516 13172 25556
rect 15052 25516 15092 25556
rect 17452 25516 17492 25556
rect 17932 25516 17972 25556
rect 19372 25516 19412 25556
rect 24556 25516 24596 25556
rect 31660 25516 31700 25556
rect 39628 25516 39668 25556
rect 41260 25516 41300 25556
rect 42412 25516 42452 25556
rect 47212 25516 47252 25556
rect 51148 25516 51188 25556
rect 1612 25432 1652 25472
rect 6700 25432 6740 25472
rect 27532 25432 27572 25472
rect 28204 25432 28244 25472
rect 29836 25432 29876 25472
rect 32524 25432 32564 25472
rect 33004 25432 33044 25472
rect 44332 25432 44372 25472
rect 22732 25348 22772 25388
rect 38476 25348 38516 25388
rect 3436 25264 3476 25304
rect 3532 25264 3572 25304
rect 3628 25264 3668 25304
rect 3820 25264 3860 25304
rect 3916 25264 3956 25304
rect 4012 25264 4052 25304
rect 4108 25264 4148 25304
rect 4300 25264 4340 25304
rect 4972 25264 5012 25304
rect 5836 25264 5876 25304
rect 6988 25264 7028 25304
rect 7852 25264 7892 25304
rect 8716 25264 8756 25304
rect 9100 25264 9140 25304
rect 9484 25264 9524 25304
rect 10348 25264 10388 25304
rect 11692 25264 11732 25304
rect 12940 25264 12980 25304
rect 13804 25264 13844 25304
rect 13996 25264 14036 25304
rect 14092 25264 14132 25304
rect 14188 25264 14228 25304
rect 14284 25264 14324 25304
rect 14668 25264 14708 25304
rect 14764 25264 14804 25304
rect 15244 25264 15284 25304
rect 16108 25264 16148 25304
rect 17164 25264 17204 25304
rect 17260 25264 17300 25304
rect 17452 25264 17492 25304
rect 17644 25264 17684 25304
rect 17740 25264 17780 25304
rect 17932 25264 17972 25304
rect 19180 25264 19220 25304
rect 20524 25264 20564 25304
rect 21388 25264 21428 25304
rect 21772 25264 21812 25304
rect 23596 25264 23636 25304
rect 24844 25264 24884 25304
rect 25132 25264 25172 25304
rect 25516 25264 25556 25304
rect 26380 25264 26420 25304
rect 27916 25264 27956 25304
rect 31180 25264 31220 25304
rect 32716 25264 32756 25304
rect 32812 25264 32852 25304
rect 33004 25264 33044 25304
rect 33868 25264 33908 25304
rect 34060 25264 34100 25304
rect 34156 25264 34196 25304
rect 34252 25264 34292 25304
rect 34348 25264 34388 25304
rect 34732 25264 34772 25304
rect 34828 25264 34868 25304
rect 34924 25264 34964 25304
rect 35212 25264 35252 25304
rect 36076 25264 36116 25304
rect 36460 25264 36500 25304
rect 37324 25264 37364 25304
rect 38943 25253 38983 25293
rect 39052 25264 39092 25304
rect 39340 25264 39380 25304
rect 40300 25264 40340 25304
rect 40492 25264 40532 25304
rect 40588 25264 40628 25304
rect 41644 25264 41684 25304
rect 41932 25264 41972 25304
rect 42316 25264 42356 25304
rect 42508 25264 42548 25304
rect 43372 25264 43412 25304
rect 43756 25264 43796 25304
rect 43852 25264 43892 25304
rect 43948 25264 43988 25304
rect 44044 25264 44084 25304
rect 44332 25264 44372 25304
rect 44524 25264 44564 25304
rect 44620 25264 44660 25304
rect 44812 25264 44852 25304
rect 45196 25264 45236 25304
rect 46060 25264 46100 25304
rect 47404 25264 47444 25304
rect 47500 25264 47540 25304
rect 47596 25264 47636 25304
rect 47884 25264 47924 25304
rect 49132 25264 49172 25304
rect 49996 25264 50036 25304
rect 12364 25180 12404 25220
rect 35020 25180 35060 25220
rect 41548 25180 41588 25220
rect 47692 25180 47732 25220
rect 48556 25180 48596 25220
rect 48748 25180 48788 25220
rect 3340 25096 3380 25136
rect 5164 25096 5204 25136
rect 14572 25092 14612 25132
rect 19084 25096 19124 25136
rect 33196 25096 33236 25136
rect 35884 25096 35924 25136
rect 40780 25096 40820 25136
rect 42700 25096 42740 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 28108 24818 28148 24858
rect 13324 24760 13364 24800
rect 16204 24760 16244 24800
rect 16876 24760 16916 24800
rect 19084 24760 19124 24800
rect 21580 24760 21620 24800
rect 25804 24760 25844 24800
rect 28396 24760 28436 24800
rect 31756 24760 31796 24800
rect 35212 24760 35252 24800
rect 35692 24760 35732 24800
rect 39820 24760 39860 24800
rect 44140 24760 44180 24800
rect 44620 24760 44660 24800
rect 45484 24760 45524 24800
rect 46348 24760 46388 24800
rect 46540 24760 46580 24800
rect 5068 24676 5108 24716
rect 10348 24676 10388 24716
rect 10828 24676 10868 24716
rect 12652 24676 12692 24716
rect 32812 24676 32852 24716
rect 38476 24676 38516 24716
rect 48940 24676 48980 24716
rect 1132 24592 1172 24632
rect 1516 24592 1556 24632
rect 2380 24592 2420 24632
rect 4204 24592 4244 24632
rect 4492 24592 4532 24632
rect 4588 24592 4628 24632
rect 5452 24592 5492 24632
rect 6316 24592 6356 24632
rect 7756 24592 7796 24632
rect 8044 24592 8084 24632
rect 8140 24592 8180 24632
rect 9292 24592 9332 24632
rect 10252 24592 10292 24632
rect 10444 24592 10484 24632
rect 10636 24592 10676 24632
rect 10732 24592 10772 24632
rect 10924 24592 10964 24632
rect 11788 24592 11828 24632
rect 12268 24592 12308 24632
rect 12556 24592 12596 24632
rect 13132 24592 13172 24632
rect 13228 24592 13268 24632
rect 13420 24592 13460 24632
rect 13612 24592 13652 24632
rect 13708 24592 13748 24632
rect 13900 24592 13940 24632
rect 14092 24592 14132 24632
rect 14188 24592 14228 24632
rect 14284 24592 14324 24632
rect 14380 24613 14420 24653
rect 14764 24592 14804 24632
rect 14860 24592 14900 24632
rect 14956 24592 14996 24632
rect 15052 24592 15092 24632
rect 15244 24592 15284 24632
rect 15532 24592 15572 24632
rect 15724 24592 15764 24632
rect 15820 24592 15860 24632
rect 15916 24592 15956 24632
rect 16012 24592 16052 24632
rect 16300 24592 16340 24632
rect 16396 24592 16436 24632
rect 16492 24592 16532 24632
rect 16684 24592 16724 24632
rect 16780 24592 16820 24632
rect 16972 24592 17012 24632
rect 17452 24592 17492 24632
rect 17548 24592 17588 24632
rect 17836 24592 17876 24632
rect 18604 24592 18644 24632
rect 18796 24592 18836 24632
rect 18892 24592 18932 24632
rect 19756 24592 19796 24632
rect 19948 24592 19988 24632
rect 22252 24592 22292 24632
rect 22444 24592 22484 24632
rect 23308 24592 23348 24632
rect 25708 24592 25748 24632
rect 25900 24592 25940 24632
rect 27916 24592 27956 24632
rect 28012 24592 28052 24632
rect 28300 24592 28340 24632
rect 28492 24592 28532 24632
rect 28588 24592 28628 24632
rect 29356 24592 29396 24632
rect 29740 24592 29780 24632
rect 30604 24592 30644 24632
rect 33196 24592 33236 24632
rect 34060 24592 34100 24632
rect 35596 24592 35636 24632
rect 35788 24592 35828 24632
rect 35884 24592 35924 24632
rect 36076 24592 36116 24632
rect 36748 24592 36788 24632
rect 36844 24592 36884 24632
rect 37804 24592 37844 24632
rect 38284 24587 38324 24627
rect 40012 24587 40052 24627
rect 40492 24592 40532 24632
rect 41452 24592 41492 24632
rect 41548 24592 41588 24632
rect 43372 24592 43412 24632
rect 43852 24592 43892 24632
rect 43948 24592 43988 24632
rect 44044 24592 44084 24632
rect 44332 24592 44372 24632
rect 44428 24592 44468 24632
rect 44524 24592 44564 24632
rect 44812 24592 44852 24632
rect 45676 24592 45716 24632
rect 47212 24592 47252 24632
rect 47404 24592 47444 24632
rect 47500 24592 47540 24632
rect 47596 24592 47636 24632
rect 47692 24592 47732 24632
rect 47980 24592 48020 24632
rect 48172 24592 48212 24632
rect 48268 24592 48308 24632
rect 48460 24592 48500 24632
rect 48652 24592 48692 24632
rect 48748 24592 48788 24632
rect 49036 24592 49076 24632
rect 49420 24592 49460 24632
rect 49804 24592 49844 24632
rect 50668 24592 50708 24632
rect 51820 24592 51860 24632
rect 3532 24508 3572 24548
rect 36172 24508 36212 24548
rect 37228 24508 37268 24548
rect 37324 24508 37364 24548
rect 40972 24508 41012 24548
rect 41068 24508 41108 24548
rect 8428 24424 8468 24464
rect 10060 24424 10100 24464
rect 15532 24424 15572 24464
rect 17164 24424 17204 24464
rect 18604 24424 18644 24464
rect 20812 24424 20852 24464
rect 21388 24424 21428 24464
rect 27628 24424 27668 24464
rect 38860 24424 38900 24464
rect 42316 24424 42356 24464
rect 48460 24424 48500 24464
rect 4876 24340 4916 24380
rect 7468 24340 7508 24380
rect 8620 24340 8660 24380
rect 11116 24340 11156 24380
rect 12940 24340 12980 24380
rect 13900 24340 13940 24380
rect 20620 24340 20660 24380
rect 22732 24340 22772 24380
rect 42988 24340 43028 24380
rect 45484 24340 45524 24380
rect 46348 24340 46388 24380
rect 46540 24340 46580 24380
rect 47980 24340 48020 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 12460 24004 12500 24044
rect 19564 24004 19604 24044
rect 22444 24004 22484 24044
rect 29452 24004 29492 24044
rect 37132 24004 37172 24044
rect 45100 24004 45140 24044
rect 47596 24004 47636 24044
rect 1708 23920 1748 23960
rect 3532 23920 3572 23960
rect 4972 23920 5012 23960
rect 6316 23920 6356 23960
rect 13612 23920 13652 23960
rect 16396 23920 16436 23960
rect 17932 23920 17972 23960
rect 23404 23920 23444 23960
rect 32428 23920 32468 23960
rect 44332 23920 44372 23960
rect 45868 23920 45908 23960
rect 49516 23920 49556 23960
rect 49900 23920 49940 23960
rect 27724 23836 27764 23876
rect 34348 23836 34388 23876
rect 34636 23836 34676 23876
rect 2284 23752 2324 23792
rect 2380 23752 2420 23792
rect 2572 23752 2612 23792
rect 2668 23752 2708 23792
rect 2860 23752 2900 23792
rect 3052 23752 3092 23792
rect 3244 23752 3284 23792
rect 3340 23752 3380 23792
rect 4204 23752 4244 23792
rect 4492 23752 4532 23792
rect 4588 23752 4628 23792
rect 4684 23752 4724 23792
rect 4876 23752 4916 23792
rect 5164 23752 5204 23792
rect 5260 23752 5300 23792
rect 5356 23752 5396 23792
rect 5452 23752 5492 23792
rect 5644 23752 5684 23792
rect 5740 23752 5780 23792
rect 5836 23752 5876 23792
rect 6508 23752 6548 23792
rect 7756 23752 7796 23792
rect 8620 23752 8660 23792
rect 10060 23752 10100 23792
rect 10444 23752 10484 23792
rect 11308 23752 11348 23792
rect 12652 23752 12692 23792
rect 12940 23752 12980 23792
rect 14476 23752 14516 23792
rect 14668 23752 14708 23792
rect 14860 23752 14900 23792
rect 15148 23752 15188 23792
rect 15244 23752 15284 23792
rect 15340 23752 15380 23792
rect 15628 23752 15668 23792
rect 15724 23752 15764 23792
rect 16108 23752 16148 23792
rect 16204 23752 16244 23792
rect 16396 23752 16436 23792
rect 16588 23752 16628 23792
rect 16684 23752 16724 23792
rect 16780 23752 16820 23792
rect 17068 23752 17108 23792
rect 19084 23752 19124 23792
rect 19180 23752 19220 23792
rect 19276 23752 19316 23792
rect 19372 23752 19412 23792
rect 19564 23752 19604 23792
rect 19756 23752 19796 23792
rect 19852 23752 19892 23792
rect 20044 23752 20084 23792
rect 20428 23752 20468 23792
rect 21292 23752 21332 23792
rect 22636 23752 22676 23792
rect 22732 23752 22772 23792
rect 22924 23752 22964 23792
rect 23404 23752 23444 23792
rect 23500 23752 23540 23792
rect 23692 23752 23732 23792
rect 23884 23752 23924 23792
rect 24652 23752 24692 23792
rect 24844 23752 24884 23792
rect 25036 23752 25076 23792
rect 25228 23752 25268 23792
rect 25324 23752 25364 23792
rect 25708 23752 25748 23792
rect 25804 23752 25844 23792
rect 25996 23752 26036 23792
rect 26092 23752 26132 23792
rect 26284 23752 26324 23792
rect 26476 23752 26516 23792
rect 26668 23752 26708 23792
rect 27148 23752 27188 23792
rect 27244 23752 27284 23792
rect 27436 23752 27476 23792
rect 27628 23752 27668 23792
rect 27820 23752 27860 23792
rect 28108 23752 28148 23792
rect 28492 23752 28532 23792
rect 28588 23752 28628 23792
rect 28684 23752 28724 23792
rect 28780 23752 28820 23792
rect 29068 23752 29108 23792
rect 29164 23752 29204 23792
rect 29260 23752 29300 23792
rect 29452 23752 29492 23792
rect 29644 23752 29684 23792
rect 29740 23752 29780 23792
rect 30796 23752 30836 23792
rect 31084 23752 31124 23792
rect 31180 23752 31220 23792
rect 31276 23752 31316 23792
rect 33100 23752 33140 23792
rect 33484 23752 33524 23792
rect 35692 23752 35732 23792
rect 36748 23752 36788 23792
rect 37228 23752 37268 23792
rect 37420 23752 37460 23792
rect 37516 23752 37556 23792
rect 37708 23752 37748 23792
rect 37900 23752 37940 23792
rect 37996 23752 38036 23792
rect 38092 23752 38132 23792
rect 38188 23752 38228 23792
rect 38764 23752 38804 23792
rect 39628 23752 39668 23792
rect 41740 23752 41780 23792
rect 41932 23752 41972 23792
rect 42316 23752 42356 23792
rect 43180 23752 43220 23792
rect 44620 23752 44660 23792
rect 45772 23752 45812 23792
rect 46156 23752 46196 23792
rect 46924 23752 46964 23792
rect 48268 23752 48308 23792
rect 48460 23752 48500 23792
rect 2764 23668 2804 23708
rect 5932 23668 5972 23708
rect 7180 23668 7220 23708
rect 7372 23668 7412 23708
rect 14764 23668 14804 23708
rect 15052 23668 15092 23708
rect 23308 23668 23348 23708
rect 23788 23668 23828 23708
rect 26572 23668 26612 23708
rect 35980 23668 36020 23708
rect 38380 23668 38420 23708
rect 3148 23584 3188 23624
rect 4396 23584 4436 23624
rect 9772 23584 9812 23624
rect 12748 23584 12788 23624
rect 13804 23584 13844 23624
rect 15916 23584 15956 23624
rect 16876 23584 16916 23624
rect 17740 23584 17780 23624
rect 22924 23584 22964 23624
rect 23116 23584 23156 23624
rect 23212 23584 23252 23624
rect 24748 23584 24788 23624
rect 25036 23584 25076 23624
rect 25516 23584 25556 23624
rect 26284 23584 26324 23624
rect 27340 23584 27380 23624
rect 28012 23584 28052 23624
rect 28300 23584 28340 23624
rect 28972 23584 29012 23624
rect 30892 23584 30932 23624
rect 31372 23584 31412 23624
rect 34828 23584 34868 23624
rect 35020 23584 35060 23624
rect 37132 23584 37172 23624
rect 37612 23584 37652 23624
rect 40780 23584 40820 23624
rect 41068 23584 41108 23624
rect 47596 23584 47636 23624
rect 49132 23584 49172 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3628 23248 3668 23288
rect 6028 23248 6068 23288
rect 7180 23248 7220 23288
rect 11116 23248 11156 23288
rect 12076 23248 12116 23288
rect 16012 23248 16052 23288
rect 19756 23248 19796 23288
rect 25900 23248 25940 23288
rect 28780 23248 28820 23288
rect 29068 23248 29108 23288
rect 30892 23248 30932 23288
rect 36556 23248 36596 23288
rect 37132 23248 37172 23288
rect 38380 23248 38420 23288
rect 43084 23248 43124 23288
rect 1228 23164 1268 23204
rect 7468 23164 7508 23204
rect 13612 23164 13652 23204
rect 17356 23164 17396 23204
rect 26284 23164 26324 23204
rect 29548 23164 29588 23204
rect 35788 23164 35828 23204
rect 47404 23164 47444 23204
rect 1612 23080 1652 23120
rect 2476 23080 2516 23120
rect 3916 23080 3956 23120
rect 4108 23080 4148 23120
rect 4204 23080 4244 23120
rect 4492 23080 4532 23120
rect 4780 23080 4820 23120
rect 4876 23080 4916 23120
rect 5452 23080 5492 23120
rect 5548 23080 5588 23120
rect 5740 23080 5780 23120
rect 6124 23080 6164 23120
rect 6700 23080 6740 23120
rect 6796 23080 6836 23120
rect 6988 23080 7028 23120
rect 7084 23080 7124 23120
rect 7276 23080 7316 23120
rect 8140 23080 8180 23120
rect 8332 23080 8372 23120
rect 8428 23080 8468 23120
rect 8524 23080 8564 23120
rect 8620 23080 8660 23120
rect 9196 23080 9236 23120
rect 9292 23080 9332 23120
rect 9388 23080 9428 23120
rect 9484 23080 9524 23120
rect 9676 23080 9716 23120
rect 9868 23080 9908 23120
rect 9964 23080 10004 23120
rect 11212 23080 11252 23120
rect 11404 23080 11444 23120
rect 12268 23080 12308 23120
rect 12364 23080 12404 23120
rect 12556 23080 12596 23120
rect 12748 23080 12788 23120
rect 13996 23080 14036 23120
rect 14860 23080 14900 23120
rect 16300 23080 16340 23120
rect 17740 23080 17780 23120
rect 18604 23080 18644 23120
rect 20620 23080 20660 23120
rect 23116 23080 23156 23120
rect 23404 23087 23444 23127
rect 23692 23080 23732 23120
rect 23788 23080 23828 23120
rect 23884 23080 23924 23120
rect 23980 23080 24020 23120
rect 24364 23080 24404 23120
rect 24460 23080 24500 23120
rect 25036 23080 25076 23120
rect 25420 23080 25460 23120
rect 25612 23080 25652 23120
rect 25708 23080 25748 23120
rect 25804 23080 25844 23120
rect 26092 23080 26132 23120
rect 26188 23080 26228 23120
rect 26380 23080 26420 23120
rect 26572 23080 26612 23120
rect 26668 23080 26708 23120
rect 26764 23080 26804 23120
rect 26860 23080 26900 23120
rect 27052 23080 27092 23120
rect 27244 23080 27284 23120
rect 27340 23080 27380 23120
rect 27724 23080 27764 23120
rect 27820 23080 27860 23120
rect 28300 23080 28340 23120
rect 28492 23080 28532 23120
rect 28588 23080 28628 23120
rect 28972 23080 29012 23120
rect 29164 23080 29204 23120
rect 29452 23080 29492 23120
rect 29644 23080 29684 23120
rect 30412 23080 30452 23120
rect 31564 23080 31604 23120
rect 31756 23080 31796 23120
rect 31852 23080 31892 23120
rect 32908 23080 32948 23120
rect 33580 23080 33620 23120
rect 33868 23080 33908 23120
rect 35020 23080 35060 23120
rect 35116 23080 35156 23120
rect 35212 23080 35252 23120
rect 35308 23080 35348 23120
rect 35884 23080 35924 23120
rect 36172 23080 36212 23120
rect 36460 23080 36500 23120
rect 36652 23080 36692 23120
rect 36748 23080 36788 23120
rect 37804 23080 37844 23120
rect 39052 23080 39092 23120
rect 39340 23080 39380 23120
rect 40300 23080 40340 23120
rect 40588 23080 40628 23120
rect 40684 23080 40724 23120
rect 41260 23080 41300 23120
rect 41356 23080 41396 23120
rect 41548 23080 41588 23120
rect 41740 23080 41780 23120
rect 41836 23080 41876 23120
rect 41932 23080 41972 23120
rect 42028 23080 42068 23120
rect 42220 23080 42260 23120
rect 43756 23080 43796 23120
rect 44812 23080 44852 23120
rect 46156 23080 46196 23120
rect 47020 23080 47060 23120
rect 48652 23080 48692 23120
rect 49900 23080 49940 23120
rect 50764 23080 50804 23120
rect 51148 23080 51188 23120
rect 652 22996 692 23036
rect 24748 22996 24788 23036
rect 25132 22996 25172 23036
rect 25324 22996 25364 23036
rect 28108 22996 28148 23036
rect 30124 22996 30164 23036
rect 37996 22996 38036 23036
rect 44140 22996 44180 23036
rect 5164 22912 5204 22952
rect 10348 22912 10388 22952
rect 12556 22912 12596 22952
rect 23404 22912 23444 22952
rect 25228 22912 25268 22952
rect 29932 22912 29972 22952
rect 32044 22912 32084 22952
rect 34156 22912 34196 22952
rect 39628 22912 39668 22952
rect 41068 22912 41108 22952
rect 41548 22912 41588 22952
rect 45004 22912 45044 22952
rect 47596 22912 47636 22952
rect 844 22828 884 22868
rect 3916 22828 3956 22868
rect 5836 22828 5876 22868
rect 9676 22828 9716 22868
rect 13420 22828 13460 22868
rect 16972 22828 17012 22868
rect 19948 22828 19988 22868
rect 24652 22828 24692 22868
rect 27052 22828 27092 22868
rect 31564 22828 31604 22868
rect 35500 22828 35540 22868
rect 37132 22828 37172 22868
rect 40012 22828 40052 22868
rect 42892 22828 42932 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4972 22492 5012 22532
rect 5644 22492 5684 22532
rect 8716 22492 8756 22532
rect 11308 22492 11348 22532
rect 12748 22492 12788 22532
rect 14860 22492 14900 22532
rect 19276 22492 19316 22532
rect 20044 22492 20084 22532
rect 23788 22492 23828 22532
rect 24460 22492 24500 22532
rect 26092 22492 26132 22532
rect 30700 22492 30740 22532
rect 33964 22492 34004 22532
rect 36844 22492 36884 22532
rect 40684 22492 40724 22532
rect 44716 22492 44756 22532
rect 45772 22492 45812 22532
rect 49132 22492 49172 22532
rect 7084 22408 7124 22448
rect 13996 22408 14036 22448
rect 15724 22408 15764 22448
rect 18508 22408 18548 22448
rect 21676 22408 21716 22448
rect 24652 22408 24692 22448
rect 37324 22408 37364 22448
rect 46156 22408 46196 22448
rect 3628 22324 3668 22364
rect 8236 22324 8276 22364
rect 29164 22324 29204 22364
rect 1228 22240 1268 22280
rect 1612 22240 1652 22280
rect 2476 22240 2516 22280
rect 3916 22240 3956 22280
rect 4012 22240 4052 22280
rect 4108 22240 4148 22280
rect 4300 22240 4340 22280
rect 5164 22240 5204 22280
rect 6028 22240 6068 22280
rect 6412 22240 6452 22280
rect 6508 22240 6548 22280
rect 6604 22240 6644 22280
rect 7372 22240 7412 22280
rect 9388 22240 9428 22280
rect 9580 22240 9620 22280
rect 10636 22240 10676 22280
rect 10924 22240 10964 22280
rect 11020 22240 11060 22280
rect 12076 22240 12116 22280
rect 12940 22240 12980 22280
rect 13516 22240 13556 22280
rect 13612 22240 13652 22280
rect 13708 22240 13748 22280
rect 13804 22240 13844 22280
rect 14572 22240 14612 22280
rect 15532 22240 15572 22280
rect 16108 22240 16148 22280
rect 17164 22240 17204 22280
rect 18124 22240 18164 22280
rect 18220 22240 18260 22280
rect 18316 22240 18356 22280
rect 18892 22240 18932 22280
rect 19180 22240 19220 22280
rect 19948 22240 19988 22280
rect 23116 22240 23156 22280
rect 23308 22240 23348 22280
rect 23500 22240 23540 22280
rect 23596 22240 23636 22280
rect 23788 22240 23828 22280
rect 23980 22240 24020 22280
rect 24172 22240 24212 22280
rect 24268 22240 24308 22280
rect 24652 22240 24692 22280
rect 24940 22240 24980 22280
rect 25036 22240 25076 22280
rect 25420 22240 25460 22280
rect 27244 22240 27284 22280
rect 27436 22240 27476 22280
rect 28588 22240 28628 22280
rect 28684 22240 28724 22280
rect 28780 22240 28820 22280
rect 28876 22240 28916 22280
rect 29932 22240 29972 22280
rect 30412 22240 30452 22280
rect 31564 22240 31604 22280
rect 31948 22240 31988 22280
rect 32812 22240 32852 22280
rect 34444 22240 34484 22280
rect 34828 22240 34868 22280
rect 35692 22240 35732 22280
rect 37516 22240 37556 22280
rect 38572 22240 38612 22280
rect 38668 22240 38708 22280
rect 38764 22240 38804 22280
rect 38956 22240 38996 22280
rect 39052 22240 39092 22280
rect 39244 22240 39284 22280
rect 40108 22240 40148 22280
rect 40396 22240 40436 22280
rect 41356 22240 41396 22280
rect 41644 22240 41684 22280
rect 41740 22240 41780 22280
rect 41836 22240 41876 22280
rect 42028 22240 42068 22280
rect 42124 22240 42164 22280
rect 42316 22240 42356 22280
rect 42700 22240 42740 22280
rect 43564 22240 43604 22280
rect 45100 22240 45140 22280
rect 46732 22240 46772 22280
rect 47116 22240 47156 22280
rect 47980 22240 48020 22280
rect 23212 22156 23252 22196
rect 652 22072 692 22112
rect 3820 22072 3860 22112
rect 6700 22072 6740 22112
rect 10252 22072 10292 22112
rect 16780 22072 16820 22112
rect 17836 22072 17876 22112
rect 18028 22072 18068 22112
rect 18988 22072 19028 22112
rect 24076 22072 24116 22112
rect 25228 22072 25268 22112
rect 26092 22072 26132 22112
rect 26572 22072 26612 22112
rect 28108 22072 28148 22112
rect 30892 22072 30932 22112
rect 38188 22072 38228 22112
rect 38476 22072 38516 22112
rect 39148 22072 39188 22112
rect 39436 22072 39476 22112
rect 41548 22072 41588 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4972 21736 5012 21776
rect 9004 21736 9044 21776
rect 9196 21736 9236 21776
rect 15436 21736 15476 21776
rect 16492 21736 16532 21776
rect 19660 21736 19700 21776
rect 25708 21736 25748 21776
rect 27340 21736 27380 21776
rect 30604 21736 30644 21776
rect 36268 21736 36308 21776
rect 36940 21736 36980 21776
rect 45292 21736 45332 21776
rect 2764 21652 2804 21692
rect 11596 21652 11636 21692
rect 13036 21652 13076 21692
rect 17260 21652 17300 21692
rect 25324 21652 25364 21692
rect 28204 21652 28244 21692
rect 39340 21652 39380 21692
rect 2668 21568 2708 21608
rect 2860 21568 2900 21608
rect 2956 21568 2996 21608
rect 3148 21568 3188 21608
rect 4108 21568 4148 21608
rect 4492 21568 4532 21608
rect 4684 21568 4724 21608
rect 4780 21568 4820 21608
rect 5068 21568 5108 21608
rect 5164 21568 5204 21608
rect 5260 21568 5300 21608
rect 5548 21568 5588 21608
rect 5740 21568 5780 21608
rect 6412 21568 6452 21608
rect 6604 21568 6644 21608
rect 6988 21568 7028 21608
rect 7852 21568 7892 21608
rect 10348 21568 10388 21608
rect 11212 21568 11252 21608
rect 13420 21568 13460 21608
rect 14284 21568 14324 21608
rect 15628 21568 15668 21608
rect 15724 21568 15764 21608
rect 16876 21568 16916 21608
rect 17644 21568 17684 21608
rect 18508 21568 18548 21608
rect 21196 21568 21236 21608
rect 21580 21568 21620 21608
rect 22444 21568 22484 21608
rect 23692 21568 23732 21608
rect 24364 21568 24404 21608
rect 24460 21568 24500 21608
rect 25228 21568 25268 21608
rect 25420 21568 25460 21608
rect 25612 21568 25652 21608
rect 25804 21568 25844 21608
rect 26092 21568 26132 21608
rect 27052 21568 27092 21608
rect 27532 21568 27572 21608
rect 27628 21568 27668 21608
rect 28588 21568 28628 21608
rect 29452 21568 29492 21608
rect 35788 21568 35828 21608
rect 38092 21568 38132 21608
rect 38956 21568 38996 21608
rect 40300 21568 40340 21608
rect 41164 21568 41204 21608
rect 41452 21568 41492 21608
rect 41644 21568 41684 21608
rect 41740 21568 41780 21608
rect 41932 21568 41972 21608
rect 42124 21568 42164 21608
rect 43276 21568 43316 21608
rect 44428 21568 44468 21608
rect 44524 21568 44564 21608
rect 44716 21568 44756 21608
rect 44812 21568 44852 21608
rect 44908 21568 44948 21608
rect 45004 21568 45044 21608
rect 45196 21568 45236 21608
rect 45388 21568 45428 21608
rect 45484 21568 45524 21608
rect 24844 21484 24884 21524
rect 1708 21400 1748 21440
rect 2188 21400 2228 21440
rect 4492 21400 4532 21440
rect 5452 21400 5492 21440
rect 11788 21400 11828 21440
rect 24172 21400 24212 21440
rect 25036 21400 25076 21440
rect 28012 21400 28052 21440
rect 34924 21400 34964 21440
rect 41932 21400 41972 21440
rect 43564 21400 43604 21440
rect 39628 21316 39668 21356
rect 40492 21316 40532 21356
rect 41356 21316 41396 21356
rect 42796 21316 42836 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4108 20980 4148 21020
rect 5932 20980 5972 21020
rect 6220 20980 6260 21020
rect 11692 20980 11732 21020
rect 16972 20980 17012 21020
rect 33772 20980 33812 21020
rect 37228 20980 37268 21020
rect 37804 20980 37844 21020
rect 38956 20980 38996 21020
rect 44620 20980 44660 21020
rect 16108 20896 16148 20936
rect 25036 20896 25076 20936
rect 27628 20896 27668 20936
rect 29068 20896 29108 20936
rect 34828 20896 34868 20936
rect 13228 20812 13268 20852
rect 17260 20812 17300 20852
rect 21292 20812 21332 20852
rect 25708 20812 25748 20852
rect 41644 20812 41684 20852
rect 1708 20728 1748 20768
rect 2092 20728 2132 20768
rect 2956 20728 2996 20768
rect 5068 20728 5108 20768
rect 5260 20728 5300 20768
rect 6892 20728 6932 20768
rect 7372 20728 7412 20768
rect 8812 20728 8852 20768
rect 9004 20728 9044 20768
rect 9292 20728 9332 20768
rect 9580 20728 9620 20768
rect 9676 20728 9716 20768
rect 9772 20728 9812 20768
rect 9868 20728 9908 20768
rect 10348 20728 10388 20768
rect 10540 20728 10580 20768
rect 10636 20728 10676 20768
rect 11500 20728 11540 20768
rect 12076 20728 12116 20768
rect 12364 20728 12404 20768
rect 13996 20728 14036 20768
rect 15148 20728 15188 20768
rect 15340 20728 15380 20768
rect 15436 20728 15476 20768
rect 15628 20728 15668 20768
rect 15724 20728 15764 20768
rect 15820 20728 15860 20768
rect 15916 20728 15956 20768
rect 16684 20728 16724 20768
rect 16780 20728 16820 20768
rect 16972 20728 17012 20768
rect 18124 20728 18164 20768
rect 19276 20728 19316 20768
rect 20140 20739 20180 20779
rect 22156 20728 22196 20768
rect 22348 20728 22388 20768
rect 22444 20728 22484 20768
rect 22540 20728 22580 20768
rect 24460 20728 24500 20768
rect 26572 20728 26612 20768
rect 26956 20728 26996 20768
rect 33292 20728 33332 20768
rect 35404 20728 35444 20768
rect 35500 20728 35540 20768
rect 35596 20728 35636 20768
rect 37132 20728 37172 20768
rect 37900 20728 37940 20768
rect 39052 20728 39092 20768
rect 39244 20728 39284 20768
rect 39628 20728 39668 20768
rect 40492 20728 40532 20768
rect 42220 20728 42260 20768
rect 42604 20728 42644 20768
rect 43468 20728 43508 20768
rect 10828 20644 10868 20684
rect 11980 20644 12020 20684
rect 18892 20644 18932 20684
rect 652 20560 692 20600
rect 4396 20560 4436 20600
rect 7852 20560 7892 20600
rect 9196 20560 9236 20600
rect 10444 20560 10484 20600
rect 15244 20560 15284 20600
rect 21484 20560 21524 20600
rect 22636 20560 22676 20600
rect 33772 20560 33812 20600
rect 35308 20560 35348 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 21100 20282 21140 20322
rect 652 20224 692 20264
rect 6508 20224 6548 20264
rect 21772 20224 21812 20264
rect 21964 20224 22004 20264
rect 4108 20140 4148 20180
rect 15628 20140 15668 20180
rect 19756 20140 19796 20180
rect 21484 20140 21524 20180
rect 26668 20140 26708 20180
rect 39724 20140 39764 20180
rect 4492 20056 4532 20096
rect 5356 20056 5396 20096
rect 6796 20056 6836 20096
rect 6988 20056 7028 20096
rect 7084 20056 7124 20096
rect 7660 20056 7700 20096
rect 9292 20056 9332 20096
rect 10156 20056 10196 20096
rect 10444 20056 10484 20096
rect 10828 20056 10868 20096
rect 11692 20056 11732 20096
rect 12940 20056 12980 20096
rect 15436 20056 15476 20096
rect 16300 20056 16340 20096
rect 16684 20056 16724 20096
rect 19276 20056 19316 20096
rect 19372 20056 19412 20096
rect 19468 20056 19508 20096
rect 19564 20056 19604 20096
rect 20428 20056 20468 20096
rect 20908 20056 20948 20096
rect 21004 20056 21044 20096
rect 21676 20056 21716 20096
rect 22156 20056 22196 20096
rect 22252 20056 22292 20096
rect 23308 20056 23348 20096
rect 24076 20056 24116 20096
rect 24268 20056 24308 20096
rect 24844 20056 24884 20096
rect 25420 20064 25460 20104
rect 25804 20056 25844 20096
rect 26092 20056 26132 20096
rect 26284 20056 26324 20096
rect 26572 20056 26612 20096
rect 26764 20056 26804 20096
rect 26956 20056 26996 20096
rect 27916 20056 27956 20096
rect 28588 20056 28628 20096
rect 28972 20056 29012 20096
rect 29836 20056 29876 20096
rect 31468 20056 31508 20096
rect 31852 20056 31892 20096
rect 32332 20056 32372 20096
rect 33292 20056 33332 20096
rect 34348 20056 34388 20096
rect 34732 20056 34772 20096
rect 35596 20056 35636 20096
rect 36844 20056 36884 20096
rect 39820 20056 39860 20096
rect 39916 20056 39956 20096
rect 40012 20056 40052 20096
rect 40204 20056 40244 20096
rect 40396 20056 40436 20096
rect 40492 20056 40532 20096
rect 33580 19972 33620 20012
rect 6796 19888 6836 19928
rect 13228 19888 13268 19928
rect 16876 19888 16916 19928
rect 18508 19888 18548 19928
rect 19084 19888 19124 19928
rect 20620 19888 20660 19928
rect 23500 19888 23540 19928
rect 24844 19888 24884 19928
rect 26284 19888 26324 19928
rect 28396 19888 28436 19928
rect 37900 19888 37940 19928
rect 39532 19888 39572 19928
rect 40204 19888 40244 19928
rect 42796 19888 42836 19928
rect 7948 19804 7988 19844
rect 14764 19804 14804 19844
rect 22636 19804 22676 19844
rect 24172 19804 24212 19844
rect 25036 19804 25076 19844
rect 25324 19804 25364 19844
rect 30988 19804 31028 19844
rect 31948 19804 31988 19844
rect 33772 19804 33812 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 5356 19468 5396 19508
rect 10348 19468 10388 19508
rect 14860 19468 14900 19508
rect 17452 19468 17492 19508
rect 20812 19468 20852 19508
rect 34924 19468 34964 19508
rect 1996 19384 2036 19424
rect 3724 19384 3764 19424
rect 5836 19384 5876 19424
rect 36364 19384 36404 19424
rect 8908 19300 8948 19340
rect 35116 19300 35156 19340
rect 3916 19216 3956 19256
rect 4012 19216 4052 19256
rect 4204 19216 4244 19256
rect 4492 19216 4532 19256
rect 5452 19216 5492 19256
rect 6028 19216 6068 19256
rect 6124 19216 6164 19256
rect 6220 19216 6260 19256
rect 6892 19216 6932 19256
rect 7756 19216 7796 19256
rect 10444 19216 10484 19256
rect 10636 19216 10676 19256
rect 11308 19216 11348 19256
rect 11692 19216 11732 19256
rect 11788 19216 11828 19256
rect 11980 19216 12020 19256
rect 12076 19216 12116 19256
rect 12268 19216 12308 19256
rect 12844 19216 12884 19256
rect 13708 19216 13748 19256
rect 15052 19216 15092 19256
rect 15436 19216 15476 19256
rect 16300 19216 16340 19256
rect 17644 19216 17684 19256
rect 17932 19216 17972 19256
rect 18508 19216 18548 19256
rect 19372 19216 19412 19256
rect 20716 19216 20756 19256
rect 21004 19216 21044 19256
rect 22156 19216 22196 19256
rect 22540 19216 22580 19256
rect 23404 19216 23444 19256
rect 24556 19216 24596 19256
rect 25612 19216 25652 19256
rect 25804 19216 25844 19256
rect 26092 19216 26132 19256
rect 26668 19216 26708 19256
rect 28012 19216 28052 19256
rect 28108 19216 28148 19256
rect 28204 19216 28244 19256
rect 28300 19216 28340 19256
rect 28684 19216 28724 19256
rect 29164 19216 29204 19256
rect 29260 19216 29300 19256
rect 29356 19216 29396 19256
rect 29548 19216 29588 19256
rect 29932 19216 29972 19256
rect 30796 19216 30836 19256
rect 31948 19216 31988 19256
rect 33196 19216 33236 19256
rect 33868 19216 33908 19256
rect 33964 19216 34004 19256
rect 34060 19216 34100 19256
rect 34252 19216 34292 19256
rect 35308 19216 35348 19256
rect 35404 19216 35444 19256
rect 36940 19216 36980 19256
rect 37324 19216 37364 19256
rect 37708 19216 37748 19256
rect 38572 19216 38612 19256
rect 39724 19216 39764 19256
rect 40684 19216 40724 19256
rect 6508 19132 6548 19172
rect 12460 19132 12500 19172
rect 18124 19132 18164 19172
rect 32428 19132 32468 19172
rect 652 19048 692 19088
rect 4108 19048 4148 19088
rect 5164 19048 5204 19088
rect 6316 19048 6356 19088
rect 12172 19048 12212 19088
rect 17836 19048 17876 19088
rect 20524 19048 20564 19088
rect 21676 19048 21716 19088
rect 25900 19048 25940 19088
rect 27148 19048 27188 19088
rect 27820 19048 27860 19088
rect 28780 19048 28820 19088
rect 29068 19048 29108 19088
rect 33772 19048 33812 19088
rect 40012 19048 40052 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 652 18712 692 18752
rect 3724 18712 3764 18752
rect 4588 18712 4628 18752
rect 4780 18712 4820 18752
rect 6796 18712 6836 18752
rect 11596 18712 11636 18752
rect 12460 18712 12500 18752
rect 13324 18712 13364 18752
rect 14956 18712 14996 18752
rect 16396 18712 16436 18752
rect 19564 18712 19604 18752
rect 20524 18712 20564 18752
rect 22060 18712 22100 18752
rect 24748 18712 24788 18752
rect 31852 18754 31892 18794
rect 26668 18712 26708 18752
rect 35404 18712 35444 18752
rect 36364 18712 36404 18752
rect 1324 18628 1364 18668
rect 23116 18628 23156 18668
rect 1708 18544 1748 18584
rect 2572 18544 2612 18584
rect 3916 18544 3956 18584
rect 4876 18544 4916 18584
rect 6604 18544 6644 18584
rect 7468 18544 7508 18584
rect 7660 18544 7700 18584
rect 7852 18544 7892 18584
rect 7948 18544 7988 18584
rect 10252 18544 10292 18584
rect 10348 18544 10388 18584
rect 10444 18544 10484 18584
rect 10540 18544 10580 18584
rect 10828 18544 10868 18584
rect 11116 18544 11156 18584
rect 11212 18544 11252 18584
rect 11308 18544 11348 18584
rect 11404 18544 11444 18584
rect 12268 18544 12308 18584
rect 13132 18544 13172 18584
rect 13996 18544 14036 18584
rect 15052 18544 15092 18584
rect 15148 18544 15188 18584
rect 15244 18544 15284 18584
rect 15436 18544 15476 18584
rect 16108 18544 16148 18584
rect 16300 18544 16340 18584
rect 20236 18544 20276 18584
rect 20620 18544 20660 18584
rect 20812 18544 20852 18584
rect 21196 18544 21236 18584
rect 21388 18544 21428 18584
rect 22252 18544 22292 18584
rect 22636 18544 22676 18584
rect 23212 18544 23252 18584
rect 23308 18544 23348 18584
rect 23404 18544 23444 18584
rect 23596 18544 23636 18584
rect 23692 18544 23732 18584
rect 23788 18544 23828 18584
rect 23884 18544 23924 18584
rect 24076 18544 24116 18584
rect 25132 18544 25172 18584
rect 26668 18544 26708 18584
rect 26764 18544 26804 18584
rect 27148 18544 27188 18584
rect 27532 18544 27572 18584
rect 28396 18544 28436 18584
rect 29548 18544 29588 18584
rect 29836 18544 29876 18584
rect 31372 18544 31412 18584
rect 31660 18544 31700 18584
rect 31852 18544 31892 18584
rect 32236 18544 32276 18584
rect 33100 18544 33140 18584
rect 33580 18544 33620 18584
rect 33676 18544 33716 18584
rect 33868 18544 33908 18584
rect 34252 18544 34292 18584
rect 34348 18544 34388 18584
rect 35020 18544 35060 18584
rect 35116 18544 35156 18584
rect 35687 18544 35727 18584
rect 35788 18544 35828 18584
rect 35884 18544 35924 18584
rect 36076 18544 36116 18584
rect 36172 18544 36212 18584
rect 37036 18544 37076 18584
rect 37228 18544 37268 18584
rect 37324 18544 37364 18584
rect 37420 18544 37460 18584
rect 37516 18544 37556 18584
rect 37900 18544 37940 18584
rect 38860 18544 38900 18584
rect 39244 18544 39284 18584
rect 40492 18544 40532 18584
rect 41452 18544 41492 18584
rect 20908 18460 20948 18500
rect 21100 18460 21140 18500
rect 22348 18460 22388 18500
rect 22540 18460 22580 18500
rect 26572 18460 26612 18500
rect 34636 18460 34676 18500
rect 5740 18376 5780 18416
rect 7660 18376 7700 18416
rect 9388 18376 9428 18416
rect 14188 18376 14228 18416
rect 18220 18376 18260 18416
rect 21004 18376 21044 18416
rect 22444 18376 22484 18416
rect 25708 18376 25748 18416
rect 26476 18376 26516 18416
rect 33868 18376 33908 18416
rect 4588 18292 4628 18332
rect 5068 18292 5108 18332
rect 5932 18292 5972 18332
rect 10924 18292 10964 18332
rect 24748 18292 24788 18332
rect 30508 18292 30548 18332
rect 30700 18292 30740 18332
rect 36172 18292 36212 18332
rect 39916 18292 39956 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 3916 17956 3956 17996
rect 11308 17956 11348 17996
rect 14956 17956 14996 17996
rect 20140 17956 20180 17996
rect 24364 17956 24404 17996
rect 26092 17956 26132 17996
rect 28972 17956 29012 17996
rect 29836 17956 29876 17996
rect 30316 17956 30356 17996
rect 34156 17956 34196 17996
rect 34636 17956 34676 17996
rect 1324 17872 1364 17912
rect 4684 17872 4724 17912
rect 8716 17872 8756 17912
rect 27244 17872 27284 17912
rect 27916 17872 27956 17912
rect 37708 17872 37748 17912
rect 31756 17788 31796 17828
rect 36652 17788 36692 17828
rect 1900 17704 1940 17744
rect 2764 17704 2804 17744
rect 4396 17704 4436 17744
rect 4492 17704 4532 17744
rect 4684 17704 4724 17744
rect 4876 17704 4916 17744
rect 5740 17704 5780 17744
rect 6124 17704 6164 17744
rect 6988 17704 7028 17744
rect 8428 17704 8468 17744
rect 8524 17704 8564 17744
rect 8716 17704 8756 17744
rect 8908 17704 8948 17744
rect 9292 17704 9332 17744
rect 10156 17704 10196 17744
rect 11692 17704 11732 17744
rect 12364 17704 12404 17744
rect 12556 17704 12596 17744
rect 12940 17704 12980 17744
rect 13804 17704 13844 17744
rect 15916 17704 15956 17744
rect 17740 17704 17780 17744
rect 18124 17704 18164 17744
rect 18988 17704 19028 17744
rect 20812 17704 20852 17744
rect 21484 17704 21524 17744
rect 21676 17704 21716 17744
rect 22540 17704 22580 17744
rect 22924 17704 22964 17744
rect 23020 17704 23060 17744
rect 23212 17704 23252 17744
rect 23404 17704 23444 17744
rect 23500 17704 23540 17744
rect 23692 17704 23732 17744
rect 23884 17704 23924 17744
rect 24076 17704 24116 17744
rect 24172 17704 24212 17744
rect 24364 17704 24404 17744
rect 24460 17704 24500 17744
rect 24652 17704 24692 17744
rect 24748 17704 24788 17744
rect 24905 17719 24945 17759
rect 26092 17704 26132 17744
rect 26284 17704 26324 17744
rect 26572 17704 26612 17744
rect 27436 17704 27476 17744
rect 27628 17704 27668 17744
rect 27916 17704 27956 17744
rect 28300 17704 28340 17744
rect 29164 17704 29204 17744
rect 30988 17704 31028 17744
rect 31372 17704 31412 17744
rect 31564 17704 31604 17744
rect 31852 17704 31892 17744
rect 33196 17704 33236 17744
rect 34156 17704 34196 17744
rect 34348 17704 34388 17744
rect 34444 17704 34484 17744
rect 34636 17704 34676 17744
rect 34732 17704 34772 17744
rect 34924 17704 34964 17744
rect 35020 17704 35060 17744
rect 35121 17704 35161 17744
rect 35404 17704 35444 17744
rect 35500 17704 35540 17744
rect 35596 17704 35636 17744
rect 35692 17704 35732 17744
rect 36556 17704 36596 17744
rect 36748 17704 36788 17744
rect 37036 17704 37076 17744
rect 37132 17683 37172 17723
rect 37228 17704 37268 17744
rect 37420 17704 37460 17744
rect 37516 17704 37556 17744
rect 37708 17704 37748 17744
rect 37900 17704 37940 17744
rect 38764 17704 38804 17744
rect 39148 17704 39188 17744
rect 40012 17704 40052 17744
rect 41260 17704 41300 17744
rect 1516 17620 1556 17660
rect 16780 17620 16820 17660
rect 23116 17620 23156 17660
rect 23596 17620 23636 17660
rect 23980 17620 24020 17660
rect 26764 17620 26804 17660
rect 27532 17620 27572 17660
rect 32428 17620 32468 17660
rect 36940 17620 36980 17660
rect 652 17536 692 17576
rect 5548 17536 5588 17576
rect 8140 17536 8180 17576
rect 26476 17536 26516 17576
rect 28108 17536 28148 17576
rect 38572 17536 38612 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 27724 17258 27764 17298
rect 652 17200 692 17240
rect 3724 17200 3764 17240
rect 4396 17200 4436 17240
rect 5836 17200 5876 17240
rect 20812 17200 20852 17240
rect 21868 17200 21908 17240
rect 23404 17200 23444 17240
rect 24172 17200 24212 17240
rect 24652 17200 24692 17240
rect 25420 17200 25460 17240
rect 26572 17200 26612 17240
rect 36652 17200 36692 17240
rect 38284 17200 38324 17240
rect 39148 17200 39188 17240
rect 4108 17116 4148 17156
rect 19372 17116 19412 17156
rect 35020 17116 35060 17156
rect 3244 17032 3284 17072
rect 3436 17032 3476 17072
rect 3628 17032 3668 17072
rect 3820 17032 3860 17072
rect 3916 17032 3956 17072
rect 4300 17032 4340 17072
rect 4684 17032 4724 17072
rect 4780 17032 4820 17072
rect 4876 17032 4916 17072
rect 4972 17032 5012 17072
rect 5644 17032 5684 17072
rect 5740 17032 5780 17072
rect 5932 17032 5972 17072
rect 6124 17032 6164 17072
rect 6796 17032 6836 17072
rect 7660 17032 7700 17072
rect 7852 17032 7892 17072
rect 7948 17032 7988 17072
rect 8044 17032 8084 17072
rect 8140 17032 8180 17072
rect 8332 17032 8372 17072
rect 8524 17032 8564 17072
rect 11212 17032 11252 17072
rect 11596 17032 11636 17072
rect 12460 17032 12500 17072
rect 12652 17032 12692 17072
rect 13612 17032 13652 17072
rect 15244 17032 15284 17072
rect 15436 17032 15476 17072
rect 16684 17032 16724 17072
rect 17548 17032 17588 17072
rect 17932 17032 17972 17072
rect 18316 17032 18356 17072
rect 20044 17032 20084 17072
rect 20332 17032 20372 17072
rect 20524 17032 20564 17072
rect 20620 17032 20660 17072
rect 20908 17032 20948 17072
rect 21004 17032 21044 17072
rect 21100 17032 21140 17072
rect 21484 17032 21524 17072
rect 22540 17032 22580 17072
rect 23500 17032 23540 17072
rect 23596 17032 23636 17072
rect 23692 17032 23732 17072
rect 23884 17032 23924 17072
rect 23980 17032 24020 17072
rect 24076 17032 24116 17072
rect 24364 17032 24404 17072
rect 24460 17032 24500 17072
rect 24556 17032 24596 17072
rect 25228 17032 25268 17072
rect 25324 17032 25364 17072
rect 25516 17032 25556 17072
rect 26476 17032 26516 17072
rect 26668 17032 26708 17072
rect 26764 17032 26804 17072
rect 27244 17032 27284 17072
rect 27340 17032 27380 17072
rect 27916 17032 27956 17072
rect 27820 16990 27860 17030
rect 28775 17032 28815 17072
rect 28876 17032 28916 17072
rect 28972 17032 29012 17072
rect 29164 17032 29204 17072
rect 29260 17032 29300 17072
rect 30412 17032 30452 17072
rect 31180 17032 31220 17072
rect 31372 17032 31412 17072
rect 31660 17032 31700 17072
rect 31948 17032 31988 17072
rect 32044 17032 32084 17072
rect 32140 17032 32180 17072
rect 32236 17032 32276 17072
rect 33388 17032 33428 17072
rect 33772 17032 33812 17072
rect 34924 17032 34964 17072
rect 35116 17032 35156 17072
rect 35884 17032 35924 17072
rect 36076 17032 36116 17072
rect 36308 17032 36348 17072
rect 36460 17032 36500 17072
rect 36556 17032 36596 17072
rect 36748 17032 36788 17072
rect 36844 17032 36884 17072
rect 37073 17032 37113 17072
rect 37228 17032 37268 17072
rect 37324 17017 37364 17057
rect 37516 17017 37556 17057
rect 37612 17032 37652 17072
rect 38188 17032 38228 17072
rect 38380 17032 38420 17072
rect 38476 17032 38516 17072
rect 39628 17032 39668 17072
rect 39916 17032 39956 17072
rect 40300 17032 40340 17072
rect 41164 17032 41204 17072
rect 3340 16948 3380 16988
rect 29548 16948 29588 16988
rect 31564 16948 31604 16988
rect 37996 16948 38036 16988
rect 9868 16864 9908 16904
rect 14380 16864 14420 16904
rect 20332 16864 20372 16904
rect 34444 16864 34484 16904
rect 5164 16780 5204 16820
rect 6988 16780 7028 16820
rect 8428 16780 8468 16820
rect 10540 16780 10580 16820
rect 14572 16780 14612 16820
rect 18988 16780 19028 16820
rect 21676 16780 21716 16820
rect 23212 16780 23252 16820
rect 27436 16780 27476 16820
rect 28204 16780 28244 16820
rect 29260 16780 29300 16820
rect 32908 16780 32948 16820
rect 34060 16780 34100 16820
rect 35980 16780 36020 16820
rect 37612 16780 37652 16820
rect 39148 16780 39188 16820
rect 42316 16780 42356 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 6412 16444 6452 16484
rect 8140 16444 8180 16484
rect 8428 16444 8468 16484
rect 11788 16444 11828 16484
rect 15628 16444 15668 16484
rect 26668 16444 26708 16484
rect 1420 16360 1460 16400
rect 5452 16360 5492 16400
rect 12076 16360 12116 16400
rect 13036 16360 13076 16400
rect 16492 16360 16532 16400
rect 20332 16360 20372 16400
rect 21388 16360 21428 16400
rect 21964 16360 22004 16400
rect 22156 16360 22196 16400
rect 37036 16360 37076 16400
rect 38476 16360 38516 16400
rect 39436 16360 39476 16400
rect 41164 16360 41204 16400
rect 6604 16276 6644 16316
rect 20236 16276 20276 16316
rect 20428 16276 20468 16316
rect 21292 16276 21332 16316
rect 21484 16276 21524 16316
rect 27724 16276 27764 16316
rect 3052 16192 3092 16232
rect 3244 16192 3284 16232
rect 3436 16192 3476 16232
rect 3628 16192 3668 16232
rect 3724 16192 3764 16232
rect 4012 16192 4052 16232
rect 4684 16192 4724 16232
rect 4972 16192 5012 16232
rect 5164 16192 5204 16232
rect 5452 16192 5492 16232
rect 5644 16192 5684 16232
rect 5740 16192 5780 16232
rect 5932 16192 5972 16232
rect 6124 16192 6164 16232
rect 6412 16192 6452 16232
rect 7084 16192 7124 16232
rect 7180 16192 7220 16232
rect 7564 16192 7604 16232
rect 7852 16192 7892 16232
rect 7948 16192 7988 16232
rect 8140 16192 8180 16232
rect 8332 16192 8372 16232
rect 8524 16192 8564 16232
rect 9388 16192 9428 16232
rect 9772 16192 9812 16232
rect 10636 16192 10676 16232
rect 12076 16192 12116 16232
rect 12268 16192 12308 16232
rect 12364 16192 12404 16232
rect 13228 16192 13268 16232
rect 14092 16192 14132 16232
rect 15340 16192 15380 16232
rect 16492 16192 16532 16232
rect 16684 16192 16724 16232
rect 18604 16192 18644 16232
rect 18892 16192 18932 16232
rect 19372 16192 19412 16232
rect 19660 16192 19700 16232
rect 20524 16192 20564 16232
rect 20140 16150 20180 16190
rect 20716 16192 20756 16232
rect 20812 16192 20852 16232
rect 20908 16192 20948 16232
rect 21004 16192 21044 16232
rect 21196 16192 21236 16232
rect 21580 16192 21620 16232
rect 21964 16192 22004 16232
rect 22348 16192 22388 16232
rect 22444 16192 22484 16232
rect 22636 16192 22676 16232
rect 22828 16192 22868 16232
rect 22924 16192 22964 16232
rect 23404 16192 23444 16232
rect 24364 16192 24404 16232
rect 24748 16192 24788 16232
rect 26188 16192 26228 16232
rect 26284 16192 26324 16232
rect 26380 16192 26420 16232
rect 26476 16192 26516 16232
rect 26668 16192 26708 16232
rect 26860 16192 26900 16232
rect 26956 16192 26996 16232
rect 27436 16192 27476 16232
rect 27532 16192 27572 16232
rect 27916 16192 27956 16232
rect 28012 16192 28052 16232
rect 28204 16192 28244 16232
rect 28396 16192 28436 16232
rect 28492 16192 28532 16232
rect 28684 16192 28724 16232
rect 28972 16192 29012 16232
rect 29068 16192 29108 16232
rect 29260 16192 29300 16232
rect 29932 16192 29972 16232
rect 30028 16192 30068 16232
rect 30124 16192 30164 16232
rect 30508 16192 30548 16232
rect 32428 16192 32468 16232
rect 32812 16192 32852 16232
rect 32908 16192 32948 16232
rect 33100 16192 33140 16232
rect 33292 16192 33332 16232
rect 33484 16192 33524 16232
rect 33580 16192 33620 16232
rect 33772 16192 33812 16232
rect 33964 16192 34004 16232
rect 34060 16192 34100 16232
rect 34636 16192 34676 16232
rect 35596 16192 35636 16232
rect 35788 16192 35828 16232
rect 35980 16192 36020 16232
rect 36076 16192 36116 16232
rect 36268 16192 36308 16232
rect 36364 16192 36404 16232
rect 36460 16192 36500 16232
rect 36556 16192 36596 16232
rect 36940 16192 36980 16232
rect 37132 16192 37172 16232
rect 37324 16192 37364 16232
rect 37420 16192 37460 16232
rect 37516 16192 37556 16232
rect 37612 16192 37652 16232
rect 38092 16192 38132 16232
rect 38188 16192 38228 16232
rect 38956 16192 38996 16232
rect 39148 16192 39188 16232
rect 39244 16192 39284 16232
rect 40108 16192 40148 16232
rect 40300 16192 40340 16232
rect 40972 16192 41012 16232
rect 3148 16108 3188 16148
rect 16204 16108 16244 16148
rect 19084 16108 19124 16148
rect 19852 16108 19892 16148
rect 24556 16108 24596 16148
rect 29164 16108 29204 16148
rect 31660 16108 31700 16148
rect 33004 16108 33044 16148
rect 35884 16108 35924 16148
rect 652 16024 692 16064
rect 3532 16024 3572 16064
rect 5068 16024 5108 16064
rect 6028 16024 6068 16064
rect 22540 16024 22580 16064
rect 23116 16024 23156 16064
rect 24844 16024 24884 16064
rect 28204 16024 28244 16064
rect 28684 16024 28724 16064
rect 29836 16024 29876 16064
rect 30892 16024 30932 16064
rect 33292 16024 33332 16064
rect 33772 16024 33812 16064
rect 37996 16020 38036 16060
rect 38956 16024 38996 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3820 15688 3860 15728
rect 4108 15688 4148 15728
rect 7660 15692 7700 15732
rect 8236 15688 8276 15728
rect 11692 15688 11732 15728
rect 19372 15688 19412 15728
rect 19852 15688 19892 15728
rect 20332 15688 20372 15728
rect 21676 15719 21716 15759
rect 23596 15688 23636 15728
rect 23884 15688 23924 15728
rect 25612 15688 25652 15728
rect 27436 15688 27476 15728
rect 27916 15688 27956 15728
rect 30508 15688 30548 15728
rect 32716 15688 32756 15728
rect 33868 15692 33908 15732
rect 35788 15688 35828 15728
rect 36844 15688 36884 15728
rect 38668 15688 38708 15728
rect 19084 15604 19124 15644
rect 19564 15604 19604 15644
rect 21004 15604 21044 15644
rect 25900 15604 25940 15644
rect 940 15520 980 15560
rect 1324 15520 1364 15560
rect 2188 15520 2228 15560
rect 4012 15520 4052 15560
rect 4300 15520 4340 15560
rect 4396 15520 4436 15560
rect 4588 15520 4628 15560
rect 4780 15520 4820 15560
rect 6316 15520 6356 15560
rect 6508 15520 6548 15560
rect 6604 15520 6644 15560
rect 7468 15520 7508 15560
rect 7564 15520 7604 15560
rect 7852 15520 7892 15560
rect 8140 15520 8180 15560
rect 8332 15520 8372 15560
rect 8524 15520 8564 15560
rect 8716 15520 8756 15560
rect 8812 15520 8852 15560
rect 9100 15520 9140 15560
rect 9292 15520 9332 15560
rect 9676 15520 9716 15560
rect 10540 15520 10580 15560
rect 12940 15520 12980 15560
rect 13324 15520 13364 15560
rect 14188 15520 14228 15560
rect 15436 15520 15476 15560
rect 16300 15520 16340 15560
rect 16684 15520 16724 15560
rect 16780 15520 16820 15560
rect 18604 15520 18644 15560
rect 18700 15520 18740 15560
rect 18892 15520 18932 15560
rect 19276 15520 19316 15560
rect 19756 15520 19796 15560
rect 20044 15520 20084 15560
rect 20140 15520 20180 15560
rect 20236 15520 20276 15560
rect 20716 15520 20756 15560
rect 20812 15520 20852 15560
rect 20908 15520 20948 15560
rect 21484 15520 21524 15560
rect 21868 15520 21908 15560
rect 6700 15436 6740 15476
rect 21580 15478 21620 15518
rect 22060 15520 22100 15560
rect 22252 15520 22292 15560
rect 22444 15520 22484 15560
rect 22540 15520 22580 15560
rect 22732 15520 22772 15560
rect 23116 15520 23156 15560
rect 23788 15520 23828 15560
rect 24076 15520 24116 15560
rect 24268 15520 24308 15560
rect 24748 15520 24788 15560
rect 25132 15520 25172 15560
rect 25324 15520 25364 15560
rect 25420 15520 25460 15560
rect 25612 15520 25652 15560
rect 26092 15520 26132 15560
rect 27628 15520 27668 15560
rect 28012 15520 28052 15560
rect 28108 15520 28148 15560
rect 28204 15520 28244 15560
rect 28396 15520 28436 15560
rect 29260 15520 29300 15560
rect 29356 15520 29396 15560
rect 29452 15520 29492 15560
rect 29548 15520 29588 15560
rect 29740 15520 29780 15560
rect 29932 15520 29972 15560
rect 30028 15520 30068 15560
rect 30604 15520 30644 15560
rect 31564 15520 31604 15560
rect 31660 15520 31700 15560
rect 31852 15520 31892 15560
rect 31948 15491 31988 15531
rect 32049 15520 32089 15560
rect 32423 15520 32463 15560
rect 32524 15520 32564 15560
rect 32620 15520 32660 15560
rect 32812 15520 32852 15560
rect 32908 15520 32948 15560
rect 33676 15520 33716 15560
rect 33772 15520 33812 15560
rect 34348 15520 34388 15560
rect 34444 15520 34484 15560
rect 34828 15520 34868 15560
rect 34924 15520 34964 15560
rect 35020 15520 35060 15560
rect 35404 15520 35444 15560
rect 35596 15520 35636 15560
rect 35884 15520 35924 15560
rect 35980 15520 36020 15560
rect 36076 15520 36116 15560
rect 36268 15501 36308 15541
rect 36364 15520 36404 15560
rect 36556 15520 36596 15560
rect 36748 15520 36788 15560
rect 36844 15520 36884 15560
rect 37516 15520 37556 15560
rect 38092 15520 38132 15560
rect 38188 15520 38228 15560
rect 38668 15520 38708 15560
rect 38860 15520 38900 15560
rect 38956 15520 38996 15560
rect 39532 15520 39572 15560
rect 40396 15520 40436 15560
rect 7948 15436 7988 15476
rect 21964 15436 22004 15476
rect 22828 15436 22868 15476
rect 23020 15436 23060 15476
rect 24844 15436 24884 15476
rect 25036 15436 25076 15476
rect 25900 15436 25940 15476
rect 34636 15436 34676 15476
rect 36940 15436 36980 15476
rect 4588 15352 4628 15392
rect 6796 15352 6836 15392
rect 6892 15352 6932 15392
rect 8812 15352 8852 15392
rect 22924 15352 22964 15392
rect 24172 15352 24212 15392
rect 24940 15352 24980 15392
rect 27628 15352 27668 15392
rect 29836 15352 29876 15392
rect 33388 15352 33428 15392
rect 35596 15352 35636 15392
rect 37036 15352 37076 15392
rect 37516 15352 37556 15392
rect 37708 15352 37748 15392
rect 39148 15352 39188 15392
rect 3340 15268 3380 15308
rect 3820 15268 3860 15308
rect 5452 15268 5492 15308
rect 5644 15268 5684 15308
rect 7180 15268 7220 15308
rect 9004 15268 9044 15308
rect 15628 15268 15668 15308
rect 16972 15268 17012 15308
rect 18892 15268 18932 15308
rect 21196 15268 21236 15308
rect 22252 15268 22292 15308
rect 29068 15268 29108 15308
rect 31564 15268 31604 15308
rect 34540 15268 34580 15308
rect 36556 15268 36596 15308
rect 38380 15268 38420 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4684 14932 4724 14972
rect 7084 14932 7124 14972
rect 9100 14932 9140 14972
rect 9292 14932 9332 14972
rect 16012 14932 16052 14972
rect 17548 14932 17588 14972
rect 20140 14932 20180 14972
rect 35692 14932 35732 14972
rect 36076 14932 36116 14972
rect 37132 14932 37172 14972
rect 41548 14932 41588 14972
rect 1516 14848 1556 14888
rect 3436 14848 3476 14888
rect 6604 14848 6644 14888
rect 10156 14848 10196 14888
rect 32332 14848 32372 14888
rect 37612 14764 37652 14804
rect 2956 14680 2996 14720
rect 3052 14680 3092 14720
rect 3244 14680 3284 14720
rect 3628 14680 3668 14720
rect 3724 14711 3764 14751
rect 4204 14680 4244 14720
rect 4300 14680 4340 14720
rect 4396 14680 4436 14720
rect 4492 14680 4532 14720
rect 5548 14680 5588 14720
rect 6412 14680 6452 14720
rect 6604 14680 6644 14720
rect 6700 14680 6740 14720
rect 6892 14680 6932 14720
rect 7756 14680 7796 14720
rect 7948 14680 7988 14720
rect 8044 14680 8084 14720
rect 8236 14680 8276 14720
rect 8812 14680 8852 14720
rect 8908 14680 8948 14720
rect 9100 14680 9140 14720
rect 9964 14680 10004 14720
rect 11404 14680 11444 14720
rect 13804 14680 13844 14720
rect 13900 14680 13940 14720
rect 13996 14680 14036 14720
rect 14380 14680 14420 14720
rect 14572 14680 14612 14720
rect 15052 14680 15092 14720
rect 15148 14680 15188 14720
rect 15820 14680 15860 14720
rect 15916 14680 15956 14720
rect 17164 14680 17204 14720
rect 17548 14680 17588 14720
rect 17644 14680 17684 14720
rect 17836 14680 17876 14720
rect 17932 14680 17972 14720
rect 18033 14680 18073 14720
rect 18316 14680 18356 14720
rect 18412 14680 18452 14720
rect 18508 14680 18548 14720
rect 18604 14680 18644 14720
rect 19852 14680 19892 14720
rect 19948 14680 19988 14720
rect 20140 14638 20180 14678
rect 20332 14680 20372 14720
rect 20620 14680 20660 14720
rect 20812 14680 20852 14720
rect 21676 14680 21716 14720
rect 22060 14680 22100 14720
rect 22924 14680 22964 14720
rect 23308 14680 23348 14720
rect 24268 14680 24308 14720
rect 24748 14680 24788 14720
rect 25612 14680 25652 14720
rect 25996 14680 26036 14720
rect 26380 14680 26420 14720
rect 26572 14680 26612 14720
rect 26860 14680 26900 14720
rect 28108 14680 28148 14720
rect 28300 14680 28340 14720
rect 28492 14680 28532 14720
rect 28588 14680 28628 14720
rect 28780 14680 28820 14720
rect 29068 14680 29108 14720
rect 29356 14680 29396 14720
rect 29548 14680 29588 14720
rect 29644 14680 29684 14720
rect 30124 14680 30164 14720
rect 31372 14680 31412 14720
rect 31468 14680 31508 14720
rect 31564 14680 31604 14720
rect 31660 14680 31700 14720
rect 31852 14680 31892 14720
rect 31948 14666 31988 14706
rect 32140 14680 32180 14720
rect 32332 14680 32372 14720
rect 32524 14680 32564 14720
rect 32620 14680 32660 14720
rect 33004 14680 33044 14720
rect 33100 14680 33140 14720
rect 33292 14680 33332 14720
rect 34348 14680 34388 14720
rect 34444 14680 34484 14720
rect 35788 14680 35828 14720
rect 36268 14680 36308 14720
rect 36364 14680 36404 14720
rect 37132 14666 37172 14706
rect 37324 14680 37364 14720
rect 37420 14680 37460 14720
rect 37900 14680 37940 14720
rect 37996 14680 38036 14720
rect 38668 14680 38708 14720
rect 38860 14680 38900 14720
rect 39148 14680 39188 14720
rect 39532 14680 39572 14720
rect 40396 14680 40436 14720
rect 14476 14596 14516 14636
rect 16396 14596 16436 14636
rect 25900 14596 25940 14636
rect 28684 14596 28724 14636
rect 29452 14596 29492 14636
rect 30316 14596 30356 14636
rect 38764 14596 38804 14636
rect 652 14512 692 14552
rect 1036 14512 1076 14552
rect 3148 14512 3188 14552
rect 3724 14512 3764 14552
rect 4876 14512 4916 14552
rect 5740 14512 5780 14552
rect 8140 14512 8180 14552
rect 11788 14512 11828 14552
rect 13708 14512 13748 14552
rect 15340 14512 15380 14552
rect 20524 14512 20564 14552
rect 25132 14512 25172 14552
rect 26668 14512 26708 14552
rect 28204 14512 28244 14552
rect 28972 14512 29012 14552
rect 30028 14512 30068 14552
rect 32044 14512 32084 14552
rect 32812 14512 32852 14552
rect 33964 14512 34004 14552
rect 34156 14512 34196 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 4780 14176 4820 14216
rect 8044 14176 8084 14216
rect 8716 14176 8756 14216
rect 15820 14176 15860 14216
rect 19852 14176 19892 14216
rect 25900 14176 25940 14216
rect 27052 14176 27092 14216
rect 27244 14176 27284 14216
rect 28588 14176 28628 14216
rect 29932 14176 29972 14216
rect 33676 14176 33716 14216
rect 35116 14176 35156 14216
rect 38956 14176 38996 14216
rect 5644 14092 5684 14132
rect 9580 14092 9620 14132
rect 13036 14092 13076 14132
rect 17836 14092 17876 14132
rect 20524 14092 20564 14132
rect 21868 14092 21908 14132
rect 29836 14092 29876 14132
rect 1036 14008 1076 14048
rect 1420 14008 1460 14048
rect 2284 14008 2324 14048
rect 3532 14008 3572 14048
rect 4588 14008 4628 14048
rect 5452 14008 5492 14048
rect 6028 14008 6068 14048
rect 6892 14008 6932 14048
rect 9388 14008 9428 14048
rect 9964 14008 10004 14048
rect 10828 14008 10868 14048
rect 12844 14008 12884 14048
rect 13708 14008 13748 14048
rect 14092 14008 14132 14048
rect 14188 14008 14228 14048
rect 14668 14008 14708 14048
rect 14764 14008 14804 14048
rect 14956 14008 14996 14048
rect 15148 14008 15188 14048
rect 15340 14008 15380 14048
rect 15532 14008 15572 14048
rect 15628 14008 15668 14048
rect 15724 14008 15764 14048
rect 16876 14008 16916 14048
rect 17260 14008 17300 14048
rect 17356 14008 17396 14048
rect 17452 14008 17492 14048
rect 17548 14008 17588 14048
rect 17740 14008 17780 14048
rect 17932 14008 17972 14048
rect 18796 14008 18836 14048
rect 18892 14008 18932 14048
rect 18988 14008 19028 14048
rect 19084 14008 19124 14048
rect 19468 14008 19508 14048
rect 19564 14008 19604 14048
rect 20044 14008 20084 14048
rect 20428 14008 20468 14048
rect 21004 14008 21044 14048
rect 21100 14008 21140 14048
rect 21292 14008 21332 14048
rect 21580 14008 21620 14048
rect 21676 14008 21716 14048
rect 21772 14008 21812 14048
rect 23020 14008 23060 14048
rect 25420 14008 25460 14048
rect 25516 14008 25556 14048
rect 25708 14008 25748 14048
rect 26092 14008 26132 14048
rect 26188 14008 26228 14048
rect 26764 14008 26804 14048
rect 26860 14008 26900 14048
rect 27436 14008 27476 14048
rect 27532 14008 27572 14048
rect 27628 14008 27668 14048
rect 27724 14008 27764 14048
rect 28204 14008 28244 14048
rect 28300 14008 28340 14048
rect 29068 14008 29108 14048
rect 29164 14008 29204 14048
rect 29644 14008 29684 14048
rect 29740 14008 29780 14048
rect 31948 14008 31988 14048
rect 34348 14008 34388 14048
rect 34636 14008 34676 14048
rect 36844 14008 36884 14048
rect 37804 14008 37844 14048
rect 38764 14008 38804 14048
rect 39148 14008 39188 14048
rect 39244 14008 39284 14048
rect 39820 14008 39860 14048
rect 40492 14008 40532 14048
rect 3916 13840 3956 13880
rect 8236 13840 8276 13880
rect 11980 13840 12020 13880
rect 25708 13840 25748 13880
rect 28972 13840 29012 13880
rect 29740 13840 29780 13880
rect 32140 13840 32180 13880
rect 33484 13840 33524 13880
rect 39628 13840 39668 13880
rect 8716 13756 8756 13796
rect 12172 13756 12212 13796
rect 13996 13756 14036 13796
rect 14764 13756 14804 13796
rect 15244 13756 15284 13796
rect 16300 13756 16340 13796
rect 21292 13756 21332 13796
rect 22540 13756 22580 13796
rect 38092 13756 38132 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 5644 13420 5684 13460
rect 6508 13420 6548 13460
rect 9580 13420 9620 13460
rect 13324 13420 13364 13460
rect 14764 13420 14804 13460
rect 15244 13420 15284 13460
rect 16300 13420 16340 13460
rect 27724 13420 27764 13460
rect 29260 13420 29300 13460
rect 36172 13420 36212 13460
rect 10060 13336 10100 13376
rect 12268 13336 12308 13376
rect 26668 13336 26708 13376
rect 28204 13336 28244 13376
rect 30220 13336 30260 13376
rect 31564 13336 31604 13376
rect 39340 13336 39380 13376
rect 11212 13252 11252 13292
rect 24844 13252 24884 13292
rect 26572 13252 26612 13292
rect 26764 13252 26804 13292
rect 3244 13168 3284 13208
rect 3628 13168 3668 13208
rect 4492 13168 4532 13208
rect 5836 13168 5876 13208
rect 6796 13168 6836 13208
rect 7180 13168 7220 13208
rect 7564 13168 7604 13208
rect 8428 13168 8468 13208
rect 12460 13168 12500 13208
rect 13036 13168 13076 13208
rect 13132 13168 13172 13208
rect 13324 13168 13364 13208
rect 13804 13168 13844 13208
rect 13900 13168 13940 13208
rect 14380 13168 14420 13208
rect 14476 13168 14516 13208
rect 14956 13168 14996 13208
rect 15052 13168 15092 13208
rect 15244 13168 15284 13208
rect 15436 13168 15476 13208
rect 15532 13168 15572 13208
rect 15628 13168 15668 13208
rect 16012 13168 16052 13208
rect 16108 13168 16148 13208
rect 16300 13168 16340 13208
rect 16972 13168 17012 13208
rect 17068 13168 17108 13208
rect 17260 13168 17300 13208
rect 17644 13168 17684 13208
rect 17740 13168 17780 13208
rect 17932 13168 17972 13208
rect 18028 13168 18068 13208
rect 18129 13168 18169 13208
rect 19084 13168 19124 13208
rect 19276 13168 19316 13208
rect 19372 13168 19412 13208
rect 19660 13168 19700 13208
rect 19756 13168 19796 13208
rect 19852 13168 19892 13208
rect 20332 13168 20372 13208
rect 20428 13168 20468 13208
rect 21100 13168 21140 13208
rect 21196 13168 21236 13208
rect 21292 13168 21332 13208
rect 21614 13183 21654 13223
rect 21772 13168 21812 13208
rect 21868 13168 21908 13208
rect 22060 13168 22100 13208
rect 22156 13168 22196 13208
rect 22444 13168 22484 13208
rect 22828 13168 22868 13208
rect 23692 13168 23732 13208
rect 26092 13168 26132 13208
rect 26860 13168 26900 13208
rect 17164 13084 17204 13124
rect 26476 13126 26516 13166
rect 27052 13168 27092 13208
rect 27148 13168 27188 13208
rect 27244 13168 27284 13208
rect 27916 13210 27956 13250
rect 27340 13168 27380 13208
rect 27724 13168 27764 13208
rect 28012 13168 28052 13208
rect 28204 13126 28244 13166
rect 28396 13168 28436 13208
rect 28492 13168 28532 13208
rect 28684 13168 28724 13208
rect 28780 13168 28820 13208
rect 28972 13168 29012 13208
rect 29452 13168 29492 13208
rect 29548 13168 29588 13208
rect 29740 13168 29780 13208
rect 29836 13168 29876 13208
rect 30220 13168 30260 13208
rect 30412 13168 30452 13208
rect 30604 13168 30644 13208
rect 30796 13168 30836 13208
rect 31372 13168 31412 13208
rect 31564 13168 31604 13208
rect 31660 13168 31700 13208
rect 32236 13168 32276 13208
rect 32428 13168 32468 13208
rect 32524 13168 32564 13208
rect 32812 13168 32852 13208
rect 33004 13168 33044 13208
rect 33100 13168 33140 13208
rect 33292 13168 33332 13208
rect 33484 13168 33524 13208
rect 33580 13168 33620 13208
rect 33772 13168 33812 13208
rect 34156 13168 34196 13208
rect 35020 13168 35060 13208
rect 36940 13168 36980 13208
rect 37324 13168 37364 13208
rect 38188 13168 38228 13208
rect 19180 13084 19220 13124
rect 28876 13084 28916 13124
rect 652 13000 692 13040
rect 12076 13000 12116 13040
rect 14092 13000 14132 13040
rect 20140 13042 20180 13082
rect 29356 13084 29396 13124
rect 32332 13084 32372 13124
rect 33388 13084 33428 13124
rect 14284 12996 14324 13036
rect 17836 13000 17876 13040
rect 19564 13000 19604 13040
rect 21388 13000 21428 13040
rect 21676 13000 21716 13040
rect 25420 13000 25460 13040
rect 29260 13000 29300 13040
rect 30028 13000 30068 13040
rect 30700 13000 30740 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 652 12664 692 12704
rect 14956 12664 14996 12704
rect 19372 12664 19412 12704
rect 27052 12664 27092 12704
rect 27244 12664 27284 12704
rect 28684 12664 28724 12704
rect 34732 12664 34772 12704
rect 36940 12664 36980 12704
rect 4300 12580 4340 12620
rect 5356 12580 5396 12620
rect 5836 12580 5876 12620
rect 9676 12580 9716 12620
rect 13804 12580 13844 12620
rect 18604 12580 18644 12620
rect 21196 12580 21236 12620
rect 27820 12580 27860 12620
rect 3724 12496 3764 12536
rect 3916 12496 3956 12536
rect 4204 12496 4244 12536
rect 4396 12496 4436 12536
rect 4492 12496 4532 12536
rect 5164 12496 5204 12536
rect 5452 12496 5492 12536
rect 5740 12496 5780 12536
rect 5932 12496 5972 12536
rect 6028 12496 6068 12536
rect 7084 12496 7124 12536
rect 8332 12496 8372 12536
rect 8620 12496 8660 12536
rect 9292 12496 9332 12536
rect 9484 12496 9524 12536
rect 9580 12496 9620 12536
rect 9772 12496 9812 12536
rect 10636 12496 10676 12536
rect 12652 12496 12692 12536
rect 13228 12496 13268 12536
rect 13324 12496 13364 12536
rect 13420 12496 13460 12536
rect 13516 12496 13556 12536
rect 13708 12496 13748 12536
rect 13900 12496 13940 12536
rect 13996 12496 14036 12536
rect 14380 12496 14420 12536
rect 14668 12496 14708 12536
rect 14764 12496 14804 12536
rect 14860 12496 14900 12536
rect 15436 12496 15476 12536
rect 15724 12496 15764 12536
rect 3820 12412 3860 12452
rect 11596 12412 11636 12452
rect 15532 12454 15572 12494
rect 15916 12496 15956 12536
rect 16012 12496 16052 12536
rect 16204 12496 16244 12536
rect 16396 12496 16436 12536
rect 16588 12496 16628 12536
rect 16684 12496 16724 12536
rect 18316 12496 18356 12536
rect 18412 12496 18452 12536
rect 18508 12517 18548 12557
rect 18796 12496 18836 12536
rect 18988 12496 19028 12536
rect 19084 12496 19124 12536
rect 19367 12496 19407 12536
rect 19468 12496 19508 12536
rect 19564 12496 19604 12536
rect 19756 12496 19796 12536
rect 19852 12496 19892 12536
rect 20044 12496 20084 12536
rect 20140 12496 20180 12536
rect 20236 12496 20276 12536
rect 20332 12496 20372 12536
rect 20620 12496 20660 12536
rect 20716 12496 20756 12536
rect 20812 12496 20852 12536
rect 20908 12496 20948 12536
rect 21100 12496 21140 12536
rect 21292 12496 21332 12536
rect 21388 12496 21428 12536
rect 21580 12496 21620 12536
rect 24748 12496 24788 12536
rect 25612 12496 25652 12536
rect 25996 12496 26036 12536
rect 26380 12496 26420 12536
rect 26668 12496 26708 12536
rect 26860 12496 26900 12536
rect 15340 12412 15380 12452
rect 26092 12412 26132 12452
rect 26764 12454 26804 12494
rect 27436 12496 27476 12536
rect 27532 12496 27572 12536
rect 27724 12496 27764 12536
rect 27916 12496 27956 12536
rect 28396 12496 28436 12536
rect 28876 12496 28916 12536
rect 28972 12496 29012 12536
rect 29164 12496 29204 12536
rect 29356 12538 29396 12578
rect 35500 12580 35540 12620
rect 36268 12580 36308 12620
rect 29548 12496 29588 12536
rect 29932 12496 29972 12536
rect 30028 12496 30068 12536
rect 30124 12496 30164 12536
rect 30220 12496 30260 12536
rect 32044 12496 32084 12536
rect 33292 12496 33332 12536
rect 34444 12496 34484 12536
rect 34540 12496 34580 12536
rect 35404 12496 35444 12536
rect 35692 12496 35732 12536
rect 35788 12496 35828 12536
rect 35980 12496 36020 12536
rect 36364 12496 36404 12536
rect 36748 12496 36788 12536
rect 37612 12496 37652 12536
rect 39052 12496 39092 12536
rect 26284 12412 26324 12452
rect 29260 12412 29300 12452
rect 29452 12412 29492 12452
rect 4684 12328 4724 12368
rect 6220 12328 6260 12368
rect 6604 12328 6644 12368
rect 6988 12328 7028 12368
rect 7468 12328 7508 12368
rect 10828 12328 10868 12368
rect 14188 12328 14228 12368
rect 14380 12328 14420 12368
rect 15148 12328 15188 12368
rect 15244 12328 15284 12368
rect 16204 12328 16244 12368
rect 22924 12328 22964 12368
rect 26188 12328 26228 12368
rect 28492 12328 28532 12368
rect 29740 12328 29780 12368
rect 33580 12328 33620 12368
rect 7660 12244 7700 12284
rect 9964 12244 10004 12284
rect 11788 12244 11828 12284
rect 11980 12244 12020 12284
rect 15724 12244 15764 12284
rect 18796 12244 18836 12284
rect 22252 12244 22292 12284
rect 32332 12244 32372 12284
rect 33772 12244 33812 12284
rect 35980 12244 36020 12284
rect 38380 12244 38420 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 8428 11908 8468 11948
rect 13708 11908 13748 11948
rect 17836 11908 17876 11948
rect 31084 11908 31124 11948
rect 33196 11908 33236 11948
rect 33964 11908 34004 11948
rect 21196 11824 21236 11864
rect 32716 11824 32756 11864
rect 33484 11824 33524 11864
rect 35020 11824 35060 11864
rect 33580 11782 33620 11822
rect 8812 11740 8852 11780
rect 15532 11740 15572 11780
rect 19276 11740 19316 11780
rect 34924 11740 34964 11780
rect 35116 11740 35156 11780
rect 6028 11656 6068 11696
rect 6412 11656 6452 11696
rect 7276 11656 7316 11696
rect 9580 11656 9620 11696
rect 10060 11656 10100 11696
rect 10444 11656 10484 11696
rect 11308 11656 11348 11696
rect 12844 11656 12884 11696
rect 13708 11656 13748 11696
rect 13900 11656 13940 11696
rect 13996 11656 14036 11696
rect 14476 11656 14516 11696
rect 14572 11656 14612 11696
rect 14668 11656 14708 11696
rect 14764 11656 14804 11696
rect 15244 11656 15284 11696
rect 15340 11656 15380 11696
rect 15724 11656 15764 11696
rect 15916 11656 15956 11696
rect 16300 11656 16340 11696
rect 16396 11656 16436 11696
rect 16588 11656 16628 11696
rect 16684 11656 16724 11696
rect 17836 11656 17876 11696
rect 17932 11656 17972 11696
rect 18076 11660 18116 11700
rect 18220 11656 18260 11696
rect 18377 11671 18417 11711
rect 19660 11656 19700 11696
rect 19756 11656 19796 11696
rect 19948 11656 19988 11696
rect 20044 11656 20084 11696
rect 20201 11671 20241 11711
rect 21772 11656 21812 11696
rect 22156 11656 22196 11696
rect 23020 11656 23060 11696
rect 24364 11656 24404 11696
rect 25801 11645 25841 11685
rect 25900 11656 25940 11696
rect 26092 11656 26132 11696
rect 26188 11656 26228 11696
rect 26284 11656 26324 11696
rect 26380 11656 26420 11696
rect 26572 11656 26612 11696
rect 26668 11656 26708 11696
rect 26764 11656 26804 11696
rect 26860 11656 26900 11696
rect 27052 11656 27092 11696
rect 27148 11656 27188 11696
rect 27244 11656 27284 11696
rect 27340 11656 27380 11696
rect 28972 11656 29012 11696
rect 29068 11656 29108 11696
rect 29164 11656 29204 11696
rect 29260 11656 29300 11696
rect 29644 11656 29684 11696
rect 29740 11656 29780 11696
rect 30124 11656 30164 11696
rect 30220 11656 30260 11696
rect 30412 11656 30452 11696
rect 31372 11656 31412 11696
rect 32332 11656 32372 11696
rect 32524 11656 32564 11696
rect 32716 11656 32756 11696
rect 32908 11656 32948 11696
rect 33196 11656 33236 11696
rect 33676 11656 33716 11696
rect 33772 11656 33812 11696
rect 33964 11656 34004 11696
rect 34252 11656 34292 11696
rect 34828 11656 34868 11696
rect 36076 11656 36116 11696
rect 36268 11656 36308 11696
rect 36940 11656 36980 11696
rect 15820 11572 15860 11612
rect 35212 11614 35252 11654
rect 37132 11656 37172 11696
rect 37516 11656 37556 11696
rect 38380 11656 38420 11696
rect 39532 11656 39572 11696
rect 652 11488 692 11528
rect 12460 11488 12500 11528
rect 13516 11488 13556 11528
rect 16108 11488 16148 11528
rect 16876 11488 16916 11528
rect 19852 11488 19892 11528
rect 24172 11488 24212 11528
rect 25036 11488 25076 11528
rect 29452 11488 29492 11528
rect 29932 11488 29972 11528
rect 32236 11488 32276 11528
rect 33676 11488 33716 11528
rect 35404 11488 35444 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 652 11152 692 11192
rect 16300 11156 16340 11196
rect 17260 11152 17300 11192
rect 25708 11152 25748 11192
rect 25996 11152 26036 11192
rect 28780 11152 28820 11192
rect 29356 11152 29396 11192
rect 30028 11152 30068 11192
rect 31468 11152 31508 11192
rect 34444 11152 34484 11192
rect 9676 11068 9716 11108
rect 27340 11068 27380 11108
rect 8428 10984 8468 11024
rect 9292 10984 9332 11024
rect 10060 10984 10100 11024
rect 10156 10984 10196 11024
rect 10348 10984 10388 11024
rect 10540 10984 10580 11024
rect 11404 10984 11444 11024
rect 11500 10984 11540 11024
rect 11596 10984 11636 11024
rect 11692 10984 11732 11024
rect 12460 10984 12500 11024
rect 12652 10984 12692 11024
rect 13900 10984 13940 11024
rect 14860 10984 14900 11024
rect 14956 10984 14996 11024
rect 16204 10984 16244 11024
rect 16967 10984 17007 11024
rect 17068 10984 17108 11024
rect 16108 10942 16148 10982
rect 17164 10984 17204 11024
rect 17356 10984 17396 11024
rect 17452 10984 17492 11024
rect 17644 10984 17684 11024
rect 18508 10984 18548 11024
rect 18892 10984 18932 11024
rect 18988 10984 19028 11024
rect 19180 10984 19220 11024
rect 19276 10984 19316 11024
rect 19377 10984 19417 11024
rect 19852 10984 19892 11024
rect 20812 10984 20852 11024
rect 21676 10984 21716 11024
rect 21868 10984 21908 11024
rect 22060 10984 22100 11024
rect 22156 10984 22196 11024
rect 23692 10984 23732 11024
rect 23788 10984 23828 11024
rect 24172 10984 24212 11024
rect 25036 10984 25076 11024
rect 25804 10984 25844 11024
rect 26092 10984 26132 11024
rect 26188 10984 26228 11024
rect 26284 10984 26324 11024
rect 26476 10984 26516 11024
rect 26668 10984 26708 11024
rect 26860 11005 26900 11045
rect 27052 10984 27092 11024
rect 27244 10984 27284 11024
rect 27436 10984 27476 11024
rect 28684 10984 28724 11024
rect 28876 10984 28916 11024
rect 29068 10984 29108 11024
rect 29164 10984 29204 11024
rect 29548 10984 29588 11024
rect 29260 10942 29300 10982
rect 29740 10984 29780 11024
rect 29644 10942 29684 10982
rect 29836 10984 29876 11024
rect 30220 10984 30260 11024
rect 30316 10984 30356 11024
rect 30508 10984 30548 11024
rect 30700 10984 30740 11024
rect 31180 10984 31220 11024
rect 31276 10984 31316 11024
rect 31468 10984 31508 11024
rect 31564 10984 31604 11024
rect 31665 10984 31705 11024
rect 32428 10984 32468 11024
rect 32716 10984 32756 11024
rect 33100 10984 33140 11024
rect 34348 10984 34388 11024
rect 34732 10984 34772 11024
rect 34828 10984 34868 11024
rect 34924 10984 34964 11024
rect 35020 10984 35060 11024
rect 35404 10984 35444 11024
rect 35788 10984 35828 11024
rect 36652 10984 36692 11024
rect 37804 10984 37844 11024
rect 38092 10984 38132 11024
rect 38764 10984 38804 11024
rect 15244 10900 15284 10940
rect 15628 10900 15668 10940
rect 23308 10900 23348 10940
rect 30604 10900 30644 10940
rect 32812 10900 32852 10940
rect 33004 10900 33044 10940
rect 10348 10816 10388 10856
rect 11884 10816 11924 10856
rect 13228 10816 13268 10856
rect 13612 10816 13652 10856
rect 18316 10816 18356 10856
rect 22348 10816 22388 10856
rect 26476 10816 26516 10856
rect 32524 10816 32564 10856
rect 32908 10816 32948 10856
rect 7276 10732 7316 10772
rect 11212 10732 11252 10772
rect 15436 10732 15476 10772
rect 15820 10732 15860 10772
rect 18892 10732 18932 10772
rect 20140 10732 20180 10772
rect 21004 10732 21044 10772
rect 21868 10732 21908 10772
rect 23500 10732 23540 10772
rect 24460 10732 24500 10772
rect 26956 10732 26996 10772
rect 35212 10732 35252 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 13516 10396 13556 10436
rect 26668 10396 26708 10436
rect 29356 10396 29396 10436
rect 30988 10396 31028 10436
rect 31276 10396 31316 10436
rect 32716 10396 32756 10436
rect 34636 10396 34676 10436
rect 35020 10396 35060 10436
rect 35308 10396 35348 10436
rect 6028 10312 6068 10352
rect 6796 10312 6836 10352
rect 9004 10312 9044 10352
rect 9964 10312 10004 10352
rect 23116 10312 23156 10352
rect 29164 10312 29204 10352
rect 20332 10228 20372 10268
rect 25132 10228 25172 10268
rect 7660 10144 7700 10184
rect 7852 10144 7892 10184
rect 9676 10144 9716 10184
rect 11116 10144 11156 10184
rect 11980 10144 12020 10184
rect 12364 10144 12404 10184
rect 12556 10144 12596 10184
rect 13228 10144 13268 10184
rect 13420 10144 13460 10184
rect 14668 10144 14708 10184
rect 15628 10144 15668 10184
rect 16108 10144 16148 10184
rect 16204 10144 16244 10184
rect 16396 10144 16436 10184
rect 16588 10144 16628 10184
rect 16780 10144 16820 10184
rect 16876 10144 16916 10184
rect 17068 10144 17108 10184
rect 18316 10144 18356 10184
rect 19180 10144 19220 10184
rect 20716 10144 20756 10184
rect 21100 10144 21140 10184
rect 21964 10144 22004 10184
rect 23308 10144 23348 10184
rect 24364 10144 24404 10184
rect 24460 10144 24500 10184
rect 24652 10144 24692 10184
rect 24748 10144 24788 10184
rect 24940 10144 24980 10184
rect 26188 10144 26228 10184
rect 26284 10144 26324 10184
rect 26380 10144 26420 10184
rect 26476 10144 26516 10184
rect 26668 10144 26708 10184
rect 26764 10144 26804 10184
rect 26956 10144 26996 10184
rect 27052 10144 27092 10184
rect 27153 10144 27193 10184
rect 28876 10144 28916 10184
rect 29068 10144 29108 10184
rect 29164 10144 29204 10184
rect 29356 10144 29396 10184
rect 29452 10144 29492 10184
rect 29644 10144 29684 10184
rect 29841 10144 29881 10184
rect 30124 10144 30164 10184
rect 6988 10060 7028 10100
rect 16684 10060 16724 10100
rect 17740 10060 17780 10100
rect 17932 10060 17972 10100
rect 23980 10060 24020 10100
rect 24844 10060 24884 10100
rect 29740 10102 29780 10142
rect 30412 10144 30452 10184
rect 30796 10144 30836 10184
rect 30995 10157 31035 10197
rect 31180 10144 31220 10184
rect 31372 10144 31412 10184
rect 32140 10144 32180 10184
rect 32236 10144 32276 10184
rect 32332 10144 32372 10184
rect 32428 10144 32468 10184
rect 32620 10144 32660 10184
rect 32812 10144 32852 10184
rect 33100 10144 33140 10184
rect 34444 10144 34484 10184
rect 34828 10144 34868 10184
rect 35020 10144 35060 10184
rect 35116 10144 35156 10184
rect 35308 10144 35348 10184
rect 35500 10144 35540 10184
rect 35596 10144 35636 10184
rect 35788 10144 35828 10184
rect 36076 10144 36116 10184
rect 36556 10144 36596 10184
rect 37228 10144 37268 10184
rect 37420 10144 37460 10184
rect 37804 10144 37844 10184
rect 38668 10144 38708 10184
rect 39820 10144 39860 10184
rect 30316 10060 30356 10100
rect 33004 10060 33044 10100
rect 36268 10060 36308 10100
rect 652 9976 692 10016
rect 8524 9976 8564 10016
rect 16396 9976 16436 10016
rect 24172 9976 24212 10016
rect 25324 9976 25364 10016
rect 34348 9976 34388 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 652 9640 692 9680
rect 9484 9640 9524 9680
rect 10060 9640 10100 9680
rect 11020 9640 11060 9680
rect 11500 9640 11540 9680
rect 13324 9640 13364 9680
rect 27340 9640 27380 9680
rect 27820 9640 27860 9680
rect 28204 9640 28244 9680
rect 29548 9640 29588 9680
rect 30604 9640 30644 9680
rect 32140 9640 32180 9680
rect 33196 9640 33236 9680
rect 35212 9640 35252 9680
rect 35596 9640 35636 9680
rect 35884 9640 35924 9680
rect 38188 9640 38228 9680
rect 5548 9556 5588 9596
rect 13804 9556 13844 9596
rect 24844 9556 24884 9596
rect 5932 9472 5972 9512
rect 6796 9472 6836 9512
rect 8140 9472 8180 9512
rect 8236 9472 8276 9512
rect 8428 9472 8468 9512
rect 9100 9472 9140 9512
rect 9292 9472 9332 9512
rect 9388 9472 9428 9512
rect 9580 9472 9620 9512
rect 9868 9472 9908 9512
rect 9964 9472 10004 9512
rect 10156 9472 10196 9512
rect 10348 9472 10388 9512
rect 10444 9472 10484 9512
rect 11116 9472 11156 9512
rect 11212 9472 11252 9512
rect 11308 9472 11348 9512
rect 11596 9472 11636 9512
rect 11692 9472 11732 9512
rect 11788 9472 11828 9512
rect 12652 9472 12692 9512
rect 12844 9472 12884 9512
rect 13036 9472 13076 9512
rect 13132 9472 13172 9512
rect 13420 9472 13460 9512
rect 13516 9472 13556 9512
rect 13612 9472 13652 9512
rect 13900 9472 13940 9512
rect 13996 9472 14036 9512
rect 14092 9472 14132 9512
rect 14284 9472 14324 9512
rect 14380 9472 14420 9512
rect 14572 9472 14612 9512
rect 14764 9472 14804 9512
rect 14860 9472 14900 9512
rect 14956 9472 14996 9512
rect 15052 9472 15092 9512
rect 15244 9472 15284 9512
rect 15340 9472 15380 9512
rect 15436 9472 15476 9512
rect 15532 9472 15572 9512
rect 15724 9493 15764 9533
rect 15820 9472 15860 9512
rect 15916 9472 15956 9512
rect 16012 9472 16052 9512
rect 16204 9472 16244 9512
rect 16300 9472 16340 9512
rect 16492 9472 16532 9512
rect 16972 9472 17012 9512
rect 17164 9472 17204 9512
rect 17260 9472 17300 9512
rect 17548 9472 17588 9512
rect 21100 9472 21140 9512
rect 21484 9472 21524 9512
rect 21676 9472 21716 9512
rect 22444 9472 22484 9512
rect 23692 9472 23732 9512
rect 24076 9472 24116 9512
rect 24172 9472 24212 9512
rect 24268 9472 24308 9512
rect 24364 9472 24404 9512
rect 24556 9472 24596 9512
rect 24652 9472 24692 9512
rect 24748 9472 24788 9512
rect 25228 9472 25268 9512
rect 27244 9472 27284 9512
rect 27436 9472 27476 9512
rect 27532 9472 27572 9512
rect 27916 9472 27956 9512
rect 28300 9472 28340 9512
rect 28396 9472 28436 9512
rect 28492 9472 28532 9512
rect 28684 9472 28724 9512
rect 28780 9472 28820 9512
rect 28876 9472 28916 9512
rect 28972 9472 29012 9512
rect 29255 9472 29295 9512
rect 29356 9472 29396 9512
rect 29452 9472 29492 9512
rect 29644 9472 29684 9512
rect 29740 9472 29780 9512
rect 29932 9472 29972 9512
rect 30316 9472 30356 9512
rect 30508 9472 30548 9512
rect 30700 9472 30740 9512
rect 31852 9472 31892 9512
rect 31948 9472 31988 9512
rect 32044 9472 32084 9512
rect 32620 9472 32660 9512
rect 32908 9472 32948 9512
rect 33004 9472 33044 9512
rect 33100 9472 33140 9512
rect 34252 9472 34292 9512
rect 34444 9472 34484 9512
rect 34636 9472 34676 9512
rect 34732 9472 34772 9512
rect 34924 9472 34964 9512
rect 35116 9472 35156 9512
rect 35212 9472 35252 9512
rect 35692 9472 35732 9512
rect 36268 9472 36308 9512
rect 37324 9472 37364 9512
rect 37996 9472 38036 9512
rect 38860 9472 38900 9512
rect 7948 9388 7988 9428
rect 22828 9388 22868 9428
rect 30028 9388 30068 9428
rect 30220 9388 30260 9428
rect 3916 9304 3956 9344
rect 12844 9304 12884 9344
rect 16492 9304 16532 9344
rect 18700 9304 18740 9344
rect 20908 9304 20948 9344
rect 23404 9304 23444 9344
rect 30124 9304 30164 9344
rect 11980 9220 12020 9260
rect 14572 9220 14612 9260
rect 16972 9220 17012 9260
rect 18220 9220 18260 9260
rect 22540 9220 22580 9260
rect 25324 9220 25364 9260
rect 32716 9220 32756 9260
rect 34156 9220 34196 9260
rect 34444 9220 34484 9260
rect 35884 9220 35924 9260
rect 36940 9220 36980 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 16300 8884 16340 8924
rect 24172 8884 24212 8924
rect 6124 8800 6164 8840
rect 18028 8800 18068 8840
rect 19756 8800 19796 8840
rect 24844 8842 24884 8882
rect 31468 8884 31508 8924
rect 32140 8884 32180 8924
rect 39052 8884 39092 8924
rect 26380 8800 26420 8840
rect 27148 8800 27188 8840
rect 30028 8800 30068 8840
rect 32524 8800 32564 8840
rect 35596 8800 35636 8840
rect 13420 8716 13460 8756
rect 24748 8716 24788 8756
rect 24940 8716 24980 8756
rect 32428 8716 32468 8756
rect 3436 8632 3476 8672
rect 3820 8632 3860 8672
rect 4684 8632 4724 8672
rect 5932 8632 5972 8672
rect 6124 8632 6164 8672
rect 6316 8632 6356 8672
rect 7084 8632 7124 8672
rect 7948 8632 7988 8672
rect 9484 8632 9524 8672
rect 10348 8632 10388 8672
rect 10444 8632 10484 8672
rect 10636 8632 10676 8672
rect 11020 8632 11060 8672
rect 11404 8632 11444 8672
rect 12268 8632 12308 8672
rect 14284 8632 14324 8672
rect 14764 8632 14804 8672
rect 14860 8632 14900 8672
rect 14956 8632 14996 8672
rect 15820 8632 15860 8672
rect 16012 8632 16052 8672
rect 16108 8632 16148 8672
rect 16300 8632 16340 8672
rect 16684 8632 16724 8672
rect 16780 8632 16820 8672
rect 16876 8632 16916 8672
rect 16972 8632 17012 8672
rect 17164 8632 17204 8672
rect 21004 8632 21044 8672
rect 22060 8632 22100 8672
rect 22348 8632 22388 8672
rect 23116 8632 23156 8672
rect 23212 8632 23252 8672
rect 23404 8632 23444 8672
rect 23500 8632 23540 8672
rect 23884 8632 23924 8672
rect 23980 8632 24020 8672
rect 24172 8632 24212 8672
rect 24652 8632 24692 8672
rect 25036 8632 25076 8672
rect 25324 8632 25364 8672
rect 25708 8674 25748 8714
rect 32620 8716 32660 8756
rect 34156 8716 34196 8756
rect 25612 8632 25652 8672
rect 25804 8632 25844 8672
rect 26092 8632 26132 8672
rect 26380 8632 26420 8672
rect 26572 8632 26612 8672
rect 26764 8632 26804 8672
rect 26860 8632 26900 8672
rect 27052 8632 27092 8672
rect 27148 8632 27188 8672
rect 27340 8632 27380 8672
rect 28780 8632 28820 8672
rect 29068 8632 29108 8672
rect 29164 8632 29204 8672
rect 29740 8632 29780 8672
rect 29836 8632 29876 8672
rect 30124 8632 30164 8672
rect 31084 8632 31124 8672
rect 31372 8632 31412 8672
rect 31468 8632 31508 8672
rect 31660 8632 31700 8672
rect 31852 8632 31892 8672
rect 31948 8632 31988 8672
rect 32140 8632 32180 8672
rect 32332 8632 32372 8672
rect 32716 8632 32756 8672
rect 32908 8632 32948 8672
rect 33004 8632 33044 8672
rect 33484 8632 33524 8672
rect 33676 8629 33716 8669
rect 33964 8632 34004 8672
rect 34252 8632 34292 8672
rect 34444 8632 34484 8672
rect 34636 8632 34676 8672
rect 34732 8657 34772 8697
rect 35308 8632 35348 8672
rect 35404 8632 35444 8672
rect 35596 8632 35636 8672
rect 35788 8632 35828 8672
rect 36460 8632 36500 8672
rect 36652 8632 36692 8672
rect 37036 8632 37076 8672
rect 37900 8632 37940 8672
rect 6700 8548 6740 8588
rect 652 8464 692 8504
rect 9100 8464 9140 8504
rect 10156 8464 10196 8504
rect 10540 8464 10580 8504
rect 13612 8464 13652 8504
rect 14668 8464 14708 8504
rect 15148 8464 15188 8504
rect 17836 8464 17876 8504
rect 20620 8464 20660 8504
rect 22252 8464 22292 8504
rect 22924 8464 22964 8504
rect 23692 8464 23732 8504
rect 25228 8464 25268 8504
rect 25900 8464 25940 8504
rect 26668 8464 26708 8504
rect 28876 8464 28916 8504
rect 29356 8464 29396 8504
rect 29548 8464 29588 8504
rect 31180 8464 31220 8504
rect 33196 8464 33236 8504
rect 34732 8422 34772 8462
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 652 8128 692 8168
rect 5644 8128 5684 8168
rect 8236 8128 8276 8168
rect 9292 8128 9332 8168
rect 13036 8128 13076 8168
rect 13612 8128 13652 8168
rect 14476 8128 14516 8168
rect 17356 8128 17396 8168
rect 20908 8128 20948 8168
rect 22828 8128 22868 8168
rect 23404 8128 23444 8168
rect 26572 8128 26612 8168
rect 26956 8128 26996 8168
rect 28396 8128 28436 8168
rect 30220 8128 30260 8168
rect 30796 8128 30836 8168
rect 32140 8128 32180 8168
rect 32716 8128 32756 8168
rect 34636 8128 34676 8168
rect 35692 8128 35732 8168
rect 14956 8044 14996 8084
rect 17548 8044 17588 8084
rect 28876 8044 28916 8084
rect 31852 8044 31892 8084
rect 4492 7960 4532 8000
rect 4684 7960 4724 8000
rect 4876 7960 4916 8000
rect 4972 7960 5012 8000
rect 5164 7960 5204 8000
rect 5260 7960 5300 8000
rect 5356 7960 5396 8000
rect 5452 7960 5492 8000
rect 5740 7960 5780 8000
rect 5836 7960 5876 8000
rect 5932 7960 5972 8000
rect 7468 7960 7508 8000
rect 7564 7960 7604 8000
rect 7756 7960 7796 8000
rect 8044 7960 8084 8000
rect 8908 7960 8948 8000
rect 9100 7960 9140 8000
rect 9196 7960 9236 8000
rect 9388 7960 9428 8000
rect 9484 7960 9524 8000
rect 9639 7960 9679 8000
rect 9964 7960 10004 8000
rect 10156 7960 10196 8000
rect 11788 7960 11828 8000
rect 12652 7960 12692 8000
rect 13132 7960 13172 8000
rect 13996 7960 14036 8000
rect 14092 7960 14132 8000
rect 14188 7960 14228 8000
rect 14284 7960 14324 8000
rect 14572 7960 14612 8000
rect 14668 7960 14708 8000
rect 14764 7960 14804 8000
rect 15340 7960 15380 8000
rect 16204 7960 16244 8000
rect 17932 7960 17972 8000
rect 18796 7960 18836 8000
rect 20236 7960 20276 8000
rect 21196 7960 21236 8000
rect 21484 7960 21524 8000
rect 21676 7960 21716 8000
rect 22540 7960 22580 8000
rect 22636 7960 22676 8000
rect 23212 7960 23252 8000
rect 23500 7960 23540 8000
rect 23788 7951 23828 7991
rect 24076 7960 24116 8000
rect 24748 7960 24788 8000
rect 25036 7960 25076 8000
rect 25228 7960 25268 8000
rect 25324 7960 25364 8000
rect 25516 7960 25556 8000
rect 25612 7960 25652 8000
rect 25767 7960 25807 8000
rect 26380 7960 26420 8000
rect 26668 7960 26708 8000
rect 27148 7960 27188 8000
rect 27436 7960 27476 8000
rect 28108 7960 28148 8000
rect 28204 7960 28244 8000
rect 28300 7960 28340 8000
rect 28588 7960 28628 8000
rect 28684 7960 28724 8000
rect 28780 7960 28820 8000
rect 29068 7960 29108 8000
rect 29452 7960 29492 8000
rect 29740 7960 29780 8000
rect 29836 7960 29876 8000
rect 30028 7960 30068 8000
rect 30124 7960 30164 8000
rect 30281 7945 30321 7985
rect 30508 7960 30548 8000
rect 30604 7960 30644 8000
rect 30700 7960 30740 8000
rect 31084 7960 31124 8000
rect 31468 7960 31508 8000
rect 31756 7960 31796 8000
rect 31948 7960 31988 8000
rect 32332 7960 32372 8000
rect 32428 7960 32468 8000
rect 32620 7960 32660 8000
rect 32908 7960 32948 8000
rect 33292 7960 33332 8000
rect 33484 7960 33524 8000
rect 33580 7960 33620 8000
rect 33772 7960 33812 8000
rect 33964 7960 34004 8000
rect 34828 7960 34868 8000
rect 36364 7960 36404 8000
rect 36556 7960 36596 8000
rect 36940 7960 36980 8000
rect 37804 7960 37844 8000
rect 6124 7901 6164 7941
rect 13804 7876 13844 7916
rect 19948 7876 19988 7916
rect 24940 7876 24980 7916
rect 29164 7876 29204 7916
rect 29356 7876 29396 7916
rect 31180 7876 31220 7916
rect 31372 7876 31412 7916
rect 2860 7792 2900 7832
rect 4684 7792 4724 7832
rect 9868 7792 9908 7832
rect 11404 7792 11444 7832
rect 29260 7792 29300 7832
rect 31276 7792 31316 7832
rect 33772 7792 33812 7832
rect 3820 7708 3860 7748
rect 6796 7708 6836 7748
rect 7756 7708 7796 7748
rect 10252 7708 10292 7748
rect 21484 7708 21524 7748
rect 22348 7708 22388 7748
rect 24076 7708 24116 7748
rect 25228 7708 25268 7748
rect 33196 7708 33236 7748
rect 35500 7708 35540 7748
rect 38956 7708 38996 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4780 7372 4820 7412
rect 5836 7372 5876 7412
rect 6988 7372 7028 7412
rect 8140 7372 8180 7412
rect 13036 7372 13076 7412
rect 22060 7372 22100 7412
rect 24172 7372 24212 7412
rect 26668 7372 26708 7412
rect 31180 7372 31220 7412
rect 31564 7372 31604 7412
rect 33772 7372 33812 7412
rect 36556 7372 36596 7412
rect 37420 7372 37460 7412
rect 10060 7288 10100 7328
rect 14476 7288 14516 7328
rect 15436 7288 15476 7328
rect 16492 7288 16532 7328
rect 29260 7288 29300 7328
rect 10732 7204 10772 7244
rect 14380 7204 14420 7244
rect 29644 7204 29684 7244
rect 2380 7120 2420 7160
rect 2764 7120 2804 7160
rect 3628 7120 3668 7160
rect 5164 7120 5204 7160
rect 6220 7120 6260 7160
rect 6508 7120 6548 7160
rect 7468 7120 7508 7160
rect 7852 7120 7892 7160
rect 8140 7120 8180 7160
rect 8332 7120 8372 7160
rect 8428 7120 8468 7160
rect 8812 7120 8852 7160
rect 8908 7120 8948 7160
rect 9100 7120 9140 7160
rect 9196 7120 9236 7160
rect 9297 7120 9337 7160
rect 9676 7120 9716 7160
rect 9772 7120 9812 7160
rect 10252 7120 10292 7160
rect 10348 7120 10388 7160
rect 11308 7120 11348 7160
rect 11404 7120 11444 7160
rect 11788 7120 11828 7160
rect 11884 7120 11924 7160
rect 12364 7120 12404 7160
rect 13612 7120 13652 7160
rect 14188 7120 14228 7160
rect 14284 7120 14324 7160
rect 14764 7120 14804 7160
rect 15052 7120 15092 7160
rect 15628 7120 15668 7160
rect 17548 7120 17588 7160
rect 17836 7120 17876 7160
rect 18988 7120 19028 7160
rect 19372 7120 19412 7160
rect 20236 7120 20276 7160
rect 22444 7120 22484 7160
rect 22924 7120 22964 7160
rect 23020 7120 23060 7160
rect 23212 7120 23252 7160
rect 23308 7120 23348 7160
rect 23465 7135 23505 7175
rect 23692 7120 23732 7160
rect 23788 7120 23828 7160
rect 24172 7120 24212 7160
rect 24268 7120 24308 7160
rect 24460 7120 24500 7160
rect 24556 7120 24596 7160
rect 24713 7135 24753 7175
rect 25228 7120 25268 7160
rect 25420 7120 25460 7160
rect 25516 7120 25556 7160
rect 25900 7120 25940 7160
rect 25996 7120 26036 7160
rect 26188 7120 26228 7160
rect 26284 7120 26324 7160
rect 26380 7120 26420 7160
rect 26668 7120 26708 7160
rect 26764 7120 26804 7160
rect 26956 7120 26996 7160
rect 27052 7120 27092 7160
rect 27207 7120 27247 7160
rect 28012 7120 28052 7160
rect 28108 7120 28148 7160
rect 28204 7120 28244 7160
rect 28684 7120 28724 7160
rect 28780 7120 28820 7160
rect 28972 7120 29012 7160
rect 29260 7120 29300 7160
rect 29452 7120 29492 7160
rect 29740 7120 29780 7160
rect 30124 7120 30164 7160
rect 30220 7120 30260 7160
rect 31276 7120 31316 7160
rect 31660 7120 31700 7160
rect 32524 7120 32564 7160
rect 34924 7120 34964 7160
rect 35788 7120 35828 7160
rect 36172 7120 36212 7160
rect 37228 7120 37268 7160
rect 38092 7120 38132 7160
rect 652 6952 692 6992
rect 5836 6952 5876 6992
rect 6028 6952 6068 6992
rect 6316 6952 6356 6992
rect 8044 6952 8084 6992
rect 8620 6952 8660 6992
rect 9292 6952 9332 6992
rect 9580 6948 9620 6988
rect 10540 6952 10580 6992
rect 11596 6952 11636 6992
rect 12076 6952 12116 6992
rect 13516 6952 13556 6992
rect 13804 6952 13844 6992
rect 14284 6952 14324 6992
rect 14956 6952 14996 6992
rect 16300 6952 16340 6992
rect 16876 6952 16916 6992
rect 17740 6952 17780 6992
rect 21388 6952 21428 6992
rect 23404 6952 23444 6992
rect 23980 6952 24020 6992
rect 25708 6952 25748 6992
rect 26476 6952 26516 6992
rect 28300 6952 28340 6992
rect 28492 6952 28532 6992
rect 29932 6952 29972 6992
rect 31852 6952 31892 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 15052 6674 15092 6714
rect 8428 6616 8468 6656
rect 8716 6616 8756 6656
rect 10060 6616 10100 6656
rect 12364 6616 12404 6656
rect 13132 6616 13172 6656
rect 13228 6616 13268 6656
rect 14188 6616 14228 6656
rect 15340 6616 15380 6656
rect 22156 6616 22196 6656
rect 23116 6616 23156 6656
rect 23500 6616 23540 6656
rect 23884 6616 23924 6656
rect 24460 6616 24500 6656
rect 25996 6616 26036 6656
rect 26572 6616 26612 6656
rect 27148 6616 27188 6656
rect 28300 6616 28340 6656
rect 35308 6616 35348 6656
rect 9964 6532 10004 6572
rect 13036 6532 13076 6572
rect 15724 6532 15764 6572
rect 21868 6532 21908 6572
rect 25900 6532 25940 6572
rect 26476 6532 26516 6572
rect 29932 6532 29972 6572
rect 3724 6448 3764 6488
rect 4108 6448 4148 6488
rect 4972 6448 5012 6488
rect 6220 6448 6260 6488
rect 6412 6435 6452 6475
rect 7468 6448 7508 6488
rect 7564 6448 7604 6488
rect 7660 6448 7700 6488
rect 7756 6448 7796 6488
rect 8236 6448 8276 6488
rect 8524 6448 8564 6488
rect 8908 6448 8948 6488
rect 9004 6448 9044 6488
rect 9196 6448 9236 6488
rect 9292 6448 9332 6488
rect 9772 6448 9812 6488
rect 9868 6448 9908 6488
rect 10348 6448 10388 6488
rect 10540 6448 10580 6488
rect 10636 6448 10676 6488
rect 10924 6448 10964 6488
rect 12556 6448 12596 6488
rect 12652 6448 12692 6488
rect 12844 6448 12884 6488
rect 12940 6448 12980 6488
rect 13708 6448 13748 6488
rect 13804 6448 13844 6488
rect 13996 6448 14036 6488
rect 14092 6448 14132 6488
rect 14193 6448 14233 6488
rect 14860 6448 14900 6488
rect 14956 6448 14996 6488
rect 15244 6448 15284 6488
rect 15436 6448 15476 6488
rect 15532 6448 15572 6488
rect 16108 6448 16148 6488
rect 16972 6448 17012 6488
rect 19564 6448 19604 6488
rect 21004 6448 21044 6488
rect 22252 6448 22292 6488
rect 22444 6448 22484 6488
rect 23692 6448 23732 6488
rect 23980 6448 24020 6488
rect 24172 6448 24212 6488
rect 24268 6448 24308 6488
rect 24652 6448 24692 6488
rect 24748 6448 24788 6488
rect 24940 6448 24980 6488
rect 25132 6448 25172 6488
rect 25516 6448 25556 6488
rect 25708 6448 25748 6488
rect 25804 6448 25844 6488
rect 26284 6448 26324 6488
rect 26380 6448 26420 6488
rect 26860 6448 26900 6488
rect 26956 6448 26996 6488
rect 28396 6448 28436 6488
rect 28588 6448 28628 6488
rect 28780 6448 28820 6488
rect 28972 6448 29012 6488
rect 29068 6448 29108 6488
rect 29260 6448 29300 6488
rect 29452 6448 29492 6488
rect 29740 6448 29780 6488
rect 30220 6448 30260 6488
rect 30892 6448 30932 6488
rect 31084 6448 31124 6488
rect 31468 6448 31508 6488
rect 32332 6448 32372 6488
rect 33484 6448 33524 6488
rect 34444 6448 34484 6488
rect 34636 6448 34676 6488
rect 35500 6448 35540 6488
rect 35884 6448 35924 6488
rect 36748 6448 36788 6488
rect 37900 6448 37940 6488
rect 9388 6364 9428 6404
rect 18796 6364 18836 6404
rect 23308 6364 23348 6404
rect 25228 6364 25268 6404
rect 25420 6364 25460 6404
rect 7084 6280 7124 6320
rect 9484 6280 9524 6320
rect 11212 6280 11252 6320
rect 14572 6280 14612 6320
rect 18124 6280 18164 6320
rect 18412 6280 18452 6320
rect 24940 6280 24980 6320
rect 25324 6280 25364 6320
rect 26572 6280 26612 6320
rect 7276 6196 7316 6236
rect 9580 6196 9620 6236
rect 10060 6196 10100 6236
rect 10540 6196 10580 6236
rect 20236 6196 20276 6236
rect 25996 6196 26036 6236
rect 28780 6196 28820 6236
rect 29260 6196 29300 6236
rect 33772 6196 33812 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4876 5860 4916 5900
rect 8236 5860 8276 5900
rect 11212 5860 11252 5900
rect 23308 5860 23348 5900
rect 28300 5860 28340 5900
rect 29356 5860 29396 5900
rect 31084 5860 31124 5900
rect 34252 5860 34292 5900
rect 4204 5776 4244 5816
rect 4684 5776 4724 5816
rect 10732 5776 10772 5816
rect 11500 5776 11540 5816
rect 11596 5776 11636 5816
rect 17452 5776 17492 5816
rect 24940 5776 24980 5816
rect 35116 5776 35156 5816
rect 11692 5692 11732 5732
rect 13708 5692 13748 5732
rect 4396 5608 4436 5648
rect 4588 5608 4628 5648
rect 4684 5608 4724 5648
rect 5548 5608 5588 5648
rect 5836 5608 5876 5648
rect 6124 5608 6164 5648
rect 6796 5608 6836 5648
rect 7180 5608 7220 5648
rect 7276 5608 7316 5648
rect 7756 5608 7796 5648
rect 7852 5608 7892 5648
rect 7948 5608 7988 5648
rect 8236 5608 8276 5648
rect 8428 5608 8468 5648
rect 8524 5608 8564 5648
rect 9388 5608 9428 5648
rect 10348 5608 10388 5648
rect 10540 5608 10580 5648
rect 10732 5608 10772 5648
rect 10828 5608 10868 5648
rect 11116 5608 11156 5648
rect 11308 5608 11348 5648
rect 11884 5650 11924 5690
rect 14092 5692 14132 5732
rect 23788 5692 23828 5732
rect 35020 5692 35060 5732
rect 35212 5692 35252 5732
rect 11788 5608 11828 5648
rect 12172 5608 12212 5648
rect 12268 5608 12308 5648
rect 13420 5608 13460 5648
rect 13612 5608 13652 5648
rect 13804 5608 13844 5648
rect 13996 5608 14036 5648
rect 14188 5608 14228 5648
rect 14380 5608 14420 5648
rect 15052 5608 15092 5648
rect 15436 5608 15476 5648
rect 15725 5625 15765 5665
rect 16012 5608 16052 5648
rect 16300 5608 16340 5648
rect 17932 5608 17972 5648
rect 18316 5608 18356 5648
rect 19180 5608 19220 5648
rect 20332 5608 20372 5648
rect 20908 5608 20948 5648
rect 21292 5608 21332 5648
rect 22156 5608 22196 5648
rect 23404 5608 23444 5648
rect 23692 5608 23732 5648
rect 23980 5608 24020 5648
rect 24268 5608 24308 5648
rect 25324 5608 25364 5648
rect 25420 5608 25460 5648
rect 25612 5608 25652 5648
rect 27143 5603 27183 5643
rect 27244 5608 27284 5648
rect 27820 5608 27860 5648
rect 27916 5608 27956 5648
rect 28108 5608 28148 5648
rect 28300 5608 28340 5648
rect 28492 5608 28532 5648
rect 30028 5608 30068 5648
rect 30892 5608 30932 5648
rect 31756 5608 31796 5648
rect 33484 5608 33524 5648
rect 33772 5608 33812 5648
rect 33964 5608 34004 5648
rect 34060 5608 34100 5648
rect 34252 5608 34292 5648
rect 34444 5608 34484 5648
rect 34636 5608 34676 5648
rect 34732 5608 34772 5648
rect 34924 5608 34964 5648
rect 35308 5608 35348 5648
rect 12748 5524 12788 5564
rect 27052 5524 27092 5564
rect 652 5440 692 5480
rect 5740 5440 5780 5480
rect 6988 5440 7028 5480
rect 8044 5440 8084 5480
rect 8716 5440 8756 5480
rect 9676 5440 9716 5480
rect 12460 5440 12500 5480
rect 15340 5440 15380 5480
rect 15820 5440 15860 5480
rect 16204 5440 16244 5480
rect 25132 5440 25172 5480
rect 26284 5440 26324 5480
rect 26860 5440 26900 5480
rect 26956 5440 26996 5480
rect 29164 5440 29204 5480
rect 30220 5440 30260 5480
rect 33676 5440 33716 5480
rect 34444 5440 34484 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 22156 5162 22196 5202
rect 652 5104 692 5144
rect 11980 5104 12020 5144
rect 12076 5104 12116 5144
rect 14764 5104 14804 5144
rect 14860 5104 14900 5144
rect 20620 5104 20660 5144
rect 26668 5104 26708 5144
rect 27340 5104 27380 5144
rect 28396 5104 28436 5144
rect 5932 5020 5972 5060
rect 11884 5020 11924 5060
rect 13804 5020 13844 5060
rect 14668 5020 14708 5060
rect 17740 5020 17780 5060
rect 20812 5020 20852 5060
rect 27436 5020 27476 5060
rect 4204 4936 4244 4976
rect 4396 4936 4436 4976
rect 4492 4936 4532 4976
rect 5356 4936 5396 4976
rect 5740 4936 5780 4976
rect 5836 4936 5876 4976
rect 6028 4936 6068 4976
rect 6220 4936 6260 4976
rect 6892 4936 6932 4976
rect 7180 4936 7220 4976
rect 7276 4936 7316 4976
rect 7372 4936 7412 4976
rect 7468 4936 7508 4976
rect 7852 4936 7892 4976
rect 8716 4936 8756 4976
rect 9100 4936 9140 4976
rect 9964 4936 10004 4976
rect 11116 4936 11156 4976
rect 11692 4936 11732 4976
rect 11788 4936 11828 4976
rect 12940 4936 12980 4976
rect 13132 4936 13172 4976
rect 13324 4936 13364 4976
rect 13420 4936 13460 4976
rect 13708 4936 13748 4976
rect 13900 4936 13940 4976
rect 14092 4936 14132 4976
rect 14284 4936 14324 4976
rect 14476 4936 14516 4976
rect 14572 4936 14612 4976
rect 15148 4936 15188 4976
rect 16012 4936 16052 4976
rect 16108 4936 16148 4976
rect 16300 4936 16340 4976
rect 16396 4936 16436 4976
rect 16588 4936 16628 4976
rect 16780 4936 16820 4976
rect 18412 4936 18452 4976
rect 19468 4936 19508 4976
rect 19948 4936 19988 4976
rect 21484 4936 21524 4976
rect 21964 4936 22004 4976
rect 22060 4936 22100 4976
rect 22348 4936 22388 4976
rect 23020 4936 23060 4976
rect 23308 4936 23348 4976
rect 24460 4936 24500 4976
rect 25324 4936 25364 4976
rect 25708 4936 25748 4976
rect 25996 4936 26036 4976
rect 26092 4936 26132 4976
rect 26476 4936 26516 4976
rect 26764 4936 26804 4976
rect 26956 4936 26996 4976
rect 27532 4936 27572 4976
rect 27628 4936 27668 4976
rect 27916 4936 27956 4976
rect 28012 4936 28052 4976
rect 28204 4936 28244 4976
rect 28588 4936 28628 4976
rect 28684 4936 28724 4976
rect 29164 4936 29204 4976
rect 29548 4936 29588 4976
rect 30412 4936 30452 4976
rect 31564 4936 31604 4976
rect 3820 4768 3860 4808
rect 4492 4768 4532 4808
rect 15820 4768 15860 4808
rect 16588 4768 16628 4808
rect 27340 4768 27380 4808
rect 4684 4684 4724 4724
rect 7660 4684 7700 4724
rect 8524 4684 8564 4724
rect 12268 4684 12308 4724
rect 13132 4684 13172 4724
rect 14188 4684 14228 4724
rect 17452 4684 17492 4724
rect 18892 4684 18932 4724
rect 21676 4684 21716 4724
rect 28204 4684 28244 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 7564 4348 7604 4388
rect 11212 4348 11252 4388
rect 19372 4348 19412 4388
rect 23308 4348 23348 4388
rect 25228 4348 25268 4388
rect 25516 4348 25556 4388
rect 8140 4264 8180 4304
rect 9196 4264 9236 4304
rect 11020 4264 11060 4304
rect 11404 4264 11444 4304
rect 14572 4264 14612 4304
rect 29068 4264 29108 4304
rect 3340 4096 3380 4136
rect 3724 4096 3764 4136
rect 4588 4096 4628 4136
rect 5836 4096 5876 4136
rect 6220 4096 6260 4136
rect 7276 4096 7316 4136
rect 7372 4096 7412 4136
rect 7852 4096 7892 4136
rect 9388 4096 9428 4136
rect 9484 4096 9524 4136
rect 9676 4096 9716 4136
rect 10444 4096 10484 4136
rect 10636 4096 10676 4136
rect 11404 4096 11444 4136
rect 11692 4096 11732 4136
rect 11788 4096 11828 4136
rect 11884 4096 11924 4136
rect 11980 4096 12020 4136
rect 12172 4096 12212 4136
rect 12556 4096 12596 4136
rect 13420 4096 13460 4136
rect 14764 4096 14804 4136
rect 14860 4096 14900 4136
rect 14956 4096 14996 4136
rect 15052 4096 15092 4136
rect 15244 4096 15284 4136
rect 16108 4096 16148 4136
rect 17356 4096 17396 4136
rect 18220 4096 18260 4136
rect 19756 4096 19796 4136
rect 20044 4096 20084 4136
rect 20716 4096 20756 4136
rect 20908 4096 20948 4136
rect 21292 4096 21332 4136
rect 22156 4096 22196 4136
rect 23596 4096 23636 4136
rect 23692 4096 23732 4136
rect 23884 4096 23924 4136
rect 25132 4096 25172 4136
rect 25708 4096 25748 4136
rect 25804 4096 25844 4136
rect 25996 4096 26036 4136
rect 26188 4096 26228 4136
rect 26476 4096 26516 4136
rect 26668 4096 26708 4136
rect 26956 4096 26996 4136
rect 28204 4096 28244 4136
rect 28396 4096 28436 4136
rect 29260 4096 29300 4136
rect 29932 4096 29972 4136
rect 30124 4096 30164 4136
rect 30508 4096 30548 4136
rect 31372 4096 31412 4136
rect 32620 4096 32660 4136
rect 10540 4012 10580 4052
rect 16972 4012 17012 4052
rect 25612 4012 25652 4052
rect 26092 4012 26132 4052
rect 652 3928 692 3968
rect 6892 3928 6932 3968
rect 7276 3928 7316 3968
rect 9676 3928 9716 3968
rect 11212 3928 11252 3968
rect 15916 3928 15956 3968
rect 16780 3928 16820 3968
rect 19564 3928 19604 3968
rect 19852 3928 19892 3968
rect 23884 3928 23924 3968
rect 25516 3928 25556 3968
rect 26764 3928 26804 3968
rect 27532 3928 27572 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 25612 3650 25652 3690
rect 652 3592 692 3632
rect 8044 3592 8084 3632
rect 9388 3592 9428 3632
rect 11404 3592 11444 3632
rect 12364 3592 12404 3632
rect 14476 3592 14516 3632
rect 15052 3592 15092 3632
rect 16300 3592 16340 3632
rect 26572 3592 26612 3632
rect 27340 3592 27380 3632
rect 27628 3592 27668 3632
rect 16780 3508 16820 3548
rect 24940 3508 24980 3548
rect 5452 3424 5492 3464
rect 5836 3424 5876 3464
rect 6700 3424 6740 3464
rect 8716 3424 8756 3464
rect 9388 3424 9428 3464
rect 9484 3424 9524 3464
rect 10540 3424 10580 3464
rect 11017 3445 11057 3485
rect 11212 3424 11252 3464
rect 12076 3424 12116 3464
rect 12268 3424 12308 3464
rect 12460 3424 12500 3464
rect 12556 3424 12596 3464
rect 14572 3424 14612 3464
rect 14956 3424 14996 3464
rect 15148 3424 15188 3464
rect 15244 3424 15284 3464
rect 15436 3424 15476 3464
rect 15820 3424 15860 3464
rect 16204 3424 16244 3464
rect 16396 3424 16436 3464
rect 16492 3424 16532 3464
rect 17164 3424 17204 3464
rect 18028 3424 18068 3464
rect 19756 3424 19796 3464
rect 20428 3424 20468 3464
rect 20620 3424 20660 3464
rect 21004 3424 21044 3464
rect 21868 3424 21908 3464
rect 23020 3424 23060 3464
rect 23308 3424 23348 3464
rect 25132 3424 25172 3464
rect 25420 3424 25460 3464
rect 25804 3424 25844 3464
rect 7852 3340 7892 3380
rect 15532 3340 15572 3380
rect 25708 3382 25748 3422
rect 26476 3424 26516 3464
rect 26668 3424 26708 3464
rect 26860 3424 26900 3464
rect 27244 3424 27284 3464
rect 28300 3424 28340 3464
rect 28492 3424 28532 3464
rect 29164 3424 29204 3464
rect 29356 3424 29396 3464
rect 29740 3424 29780 3464
rect 30604 3424 30644 3464
rect 31852 3424 31892 3464
rect 15724 3340 15764 3380
rect 12748 3256 12788 3296
rect 13324 3256 13364 3296
rect 15628 3256 15668 3296
rect 9676 3172 9716 3212
rect 9868 3172 9908 3212
rect 11116 3172 11156 3212
rect 14764 3172 14804 3212
rect 19180 3172 19220 3212
rect 23980 3172 24020 3212
rect 26092 3172 26132 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 6700 2836 6740 2876
rect 9388 2836 9428 2876
rect 11980 2836 12020 2876
rect 15244 2836 15284 2876
rect 16876 2836 16916 2876
rect 21388 2836 21428 2876
rect 26380 2836 26420 2876
rect 26572 2836 26612 2876
rect 29836 2836 29876 2876
rect 30220 2836 30260 2876
rect 6892 2752 6932 2792
rect 9196 2752 9236 2792
rect 17260 2752 17300 2792
rect 25516 2752 25556 2792
rect 844 2668 884 2708
rect 6124 2668 6164 2708
rect 8524 2668 8564 2708
rect 19948 2668 19988 2708
rect 21964 2668 22004 2708
rect 24556 2668 24596 2708
rect 6028 2584 6068 2624
rect 6220 2584 6260 2624
rect 6412 2584 6452 2624
rect 6508 2584 6548 2624
rect 6700 2584 6740 2624
rect 8044 2584 8084 2624
rect 8140 2584 8180 2624
rect 8236 2584 8276 2624
rect 8428 2584 8468 2624
rect 8620 2584 8660 2624
rect 9196 2584 9236 2624
rect 9580 2584 9620 2624
rect 9964 2584 10004 2624
rect 10828 2584 10868 2624
rect 12076 2584 12116 2624
rect 12844 2584 12884 2624
rect 13228 2584 13268 2624
rect 14092 2584 14132 2624
rect 15724 2584 15764 2624
rect 15916 2584 15956 2624
rect 16108 2584 16148 2624
rect 16300 2584 16340 2624
rect 16492 2584 16532 2624
rect 16684 2584 16724 2624
rect 16972 2584 17012 2624
rect 18700 2584 18740 2624
rect 20236 2584 20276 2624
rect 20332 2584 20372 2624
rect 20716 2584 20756 2624
rect 23116 2584 23156 2624
rect 23980 2584 24020 2624
rect 24364 2584 24404 2624
rect 25228 2584 25268 2624
rect 25420 2584 25460 2624
rect 25708 2584 25748 2624
rect 27244 2584 27284 2624
rect 27436 2584 27476 2624
rect 27820 2584 27860 2624
rect 28684 2584 28724 2624
rect 30892 2584 30932 2624
rect 16204 2500 16244 2540
rect 16588 2500 16628 2540
rect 18028 2500 18068 2540
rect 652 2416 692 2456
rect 26380 2416 26420 2456
rect 26572 2416 26612 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 20812 2080 20852 2120
rect 22060 2080 22100 2120
rect 29356 2080 29396 2120
rect 15052 1996 15092 2036
rect 9676 1912 9716 1952
rect 9772 1912 9812 1952
rect 9964 1912 10004 1952
rect 10732 1912 10772 1952
rect 11116 1912 11156 1952
rect 11980 1912 12020 1952
rect 13132 1912 13172 1952
rect 15436 1912 15476 1952
rect 16300 1912 16340 1952
rect 21004 1912 21044 1952
rect 21292 1912 21332 1952
rect 22540 1912 22580 1952
rect 23596 1912 23636 1952
rect 23980 1912 24020 1952
rect 24844 1912 24884 1952
rect 25996 1912 26036 1952
rect 26284 1912 26324 1952
rect 26668 1912 26708 1952
rect 27532 1912 27572 1952
rect 28780 1912 28820 1952
rect 29452 1912 29492 1952
rect 9964 1744 10004 1784
rect 10156 1744 10196 1784
rect 17452 1660 17492 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 26284 1324 26324 1364
rect 10156 1240 10196 1280
rect 11212 1240 11252 1280
rect 15532 1240 15572 1280
rect 24364 1240 24404 1280
rect 25228 1156 25268 1196
rect 10252 1072 10292 1112
rect 11884 1072 11924 1112
rect 23308 1072 23348 1112
rect 23980 1072 24020 1112
rect 25036 1072 25076 1112
rect 25516 1072 25556 1112
rect 25612 1072 25652 1112
rect 26092 1072 26132 1112
rect 26476 1072 26516 1112
rect 26668 1072 26708 1112
rect 26764 1072 26804 1112
rect 25996 904 26036 944
rect 26476 904 26516 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 267 37568 309 37577
rect 267 37528 268 37568
rect 308 37528 309 37568
rect 267 37519 309 37528
rect 27435 37568 27477 37577
rect 27435 37528 27436 37568
rect 27476 37528 27477 37568
rect 27435 37519 27477 37528
rect 27819 37568 27861 37577
rect 27819 37528 27820 37568
rect 27860 37528 27861 37568
rect 27819 37519 27861 37528
rect 268 20945 308 37519
rect 26571 37232 26613 37241
rect 26571 37192 26572 37232
rect 26612 37192 26613 37232
rect 26571 37183 26613 37192
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 25708 36856 26420 36896
rect 12556 36728 12596 36737
rect 9964 36560 10004 36569
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 9868 35888 9908 35897
rect 9964 35888 10004 36520
rect 12556 36140 12596 36688
rect 12652 36728 12692 36737
rect 12844 36728 12884 36737
rect 13708 36728 13748 36737
rect 12652 36485 12692 36688
rect 12748 36688 12844 36728
rect 12651 36476 12693 36485
rect 12651 36436 12652 36476
rect 12692 36436 12693 36476
rect 12651 36427 12693 36436
rect 12556 36091 12596 36100
rect 12748 36056 12788 36688
rect 12844 36679 12884 36688
rect 12940 36688 13708 36728
rect 12844 36560 12884 36569
rect 12940 36560 12980 36688
rect 13708 36679 13748 36688
rect 16108 36728 16148 36737
rect 25612 36728 25652 36737
rect 16148 36688 16436 36728
rect 16108 36679 16148 36688
rect 12884 36520 12980 36560
rect 13131 36560 13173 36569
rect 13131 36520 13132 36560
rect 13172 36520 13173 36560
rect 12844 36511 12884 36520
rect 13131 36511 13173 36520
rect 13899 36560 13941 36569
rect 13899 36520 13900 36560
rect 13940 36520 13941 36560
rect 13899 36511 13941 36520
rect 16300 36560 16340 36569
rect 13036 36476 13076 36485
rect 12652 36016 12788 36056
rect 12940 36436 13036 36476
rect 9908 35848 10004 35888
rect 10732 35888 10772 35897
rect 12460 35888 12500 35897
rect 9868 35839 9908 35848
rect 9484 35804 9524 35813
rect 9004 35764 9484 35804
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 9004 35384 9044 35764
rect 9484 35755 9524 35764
rect 9004 35335 9044 35344
rect 5931 35300 5973 35309
rect 5931 35260 5932 35300
rect 5972 35260 5973 35300
rect 5931 35251 5973 35260
rect 6987 35300 7029 35309
rect 6987 35260 6988 35300
rect 7028 35260 7029 35300
rect 6987 35251 7029 35260
rect 4779 35216 4821 35225
rect 4779 35176 4780 35216
rect 4820 35176 4821 35216
rect 4779 35167 4821 35176
rect 5355 35216 5397 35225
rect 5355 35176 5356 35216
rect 5396 35176 5397 35216
rect 5355 35167 5397 35176
rect 5452 35216 5492 35227
rect 4492 35048 4532 35057
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 2572 34544 2612 34553
rect 1996 33704 2036 33713
rect 1323 33116 1365 33125
rect 1323 33076 1324 33116
rect 1364 33076 1365 33116
rect 1323 33067 1365 33076
rect 1324 32276 1364 33067
rect 1324 32227 1364 32236
rect 1708 33032 1748 33041
rect 1708 32192 1748 32992
rect 1996 32957 2036 33664
rect 2380 33704 2420 33713
rect 2572 33704 2612 34504
rect 3627 34376 3669 34385
rect 3627 34336 3628 34376
rect 3668 34336 3669 34376
rect 3627 34327 3669 34336
rect 4012 34376 4052 34385
rect 4492 34376 4532 35008
rect 4052 34336 4532 34376
rect 4012 34327 4052 34336
rect 3628 34242 3668 34327
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3243 33956 3285 33965
rect 3243 33916 3244 33956
rect 3284 33916 3285 33956
rect 3243 33907 3285 33916
rect 2420 33664 2612 33704
rect 3244 33704 3284 33907
rect 4588 33872 4628 33881
rect 4780 33872 4820 35167
rect 5356 35082 5396 35167
rect 5452 35141 5492 35176
rect 5644 35216 5684 35225
rect 5836 35216 5876 35225
rect 5684 35176 5780 35216
rect 5644 35167 5684 35176
rect 5451 35132 5493 35141
rect 5451 35092 5452 35132
rect 5492 35092 5493 35132
rect 5451 35083 5493 35092
rect 5644 34964 5684 34973
rect 5644 34385 5684 34924
rect 4876 34376 4916 34385
rect 4876 34049 4916 34336
rect 5643 34376 5685 34385
rect 5643 34336 5644 34376
rect 5684 34336 5685 34376
rect 5643 34327 5685 34336
rect 4971 34124 5013 34133
rect 4971 34084 4972 34124
rect 5012 34084 5013 34124
rect 4971 34075 5013 34084
rect 4875 34040 4917 34049
rect 4875 34000 4876 34040
rect 4916 34000 4917 34040
rect 4875 33991 4917 34000
rect 4972 33872 5012 34075
rect 5740 34049 5780 35176
rect 5836 34133 5876 35176
rect 5932 35166 5972 35251
rect 6028 35216 6068 35225
rect 6028 35141 6068 35176
rect 6124 35216 6164 35225
rect 6027 35132 6069 35141
rect 6027 35092 6028 35132
rect 6068 35092 6069 35132
rect 6027 35083 6069 35092
rect 6028 34796 6068 35083
rect 5932 34756 6068 34796
rect 5835 34124 5877 34133
rect 5835 34084 5836 34124
rect 5876 34084 5877 34124
rect 5835 34075 5877 34084
rect 5739 34040 5781 34049
rect 5739 34000 5740 34040
rect 5780 34000 5781 34040
rect 5739 33991 5781 34000
rect 4628 33832 4820 33872
rect 4876 33832 5012 33872
rect 5067 33872 5109 33881
rect 5067 33832 5068 33872
rect 5108 33832 5109 33872
rect 4588 33823 4628 33832
rect 4876 33788 4916 33832
rect 5067 33823 5109 33832
rect 4876 33739 4916 33748
rect 2380 33655 2420 33664
rect 3244 33655 3284 33664
rect 4683 33704 4725 33713
rect 4683 33664 4684 33704
rect 4724 33664 4725 33704
rect 4683 33655 4725 33664
rect 4972 33704 5012 33713
rect 2763 33620 2805 33629
rect 2763 33580 2764 33620
rect 2804 33580 2805 33620
rect 2763 33571 2805 33580
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 2380 33041 2420 33126
rect 2379 33032 2421 33041
rect 2379 32992 2380 33032
rect 2420 32992 2421 33032
rect 2379 32983 2421 32992
rect 1995 32948 2037 32957
rect 1995 32908 1996 32948
rect 2036 32908 2037 32948
rect 1995 32899 2037 32908
rect 2188 32873 2228 32958
rect 1708 32143 1748 32152
rect 2092 32864 2132 32873
rect 2092 31529 2132 32824
rect 2187 32864 2229 32873
rect 2187 32824 2188 32864
rect 2228 32824 2229 32864
rect 2187 32815 2229 32824
rect 2380 32864 2420 32873
rect 2572 32864 2612 32873
rect 2420 32824 2572 32864
rect 2380 32815 2420 32824
rect 2572 32815 2612 32824
rect 2668 32864 2708 32875
rect 2668 32789 2708 32824
rect 2764 32864 2804 33571
rect 4203 33536 4245 33545
rect 4203 33496 4204 33536
rect 4244 33496 4245 33536
rect 4203 33487 4245 33496
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 3723 33032 3765 33041
rect 3723 32992 3724 33032
rect 3764 32992 3765 33032
rect 3723 32983 3765 32992
rect 3051 32948 3093 32957
rect 3051 32908 3052 32948
rect 3092 32908 3093 32948
rect 3051 32899 3093 32908
rect 2764 32815 2804 32824
rect 2859 32864 2901 32873
rect 2859 32824 2860 32864
rect 2900 32824 2901 32864
rect 2859 32815 2901 32824
rect 2667 32780 2709 32789
rect 2667 32740 2668 32780
rect 2708 32740 2709 32780
rect 2667 32731 2709 32740
rect 2860 32730 2900 32815
rect 3052 32814 3092 32899
rect 3724 32864 3764 32983
rect 3724 32815 3764 32824
rect 4011 32864 4053 32873
rect 4011 32824 4012 32864
rect 4052 32824 4053 32864
rect 4011 32815 4053 32824
rect 4108 32864 4148 32873
rect 4012 32730 4052 32815
rect 4108 32360 4148 32824
rect 4204 32864 4244 33487
rect 4396 33486 4436 33571
rect 4684 33570 4724 33655
rect 4972 33545 5012 33664
rect 5068 33704 5108 33823
rect 5163 33788 5205 33797
rect 5163 33748 5164 33788
rect 5204 33748 5205 33788
rect 5163 33739 5205 33748
rect 5068 33655 5108 33664
rect 5164 33704 5204 33739
rect 5932 33713 5972 34756
rect 6027 34628 6069 34637
rect 6027 34588 6028 34628
rect 6068 34588 6069 34628
rect 6027 34579 6069 34588
rect 6028 34494 6068 34579
rect 5164 33653 5204 33664
rect 5355 33704 5397 33713
rect 5355 33664 5356 33704
rect 5396 33664 5397 33704
rect 5355 33655 5397 33664
rect 5931 33704 5973 33713
rect 5931 33664 5932 33704
rect 5972 33664 5973 33704
rect 5931 33655 5973 33664
rect 6028 33704 6068 33715
rect 5356 33570 5396 33655
rect 6028 33629 6068 33664
rect 6027 33620 6069 33629
rect 6027 33580 6028 33620
rect 6068 33580 6069 33620
rect 6027 33571 6069 33580
rect 4971 33536 5013 33545
rect 4971 33496 4972 33536
rect 5012 33496 5013 33536
rect 4971 33487 5013 33496
rect 4491 33116 4533 33125
rect 4491 33076 4492 33116
rect 4532 33076 4533 33116
rect 4491 33067 4533 33076
rect 4779 33116 4821 33125
rect 4779 33076 4780 33116
rect 4820 33076 4821 33116
rect 4779 33067 4821 33076
rect 4492 32982 4532 33067
rect 4204 32789 4244 32824
rect 4300 32864 4340 32873
rect 4492 32864 4532 32873
rect 4340 32824 4492 32864
rect 4300 32815 4340 32824
rect 4492 32815 4532 32824
rect 4683 32864 4725 32873
rect 4683 32824 4684 32864
rect 4724 32824 4725 32864
rect 4683 32815 4725 32824
rect 4780 32864 4820 33067
rect 4780 32815 4820 32824
rect 5164 33032 5204 33041
rect 4203 32780 4245 32789
rect 4203 32740 4204 32780
rect 4244 32740 4245 32780
rect 4203 32731 4245 32740
rect 4108 32311 4148 32320
rect 2572 32192 2612 32201
rect 1900 31520 1940 31529
rect 1227 31184 1269 31193
rect 1227 31144 1228 31184
rect 1268 31144 1269 31184
rect 1227 31135 1269 31144
rect 1035 30008 1077 30017
rect 1035 29968 1036 30008
rect 1076 29968 1077 30008
rect 1035 29959 1077 29968
rect 1036 29874 1076 29959
rect 1228 29840 1268 31135
rect 1228 29791 1268 29800
rect 1324 30680 1364 30689
rect 1324 29009 1364 30640
rect 1708 30680 1748 30689
rect 1900 30680 1940 31480
rect 2091 31520 2133 31529
rect 2091 31480 2092 31520
rect 2132 31480 2133 31520
rect 2091 31471 2133 31480
rect 1748 30640 1940 30680
rect 2572 30680 2612 32152
rect 3723 32192 3765 32201
rect 3723 32152 3724 32192
rect 3764 32152 3765 32192
rect 3723 32143 3765 32152
rect 3724 32108 3764 32143
rect 3724 32057 3764 32068
rect 3531 31940 3573 31949
rect 3531 31900 3532 31940
rect 3572 31900 3573 31940
rect 3531 31891 3573 31900
rect 4107 31940 4149 31949
rect 4107 31900 4108 31940
rect 4148 31900 4149 31940
rect 4107 31891 4149 31900
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3435 31520 3477 31529
rect 3435 31480 3436 31520
rect 3476 31480 3477 31520
rect 3435 31471 3477 31480
rect 2667 31436 2709 31445
rect 2667 31396 2668 31436
rect 2708 31396 2709 31436
rect 2667 31387 2709 31396
rect 1708 30631 1748 30640
rect 1611 30008 1653 30017
rect 1611 29968 1612 30008
rect 1652 29968 1653 30008
rect 1611 29959 1653 29968
rect 1612 29840 1652 29959
rect 1612 29791 1652 29800
rect 2476 29840 2516 29849
rect 2572 29840 2612 30640
rect 2516 29800 2612 29840
rect 2476 29791 2516 29800
rect 2572 29177 2612 29800
rect 2571 29168 2613 29177
rect 2571 29128 2572 29168
rect 2612 29128 2613 29168
rect 2571 29119 2613 29128
rect 1323 29000 1365 29009
rect 1323 28960 1324 29000
rect 1364 28960 1365 29000
rect 1323 28951 1365 28960
rect 1804 29000 1844 29009
rect 1708 28328 1748 28337
rect 1804 28328 1844 28960
rect 2572 28328 2612 29119
rect 1748 28288 1844 28328
rect 2476 28288 2572 28328
rect 1708 28279 1748 28288
rect 1323 28244 1365 28253
rect 1323 28204 1324 28244
rect 1364 28204 1365 28244
rect 1323 28195 1365 28204
rect 1324 28110 1364 28195
rect 1708 27488 1748 27497
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1612 26816 1652 26825
rect 1708 26816 1748 27448
rect 1652 26776 1748 26816
rect 2476 26816 2516 28288
rect 2572 28193 2612 28288
rect 2668 27740 2708 31387
rect 3436 31386 3476 31471
rect 3532 31352 3572 31891
rect 4108 31806 4148 31891
rect 4011 31520 4053 31529
rect 4011 31480 4012 31520
rect 4052 31480 4053 31520
rect 4011 31471 4053 31480
rect 3532 31303 3572 31312
rect 3820 31352 3860 31361
rect 4012 31352 4052 31471
rect 3860 31312 3956 31352
rect 3820 31303 3860 31312
rect 3724 31184 3764 31193
rect 3532 31144 3724 31184
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3532 30092 3572 31144
rect 3724 31135 3764 31144
rect 3916 30848 3956 31312
rect 4012 31016 4052 31312
rect 4107 31352 4149 31361
rect 4107 31312 4108 31352
rect 4148 31312 4149 31352
rect 4107 31303 4149 31312
rect 4204 31352 4244 32731
rect 4684 32730 4724 32815
rect 4971 32780 5013 32789
rect 4971 32740 4972 32780
rect 5012 32740 5013 32780
rect 4971 32731 5013 32740
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4780 32217 4820 32287
rect 4972 32276 5012 32731
rect 4972 32227 5012 32236
rect 4779 32152 4780 32201
rect 4820 32152 4821 32201
rect 5164 32192 5204 32992
rect 6124 32957 6164 35176
rect 6988 35216 7028 35251
rect 6988 35165 7028 35176
rect 8332 35216 8372 35225
rect 7180 35048 7220 35057
rect 6316 34964 6356 34973
rect 6220 34376 6260 34385
rect 6316 34376 6356 34924
rect 6507 34964 6549 34973
rect 6507 34924 6508 34964
rect 6548 34924 6549 34964
rect 6507 34915 6549 34924
rect 6260 34336 6356 34376
rect 6220 34327 6260 34336
rect 6315 34040 6357 34049
rect 6315 34000 6316 34040
rect 6356 34000 6357 34040
rect 6315 33991 6357 34000
rect 6316 33872 6356 33991
rect 6316 33823 6356 33832
rect 6411 33788 6453 33797
rect 6411 33748 6412 33788
rect 6452 33748 6453 33788
rect 6411 33739 6453 33748
rect 6412 33704 6452 33739
rect 6412 33545 6452 33664
rect 6508 33704 6548 34915
rect 6604 34376 6644 34385
rect 7180 34376 7220 35008
rect 7659 34964 7701 34973
rect 7659 34924 7660 34964
rect 7700 34924 7701 34964
rect 7659 34915 7701 34924
rect 7660 34830 7700 34915
rect 8332 34637 8372 35176
rect 8811 35216 8853 35225
rect 8811 35176 8812 35216
rect 8852 35176 8853 35216
rect 8811 35167 8853 35176
rect 8908 35216 8948 35227
rect 8812 35082 8852 35167
rect 8908 35141 8948 35176
rect 9100 35216 9140 35225
rect 8907 35132 8949 35141
rect 8907 35092 8908 35132
rect 8948 35092 8949 35132
rect 8907 35083 8949 35092
rect 8811 34964 8853 34973
rect 8811 34924 8812 34964
rect 8852 34924 8853 34964
rect 8811 34915 8853 34924
rect 8331 34628 8373 34637
rect 8331 34588 8332 34628
rect 8372 34588 8373 34628
rect 8331 34579 8373 34588
rect 6644 34336 7220 34376
rect 7468 34376 7508 34385
rect 6604 34327 6644 34336
rect 7468 33965 7508 34336
rect 8332 34049 8372 34579
rect 8812 34376 8852 34915
rect 9100 34637 9140 35176
rect 9292 35216 9332 35225
rect 9195 35132 9237 35141
rect 9195 35092 9196 35132
rect 9236 35092 9237 35132
rect 9195 35083 9237 35092
rect 9099 34628 9141 34637
rect 9099 34588 9100 34628
rect 9140 34588 9141 34628
rect 9099 34579 9141 34588
rect 8812 34327 8852 34336
rect 8908 34376 8948 34385
rect 9100 34376 9140 34385
rect 8948 34336 9100 34376
rect 8908 34327 8948 34336
rect 9100 34327 9140 34336
rect 9196 34376 9236 35083
rect 9292 34628 9332 35176
rect 9676 35216 9716 35225
rect 9388 34628 9428 34637
rect 9292 34588 9388 34628
rect 9388 34579 9428 34588
rect 9676 34553 9716 35176
rect 10540 35216 10580 35225
rect 10732 35216 10772 35848
rect 12268 35848 12460 35888
rect 11883 35720 11925 35729
rect 11883 35680 11884 35720
rect 11924 35680 11925 35720
rect 11883 35671 11925 35680
rect 11884 35586 11924 35671
rect 12268 35384 12308 35848
rect 12460 35839 12500 35848
rect 12268 35335 12308 35344
rect 10580 35176 10772 35216
rect 10923 35216 10965 35225
rect 10923 35176 10924 35216
rect 10964 35176 10965 35216
rect 9675 34544 9717 34553
rect 9675 34504 9676 34544
rect 9716 34504 9717 34544
rect 9675 34495 9717 34504
rect 10443 34544 10485 34553
rect 10443 34504 10444 34544
rect 10484 34504 10485 34544
rect 10443 34495 10485 34504
rect 10444 34410 10484 34495
rect 8620 34208 8660 34217
rect 8331 34040 8373 34049
rect 8331 34000 8332 34040
rect 8372 34000 8373 34040
rect 8331 33991 8373 34000
rect 6699 33956 6741 33965
rect 6699 33916 6700 33956
rect 6740 33916 6741 33956
rect 6699 33907 6741 33916
rect 7467 33956 7509 33965
rect 7467 33916 7468 33956
rect 7508 33916 7509 33956
rect 7467 33907 7509 33916
rect 6508 33655 6548 33664
rect 6603 33704 6645 33713
rect 6603 33664 6604 33704
rect 6644 33664 6645 33704
rect 6603 33655 6645 33664
rect 6604 33570 6644 33655
rect 6411 33536 6453 33545
rect 6411 33496 6412 33536
rect 6452 33496 6453 33536
rect 6411 33487 6453 33496
rect 6411 33368 6453 33377
rect 6411 33328 6412 33368
rect 6452 33328 6453 33368
rect 6411 33319 6453 33328
rect 6123 32948 6165 32957
rect 6123 32908 6124 32948
rect 6164 32908 6165 32948
rect 6123 32899 6165 32908
rect 5451 32864 5493 32873
rect 6028 32864 6068 32873
rect 5451 32824 5452 32864
rect 5492 32824 5493 32864
rect 5451 32815 5493 32824
rect 5548 32824 6028 32864
rect 5355 32780 5397 32789
rect 5355 32740 5356 32780
rect 5396 32740 5397 32780
rect 5355 32731 5397 32740
rect 5356 32646 5396 32731
rect 5356 32192 5396 32201
rect 5164 32152 5356 32192
rect 4779 32143 4821 32152
rect 5356 32143 5396 32152
rect 4587 31520 4629 31529
rect 4779 31520 4821 31529
rect 4587 31480 4588 31520
rect 4628 31480 4724 31520
rect 4587 31471 4629 31480
rect 4108 31218 4148 31303
rect 4012 30976 4148 31016
rect 4012 30848 4052 30857
rect 3916 30808 4012 30848
rect 4012 30799 4052 30808
rect 3723 30596 3765 30605
rect 3723 30556 3724 30596
rect 3764 30556 3765 30596
rect 3723 30547 3765 30556
rect 3724 30462 3764 30547
rect 4108 30512 4148 30976
rect 4204 30596 4244 31312
rect 4300 31352 4340 31361
rect 4492 31352 4532 31361
rect 4340 31312 4492 31352
rect 4300 31303 4340 31312
rect 4492 31303 4532 31312
rect 4684 31352 4724 31480
rect 4779 31480 4780 31520
rect 4820 31480 4821 31520
rect 4779 31471 4821 31480
rect 4684 31303 4724 31312
rect 4780 31352 4820 31471
rect 4780 31303 4820 31312
rect 4971 31352 5013 31361
rect 4971 31312 4972 31352
rect 5012 31312 5013 31352
rect 4971 31303 5013 31312
rect 5068 31352 5108 31361
rect 5260 31352 5300 31361
rect 5108 31312 5260 31352
rect 5068 31303 5108 31312
rect 5260 31303 5300 31312
rect 5356 31352 5396 31361
rect 5452 31352 5492 32815
rect 5548 31520 5588 32824
rect 6028 32815 6068 32824
rect 6412 32864 6452 33319
rect 6412 32815 6452 32824
rect 6508 32864 6548 32875
rect 6508 32789 6548 32824
rect 6603 32864 6645 32873
rect 6603 32824 6604 32864
rect 6644 32824 6645 32864
rect 6603 32815 6645 32824
rect 6507 32780 6549 32789
rect 6507 32740 6508 32780
rect 6548 32740 6549 32780
rect 6507 32731 6549 32740
rect 6604 32730 6644 32815
rect 5643 32696 5685 32705
rect 5643 32656 5644 32696
rect 5684 32656 5685 32696
rect 5643 32647 5685 32656
rect 6315 32696 6357 32705
rect 6315 32656 6316 32696
rect 6356 32656 6357 32696
rect 6315 32647 6357 32656
rect 5548 31471 5588 31480
rect 5396 31312 5492 31352
rect 5548 31352 5588 31361
rect 5644 31352 5684 32647
rect 6316 32562 6356 32647
rect 6700 32201 6740 33907
rect 8620 33881 8660 34168
rect 8907 34040 8949 34049
rect 8907 34000 8908 34040
rect 8948 34000 8949 34040
rect 8907 33991 8949 34000
rect 8619 33872 8661 33881
rect 8619 33832 8620 33872
rect 8660 33832 8661 33872
rect 8619 33823 8661 33832
rect 6987 33788 7029 33797
rect 6987 33748 6988 33788
rect 7028 33748 7029 33788
rect 6987 33739 7029 33748
rect 6988 33654 7028 33739
rect 7852 33704 7892 33713
rect 7179 33620 7221 33629
rect 7179 33580 7180 33620
rect 7220 33580 7221 33620
rect 7179 33571 7221 33580
rect 6891 33200 6933 33209
rect 6891 33160 6892 33200
rect 6932 33160 6933 33200
rect 6891 33151 6933 33160
rect 6892 32873 6932 33151
rect 7084 33041 7124 33126
rect 7083 33032 7125 33041
rect 7083 32992 7084 33032
rect 7124 32992 7125 33032
rect 7083 32983 7125 32992
rect 6796 32864 6836 32873
rect 6219 32192 6261 32201
rect 6219 32152 6220 32192
rect 6260 32152 6261 32192
rect 6219 32143 6261 32152
rect 6699 32192 6741 32201
rect 6699 32152 6700 32192
rect 6740 32152 6741 32192
rect 6699 32143 6741 32152
rect 6220 32058 6260 32143
rect 6700 31520 6740 32143
rect 6796 31529 6836 32824
rect 6891 32864 6933 32873
rect 6891 32824 6892 32864
rect 6932 32824 6933 32864
rect 6891 32815 6933 32824
rect 7083 32864 7125 32873
rect 7083 32824 7084 32864
rect 7124 32824 7125 32864
rect 7083 32815 7125 32824
rect 6892 32730 6932 32815
rect 7084 32730 7124 32815
rect 6700 31471 6740 31480
rect 6795 31520 6837 31529
rect 6795 31480 6796 31520
rect 6836 31480 6837 31520
rect 6795 31471 6837 31480
rect 6891 31436 6933 31445
rect 6891 31396 6892 31436
rect 6932 31396 6933 31436
rect 6891 31387 6933 31396
rect 5588 31312 5684 31352
rect 6124 31352 6164 31361
rect 6164 31312 6260 31352
rect 5356 31303 5396 31312
rect 5548 31303 5588 31312
rect 6124 31303 6164 31312
rect 4588 31193 4628 31278
rect 4587 31184 4629 31193
rect 4587 31144 4588 31184
rect 4628 31144 4629 31184
rect 4587 31135 4629 31144
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4876 30848 4916 30857
rect 4972 30848 5012 31303
rect 4916 30808 5012 30848
rect 4876 30799 4916 30808
rect 4684 30680 4724 30689
rect 5548 30680 5588 30689
rect 4724 30640 4820 30680
rect 4684 30631 4724 30640
rect 4204 30556 4436 30596
rect 4108 30472 4340 30512
rect 4012 30428 4052 30437
rect 4052 30388 4244 30428
rect 4012 30379 4052 30388
rect 3723 30344 3765 30353
rect 3723 30304 3724 30344
rect 3764 30304 3765 30344
rect 3723 30295 3765 30304
rect 3052 30052 3572 30092
rect 2764 29261 2804 29305
rect 2763 29252 2805 29261
rect 2763 29212 2764 29252
rect 2804 29212 2805 29252
rect 2763 29210 2805 29212
rect 2763 29203 2764 29210
rect 2804 29203 2805 29210
rect 2764 29161 2804 29170
rect 2956 29168 2996 29179
rect 2956 29093 2996 29128
rect 3052 29168 3092 30052
rect 3339 29924 3381 29933
rect 3339 29884 3340 29924
rect 3380 29884 3381 29924
rect 3339 29875 3381 29884
rect 3627 29924 3669 29933
rect 3627 29884 3628 29924
rect 3668 29884 3669 29924
rect 3627 29875 3669 29884
rect 3243 29252 3285 29261
rect 3243 29212 3244 29252
rect 3284 29212 3285 29252
rect 3243 29203 3285 29212
rect 3052 29119 3092 29128
rect 3244 29118 3284 29203
rect 3340 29168 3380 29875
rect 3628 29790 3668 29875
rect 3724 29672 3764 30295
rect 4107 30008 4149 30017
rect 4107 29968 4108 30008
rect 4148 29968 4149 30008
rect 4107 29959 4149 29968
rect 3819 29840 3861 29849
rect 3819 29800 3820 29840
rect 3860 29800 3861 29840
rect 3819 29791 3861 29800
rect 4108 29840 4148 29959
rect 3340 29119 3380 29128
rect 3436 29632 3764 29672
rect 3436 29168 3476 29632
rect 3531 29252 3573 29261
rect 3531 29212 3532 29252
rect 3572 29212 3573 29252
rect 3531 29203 3573 29212
rect 3436 29119 3476 29128
rect 3532 29168 3572 29203
rect 3724 29177 3764 29262
rect 3532 29117 3572 29128
rect 3723 29168 3765 29177
rect 3723 29128 3724 29168
rect 3764 29128 3765 29168
rect 3723 29119 3765 29128
rect 2955 29084 2997 29093
rect 2955 29044 2956 29084
rect 2996 29044 2997 29084
rect 2955 29035 2997 29044
rect 2763 29000 2805 29009
rect 3820 29000 3860 29791
rect 4012 29672 4052 29681
rect 3915 29168 3957 29177
rect 3915 29128 3916 29168
rect 3956 29128 3957 29168
rect 3915 29119 3957 29128
rect 2763 28960 2764 29000
rect 2804 28960 2805 29000
rect 2763 28951 2805 28960
rect 3724 28960 3860 29000
rect 2764 28866 2804 28951
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3724 28580 3764 28960
rect 3724 28531 3764 28540
rect 3819 28496 3861 28505
rect 3819 28456 3820 28496
rect 3860 28456 3861 28496
rect 3819 28447 3861 28456
rect 3820 27824 3860 28447
rect 3916 28160 3956 29119
rect 4012 28328 4052 29632
rect 4108 29429 4148 29800
rect 4204 29840 4244 30388
rect 4204 29791 4244 29800
rect 4300 29840 4340 30472
rect 4396 30017 4436 30556
rect 4683 30512 4725 30521
rect 4683 30472 4684 30512
rect 4724 30472 4725 30512
rect 4683 30463 4725 30472
rect 4395 30008 4437 30017
rect 4395 29968 4396 30008
rect 4436 29968 4437 30008
rect 4395 29959 4437 29968
rect 4300 29672 4340 29800
rect 4588 29840 4628 29849
rect 4588 29681 4628 29800
rect 4684 29840 4724 30463
rect 4780 29849 4820 30640
rect 5548 30017 5588 30640
rect 6123 30512 6165 30521
rect 6123 30472 6124 30512
rect 6164 30472 6165 30512
rect 6123 30463 6165 30472
rect 5932 30428 5972 30439
rect 5932 30353 5972 30388
rect 5931 30344 5973 30353
rect 5931 30304 5932 30344
rect 5972 30304 5973 30344
rect 5931 30295 5973 30304
rect 5547 30008 5589 30017
rect 5547 29968 5548 30008
rect 5588 29968 5589 30008
rect 5547 29959 5589 29968
rect 5835 30008 5877 30017
rect 5835 29968 5836 30008
rect 5876 29968 5877 30008
rect 5835 29959 5877 29968
rect 5067 29924 5109 29933
rect 5067 29884 5068 29924
rect 5108 29884 5109 29924
rect 5067 29875 5109 29884
rect 4684 29791 4724 29800
rect 4779 29840 4821 29849
rect 4779 29800 4780 29840
rect 4820 29800 4821 29840
rect 4779 29791 4821 29800
rect 5068 29790 5108 29875
rect 5163 29840 5205 29849
rect 5163 29800 5164 29840
rect 5204 29800 5205 29840
rect 5163 29791 5205 29800
rect 5643 29840 5685 29849
rect 5643 29800 5644 29840
rect 5684 29800 5685 29840
rect 5643 29791 5685 29800
rect 5164 29706 5204 29791
rect 5644 29706 5684 29791
rect 4204 29632 4340 29672
rect 4587 29672 4629 29681
rect 4587 29632 4588 29672
rect 4628 29632 4629 29672
rect 4107 29420 4149 29429
rect 4107 29380 4108 29420
rect 4148 29380 4149 29420
rect 4107 29371 4149 29380
rect 4204 29261 4244 29632
rect 4587 29623 4629 29632
rect 5259 29672 5301 29681
rect 5259 29632 5260 29672
rect 5300 29632 5301 29672
rect 5259 29623 5301 29632
rect 4352 29504 4720 29513
rect 5260 29504 5300 29623
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 5255 29464 5300 29504
rect 5255 29261 5295 29464
rect 5643 29420 5685 29429
rect 5643 29380 5644 29420
rect 5684 29380 5685 29420
rect 5643 29371 5685 29380
rect 5355 29336 5397 29345
rect 5355 29296 5356 29336
rect 5396 29296 5397 29336
rect 5355 29287 5397 29296
rect 5547 29336 5589 29345
rect 5547 29296 5548 29336
rect 5588 29296 5589 29336
rect 5547 29287 5589 29296
rect 4203 29252 4245 29261
rect 4203 29212 4204 29252
rect 4244 29212 4245 29252
rect 4203 29203 4245 29212
rect 5163 29252 5205 29261
rect 5163 29212 5164 29252
rect 5204 29212 5205 29252
rect 5255 29252 5300 29261
rect 5255 29212 5260 29252
rect 5163 29203 5205 29212
rect 5260 29203 5300 29212
rect 4204 28505 4244 29203
rect 4683 29168 4725 29177
rect 4683 29128 4684 29168
rect 4724 29128 4725 29168
rect 4683 29119 4725 29128
rect 5068 29168 5108 29177
rect 4684 29034 4724 29119
rect 4203 28496 4245 28505
rect 4203 28456 4204 28496
rect 4244 28456 4245 28496
rect 4203 28447 4245 28456
rect 4875 28496 4917 28505
rect 4875 28456 4876 28496
rect 4916 28456 4917 28496
rect 4875 28447 4917 28456
rect 4012 28279 4052 28288
rect 4204 28328 4244 28447
rect 4300 28337 4340 28422
rect 4204 28279 4244 28288
rect 4299 28328 4341 28337
rect 4299 28288 4300 28328
rect 4340 28288 4341 28328
rect 4299 28279 4341 28288
rect 4107 28244 4149 28253
rect 4107 28204 4108 28244
rect 4148 28204 4149 28244
rect 4107 28195 4149 28204
rect 3916 28120 4052 28160
rect 3628 27784 3860 27824
rect 2668 27691 2708 27700
rect 3051 27740 3093 27749
rect 3051 27700 3052 27740
rect 3092 27700 3093 27740
rect 3051 27691 3093 27700
rect 2764 27656 2804 27665
rect 2764 27329 2804 27616
rect 3052 27656 3092 27691
rect 3340 27665 3380 27750
rect 3052 27605 3092 27616
rect 3339 27656 3381 27665
rect 3339 27616 3340 27656
rect 3380 27616 3381 27656
rect 3339 27607 3381 27616
rect 3532 27656 3572 27665
rect 3244 27488 3284 27497
rect 3532 27488 3572 27616
rect 3284 27448 3572 27488
rect 3628 27656 3668 27784
rect 3244 27439 3284 27448
rect 2955 27404 2997 27413
rect 2955 27364 2956 27404
rect 2996 27364 2997 27404
rect 2955 27355 2997 27364
rect 2763 27320 2805 27329
rect 2763 27280 2764 27320
rect 2804 27280 2805 27320
rect 2763 27271 2805 27280
rect 2956 27270 2996 27355
rect 3628 27245 3668 27616
rect 3723 27656 3765 27665
rect 3723 27616 3724 27656
rect 3764 27616 3765 27656
rect 3723 27607 3765 27616
rect 3820 27656 3860 27665
rect 4012 27656 4052 28120
rect 4108 28110 4148 28195
rect 4492 28160 4532 28169
rect 4204 28120 4492 28160
rect 4204 27833 4244 28120
rect 4492 28111 4532 28120
rect 4779 28076 4821 28085
rect 4779 28036 4780 28076
rect 4820 28036 4821 28076
rect 4779 28027 4821 28036
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4203 27824 4245 27833
rect 4203 27784 4204 27824
rect 4244 27784 4245 27824
rect 4203 27775 4245 27784
rect 4683 27824 4725 27833
rect 4683 27784 4684 27824
rect 4724 27784 4725 27824
rect 4683 27775 4725 27784
rect 4684 27690 4724 27775
rect 4204 27656 4244 27665
rect 3860 27616 3956 27656
rect 4012 27616 4204 27656
rect 3820 27607 3860 27616
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3627 27236 3669 27245
rect 3627 27196 3628 27236
rect 3668 27196 3669 27236
rect 3627 27187 3669 27196
rect 3627 27068 3669 27077
rect 3627 27028 3628 27068
rect 3668 27028 3669 27068
rect 3627 27019 3669 27028
rect 3628 26934 3668 27019
rect 1612 26767 1652 26776
rect 1228 26682 1268 26767
rect 1227 26228 1269 26237
rect 1227 26188 1228 26228
rect 1268 26188 1269 26228
rect 1227 26179 1269 26188
rect 1228 26094 1268 26179
rect 1612 26144 1652 26153
rect 1612 25985 1652 26104
rect 2476 26144 2516 26776
rect 3724 26648 3764 27607
rect 3820 27404 3860 27413
rect 3820 26825 3860 27364
rect 3819 26816 3861 26825
rect 3819 26776 3820 26816
rect 3860 26776 3861 26816
rect 3819 26767 3861 26776
rect 3820 26648 3860 26657
rect 3724 26608 3820 26648
rect 3627 26312 3669 26321
rect 3627 26272 3628 26312
rect 3668 26272 3669 26312
rect 3627 26263 3669 26272
rect 3628 26178 3668 26263
rect 3724 26144 3764 26608
rect 3820 26599 3860 26608
rect 3916 26480 3956 27616
rect 4204 27607 4244 27616
rect 4011 27488 4053 27497
rect 4011 27448 4012 27488
rect 4052 27448 4053 27488
rect 4011 27439 4053 27448
rect 3820 26440 3956 26480
rect 3820 26312 3860 26440
rect 3820 26263 3860 26272
rect 4012 26165 4052 27439
rect 4107 27236 4149 27245
rect 4107 27196 4108 27236
rect 4148 27196 4149 27236
rect 4107 27187 4149 27196
rect 3724 26104 3860 26144
rect 4012 26116 4052 26125
rect 4108 26144 4148 27187
rect 4684 27068 4724 27077
rect 4780 27068 4820 28027
rect 4876 27833 4916 28447
rect 4875 27824 4917 27833
rect 4875 27784 4876 27824
rect 4916 27784 4917 27824
rect 4875 27775 4917 27784
rect 5068 27413 5108 29128
rect 5164 29168 5204 29203
rect 5164 29117 5204 29128
rect 5356 29168 5396 29287
rect 5548 29202 5588 29287
rect 5356 29119 5396 29128
rect 5644 29168 5684 29371
rect 5739 29336 5781 29345
rect 5739 29296 5740 29336
rect 5780 29296 5781 29336
rect 5739 29287 5781 29296
rect 5644 29119 5684 29128
rect 5740 29168 5780 29287
rect 5836 29261 5876 29959
rect 6124 29854 6164 30463
rect 6124 29805 6164 29814
rect 6027 29336 6069 29345
rect 6027 29296 6028 29336
rect 6068 29296 6069 29336
rect 6027 29287 6069 29296
rect 5835 29252 5877 29261
rect 5835 29212 5836 29252
rect 5876 29212 5877 29252
rect 5835 29203 5877 29212
rect 5740 29119 5780 29128
rect 5836 29168 5876 29203
rect 6028 29202 6068 29287
rect 6220 29177 6260 31312
rect 6604 30680 6644 30691
rect 6604 30605 6644 30640
rect 6892 30680 6932 31387
rect 6988 31352 7028 31361
rect 7028 31312 7124 31352
rect 6988 31303 7028 31312
rect 6892 30631 6932 30640
rect 6987 30680 7029 30689
rect 6987 30640 6988 30680
rect 7028 30640 7029 30680
rect 6987 30631 7029 30640
rect 6603 30596 6645 30605
rect 6603 30556 6604 30596
rect 6644 30556 6645 30596
rect 6603 30547 6645 30556
rect 6988 30546 7028 30631
rect 6508 29840 6548 29849
rect 6508 29681 6548 29800
rect 6316 29672 6356 29681
rect 6316 29513 6356 29632
rect 6507 29672 6549 29681
rect 6507 29632 6508 29672
rect 6548 29632 6549 29672
rect 6507 29623 6549 29632
rect 6315 29504 6357 29513
rect 6315 29464 6316 29504
rect 6356 29464 6357 29504
rect 6315 29455 6357 29464
rect 7084 29420 7124 31312
rect 7180 30689 7220 33571
rect 7852 33377 7892 33664
rect 8620 33704 8660 33713
rect 8908 33704 8948 33991
rect 9003 33872 9045 33881
rect 9003 33832 9004 33872
rect 9044 33832 9045 33872
rect 9003 33823 9045 33832
rect 9196 33872 9236 34336
rect 9388 34376 9428 34385
rect 9388 34217 9428 34336
rect 9580 34376 9620 34385
rect 9387 34208 9429 34217
rect 9387 34168 9388 34208
rect 9428 34168 9429 34208
rect 9387 34159 9429 34168
rect 9580 33881 9620 34336
rect 10251 34376 10293 34385
rect 10251 34336 10252 34376
rect 10292 34336 10293 34376
rect 10251 34327 10293 34336
rect 10252 34242 10292 34327
rect 9484 33872 9524 33881
rect 9196 33832 9484 33872
rect 9004 33788 9044 33823
rect 9004 33737 9044 33748
rect 9196 33713 9236 33832
rect 9484 33823 9524 33832
rect 9579 33872 9621 33881
rect 9579 33832 9580 33872
rect 9620 33832 9621 33872
rect 9579 33823 9621 33832
rect 10540 33713 10580 35176
rect 10923 35167 10965 35176
rect 10924 34628 10964 35167
rect 11691 35132 11733 35141
rect 11691 35092 11692 35132
rect 11732 35092 11733 35132
rect 11691 35083 11733 35092
rect 11692 34998 11732 35083
rect 12076 35057 12116 35142
rect 12075 35048 12117 35057
rect 12075 35008 12076 35048
rect 12116 35008 12117 35048
rect 12652 35048 12692 36016
rect 12748 35888 12788 35897
rect 12940 35888 12980 36436
rect 13036 36427 13076 36436
rect 12788 35848 12980 35888
rect 13132 35888 13172 36511
rect 13227 36476 13269 36485
rect 13227 36436 13228 36476
rect 13268 36436 13269 36476
rect 13227 36427 13269 36436
rect 12748 35839 12788 35848
rect 13132 35839 13172 35848
rect 12939 35720 12981 35729
rect 12939 35680 12940 35720
rect 12980 35680 12981 35720
rect 12939 35671 12981 35680
rect 12940 35309 12980 35671
rect 12939 35300 12981 35309
rect 12939 35260 12940 35300
rect 12980 35260 12981 35300
rect 12939 35251 12981 35260
rect 12940 35216 12980 35251
rect 12940 35166 12980 35176
rect 12652 35008 12980 35048
rect 12075 34999 12117 35008
rect 11595 34964 11637 34973
rect 12268 34964 12308 34973
rect 11595 34924 11596 34964
rect 11636 34924 11637 34964
rect 11595 34915 11637 34924
rect 12172 34924 12268 34964
rect 10924 34579 10964 34588
rect 10827 34376 10869 34385
rect 10827 34336 10828 34376
rect 10868 34336 10869 34376
rect 10827 34327 10869 34336
rect 11211 34376 11253 34385
rect 11211 34336 11212 34376
rect 11252 34336 11253 34376
rect 11211 34327 11253 34336
rect 11500 34376 11540 34385
rect 10828 34242 10868 34327
rect 11212 34242 11252 34327
rect 11500 34301 11540 34336
rect 11596 34376 11636 34915
rect 12172 34880 12212 34924
rect 12268 34915 12308 34924
rect 12076 34840 12212 34880
rect 11883 34628 11925 34637
rect 11883 34588 11884 34628
rect 11924 34588 11925 34628
rect 11883 34579 11925 34588
rect 11691 34460 11733 34469
rect 11691 34420 11692 34460
rect 11732 34420 11733 34460
rect 11691 34411 11733 34420
rect 11596 34327 11636 34336
rect 11692 34376 11732 34411
rect 11499 34292 11541 34301
rect 11499 34252 11500 34292
rect 11540 34252 11541 34292
rect 11499 34243 11541 34252
rect 11116 34208 11156 34217
rect 10635 34124 10677 34133
rect 10635 34084 10636 34124
rect 10676 34084 10677 34124
rect 10635 34075 10677 34084
rect 8660 33664 8756 33704
rect 8620 33655 8660 33664
rect 7851 33368 7893 33377
rect 7851 33328 7852 33368
rect 7892 33328 7893 33368
rect 7851 33319 7893 33328
rect 7563 32948 7605 32957
rect 7563 32908 7564 32948
rect 7604 32908 7605 32948
rect 7563 32899 7605 32908
rect 7276 32864 7316 32873
rect 7276 32789 7316 32824
rect 7275 32780 7317 32789
rect 7275 32740 7276 32780
rect 7316 32740 7317 32780
rect 7275 32731 7317 32740
rect 7276 32360 7316 32731
rect 7372 32360 7412 32369
rect 7276 32320 7372 32360
rect 7372 32311 7412 32320
rect 7564 32360 7604 32899
rect 7659 32696 7701 32705
rect 7659 32656 7660 32696
rect 7700 32656 7701 32696
rect 7659 32647 7701 32656
rect 7564 32311 7604 32320
rect 7660 32192 7700 32647
rect 7852 32192 7892 33319
rect 8235 33200 8277 33209
rect 8235 33160 8236 33200
rect 8276 33160 8277 33200
rect 8235 33151 8277 33160
rect 8139 33032 8181 33041
rect 8139 32992 8140 33032
rect 8180 32992 8181 33032
rect 8139 32983 8181 32992
rect 8043 32864 8085 32873
rect 8043 32824 8044 32864
rect 8084 32824 8085 32864
rect 8043 32815 8085 32824
rect 8140 32864 8180 32983
rect 8236 32873 8276 33151
rect 8140 32815 8180 32824
rect 8235 32864 8277 32873
rect 8235 32824 8236 32864
rect 8276 32824 8277 32864
rect 8235 32815 8277 32824
rect 7947 32696 7989 32705
rect 7947 32656 7948 32696
rect 7988 32656 7989 32696
rect 7947 32647 7989 32656
rect 7948 32562 7988 32647
rect 7948 32360 7988 32369
rect 8044 32360 8084 32815
rect 7988 32320 8084 32360
rect 7948 32311 7988 32320
rect 8044 32192 8084 32201
rect 7852 32152 8044 32192
rect 7660 32143 7700 32152
rect 8044 32143 8084 32152
rect 8139 32192 8181 32201
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8236 32192 8276 32815
rect 8427 32780 8469 32789
rect 8427 32740 8428 32780
rect 8468 32740 8469 32780
rect 8427 32731 8469 32740
rect 8428 32276 8468 32731
rect 8428 32227 8468 32236
rect 8236 32143 8276 32152
rect 8140 32058 8180 32143
rect 7372 31940 7412 31949
rect 7412 31900 7508 31940
rect 7372 31891 7412 31900
rect 7372 31520 7412 31529
rect 7276 31480 7372 31520
rect 7179 30680 7221 30689
rect 7179 30640 7180 30680
rect 7220 30640 7221 30680
rect 7179 30631 7221 30640
rect 7179 29672 7221 29681
rect 7179 29632 7180 29672
rect 7220 29632 7221 29672
rect 7179 29623 7221 29632
rect 7180 29538 7220 29623
rect 7084 29380 7220 29420
rect 5836 29118 5876 29128
rect 6219 29168 6261 29177
rect 6219 29128 6220 29168
rect 6260 29128 6261 29168
rect 6219 29119 6261 29128
rect 7180 29168 7220 29380
rect 7276 29177 7316 31480
rect 7372 31471 7412 31480
rect 7468 31352 7508 31900
rect 7659 31520 7701 31529
rect 7659 31480 7660 31520
rect 7700 31480 7701 31520
rect 7659 31471 7701 31480
rect 7852 31520 7892 31529
rect 8331 31520 8373 31529
rect 7892 31480 8276 31520
rect 7852 31471 7892 31480
rect 7660 31386 7700 31471
rect 7372 31312 7508 31352
rect 7564 31352 7604 31361
rect 7372 30680 7412 31312
rect 7372 30631 7412 30640
rect 7467 30596 7509 30605
rect 7467 30556 7468 30596
rect 7508 30556 7509 30596
rect 7467 30547 7509 30556
rect 7468 30462 7508 30547
rect 7564 30353 7604 31312
rect 7948 31352 7988 31361
rect 7948 30848 7988 31312
rect 8236 31268 8276 31480
rect 8331 31480 8332 31520
rect 8372 31480 8373 31520
rect 8331 31471 8373 31480
rect 8332 31386 8372 31471
rect 8716 31445 8756 33664
rect 8908 33655 8948 33664
rect 9195 33704 9237 33713
rect 9195 33664 9196 33704
rect 9236 33664 9237 33704
rect 9195 33655 9237 33664
rect 10444 33704 10484 33713
rect 9676 33620 9716 33629
rect 9292 33452 9332 33461
rect 9292 32957 9332 33412
rect 9291 32948 9333 32957
rect 9291 32908 9292 32948
rect 9332 32908 9333 32948
rect 9291 32899 9333 32908
rect 9676 32873 9716 33580
rect 9867 33116 9909 33125
rect 9867 33076 9868 33116
rect 9908 33076 9909 33116
rect 9867 33067 9909 33076
rect 9003 32864 9045 32873
rect 9003 32824 9004 32864
rect 9044 32824 9045 32864
rect 9003 32815 9045 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9675 32815 9717 32824
rect 8811 32780 8853 32789
rect 8811 32740 8812 32780
rect 8852 32740 8853 32780
rect 8811 32731 8853 32740
rect 8812 32646 8852 32731
rect 9004 32730 9044 32815
rect 8812 32192 8852 32201
rect 8812 31529 8852 32152
rect 9676 32192 9716 32201
rect 9676 31781 9716 32152
rect 9675 31772 9717 31781
rect 9675 31732 9676 31772
rect 9716 31732 9717 31772
rect 9675 31723 9717 31732
rect 8811 31520 8853 31529
rect 8811 31480 8812 31520
rect 8852 31480 8853 31520
rect 9868 31520 9908 33067
rect 10444 32873 10484 33664
rect 10539 33704 10581 33713
rect 10539 33664 10540 33704
rect 10580 33664 10581 33704
rect 10539 33655 10581 33664
rect 10636 33704 10676 34075
rect 10636 33655 10676 33664
rect 10924 33452 10964 33461
rect 9963 32864 10005 32873
rect 9963 32824 9964 32864
rect 10004 32824 10005 32864
rect 9963 32815 10005 32824
rect 10252 32864 10292 32873
rect 10443 32864 10485 32873
rect 10292 32824 10388 32864
rect 10252 32815 10292 32824
rect 9964 32730 10004 32815
rect 9964 31520 10004 31529
rect 9868 31480 9964 31520
rect 8811 31471 8853 31480
rect 9964 31471 10004 31480
rect 8715 31436 8757 31445
rect 8715 31396 8716 31436
rect 8756 31396 8757 31436
rect 8715 31387 8757 31396
rect 8524 31352 8564 31361
rect 8524 31268 8564 31312
rect 8236 31228 8564 31268
rect 8620 31352 8660 31361
rect 8331 31016 8373 31025
rect 8331 30976 8332 31016
rect 8372 30976 8373 31016
rect 8331 30967 8373 30976
rect 7948 30808 8084 30848
rect 7948 30680 7988 30689
rect 7563 30344 7605 30353
rect 7563 30304 7564 30344
rect 7604 30304 7605 30344
rect 7563 30295 7605 30304
rect 7851 30260 7893 30269
rect 7851 30220 7852 30260
rect 7892 30220 7893 30260
rect 7851 30211 7893 30220
rect 7563 30008 7605 30017
rect 7563 29968 7564 30008
rect 7604 29968 7605 30008
rect 7563 29959 7605 29968
rect 7564 29840 7604 29959
rect 7564 29791 7604 29800
rect 7659 29840 7701 29849
rect 7659 29800 7660 29840
rect 7700 29800 7701 29840
rect 7659 29791 7701 29800
rect 7756 29840 7796 29849
rect 7660 29706 7700 29791
rect 6123 29084 6165 29093
rect 6123 29044 6124 29084
rect 6164 29044 6165 29084
rect 6123 29035 6165 29044
rect 5163 28328 5205 28337
rect 5163 28288 5164 28328
rect 5204 28288 5205 28328
rect 5163 28279 5205 28288
rect 5356 28328 5396 28337
rect 5067 27404 5109 27413
rect 5067 27364 5068 27404
rect 5108 27364 5109 27404
rect 5067 27355 5109 27364
rect 5164 27077 5204 28279
rect 5356 28085 5396 28288
rect 6027 28160 6069 28169
rect 6027 28120 6028 28160
rect 6068 28120 6069 28160
rect 6027 28111 6069 28120
rect 5355 28076 5397 28085
rect 5355 28036 5356 28076
rect 5396 28036 5397 28076
rect 5355 28027 5397 28036
rect 6028 28026 6068 28111
rect 5931 27656 5973 27665
rect 5931 27616 5932 27656
rect 5972 27616 5973 27656
rect 5931 27607 5973 27616
rect 5644 27572 5684 27581
rect 5452 27404 5492 27413
rect 4724 27028 4820 27068
rect 5163 27068 5205 27077
rect 5163 27028 5164 27068
rect 5204 27028 5205 27068
rect 4684 27019 4724 27028
rect 5163 27019 5205 27028
rect 4492 26816 4532 26825
rect 4532 26776 4820 26816
rect 4492 26767 4532 26776
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4587 26312 4629 26321
rect 4587 26272 4588 26312
rect 4628 26272 4629 26312
rect 4587 26263 4629 26272
rect 4395 26228 4437 26237
rect 4395 26188 4396 26228
rect 4436 26188 4437 26228
rect 4395 26179 4437 26188
rect 4300 26144 4340 26153
rect 2476 26095 2516 26104
rect 1035 25976 1077 25985
rect 1035 25936 1036 25976
rect 1076 25936 1077 25976
rect 1035 25927 1077 25936
rect 1611 25976 1653 25985
rect 1611 25936 1612 25976
rect 1652 25936 1653 25976
rect 3820 25976 3860 26104
rect 3916 26102 3956 26111
rect 4108 26095 4148 26104
rect 4204 26104 4300 26144
rect 3916 26060 3956 26062
rect 3916 26020 4052 26060
rect 3820 25936 3956 25976
rect 1611 25927 1653 25936
rect 1036 25842 1076 25927
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 1612 25472 1652 25481
rect 1131 24632 1173 24641
rect 1131 24592 1132 24632
rect 1172 24592 1173 24632
rect 1131 24583 1173 24592
rect 1516 24632 1556 24641
rect 1612 24632 1652 25432
rect 3435 25388 3477 25397
rect 3435 25348 3436 25388
rect 3476 25348 3477 25388
rect 3435 25339 3477 25348
rect 3436 25304 3476 25339
rect 3436 25253 3476 25264
rect 3531 25304 3573 25313
rect 3531 25264 3532 25304
rect 3572 25264 3573 25304
rect 3531 25255 3573 25264
rect 3628 25304 3668 25315
rect 2667 25220 2709 25229
rect 2667 25180 2668 25220
rect 2708 25180 2709 25220
rect 2667 25171 2709 25180
rect 1556 24592 1652 24632
rect 2380 24632 2420 24641
rect 2420 24592 2516 24632
rect 1516 24583 1556 24592
rect 2380 24583 2420 24592
rect 1132 24498 1172 24583
rect 1708 23960 1748 23969
rect 1612 23920 1708 23960
rect 1227 23204 1269 23213
rect 1227 23164 1228 23204
rect 1268 23164 1269 23204
rect 1227 23155 1269 23164
rect 1228 23070 1268 23155
rect 1612 23120 1652 23920
rect 1708 23911 1748 23920
rect 2379 23876 2421 23885
rect 2379 23836 2380 23876
rect 2420 23836 2421 23876
rect 2379 23827 2421 23836
rect 2283 23792 2325 23801
rect 2283 23752 2284 23792
rect 2324 23752 2325 23792
rect 2283 23743 2325 23752
rect 2380 23792 2420 23827
rect 2284 23658 2324 23743
rect 2380 23741 2420 23752
rect 1612 23071 1652 23080
rect 2476 23120 2516 24592
rect 2571 23792 2613 23801
rect 2571 23752 2572 23792
rect 2612 23752 2613 23792
rect 2571 23743 2613 23752
rect 2668 23792 2708 25171
rect 3532 25170 3572 25255
rect 3628 25229 3668 25264
rect 3820 25304 3860 25313
rect 3627 25220 3669 25229
rect 3627 25180 3628 25220
rect 3668 25180 3669 25220
rect 3627 25171 3669 25180
rect 3340 25136 3380 25145
rect 2860 25096 3340 25136
rect 2763 24632 2805 24641
rect 2763 24592 2764 24632
rect 2804 24592 2805 24632
rect 2763 24583 2805 24592
rect 2668 23743 2708 23752
rect 2572 23658 2612 23743
rect 2764 23708 2804 24583
rect 2860 23792 2900 25096
rect 3340 25087 3380 25096
rect 3531 24548 3573 24557
rect 3531 24508 3532 24548
rect 3572 24508 3573 24548
rect 3531 24499 3573 24508
rect 3532 24414 3572 24499
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3531 23960 3573 23969
rect 3531 23920 3532 23960
rect 3572 23920 3573 23960
rect 3531 23911 3573 23920
rect 3532 23826 3572 23911
rect 3820 23885 3860 25264
rect 3916 25304 3956 25936
rect 4012 25733 4052 26020
rect 4011 25724 4053 25733
rect 4011 25684 4012 25724
rect 4052 25684 4053 25724
rect 4011 25675 4053 25684
rect 4012 25397 4052 25675
rect 4011 25388 4053 25397
rect 4011 25348 4012 25388
rect 4052 25348 4053 25388
rect 4011 25339 4053 25348
rect 3916 25255 3956 25264
rect 4012 25304 4052 25339
rect 4012 24053 4052 25264
rect 4108 25304 4148 25313
rect 4204 25304 4244 26104
rect 4300 26095 4340 26104
rect 4396 26094 4436 26179
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 4588 26144 4628 26263
rect 4780 26237 4820 26776
rect 4779 26228 4821 26237
rect 4779 26188 4780 26228
rect 4820 26188 4821 26228
rect 4779 26179 4821 26188
rect 5452 26153 5492 27364
rect 5644 26741 5684 27532
rect 5932 27522 5972 27607
rect 5836 27404 5876 27413
rect 5740 27364 5836 27404
rect 5643 26732 5685 26741
rect 5643 26692 5644 26732
rect 5684 26692 5685 26732
rect 5643 26683 5685 26692
rect 5740 26321 5780 27364
rect 5836 27355 5876 27364
rect 5836 26816 5876 26825
rect 6124 26816 6164 29035
rect 6220 29000 6260 29119
rect 7180 29093 7220 29128
rect 7275 29168 7317 29177
rect 7275 29128 7276 29168
rect 7316 29128 7317 29168
rect 7275 29119 7317 29128
rect 7179 29084 7221 29093
rect 7179 29044 7180 29084
rect 7220 29044 7221 29084
rect 7179 29035 7221 29044
rect 7371 29084 7413 29093
rect 7371 29044 7372 29084
rect 7412 29044 7413 29084
rect 7371 29035 7413 29044
rect 7180 29004 7220 29035
rect 6220 28960 6356 29000
rect 5876 26776 6164 26816
rect 5836 26767 5876 26776
rect 5739 26312 5781 26321
rect 5739 26272 5740 26312
rect 5780 26272 5781 26312
rect 5739 26263 5781 26272
rect 4972 26144 5012 26153
rect 4588 26095 4628 26104
rect 4876 26104 4972 26144
rect 4395 25388 4437 25397
rect 4395 25348 4396 25388
rect 4436 25348 4437 25388
rect 4395 25339 4437 25348
rect 4148 25264 4244 25304
rect 4300 25304 4340 25313
rect 4108 25255 4148 25264
rect 4300 25136 4340 25264
rect 4396 25145 4436 25339
rect 4492 25229 4532 26095
rect 4779 25304 4821 25313
rect 4779 25264 4780 25304
rect 4820 25264 4821 25304
rect 4779 25255 4821 25264
rect 4491 25220 4533 25229
rect 4491 25180 4492 25220
rect 4532 25180 4533 25220
rect 4491 25171 4533 25180
rect 4108 25096 4340 25136
rect 4395 25136 4437 25145
rect 4395 25096 4396 25136
rect 4436 25096 4437 25136
rect 4108 24557 4148 25096
rect 4395 25087 4437 25096
rect 4203 24968 4245 24977
rect 4203 24928 4204 24968
rect 4244 24928 4245 24968
rect 4203 24919 4245 24928
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4204 24632 4244 24919
rect 4107 24548 4149 24557
rect 4107 24508 4108 24548
rect 4148 24508 4149 24548
rect 4107 24499 4149 24508
rect 4204 24380 4244 24592
rect 4492 24632 4532 24643
rect 4492 24557 4532 24592
rect 4588 24632 4628 24641
rect 4491 24548 4533 24557
rect 4491 24508 4492 24548
rect 4532 24508 4533 24548
rect 4491 24499 4533 24508
rect 4108 24340 4244 24380
rect 4011 24044 4053 24053
rect 4011 24004 4012 24044
rect 4052 24004 4053 24044
rect 4011 23995 4053 24004
rect 3819 23876 3861 23885
rect 3819 23836 3820 23876
rect 3860 23836 3861 23876
rect 3819 23827 3861 23836
rect 2860 23743 2900 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3051 23743 3093 23752
rect 3244 23792 3284 23801
rect 2764 23659 2804 23668
rect 3052 23658 3092 23743
rect 3148 23624 3188 23633
rect 3148 23213 3188 23584
rect 3147 23204 3189 23213
rect 3147 23164 3148 23204
rect 3188 23164 3189 23204
rect 3147 23155 3189 23164
rect 652 23036 692 23045
rect 652 22457 692 22996
rect 844 22868 884 22877
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 652 22112 692 22121
rect 652 21617 692 22072
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 267 20936 309 20945
rect 267 20896 268 20936
rect 308 20896 309 20936
rect 267 20887 309 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 652 20600 692 20719
rect 652 20551 692 20560
rect 652 20264 692 20273
rect 652 19937 692 20224
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18954 692 19039
rect 652 18752 692 18761
rect 652 18257 692 18712
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17576 692 17585
rect 652 17417 692 17536
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 17240 692 17249
rect 652 16577 692 17200
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16064 692 16073
rect 652 15737 692 16024
rect 844 15821 884 22828
rect 1227 22868 1269 22877
rect 1227 22828 1228 22868
rect 1268 22828 1269 22868
rect 1227 22819 1269 22828
rect 1228 22280 1268 22819
rect 2476 22289 2516 23080
rect 3244 23036 3284 23752
rect 3340 23792 3380 23801
rect 3340 23297 3380 23752
rect 3627 23792 3669 23801
rect 3627 23752 3628 23792
rect 3668 23752 3669 23792
rect 3627 23743 3669 23752
rect 3339 23288 3381 23297
rect 3339 23248 3340 23288
rect 3380 23248 3381 23288
rect 3339 23239 3381 23248
rect 3628 23288 3668 23743
rect 4012 23708 4052 23995
rect 3628 23239 3668 23248
rect 3820 23668 4052 23708
rect 2956 22996 3284 23036
rect 1228 22231 1268 22240
rect 1612 22280 1652 22289
rect 1612 21440 1652 22240
rect 2475 22280 2517 22289
rect 2475 22240 2476 22280
rect 2516 22240 2517 22280
rect 2475 22231 2517 22240
rect 2476 22146 2516 22231
rect 2859 22196 2901 22205
rect 2956 22196 2996 22996
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3628 22364 3668 22375
rect 3628 22289 3668 22324
rect 3147 22280 3189 22289
rect 3147 22240 3148 22280
rect 3188 22240 3189 22280
rect 3147 22231 3189 22240
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3820 22280 3860 23668
rect 3915 23540 3957 23549
rect 4108 23540 4148 24340
rect 4588 24296 4628 24592
rect 4300 24256 4628 24296
rect 4204 23801 4244 23886
rect 4203 23792 4245 23801
rect 4300 23792 4340 24256
rect 4780 24128 4820 25255
rect 4876 24884 4916 26104
rect 4972 26095 5012 26104
rect 5067 26144 5109 26153
rect 5260 26144 5300 26153
rect 5067 26104 5068 26144
rect 5108 26104 5109 26144
rect 5067 26095 5109 26104
rect 5164 26104 5260 26144
rect 5068 26010 5108 26095
rect 4971 25304 5013 25313
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 5164 25304 5204 26104
rect 5260 26095 5300 26104
rect 5451 26144 5493 26153
rect 5451 26104 5452 26144
rect 5492 26104 5493 26144
rect 5451 26095 5493 26104
rect 5548 26104 5876 26144
rect 5260 25976 5300 25985
rect 5548 25976 5588 26104
rect 5300 25936 5588 25976
rect 5644 25976 5684 25985
rect 5260 25927 5300 25936
rect 5164 25264 5300 25304
rect 4971 25255 5013 25264
rect 4972 25170 5012 25255
rect 5164 25136 5204 25145
rect 4876 24844 5012 24884
rect 4875 24380 4917 24389
rect 4875 24340 4876 24380
rect 4916 24340 4917 24380
rect 4875 24331 4917 24340
rect 4876 24246 4916 24331
rect 4780 24088 4916 24128
rect 4395 24044 4437 24053
rect 4395 24004 4396 24044
rect 4436 24004 4437 24044
rect 4395 23995 4437 24004
rect 4396 23876 4436 23995
rect 4683 23876 4725 23885
rect 4396 23836 4532 23876
rect 4203 23752 4204 23792
rect 4244 23752 4245 23792
rect 4203 23743 4245 23752
rect 4299 23752 4340 23792
rect 4492 23792 4532 23836
rect 4683 23836 4684 23876
rect 4724 23836 4725 23876
rect 4683 23827 4725 23836
rect 4299 23708 4339 23752
rect 4492 23743 4532 23752
rect 4588 23792 4628 23801
rect 4299 23668 4340 23708
rect 4300 23624 4340 23668
rect 4396 23633 4436 23718
rect 4588 23633 4628 23752
rect 4684 23792 4724 23827
rect 4684 23741 4724 23752
rect 4779 23792 4821 23801
rect 4779 23752 4780 23792
rect 4820 23752 4821 23792
rect 4779 23743 4821 23752
rect 4876 23792 4916 24088
rect 4972 23960 5012 24844
rect 5068 24716 5108 24725
rect 5164 24716 5204 25096
rect 5108 24676 5204 24716
rect 5068 24667 5108 24676
rect 5260 24632 5300 25264
rect 5355 25220 5397 25229
rect 5355 25180 5356 25220
rect 5396 25180 5397 25220
rect 5355 25171 5397 25180
rect 4972 23911 5012 23920
rect 5164 24592 5300 24632
rect 4876 23743 4916 23752
rect 5164 23792 5204 24592
rect 5356 24464 5396 25171
rect 5452 24632 5492 24641
rect 5644 24632 5684 25936
rect 5836 25304 5876 26104
rect 6316 25976 6356 28960
rect 6412 28496 6452 28505
rect 6412 26816 6452 28456
rect 6604 28328 6644 28337
rect 6604 27833 6644 28288
rect 6700 28328 6740 28337
rect 6700 28085 6740 28288
rect 6796 28328 6836 28337
rect 6699 28076 6741 28085
rect 6699 28036 6700 28076
rect 6740 28036 6741 28076
rect 6699 28027 6741 28036
rect 6796 28001 6836 28288
rect 6892 28328 6932 28337
rect 7084 28328 7124 28337
rect 6932 28288 7084 28328
rect 6892 28279 6932 28288
rect 7084 28279 7124 28288
rect 7275 28328 7317 28337
rect 7275 28288 7276 28328
rect 7316 28288 7317 28328
rect 7275 28279 7317 28288
rect 7372 28328 7412 29035
rect 7467 28412 7509 28421
rect 7467 28372 7468 28412
rect 7508 28372 7509 28412
rect 7467 28363 7509 28372
rect 7372 28279 7412 28288
rect 7179 28244 7221 28253
rect 7179 28204 7180 28244
rect 7220 28204 7221 28244
rect 7179 28195 7221 28204
rect 7180 28110 7220 28195
rect 7276 28194 7316 28279
rect 7371 28160 7413 28169
rect 7371 28120 7372 28160
rect 7412 28120 7413 28160
rect 7371 28111 7413 28120
rect 7275 28076 7317 28085
rect 7275 28036 7276 28076
rect 7316 28036 7317 28076
rect 7275 28027 7317 28036
rect 6795 27992 6837 28001
rect 6795 27952 6796 27992
rect 6836 27952 6837 27992
rect 6795 27943 6837 27952
rect 6603 27824 6645 27833
rect 6603 27784 6604 27824
rect 6644 27784 6645 27824
rect 6603 27775 6645 27784
rect 7083 27740 7125 27749
rect 7083 27700 7084 27740
rect 7124 27700 7125 27740
rect 7083 27691 7125 27700
rect 6988 27656 7028 27665
rect 6796 27404 6836 27413
rect 6700 26816 6740 26825
rect 6412 26776 6700 26816
rect 6700 26767 6740 26776
rect 6412 25976 6452 25985
rect 6316 25936 6412 25976
rect 6412 25927 6452 25936
rect 6796 25733 6836 27364
rect 6988 27245 7028 27616
rect 6987 27236 7029 27245
rect 6987 27196 6988 27236
rect 7028 27196 7029 27236
rect 6987 27187 7029 27196
rect 7084 26816 7124 27691
rect 7276 27488 7316 28027
rect 7372 27656 7412 28111
rect 7468 27740 7508 28363
rect 7564 28160 7604 28169
rect 7564 27749 7604 28120
rect 7756 27833 7796 29800
rect 7852 29840 7892 30211
rect 7852 29791 7892 29800
rect 7948 29345 7988 30640
rect 8044 30092 8084 30808
rect 8044 30043 8084 30052
rect 8139 30008 8181 30017
rect 8139 29968 8140 30008
rect 8180 29968 8181 30008
rect 8139 29959 8181 29968
rect 7947 29336 7989 29345
rect 7947 29296 7948 29336
rect 7988 29296 7989 29336
rect 7947 29287 7989 29296
rect 8044 29177 8084 29262
rect 8043 29168 8085 29177
rect 8043 29128 8044 29168
rect 8084 29128 8085 29168
rect 8043 29119 8085 29128
rect 8140 29000 8180 29959
rect 8044 28960 8180 29000
rect 7851 27992 7893 28001
rect 7851 27952 7852 27992
rect 7892 27952 7893 27992
rect 7851 27943 7893 27952
rect 7755 27824 7797 27833
rect 7755 27784 7756 27824
rect 7796 27784 7797 27824
rect 7755 27775 7797 27784
rect 7468 27691 7508 27700
rect 7563 27740 7605 27749
rect 7563 27700 7564 27740
rect 7604 27700 7605 27740
rect 7563 27691 7605 27700
rect 7372 27607 7412 27616
rect 7660 27656 7700 27667
rect 7660 27581 7700 27616
rect 7756 27656 7796 27665
rect 7659 27572 7701 27581
rect 7659 27532 7660 27572
rect 7700 27532 7701 27572
rect 7659 27523 7701 27532
rect 7756 27497 7796 27616
rect 7852 27656 7892 27943
rect 7755 27488 7797 27497
rect 7276 27448 7604 27488
rect 7084 26767 7124 26776
rect 6988 26144 7028 26153
rect 6795 25724 6837 25733
rect 6795 25684 6796 25724
rect 6836 25684 6837 25724
rect 6795 25675 6837 25684
rect 6700 25472 6740 25481
rect 6740 25432 6932 25472
rect 6700 25423 6740 25432
rect 5836 25255 5876 25264
rect 5492 24592 5684 24632
rect 6316 24632 6356 24641
rect 6356 24592 6452 24632
rect 5452 24583 5492 24592
rect 6316 24583 6356 24592
rect 5356 24424 5492 24464
rect 5355 24296 5397 24305
rect 5355 24256 5356 24296
rect 5396 24256 5397 24296
rect 5355 24247 5397 24256
rect 5259 24044 5301 24053
rect 5259 24004 5260 24044
rect 5300 24004 5301 24044
rect 5259 23995 5301 24004
rect 5164 23743 5204 23752
rect 5260 23792 5300 23995
rect 5260 23743 5300 23752
rect 5356 23792 5396 24247
rect 5356 23743 5396 23752
rect 5452 23792 5492 24424
rect 5835 24044 5877 24053
rect 5835 24004 5836 24044
rect 5876 24004 5877 24044
rect 5835 23995 5877 24004
rect 5739 23960 5781 23969
rect 5739 23920 5740 23960
rect 5780 23920 5781 23960
rect 5644 23885 5684 23916
rect 5739 23911 5781 23920
rect 5643 23876 5685 23885
rect 5643 23836 5644 23876
rect 5684 23836 5685 23876
rect 5643 23827 5685 23836
rect 5452 23743 5492 23752
rect 5644 23792 5684 23827
rect 4252 23584 4340 23624
rect 4395 23624 4437 23633
rect 4395 23584 4396 23624
rect 4436 23584 4437 23624
rect 4252 23540 4292 23584
rect 4395 23575 4437 23584
rect 4587 23624 4629 23633
rect 4587 23584 4588 23624
rect 4628 23584 4629 23624
rect 4587 23575 4629 23584
rect 3915 23500 3916 23540
rect 3956 23500 3957 23540
rect 3915 23491 3957 23500
rect 4012 23500 4148 23540
rect 4204 23500 4292 23540
rect 3916 23120 3956 23491
rect 3916 23071 3956 23080
rect 4012 22961 4052 23500
rect 4204 23288 4244 23500
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 4204 23248 4340 23288
rect 4108 23120 4148 23129
rect 4011 22952 4053 22961
rect 4011 22912 4012 22952
rect 4052 22912 4053 22952
rect 4011 22903 4053 22912
rect 3915 22868 3957 22877
rect 3915 22828 3916 22868
rect 3956 22828 3957 22868
rect 3915 22819 3957 22828
rect 3916 22734 3956 22819
rect 3916 22280 3956 22289
rect 3820 22240 3916 22280
rect 3627 22231 3669 22240
rect 2859 22156 2860 22196
rect 2900 22156 2996 22196
rect 2859 22147 2901 22156
rect 1803 21692 1845 21701
rect 1803 21652 1804 21692
rect 1844 21652 1845 21692
rect 1803 21643 1845 21652
rect 2763 21692 2805 21701
rect 2763 21652 2764 21692
rect 2804 21652 2805 21692
rect 2763 21643 2805 21652
rect 1708 21440 1748 21449
rect 1612 21400 1708 21440
rect 1708 21391 1748 21400
rect 1708 20768 1748 20777
rect 1804 20768 1844 21643
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 2668 21474 2708 21559
rect 2764 21558 2804 21643
rect 2860 21608 2900 22147
rect 2955 21692 2997 21701
rect 2955 21652 2956 21692
rect 2996 21652 2997 21692
rect 2955 21643 2997 21652
rect 2860 21559 2900 21568
rect 2956 21608 2996 21643
rect 3148 21608 3188 22231
rect 3820 22112 3860 22121
rect 3820 21617 3860 22072
rect 3916 21869 3956 22240
rect 4012 22280 4052 22289
rect 3915 21860 3957 21869
rect 3915 21820 3916 21860
rect 3956 21820 3957 21860
rect 3915 21811 3957 21820
rect 2956 21557 2996 21568
rect 3052 21568 3148 21608
rect 3052 21524 3092 21568
rect 3148 21559 3188 21568
rect 3819 21608 3861 21617
rect 3819 21568 3820 21608
rect 3860 21568 3861 21608
rect 3819 21559 3861 21568
rect 4012 21533 4052 22240
rect 4108 22280 4148 23080
rect 4203 23120 4245 23129
rect 4203 23080 4204 23120
rect 4244 23080 4245 23120
rect 4203 23071 4245 23080
rect 4204 22986 4244 23071
rect 4300 22448 4340 23248
rect 4492 23120 4532 23129
rect 4492 22961 4532 23080
rect 4780 23120 4820 23743
rect 4971 23624 5013 23633
rect 4971 23584 4972 23624
rect 5012 23584 5013 23624
rect 4971 23575 5013 23584
rect 4972 23213 5012 23575
rect 5163 23456 5205 23465
rect 5163 23416 5164 23456
rect 5204 23416 5205 23456
rect 5163 23407 5205 23416
rect 4971 23204 5013 23213
rect 4971 23164 4972 23204
rect 5012 23164 5013 23204
rect 4971 23155 5013 23164
rect 4780 23071 4820 23080
rect 4876 23120 4916 23129
rect 4491 22952 4533 22961
rect 4491 22912 4492 22952
rect 4532 22912 4533 22952
rect 4491 22903 4533 22912
rect 4108 22205 4148 22240
rect 4204 22408 4340 22448
rect 4107 22196 4149 22205
rect 4107 22156 4108 22196
rect 4148 22156 4149 22196
rect 4107 22147 4149 22156
rect 4107 21608 4149 21617
rect 4107 21568 4108 21608
rect 4148 21568 4149 21608
rect 4107 21559 4149 21568
rect 3044 21484 3092 21524
rect 4011 21524 4053 21533
rect 4011 21484 4012 21524
rect 4052 21484 4053 21524
rect 2188 21440 2228 21449
rect 3044 21440 3084 21484
rect 4011 21475 4053 21484
rect 4108 21474 4148 21559
rect 1748 20728 1844 20768
rect 2092 20768 2132 20777
rect 2188 20768 2228 21400
rect 2132 20728 2228 20768
rect 2956 21400 3084 21440
rect 2956 20768 2996 21400
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4108 21020 4148 21029
rect 4204 21020 4244 22408
rect 4876 22289 4916 23080
rect 4972 22532 5012 23155
rect 5164 22952 5204 23407
rect 5451 23120 5493 23129
rect 5451 23080 5452 23120
rect 5492 23080 5493 23120
rect 5451 23071 5493 23080
rect 5548 23120 5588 23129
rect 5452 22986 5492 23071
rect 5164 22903 5204 22912
rect 5548 22709 5588 23080
rect 5547 22700 5589 22709
rect 5547 22660 5548 22700
rect 5588 22660 5589 22700
rect 5547 22651 5589 22660
rect 4972 22483 5012 22492
rect 5644 22532 5684 23752
rect 5740 23792 5780 23911
rect 5740 23743 5780 23752
rect 5836 23792 5876 23995
rect 6315 23960 6357 23969
rect 6315 23920 6316 23960
rect 6356 23920 6357 23960
rect 6315 23911 6357 23920
rect 6316 23826 6356 23911
rect 5836 23743 5876 23752
rect 5931 23708 5973 23717
rect 5931 23668 5932 23708
rect 5972 23668 5973 23708
rect 5931 23659 5973 23668
rect 5932 23574 5972 23659
rect 6027 23288 6069 23297
rect 6027 23248 6028 23288
rect 6068 23248 6069 23288
rect 6027 23239 6069 23248
rect 5739 23204 5781 23213
rect 5739 23164 5740 23204
rect 5780 23164 5781 23204
rect 5739 23155 5781 23164
rect 5740 23120 5780 23155
rect 6028 23154 6068 23239
rect 6123 23204 6165 23213
rect 6123 23164 6124 23204
rect 6164 23164 6165 23204
rect 6123 23155 6165 23164
rect 5740 23069 5780 23080
rect 6124 23120 6164 23155
rect 6124 23069 6164 23080
rect 6315 23036 6357 23045
rect 6315 22996 6316 23036
rect 6356 22996 6357 23036
rect 6315 22987 6357 22996
rect 5644 22483 5684 22492
rect 5836 22868 5876 22877
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4875 22280 4917 22289
rect 4875 22240 4876 22280
rect 4916 22240 4917 22280
rect 4875 22231 4917 22240
rect 5164 22280 5204 22291
rect 4300 22146 4340 22231
rect 5164 22205 5204 22240
rect 5163 22196 5205 22205
rect 5163 22156 5164 22196
rect 5204 22156 5300 22196
rect 5163 22147 5205 22156
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 5067 21860 5109 21869
rect 5067 21820 5068 21860
rect 5108 21820 5109 21860
rect 5067 21811 5109 21820
rect 4972 21776 5012 21785
rect 4492 21736 4972 21776
rect 4492 21608 4532 21736
rect 4972 21727 5012 21736
rect 4492 21559 4532 21568
rect 4684 21608 4724 21617
rect 4491 21440 4533 21449
rect 4491 21400 4492 21440
rect 4532 21400 4533 21440
rect 4491 21391 4533 21400
rect 4492 21306 4532 21391
rect 4148 20980 4244 21020
rect 4108 20971 4148 20980
rect 4204 20777 4244 20980
rect 4684 20852 4724 21568
rect 4780 21608 4820 21617
rect 4780 21440 4820 21568
rect 5068 21608 5108 21811
rect 5163 21776 5205 21785
rect 5163 21736 5164 21776
rect 5204 21736 5205 21776
rect 5163 21727 5205 21736
rect 5068 21559 5108 21568
rect 5164 21608 5204 21727
rect 5164 21559 5204 21568
rect 5260 21608 5300 22156
rect 5836 21701 5876 22828
rect 6316 22364 6356 22987
rect 6412 22457 6452 24592
rect 6795 24044 6837 24053
rect 6795 24004 6796 24044
rect 6836 24004 6837 24044
rect 6795 23995 6837 24004
rect 6508 23792 6548 23801
rect 6508 23297 6548 23752
rect 6507 23288 6549 23297
rect 6507 23248 6508 23288
rect 6548 23248 6549 23288
rect 6507 23239 6549 23248
rect 6699 23120 6741 23129
rect 6699 23080 6700 23120
rect 6740 23080 6741 23120
rect 6699 23071 6741 23080
rect 6796 23120 6836 23995
rect 6796 23071 6836 23080
rect 6700 22986 6740 23071
rect 6411 22448 6453 22457
rect 6411 22408 6412 22448
rect 6452 22408 6453 22448
rect 6411 22399 6453 22408
rect 6028 22324 6356 22364
rect 6028 22280 6068 22324
rect 6316 22280 6356 22324
rect 6412 22280 6452 22289
rect 6316 22240 6412 22280
rect 6028 22231 6068 22240
rect 6412 22231 6452 22240
rect 6507 22280 6549 22289
rect 6507 22240 6508 22280
rect 6548 22240 6549 22280
rect 6507 22231 6549 22240
rect 6604 22280 6644 22291
rect 6123 22196 6165 22205
rect 6123 22156 6124 22196
rect 6164 22156 6165 22196
rect 6123 22147 6165 22156
rect 5835 21692 5877 21701
rect 5835 21652 5836 21692
rect 5876 21652 5877 21692
rect 5835 21643 5877 21652
rect 5260 21559 5300 21568
rect 5548 21608 5588 21617
rect 5355 21524 5397 21533
rect 5355 21484 5356 21524
rect 5396 21484 5397 21524
rect 5355 21475 5397 21484
rect 4780 21400 5204 21440
rect 5067 21272 5109 21281
rect 5067 21232 5068 21272
rect 5108 21232 5109 21272
rect 5067 21223 5109 21232
rect 4684 20812 4820 20852
rect 1708 20719 1748 20728
rect 2092 20719 2132 20728
rect 1996 19424 2036 19433
rect 1323 19088 1365 19097
rect 1323 19048 1324 19088
rect 1364 19048 1365 19088
rect 1323 19039 1365 19048
rect 1324 18668 1364 19039
rect 1324 18619 1364 18628
rect 1708 18584 1748 18593
rect 1420 18544 1708 18584
rect 1324 17912 1364 17921
rect 1420 17912 1460 18544
rect 1708 18535 1748 18544
rect 1364 17872 1460 17912
rect 1324 17863 1364 17872
rect 1900 17744 1940 17753
rect 1996 17744 2036 19384
rect 2956 18593 2996 20728
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4396 20600 4436 20609
rect 4204 20560 4396 20600
rect 4108 20180 4148 20189
rect 4204 20180 4244 20560
rect 4396 20551 4436 20560
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4148 20140 4244 20180
rect 4108 20131 4148 20140
rect 4492 20096 4532 20105
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4492 19433 4532 20056
rect 3723 19424 3765 19433
rect 3723 19384 3724 19424
rect 3764 19384 3765 19424
rect 3723 19375 3765 19384
rect 4491 19424 4533 19433
rect 4491 19384 4492 19424
rect 4532 19384 4533 19424
rect 4491 19375 4533 19384
rect 3724 19290 3764 19375
rect 4203 19340 4245 19349
rect 4203 19300 4204 19340
rect 4244 19300 4245 19340
rect 4203 19291 4245 19300
rect 3916 19256 3956 19265
rect 3820 19216 3916 19256
rect 3723 19172 3765 19181
rect 3723 19132 3724 19172
rect 3764 19132 3765 19172
rect 3723 19123 3765 19132
rect 3724 18752 3764 19123
rect 3724 18703 3764 18712
rect 3820 18593 3860 19216
rect 3916 19207 3956 19216
rect 4012 19256 4052 19265
rect 2571 18584 2613 18593
rect 2571 18544 2572 18584
rect 2612 18544 2613 18584
rect 2571 18535 2613 18544
rect 2763 18584 2805 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 2955 18584 2997 18593
rect 2955 18544 2956 18584
rect 2996 18544 2997 18584
rect 2955 18535 2997 18544
rect 3819 18584 3861 18593
rect 3819 18544 3820 18584
rect 3860 18544 3861 18584
rect 3819 18535 3861 18544
rect 3916 18584 3956 18593
rect 2572 18450 2612 18535
rect 1940 17704 2036 17744
rect 2764 17744 2804 18535
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 1900 17695 1940 17704
rect 2764 17695 2804 17704
rect 1516 17660 1556 17669
rect 1516 17249 1556 17620
rect 3627 17576 3669 17585
rect 3627 17536 3628 17576
rect 3668 17536 3669 17576
rect 3627 17527 3669 17536
rect 1515 17240 1557 17249
rect 1515 17200 1516 17240
rect 1556 17200 1557 17240
rect 1515 17191 1557 17200
rect 3531 17156 3573 17165
rect 3436 17116 3532 17156
rect 3572 17116 3573 17156
rect 3243 17072 3285 17081
rect 3243 17032 3244 17072
rect 3284 17032 3285 17072
rect 3243 17023 3285 17032
rect 3436 17072 3476 17116
rect 3531 17107 3573 17116
rect 3436 17023 3476 17032
rect 3628 17072 3668 17527
rect 3820 17333 3860 18535
rect 3916 17996 3956 18544
rect 3916 17947 3956 17956
rect 4012 17669 4052 19216
rect 4204 19256 4244 19291
rect 4204 19205 4244 19216
rect 4491 19256 4533 19265
rect 4491 19216 4492 19256
rect 4532 19216 4533 19256
rect 4491 19207 4533 19216
rect 4492 19122 4532 19207
rect 4780 19181 4820 20812
rect 5068 20768 5108 21223
rect 5068 20719 5108 20728
rect 5164 20180 5204 21400
rect 5356 21020 5396 21475
rect 5451 21440 5493 21449
rect 5451 21400 5452 21440
rect 5492 21400 5493 21440
rect 5451 21391 5493 21400
rect 5452 21306 5492 21391
rect 5548 21029 5588 21568
rect 5740 21608 5780 21617
rect 5547 21020 5589 21029
rect 5356 20980 5492 21020
rect 5259 20768 5301 20777
rect 5259 20728 5260 20768
rect 5300 20728 5301 20768
rect 5259 20719 5301 20728
rect 5260 20634 5300 20719
rect 5164 20140 5300 20180
rect 5260 19508 5300 20140
rect 5355 20096 5397 20105
rect 5355 20056 5356 20096
rect 5396 20056 5397 20096
rect 5355 20047 5397 20056
rect 5356 19962 5396 20047
rect 5356 19508 5396 19517
rect 5260 19468 5356 19508
rect 5356 19459 5396 19468
rect 5452 19256 5492 20980
rect 5547 20980 5548 21020
rect 5588 20980 5589 21020
rect 5547 20971 5589 20980
rect 5740 19937 5780 21568
rect 5931 21524 5973 21533
rect 5931 21484 5932 21524
rect 5972 21484 5973 21524
rect 5931 21475 5973 21484
rect 5932 21020 5972 21475
rect 5932 20971 5972 20980
rect 6124 20180 6164 22147
rect 6508 22146 6548 22231
rect 6604 22205 6644 22240
rect 6603 22196 6645 22205
rect 6603 22156 6604 22196
rect 6644 22156 6645 22196
rect 6603 22147 6645 22156
rect 6700 22112 6740 22121
rect 6412 21608 6452 21617
rect 6604 21608 6644 21617
rect 6452 21568 6604 21608
rect 6412 21559 6452 21568
rect 6604 21559 6644 21568
rect 6219 21020 6261 21029
rect 6219 20980 6220 21020
rect 6260 20980 6261 21020
rect 6219 20971 6261 20980
rect 6220 20886 6260 20971
rect 6508 20273 6548 20358
rect 6507 20264 6549 20273
rect 6507 20224 6508 20264
rect 6548 20224 6549 20264
rect 6507 20215 6549 20224
rect 6124 20140 6260 20180
rect 5739 19928 5781 19937
rect 5739 19888 5740 19928
rect 5780 19888 5781 19928
rect 5739 19879 5781 19888
rect 5835 19424 5877 19433
rect 5835 19384 5836 19424
rect 5876 19384 5877 19424
rect 5835 19375 5877 19384
rect 5836 19290 5876 19375
rect 5452 19207 5492 19216
rect 6028 19256 6068 19267
rect 6028 19181 6068 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6220 19256 6260 20140
rect 6700 20096 6740 22072
rect 6795 21692 6837 21701
rect 6795 21652 6796 21692
rect 6836 21652 6837 21692
rect 6795 21643 6837 21652
rect 6796 20768 6836 21643
rect 6892 21617 6932 25432
rect 6988 25304 7028 26104
rect 7468 26144 7508 26153
rect 7564 26144 7604 27448
rect 7755 27448 7756 27488
rect 7796 27448 7797 27488
rect 7755 27439 7797 27448
rect 7852 27068 7892 27616
rect 7852 27019 7892 27028
rect 7948 27656 7988 27665
rect 7948 26489 7988 27616
rect 8044 27581 8084 28960
rect 8332 28925 8372 30967
rect 8620 30932 8660 31312
rect 8812 31352 8852 31361
rect 8715 31268 8757 31277
rect 8715 31228 8716 31268
rect 8756 31228 8757 31268
rect 8715 31219 8757 31228
rect 8716 31134 8756 31219
rect 8620 30892 8756 30932
rect 8620 30764 8660 30773
rect 8524 30724 8620 30764
rect 8428 30666 8468 30675
rect 8428 30521 8468 30626
rect 8427 30512 8469 30521
rect 8427 30472 8428 30512
rect 8468 30472 8469 30512
rect 8427 30463 8469 30472
rect 8427 29672 8469 29681
rect 8427 29632 8428 29672
rect 8468 29632 8469 29672
rect 8427 29623 8469 29632
rect 8428 29252 8468 29623
rect 8428 29203 8468 29212
rect 8331 28916 8373 28925
rect 8331 28876 8332 28916
rect 8372 28876 8373 28916
rect 8331 28867 8373 28876
rect 8236 28328 8276 28339
rect 8236 28253 8276 28288
rect 8235 28244 8277 28253
rect 8235 28204 8236 28244
rect 8276 28204 8277 28244
rect 8235 28195 8277 28204
rect 8139 27656 8181 27665
rect 8139 27616 8140 27656
rect 8180 27616 8181 27656
rect 8139 27607 8181 27616
rect 8043 27572 8085 27581
rect 8043 27532 8044 27572
rect 8084 27532 8085 27572
rect 8043 27523 8085 27532
rect 8140 27522 8180 27607
rect 8044 26648 8084 26657
rect 7947 26480 7989 26489
rect 7947 26440 7948 26480
rect 7988 26440 7989 26480
rect 7947 26431 7989 26440
rect 7851 26228 7893 26237
rect 7851 26188 7852 26228
rect 7892 26188 7893 26228
rect 7851 26179 7893 26188
rect 7756 26144 7796 26153
rect 7564 26104 7756 26144
rect 7468 25397 7508 26104
rect 7756 26095 7796 26104
rect 7852 26094 7892 26179
rect 7467 25388 7509 25397
rect 7467 25348 7468 25388
rect 7508 25348 7509 25388
rect 7467 25339 7509 25348
rect 7851 25388 7893 25397
rect 7851 25348 7852 25388
rect 7892 25348 7893 25388
rect 7851 25339 7893 25348
rect 6988 25229 7028 25264
rect 7852 25304 7892 25339
rect 6987 25220 7029 25229
rect 6987 25180 6988 25220
rect 7028 25180 7029 25220
rect 6987 25171 7029 25180
rect 7756 24632 7796 24641
rect 7852 24632 7892 25264
rect 8044 24800 8084 26608
rect 8140 25892 8180 25901
rect 8140 24809 8180 25852
rect 8235 25892 8277 25901
rect 8235 25852 8236 25892
rect 8276 25852 8277 25892
rect 8235 25843 8277 25852
rect 7796 24592 7892 24632
rect 7948 24760 8084 24800
rect 8139 24800 8181 24809
rect 8139 24760 8140 24800
rect 8180 24760 8181 24800
rect 7756 24583 7796 24592
rect 7468 24380 7508 24391
rect 7468 24305 7508 24340
rect 7467 24296 7509 24305
rect 7467 24256 7468 24296
rect 7508 24256 7509 24296
rect 7467 24247 7509 24256
rect 7755 23960 7797 23969
rect 7755 23920 7756 23960
rect 7796 23920 7797 23960
rect 7755 23911 7797 23920
rect 7756 23792 7796 23911
rect 7756 23743 7796 23752
rect 7180 23708 7220 23717
rect 7372 23708 7412 23717
rect 7220 23668 7372 23708
rect 7180 23659 7220 23668
rect 7372 23659 7412 23668
rect 7179 23288 7221 23297
rect 7179 23248 7180 23288
rect 7220 23248 7221 23288
rect 7179 23239 7221 23248
rect 7180 23154 7220 23239
rect 7467 23204 7509 23213
rect 7467 23164 7468 23204
rect 7508 23164 7509 23204
rect 7467 23155 7509 23164
rect 6987 23120 7029 23129
rect 6987 23080 6988 23120
rect 7028 23080 7029 23120
rect 6987 23071 7029 23080
rect 7084 23120 7124 23131
rect 6988 22986 7028 23071
rect 7084 23045 7124 23080
rect 7275 23120 7317 23129
rect 7275 23080 7276 23120
rect 7316 23080 7317 23120
rect 7275 23071 7317 23080
rect 7083 23036 7125 23045
rect 7083 22996 7084 23036
rect 7124 22996 7125 23036
rect 7083 22987 7125 22996
rect 7276 22986 7316 23071
rect 7468 23070 7508 23155
rect 7084 22448 7124 22457
rect 6988 22408 7084 22448
rect 6891 21608 6933 21617
rect 6891 21568 6892 21608
rect 6932 21568 6933 21608
rect 6891 21559 6933 21568
rect 6988 21608 7028 22408
rect 7084 22399 7124 22408
rect 7755 22448 7797 22457
rect 7755 22408 7756 22448
rect 7796 22408 7797 22448
rect 7755 22399 7797 22408
rect 6988 21559 7028 21568
rect 7372 22280 7412 22289
rect 6892 20768 6932 20777
rect 6796 20728 6892 20768
rect 6796 20273 6836 20728
rect 6892 20719 6932 20728
rect 7372 20768 7412 22240
rect 7659 21608 7701 21617
rect 7659 21568 7660 21608
rect 7700 21568 7701 21608
rect 7756 21608 7796 22399
rect 7948 22205 7988 24760
rect 8139 24751 8181 24760
rect 8043 24632 8085 24641
rect 8043 24592 8044 24632
rect 8084 24592 8085 24632
rect 8043 24583 8085 24592
rect 8140 24632 8180 24641
rect 8044 24305 8084 24583
rect 8043 24296 8085 24305
rect 8043 24256 8044 24296
rect 8084 24256 8085 24296
rect 8043 24247 8085 24256
rect 8140 23288 8180 24592
rect 8236 24464 8276 25843
rect 8332 25304 8372 28867
rect 8427 27740 8469 27749
rect 8427 27700 8428 27740
rect 8468 27700 8469 27740
rect 8427 27691 8469 27700
rect 8428 27245 8468 27691
rect 8427 27236 8469 27245
rect 8427 27196 8428 27236
rect 8468 27196 8469 27236
rect 8427 27187 8469 27196
rect 8428 26816 8468 27187
rect 8428 26767 8468 26776
rect 8524 26405 8564 30724
rect 8620 30715 8660 30724
rect 8716 30017 8756 30892
rect 8812 30269 8852 31312
rect 9676 31352 9716 31363
rect 9676 31277 9716 31312
rect 10059 31352 10101 31361
rect 10059 31312 10060 31352
rect 10100 31312 10101 31352
rect 10059 31303 10101 31312
rect 9675 31268 9717 31277
rect 9675 31228 9676 31268
rect 9716 31228 9717 31268
rect 9675 31219 9717 31228
rect 10060 31218 10100 31303
rect 9004 31184 9044 31193
rect 8908 31144 9004 31184
rect 8811 30260 8853 30269
rect 8811 30220 8812 30260
rect 8852 30220 8853 30260
rect 8811 30211 8853 30220
rect 8715 30008 8757 30017
rect 8715 29968 8716 30008
rect 8756 29968 8757 30008
rect 8715 29959 8757 29968
rect 8716 29840 8756 29849
rect 8716 29345 8756 29800
rect 8908 29840 8948 31144
rect 9004 31135 9044 31144
rect 9675 30680 9717 30689
rect 9675 30640 9676 30680
rect 9716 30640 9717 30680
rect 9675 30631 9717 30640
rect 9676 30546 9716 30631
rect 9868 30512 9908 30521
rect 8908 29791 8948 29800
rect 9004 30428 9044 30437
rect 9004 29672 9044 30388
rect 9099 30092 9141 30101
rect 9099 30052 9100 30092
rect 9140 30052 9141 30092
rect 9099 30043 9141 30052
rect 8908 29632 9044 29672
rect 8715 29336 8757 29345
rect 8715 29296 8716 29336
rect 8756 29296 8757 29336
rect 8715 29287 8757 29296
rect 8620 29093 8660 29178
rect 8715 29168 8757 29177
rect 8715 29128 8716 29168
rect 8756 29128 8757 29168
rect 8715 29119 8757 29128
rect 8619 29084 8661 29093
rect 8619 29044 8620 29084
rect 8660 29044 8661 29084
rect 8619 29035 8661 29044
rect 8716 29034 8756 29119
rect 8908 29000 8948 29632
rect 9100 29597 9140 30043
rect 9292 29840 9332 29849
rect 9868 29840 9908 30472
rect 9963 29924 10005 29933
rect 9963 29884 9964 29924
rect 10004 29884 10005 29924
rect 9963 29875 10005 29884
rect 9332 29800 9908 29840
rect 9292 29791 9332 29800
rect 9099 29588 9141 29597
rect 9099 29548 9100 29588
rect 9140 29548 9141 29588
rect 9099 29539 9141 29548
rect 9100 29168 9140 29539
rect 9100 29119 9140 29128
rect 9964 29168 10004 29875
rect 10156 29840 10196 29849
rect 10156 29177 10196 29800
rect 9964 29119 10004 29128
rect 10155 29168 10197 29177
rect 10155 29128 10156 29168
rect 10196 29128 10197 29168
rect 10155 29119 10197 29128
rect 8812 28960 8948 29000
rect 10156 29000 10196 29119
rect 10156 28960 10292 29000
rect 8715 28328 8757 28337
rect 8715 28288 8716 28328
rect 8756 28288 8757 28328
rect 8715 28279 8757 28288
rect 8716 28169 8756 28279
rect 8715 28160 8757 28169
rect 8715 28120 8716 28160
rect 8756 28120 8757 28160
rect 8715 28111 8757 28120
rect 8812 27824 8852 28960
rect 9291 28916 9333 28925
rect 9291 28876 9292 28916
rect 9332 28876 9333 28916
rect 9291 28867 9333 28876
rect 9292 28782 9332 28867
rect 8620 27784 8852 27824
rect 8908 28496 8948 28505
rect 8620 27329 8660 27784
rect 8800 27665 8840 27684
rect 8800 27656 8852 27665
rect 8716 27616 8812 27656
rect 8716 27497 8756 27616
rect 8812 27607 8852 27616
rect 8908 27581 8948 28456
rect 10155 28328 10197 28337
rect 10155 28288 10156 28328
rect 10196 28288 10197 28328
rect 10155 28279 10197 28288
rect 10156 28194 10196 28279
rect 10060 28160 10100 28169
rect 9292 28120 10060 28160
rect 9004 27656 9044 27665
rect 9044 27616 9236 27656
rect 9004 27607 9044 27616
rect 8907 27572 8949 27581
rect 8907 27532 8908 27572
rect 8948 27532 8949 27572
rect 8907 27523 8949 27532
rect 8715 27488 8757 27497
rect 8715 27448 8716 27488
rect 8756 27448 8757 27488
rect 8715 27439 8757 27448
rect 8619 27320 8661 27329
rect 8619 27280 8620 27320
rect 8660 27280 8661 27320
rect 8619 27271 8661 27280
rect 8908 26993 8948 27523
rect 9196 27068 9236 27616
rect 9292 27152 9332 28120
rect 10060 28111 10100 28120
rect 9388 27656 9428 27665
rect 10252 27656 10292 28960
rect 10348 28169 10388 32824
rect 10443 32824 10444 32864
rect 10484 32824 10485 32864
rect 10443 32815 10485 32824
rect 10444 32730 10484 32815
rect 10827 32192 10869 32201
rect 10827 32152 10828 32192
rect 10868 32152 10869 32192
rect 10827 32143 10869 32152
rect 10828 32108 10868 32143
rect 10828 32057 10868 32068
rect 10827 31772 10869 31781
rect 10827 31732 10828 31772
rect 10868 31732 10869 31772
rect 10827 31723 10869 31732
rect 10443 31688 10485 31697
rect 10443 31648 10444 31688
rect 10484 31648 10485 31688
rect 10443 31639 10485 31648
rect 10444 31520 10484 31639
rect 10444 31471 10484 31480
rect 10828 31436 10868 31723
rect 10828 31387 10868 31396
rect 10924 31361 10964 33412
rect 11116 33125 11156 34168
rect 11403 34208 11445 34217
rect 11403 34168 11404 34208
rect 11444 34168 11445 34208
rect 11403 34159 11445 34168
rect 11404 34074 11444 34159
rect 11211 33704 11253 33713
rect 11211 33664 11212 33704
rect 11252 33664 11253 33704
rect 11211 33655 11253 33664
rect 11115 33116 11157 33125
rect 11115 33076 11116 33116
rect 11156 33076 11157 33116
rect 11115 33067 11157 33076
rect 11115 32864 11157 32873
rect 11115 32824 11116 32864
rect 11156 32824 11157 32864
rect 11115 32815 11157 32824
rect 11116 32730 11156 32815
rect 11019 32192 11061 32201
rect 11019 32152 11020 32192
rect 11060 32152 11061 32192
rect 11019 32143 11061 32152
rect 11020 31865 11060 32143
rect 11019 31856 11061 31865
rect 11019 31816 11020 31856
rect 11060 31816 11061 31856
rect 11019 31807 11061 31816
rect 11212 31781 11252 33655
rect 11500 33377 11540 34243
rect 11692 34133 11732 34336
rect 11884 34376 11924 34579
rect 11884 34327 11924 34336
rect 11980 34376 12020 34387
rect 11980 34301 12020 34336
rect 12076 34376 12116 34840
rect 12171 34460 12213 34469
rect 12171 34420 12172 34460
rect 12212 34420 12213 34460
rect 12171 34411 12213 34420
rect 12076 34327 12116 34336
rect 12172 34376 12212 34411
rect 12172 34325 12212 34336
rect 12364 34376 12404 34385
rect 11979 34292 12021 34301
rect 11979 34252 11980 34292
rect 12020 34252 12021 34292
rect 11979 34243 12021 34252
rect 12364 34217 12404 34336
rect 12460 34376 12500 34385
rect 12363 34208 12405 34217
rect 12363 34168 12364 34208
rect 12404 34168 12405 34208
rect 12363 34159 12405 34168
rect 11691 34124 11733 34133
rect 11691 34084 11692 34124
rect 11732 34084 11733 34124
rect 11691 34075 11733 34084
rect 11979 34124 12021 34133
rect 11979 34084 11980 34124
rect 12020 34084 12021 34124
rect 11979 34075 12021 34084
rect 11787 33872 11829 33881
rect 11787 33832 11788 33872
rect 11828 33832 11829 33872
rect 11787 33823 11829 33832
rect 11788 33738 11828 33823
rect 11596 33704 11636 33713
rect 11596 33452 11636 33664
rect 11788 33452 11828 33461
rect 11596 33412 11788 33452
rect 11499 33368 11541 33377
rect 11499 33328 11500 33368
rect 11540 33328 11541 33368
rect 11499 33319 11541 33328
rect 11211 31772 11253 31781
rect 11211 31732 11212 31772
rect 11252 31732 11253 31772
rect 11211 31723 11253 31732
rect 11500 31604 11540 33319
rect 11691 31940 11733 31949
rect 11691 31900 11692 31940
rect 11732 31900 11733 31940
rect 11691 31891 11733 31900
rect 11692 31806 11732 31891
rect 11500 31555 11540 31564
rect 11691 31520 11733 31529
rect 11691 31480 11692 31520
rect 11732 31480 11733 31520
rect 11691 31471 11733 31480
rect 11692 31386 11732 31471
rect 10923 31352 10965 31361
rect 10923 31312 10924 31352
rect 10964 31312 10965 31352
rect 10923 31303 10965 31312
rect 11019 30848 11061 30857
rect 11019 30808 11020 30848
rect 11060 30808 11061 30848
rect 11019 30799 11061 30808
rect 10923 30680 10965 30689
rect 10923 30640 10924 30680
rect 10964 30640 10965 30680
rect 10923 30631 10965 30640
rect 11020 30680 11060 30799
rect 11020 30631 11060 30640
rect 11116 30680 11156 30691
rect 10924 30546 10964 30631
rect 11116 30605 11156 30640
rect 11212 30680 11252 30689
rect 11115 30596 11157 30605
rect 11115 30556 11116 30596
rect 11156 30556 11157 30596
rect 11115 30547 11157 30556
rect 10923 30428 10965 30437
rect 10923 30388 10924 30428
rect 10964 30388 10965 30428
rect 10923 30379 10965 30388
rect 10924 29252 10964 30379
rect 11116 30269 11156 30547
rect 11212 30353 11252 30640
rect 11499 30680 11541 30689
rect 11691 30680 11733 30689
rect 11499 30640 11500 30680
rect 11540 30640 11541 30680
rect 11499 30631 11541 30640
rect 11596 30640 11692 30680
rect 11732 30640 11733 30680
rect 11403 30428 11445 30437
rect 11403 30388 11404 30428
rect 11444 30388 11445 30428
rect 11403 30379 11445 30388
rect 11211 30344 11253 30353
rect 11211 30304 11212 30344
rect 11252 30304 11253 30344
rect 11211 30295 11253 30304
rect 11404 30294 11444 30379
rect 11115 30260 11157 30269
rect 11115 30220 11116 30260
rect 11156 30220 11157 30260
rect 11115 30211 11157 30220
rect 11308 30017 11348 30048
rect 11307 30008 11349 30017
rect 11307 29968 11308 30008
rect 11348 29968 11349 30008
rect 11307 29959 11349 29968
rect 11308 29924 11348 29959
rect 11308 29849 11348 29884
rect 11307 29840 11349 29849
rect 11307 29800 11308 29840
rect 11348 29800 11349 29840
rect 11500 29840 11540 30631
rect 11596 30092 11636 30640
rect 11691 30631 11733 30640
rect 11691 30344 11733 30353
rect 11691 30304 11692 30344
rect 11732 30304 11733 30344
rect 11691 30295 11733 30304
rect 11596 30043 11636 30052
rect 11596 29840 11636 29849
rect 11500 29800 11596 29840
rect 11692 29840 11732 30295
rect 11788 30185 11828 33412
rect 11980 32948 12020 34075
rect 12460 33881 12500 34336
rect 12556 34376 12596 34387
rect 12556 34301 12596 34336
rect 12940 34376 12980 35008
rect 13131 34964 13173 34973
rect 13131 34924 13132 34964
rect 13172 34924 13173 34964
rect 13131 34915 13173 34924
rect 13132 34830 13172 34915
rect 13228 34889 13268 36427
rect 13900 36426 13940 36511
rect 15436 36476 15476 36485
rect 13996 35888 14036 35897
rect 13900 35848 13996 35888
rect 13611 35300 13653 35309
rect 13611 35260 13612 35300
rect 13652 35260 13653 35300
rect 13611 35251 13653 35260
rect 13227 34880 13269 34889
rect 13227 34840 13228 34880
rect 13268 34840 13269 34880
rect 13227 34831 13269 34840
rect 13131 34628 13173 34637
rect 13131 34588 13132 34628
rect 13172 34588 13173 34628
rect 13131 34579 13173 34588
rect 12940 34327 12980 34336
rect 13036 34376 13076 34387
rect 13036 34301 13076 34336
rect 13132 34376 13172 34579
rect 13228 34469 13268 34831
rect 13227 34460 13269 34469
rect 13227 34420 13228 34460
rect 13268 34420 13269 34460
rect 13227 34411 13269 34420
rect 13132 34327 13172 34336
rect 13228 34376 13268 34411
rect 13516 34376 13556 34385
rect 12555 34292 12597 34301
rect 12555 34252 12556 34292
rect 12596 34252 12597 34292
rect 12555 34243 12597 34252
rect 13035 34292 13077 34301
rect 13035 34252 13036 34292
rect 13076 34252 13077 34292
rect 13035 34243 13077 34252
rect 12652 34208 12692 34217
rect 12459 33872 12501 33881
rect 12459 33832 12460 33872
rect 12500 33832 12501 33872
rect 12459 33823 12501 33832
rect 12020 32908 12500 32948
rect 11980 32899 12020 32908
rect 11884 32192 11924 32201
rect 12268 32192 12308 32201
rect 11924 32152 12116 32192
rect 11884 32143 11924 32152
rect 12076 31604 12116 32152
rect 12268 31781 12308 32152
rect 12363 31856 12405 31865
rect 12363 31816 12364 31856
rect 12404 31816 12405 31856
rect 12363 31807 12405 31816
rect 12267 31772 12309 31781
rect 12267 31732 12268 31772
rect 12308 31732 12309 31772
rect 12267 31723 12309 31732
rect 12268 31604 12308 31613
rect 12076 31564 12268 31604
rect 12268 31555 12308 31564
rect 12171 31436 12213 31445
rect 12171 31396 12172 31436
rect 12212 31396 12213 31436
rect 12171 31387 12213 31396
rect 11884 31352 11924 31361
rect 11884 30857 11924 31312
rect 11883 30848 11925 30857
rect 11883 30808 11884 30848
rect 11924 30808 11925 30848
rect 11883 30799 11925 30808
rect 11883 30680 11925 30689
rect 12076 30680 12116 30689
rect 11883 30640 11884 30680
rect 11924 30640 12076 30680
rect 11883 30631 11925 30640
rect 12076 30631 12116 30640
rect 11979 30512 12021 30521
rect 11979 30472 11980 30512
rect 12020 30472 12021 30512
rect 11979 30463 12021 30472
rect 11883 30260 11925 30269
rect 11883 30220 11884 30260
rect 11924 30220 11925 30260
rect 11883 30211 11925 30220
rect 11787 30176 11829 30185
rect 11787 30136 11788 30176
rect 11828 30136 11829 30176
rect 11787 30127 11829 30136
rect 11787 29840 11829 29849
rect 11692 29800 11788 29840
rect 11828 29800 11829 29840
rect 11307 29791 11349 29800
rect 11596 29791 11636 29800
rect 11787 29791 11829 29800
rect 11884 29840 11924 30211
rect 11884 29791 11924 29800
rect 11788 29706 11828 29791
rect 10924 29203 10964 29212
rect 11320 29177 11360 29196
rect 11308 29168 11360 29177
rect 11348 29128 11444 29168
rect 11308 29119 11348 29128
rect 11404 28496 11444 29128
rect 11980 28496 12020 30463
rect 12172 30260 12212 31387
rect 12267 31352 12309 31361
rect 12267 31312 12268 31352
rect 12308 31312 12309 31352
rect 12267 31303 12309 31312
rect 12268 31218 12308 31303
rect 12076 30220 12212 30260
rect 12268 30680 12308 30689
rect 12076 29849 12116 30220
rect 12171 30092 12213 30101
rect 12171 30052 12172 30092
rect 12212 30052 12213 30092
rect 12171 30043 12213 30052
rect 12075 29840 12117 29849
rect 12075 29800 12076 29840
rect 12116 29800 12117 29840
rect 12075 29791 12117 29800
rect 12172 29840 12212 30043
rect 12268 30017 12308 30640
rect 12267 30008 12309 30017
rect 12267 29968 12268 30008
rect 12308 29968 12309 30008
rect 12267 29959 12309 29968
rect 12364 29840 12404 31807
rect 12460 31445 12500 32908
rect 12652 32873 12692 34168
rect 13228 34049 13268 34336
rect 13420 34336 13516 34376
rect 13227 34040 13269 34049
rect 13227 34000 13228 34040
rect 13268 34000 13269 34040
rect 13227 33991 13269 34000
rect 12939 33704 12981 33713
rect 12939 33664 12940 33704
rect 12980 33664 12981 33704
rect 12939 33655 12981 33664
rect 12940 33116 12980 33655
rect 12980 33076 13172 33116
rect 12940 33067 12980 33076
rect 12747 32948 12789 32957
rect 12747 32908 12748 32948
rect 12788 32908 12789 32948
rect 12747 32899 12789 32908
rect 12651 32864 12693 32873
rect 12651 32824 12652 32864
rect 12692 32824 12693 32864
rect 12651 32815 12693 32824
rect 12748 32696 12788 32899
rect 12652 32656 12788 32696
rect 12939 32696 12981 32705
rect 12939 32656 12940 32696
rect 12980 32656 12981 32696
rect 12459 31436 12501 31445
rect 12459 31396 12460 31436
rect 12500 31396 12501 31436
rect 12459 31387 12501 31396
rect 12460 31352 12500 31387
rect 12460 31302 12500 31312
rect 12556 31352 12596 31363
rect 12556 31277 12596 31312
rect 12555 31268 12597 31277
rect 12555 31228 12556 31268
rect 12596 31228 12597 31268
rect 12555 31219 12597 31228
rect 12555 30008 12597 30017
rect 12555 29968 12556 30008
rect 12596 29968 12597 30008
rect 12555 29959 12597 29968
rect 12460 29840 12500 29849
rect 12364 29800 12460 29840
rect 12172 29791 12212 29800
rect 12460 29791 12500 29800
rect 12556 29840 12596 29959
rect 12556 29791 12596 29800
rect 12171 29168 12213 29177
rect 12171 29128 12172 29168
rect 12212 29128 12213 29168
rect 12171 29119 12213 29128
rect 12172 29034 12212 29119
rect 11980 28456 12212 28496
rect 11404 28447 11444 28456
rect 11884 28328 11924 28337
rect 10347 28160 10389 28169
rect 10347 28120 10348 28160
rect 10388 28120 10389 28160
rect 10347 28111 10389 28120
rect 9428 27616 10100 27656
rect 9388 27607 9428 27616
rect 9292 27112 9428 27152
rect 9196 27019 9236 27028
rect 8907 26984 8949 26993
rect 8907 26944 8908 26984
rect 8948 26944 8949 26984
rect 8907 26935 8949 26944
rect 9291 26984 9333 26993
rect 9291 26944 9292 26984
rect 9332 26944 9333 26984
rect 9291 26935 9333 26944
rect 9099 26480 9141 26489
rect 9099 26440 9100 26480
rect 9140 26440 9141 26480
rect 9099 26431 9141 26440
rect 8523 26396 8565 26405
rect 8523 26356 8524 26396
rect 8564 26356 8565 26396
rect 8523 26347 8565 26356
rect 9100 26144 9140 26431
rect 9195 26312 9237 26321
rect 9195 26272 9196 26312
rect 9236 26272 9237 26312
rect 9195 26263 9237 26272
rect 9196 26178 9236 26263
rect 9100 26095 9140 26104
rect 9292 26144 9332 26935
rect 9292 26095 9332 26104
rect 9388 26144 9428 27112
rect 10060 26984 10100 27616
rect 10060 26935 10100 26944
rect 9868 26816 9908 26825
rect 9868 26321 9908 26776
rect 10059 26732 10101 26741
rect 10059 26692 10060 26732
rect 10100 26692 10101 26732
rect 10059 26683 10101 26692
rect 9867 26312 9909 26321
rect 9867 26272 9868 26312
rect 9908 26272 9909 26312
rect 9867 26263 9909 26272
rect 9388 26095 9428 26104
rect 9675 26060 9717 26069
rect 10060 26060 10100 26683
rect 10252 26153 10292 27616
rect 11692 27656 11732 27665
rect 11403 27404 11445 27413
rect 11403 27364 11404 27404
rect 11444 27364 11445 27404
rect 11403 27355 11445 27364
rect 11595 27404 11637 27413
rect 11595 27364 11596 27404
rect 11636 27364 11637 27404
rect 11595 27355 11637 27364
rect 11404 27270 11444 27355
rect 10539 26984 10581 26993
rect 10539 26944 10540 26984
rect 10580 26944 10581 26984
rect 10539 26935 10581 26944
rect 10540 26816 10580 26935
rect 10828 26825 10868 26910
rect 10540 26767 10580 26776
rect 10732 26816 10772 26825
rect 10444 26648 10484 26657
rect 10732 26648 10772 26776
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 11019 26816 11061 26825
rect 11308 26816 11348 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 11212 26776 11308 26816
rect 11020 26682 11060 26767
rect 10924 26648 10964 26657
rect 10484 26608 10772 26648
rect 10828 26608 10924 26648
rect 10444 26599 10484 26608
rect 10251 26144 10293 26153
rect 10251 26104 10252 26144
rect 10292 26104 10293 26144
rect 10251 26095 10293 26104
rect 10732 26144 10772 26153
rect 10828 26144 10868 26608
rect 10924 26599 10964 26608
rect 10924 26237 10964 26268
rect 10923 26228 10965 26237
rect 10923 26188 10924 26228
rect 10964 26188 10965 26228
rect 10923 26179 10965 26188
rect 10772 26104 10868 26144
rect 10924 26144 10964 26179
rect 10732 26095 10772 26104
rect 9675 26020 9676 26060
rect 9716 26020 9717 26060
rect 9675 26011 9717 26020
rect 9964 26020 10100 26060
rect 10155 26060 10197 26069
rect 10155 26020 10156 26060
rect 10196 26020 10197 26060
rect 8908 25976 8948 25985
rect 8908 25640 8948 25936
rect 9676 25926 9716 26011
rect 8908 25600 9236 25640
rect 8716 25304 8756 25313
rect 8332 25264 8716 25304
rect 8716 25255 8756 25264
rect 9099 25304 9141 25313
rect 9099 25264 9100 25304
rect 9140 25264 9141 25304
rect 9196 25304 9236 25600
rect 9484 25304 9524 25313
rect 9196 25264 9484 25304
rect 9099 25255 9141 25264
rect 9484 25255 9524 25264
rect 9100 25170 9140 25255
rect 9291 24632 9333 24641
rect 9291 24592 9292 24632
rect 9332 24592 9333 24632
rect 9291 24583 9333 24592
rect 9292 24498 9332 24583
rect 8428 24464 8468 24473
rect 8236 24424 8428 24464
rect 8428 24415 8468 24424
rect 8620 24380 8660 24389
rect 8620 24053 8660 24340
rect 8619 24044 8661 24053
rect 8619 24004 8620 24044
rect 8660 24004 8661 24044
rect 8619 23995 8661 24004
rect 9964 23960 10004 26020
rect 10155 26011 10197 26020
rect 10060 25892 10100 25901
rect 10060 25313 10100 25852
rect 10059 25304 10101 25313
rect 10059 25264 10060 25304
rect 10100 25264 10101 25304
rect 10059 25255 10101 25264
rect 10156 25304 10196 26011
rect 10924 25985 10964 26104
rect 11116 26144 11156 26153
rect 11019 26060 11061 26069
rect 11019 26020 11020 26060
rect 11060 26020 11061 26060
rect 11019 26011 11061 26020
rect 10443 25976 10485 25985
rect 10443 25936 10444 25976
rect 10484 25936 10485 25976
rect 10443 25927 10485 25936
rect 10923 25976 10965 25985
rect 10923 25936 10924 25976
rect 10964 25936 10965 25976
rect 10923 25927 10965 25936
rect 10348 25304 10388 25313
rect 10156 25264 10348 25304
rect 10059 24464 10101 24473
rect 10059 24424 10060 24464
rect 10100 24424 10101 24464
rect 10059 24415 10101 24424
rect 10060 24330 10100 24415
rect 10059 24044 10101 24053
rect 10059 24004 10060 24044
rect 10100 24004 10101 24044
rect 10059 23995 10101 24004
rect 9868 23920 10004 23960
rect 8619 23792 8661 23801
rect 8619 23752 8620 23792
rect 8660 23752 8661 23792
rect 8619 23743 8661 23752
rect 8523 23708 8565 23717
rect 8523 23668 8524 23708
rect 8564 23668 8565 23708
rect 8523 23659 8565 23668
rect 8044 23248 8180 23288
rect 7947 22196 7989 22205
rect 7947 22156 7948 22196
rect 7988 22156 7989 22196
rect 7947 22147 7989 22156
rect 8044 21701 8084 23248
rect 8235 23204 8277 23213
rect 8235 23164 8236 23204
rect 8276 23164 8277 23204
rect 8235 23155 8277 23164
rect 8140 23120 8180 23129
rect 8140 22289 8180 23080
rect 8236 23045 8276 23155
rect 8331 23120 8373 23129
rect 8331 23080 8332 23120
rect 8372 23080 8373 23120
rect 8331 23071 8373 23080
rect 8428 23120 8468 23129
rect 8235 23036 8277 23045
rect 8235 22996 8236 23036
rect 8276 22996 8277 23036
rect 8235 22987 8277 22996
rect 8236 22364 8276 22987
rect 8332 22986 8372 23071
rect 8428 22625 8468 23080
rect 8524 23120 8564 23659
rect 8620 23658 8660 23743
rect 9771 23708 9813 23717
rect 9771 23668 9772 23708
rect 9812 23668 9813 23708
rect 9771 23659 9813 23668
rect 9772 23624 9812 23659
rect 9772 23573 9812 23584
rect 9868 23213 9908 23920
rect 10060 23792 10100 23995
rect 10156 23801 10196 25264
rect 10348 25255 10388 25264
rect 10347 24884 10389 24893
rect 10347 24844 10348 24884
rect 10388 24844 10389 24884
rect 10347 24835 10389 24844
rect 10251 24800 10293 24809
rect 10251 24760 10252 24800
rect 10292 24760 10293 24800
rect 10251 24751 10293 24760
rect 10252 24632 10292 24751
rect 10348 24716 10388 24835
rect 10348 24667 10388 24676
rect 10252 24583 10292 24592
rect 10444 24632 10484 25927
rect 11020 25926 11060 26011
rect 11116 25313 11156 26104
rect 11212 25388 11252 26776
rect 11308 26767 11348 26776
rect 11596 26816 11636 27355
rect 11692 27245 11732 27616
rect 11691 27236 11733 27245
rect 11691 27196 11692 27236
rect 11732 27196 11733 27236
rect 11691 27187 11733 27196
rect 11596 26767 11636 26776
rect 11692 26732 11732 26741
rect 11307 26144 11349 26153
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 11308 26010 11348 26095
rect 11500 25556 11540 25565
rect 11692 25556 11732 26692
rect 11540 25516 11732 25556
rect 11500 25507 11540 25516
rect 11307 25388 11349 25397
rect 11212 25348 11308 25388
rect 11348 25348 11349 25388
rect 11307 25339 11349 25348
rect 11115 25304 11157 25313
rect 11115 25264 11116 25304
rect 11156 25264 11157 25304
rect 11115 25255 11157 25264
rect 11308 25145 11348 25339
rect 11595 25304 11637 25313
rect 11595 25264 11596 25304
rect 11636 25264 11637 25304
rect 11595 25255 11637 25264
rect 11692 25304 11732 25516
rect 11692 25255 11732 25264
rect 11307 25136 11349 25145
rect 11307 25096 11308 25136
rect 11348 25096 11349 25136
rect 11596 25136 11636 25255
rect 11596 25096 11732 25136
rect 11307 25087 11349 25096
rect 11211 25052 11253 25061
rect 11211 25012 11212 25052
rect 11252 25012 11253 25052
rect 11211 25003 11253 25012
rect 10827 24716 10869 24725
rect 10827 24676 10828 24716
rect 10868 24676 10869 24716
rect 10827 24667 10869 24676
rect 10444 24583 10484 24592
rect 10636 24632 10676 24641
rect 10443 24464 10485 24473
rect 10443 24424 10444 24464
rect 10484 24424 10485 24464
rect 10443 24415 10485 24424
rect 10060 23743 10100 23752
rect 10155 23792 10197 23801
rect 10155 23752 10156 23792
rect 10196 23752 10197 23792
rect 10155 23743 10197 23752
rect 10444 23792 10484 24415
rect 10636 23792 10676 24592
rect 10732 24632 10772 24641
rect 10732 24305 10772 24592
rect 10828 24582 10868 24667
rect 10923 24632 10965 24641
rect 10923 24592 10924 24632
rect 10964 24592 10965 24632
rect 10923 24583 10965 24592
rect 10924 24498 10964 24583
rect 11116 24380 11156 24389
rect 10731 24296 10773 24305
rect 10731 24256 10732 24296
rect 10772 24256 10773 24296
rect 10731 24247 10773 24256
rect 11116 24053 11156 24340
rect 11115 24044 11157 24053
rect 11115 24004 11116 24044
rect 11156 24004 11157 24044
rect 11115 23995 11157 24004
rect 10636 23752 11156 23792
rect 10444 23743 10484 23752
rect 11116 23288 11156 23752
rect 11116 23239 11156 23248
rect 8619 23204 8661 23213
rect 8619 23164 8620 23204
rect 8660 23164 8661 23204
rect 8619 23155 8661 23164
rect 9867 23204 9909 23213
rect 9867 23164 9868 23204
rect 9908 23164 9909 23204
rect 9867 23155 9909 23164
rect 8524 23071 8564 23080
rect 8620 23120 8660 23155
rect 9196 23120 9236 23129
rect 8620 23069 8660 23080
rect 9100 23080 9196 23120
rect 8715 22700 8757 22709
rect 8715 22660 8716 22700
rect 8756 22660 8757 22700
rect 8715 22651 8757 22660
rect 8427 22616 8469 22625
rect 8427 22576 8428 22616
rect 8468 22576 8469 22616
rect 8427 22567 8469 22576
rect 8236 22315 8276 22324
rect 8139 22280 8181 22289
rect 8139 22240 8140 22280
rect 8180 22240 8181 22280
rect 8139 22231 8181 22240
rect 8140 21785 8180 22231
rect 8428 22205 8468 22567
rect 8716 22532 8756 22651
rect 8716 22483 8756 22492
rect 8427 22196 8469 22205
rect 8427 22156 8428 22196
rect 8468 22156 8469 22196
rect 8427 22147 8469 22156
rect 8139 21776 8181 21785
rect 8139 21736 8140 21776
rect 8180 21736 8181 21776
rect 8139 21727 8181 21736
rect 9003 21776 9045 21785
rect 9003 21736 9004 21776
rect 9044 21736 9045 21776
rect 9003 21727 9045 21736
rect 8043 21692 8085 21701
rect 8043 21652 8044 21692
rect 8084 21652 8085 21692
rect 8043 21643 8085 21652
rect 9004 21642 9044 21727
rect 7852 21608 7892 21617
rect 7756 21568 7852 21608
rect 7892 21568 7988 21608
rect 7659 21559 7701 21568
rect 7852 21559 7892 21568
rect 6795 20264 6837 20273
rect 6795 20224 6796 20264
rect 6836 20224 6837 20264
rect 6795 20215 6837 20224
rect 7372 20180 7412 20728
rect 7372 20140 7508 20180
rect 6796 20096 6836 20105
rect 6700 20056 6796 20096
rect 6796 20047 6836 20056
rect 6988 20096 7028 20107
rect 6988 20021 7028 20056
rect 7084 20096 7124 20105
rect 6987 20012 7029 20021
rect 6987 19972 6988 20012
rect 7028 19972 7029 20012
rect 6987 19963 7029 19972
rect 7084 19937 7124 20056
rect 7468 20021 7508 20140
rect 7660 20096 7700 21559
rect 7660 20047 7700 20056
rect 7852 20600 7892 20609
rect 7467 20012 7509 20021
rect 7467 19972 7468 20012
rect 7508 19972 7509 20012
rect 7467 19963 7509 19972
rect 6795 19928 6837 19937
rect 6795 19888 6796 19928
rect 6836 19888 6837 19928
rect 6795 19879 6837 19888
rect 7083 19928 7125 19937
rect 7852 19928 7892 20560
rect 7948 20105 7988 21568
rect 8043 21440 8085 21449
rect 8043 21400 8044 21440
rect 8084 21400 8085 21440
rect 8043 21391 8085 21400
rect 7947 20096 7989 20105
rect 7947 20056 7948 20096
rect 7988 20056 7989 20096
rect 7947 20047 7989 20056
rect 7083 19888 7084 19928
rect 7124 19888 7125 19928
rect 7083 19879 7125 19888
rect 7849 19888 7892 19928
rect 6796 19794 6836 19879
rect 7849 19844 7889 19888
rect 7948 19844 7988 20047
rect 7849 19804 7892 19844
rect 6891 19424 6933 19433
rect 6891 19384 6892 19424
rect 6932 19384 6933 19424
rect 6891 19375 6933 19384
rect 6220 19207 6260 19216
rect 6892 19256 6932 19375
rect 6892 19207 6932 19216
rect 7756 19256 7796 19265
rect 4779 19172 4821 19181
rect 4779 19132 4780 19172
rect 4820 19132 4821 19172
rect 4779 19123 4821 19132
rect 6027 19172 6069 19181
rect 6027 19132 6028 19172
rect 6068 19132 6069 19172
rect 6027 19123 6069 19132
rect 6124 19122 6164 19207
rect 6508 19172 6548 19181
rect 6548 19132 6836 19172
rect 6508 19123 6548 19132
rect 4107 19088 4149 19097
rect 4107 19048 4108 19088
rect 4148 19048 4149 19088
rect 4107 19039 4149 19048
rect 5164 19088 5204 19097
rect 4108 18954 4148 19039
rect 4203 19004 4245 19013
rect 4203 18964 4204 19004
rect 4244 18964 4245 19004
rect 4203 18955 4245 18964
rect 4011 17660 4053 17669
rect 4204 17660 4244 18955
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4588 18752 4628 18761
rect 4780 18752 4820 18761
rect 4628 18712 4780 18752
rect 4588 18703 4628 18712
rect 4780 18703 4820 18712
rect 4875 18584 4917 18593
rect 4875 18544 4876 18584
rect 4916 18544 4917 18584
rect 4875 18535 4917 18544
rect 4876 18450 4916 18535
rect 4588 18332 4628 18341
rect 4492 18292 4588 18332
rect 4396 17753 4436 17838
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4492 17744 4532 18292
rect 4588 18283 4628 18292
rect 5068 18332 5108 18341
rect 4684 17921 4724 18006
rect 4683 17912 4725 17921
rect 4683 17872 4684 17912
rect 4724 17872 4725 17912
rect 4683 17863 4725 17872
rect 4684 17744 4724 17753
rect 4876 17744 4916 17753
rect 4011 17620 4012 17660
rect 4052 17620 4053 17660
rect 4011 17611 4053 17620
rect 4108 17620 4244 17660
rect 3915 17492 3957 17501
rect 3915 17452 3916 17492
rect 3956 17452 3957 17492
rect 3915 17443 3957 17452
rect 3819 17324 3861 17333
rect 3819 17284 3820 17324
rect 3860 17284 3861 17324
rect 3819 17275 3861 17284
rect 3723 17240 3765 17249
rect 3723 17200 3724 17240
rect 3764 17200 3765 17240
rect 3723 17191 3765 17200
rect 3724 17106 3764 17191
rect 3244 16938 3284 17023
rect 3339 16988 3381 16997
rect 3339 16948 3340 16988
rect 3380 16948 3381 16988
rect 3339 16939 3381 16948
rect 3340 16854 3380 16939
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 3628 16577 3668 17032
rect 3820 17072 3860 17083
rect 3820 16997 3860 17032
rect 3916 17072 3956 17443
rect 4108 17324 4148 17620
rect 4492 17576 4532 17704
rect 4588 17704 4684 17744
rect 4588 17585 4628 17704
rect 4684 17695 4724 17704
rect 4780 17704 4876 17744
rect 3916 17023 3956 17032
rect 4012 17284 4148 17324
rect 4204 17536 4532 17576
rect 4587 17576 4629 17585
rect 4587 17536 4588 17576
rect 4628 17536 4629 17576
rect 3819 16988 3861 16997
rect 3819 16948 3820 16988
rect 3860 16948 3861 16988
rect 3819 16939 3861 16948
rect 4012 16904 4052 17284
rect 4107 17156 4149 17165
rect 4107 17116 4108 17156
rect 4148 17116 4149 17156
rect 4107 17107 4149 17116
rect 4108 17022 4148 17107
rect 4204 17081 4244 17536
rect 4587 17527 4629 17536
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4395 17240 4437 17249
rect 4780 17240 4820 17704
rect 4876 17695 4916 17704
rect 4971 17744 5013 17753
rect 4971 17704 4972 17744
rect 5012 17704 5013 17744
rect 4971 17695 5013 17704
rect 4395 17200 4396 17240
rect 4436 17200 4437 17240
rect 4395 17191 4437 17200
rect 4588 17200 4820 17240
rect 4875 17240 4917 17249
rect 4972 17240 5012 17695
rect 5068 17501 5108 18292
rect 5164 17753 5204 19048
rect 6316 19088 6356 19097
rect 6316 18845 6356 19048
rect 6315 18836 6357 18845
rect 6315 18796 6316 18836
rect 6356 18796 6357 18836
rect 6315 18787 6357 18796
rect 6796 18752 6836 19132
rect 7756 18929 7796 19216
rect 7852 19181 7892 19804
rect 7851 19172 7893 19181
rect 7851 19132 7852 19172
rect 7892 19132 7893 19172
rect 7851 19123 7893 19132
rect 6987 18920 7029 18929
rect 6987 18880 6988 18920
rect 7028 18880 7029 18920
rect 6987 18871 7029 18880
rect 7755 18920 7797 18929
rect 7755 18880 7756 18920
rect 7796 18880 7797 18920
rect 7755 18871 7797 18880
rect 6796 18703 6836 18712
rect 6604 18584 6644 18593
rect 5740 18460 6164 18500
rect 5740 18416 5780 18460
rect 5740 18367 5780 18376
rect 5932 18332 5972 18341
rect 5836 18292 5932 18332
rect 5163 17744 5205 17753
rect 5163 17704 5164 17744
rect 5204 17704 5205 17744
rect 5163 17695 5205 17704
rect 5740 17744 5780 17753
rect 5836 17744 5876 18292
rect 5932 18283 5972 18292
rect 5931 18164 5973 18173
rect 5931 18124 5932 18164
rect 5972 18124 5973 18164
rect 5931 18115 5973 18124
rect 5780 17704 5876 17744
rect 5740 17695 5780 17704
rect 5259 17660 5301 17669
rect 5259 17620 5260 17660
rect 5300 17620 5301 17660
rect 5259 17611 5301 17620
rect 5163 17576 5205 17585
rect 5163 17536 5164 17576
rect 5204 17536 5205 17576
rect 5163 17527 5205 17536
rect 5067 17492 5109 17501
rect 5067 17452 5068 17492
rect 5108 17452 5109 17492
rect 5067 17443 5109 17452
rect 4875 17200 4876 17240
rect 4916 17200 5108 17240
rect 4396 17106 4436 17191
rect 4203 17072 4245 17081
rect 4203 17032 4204 17072
rect 4244 17032 4245 17072
rect 4203 17023 4245 17032
rect 4300 17072 4340 17081
rect 4300 16913 4340 17032
rect 4299 16904 4341 16913
rect 4012 16864 4300 16904
rect 4340 16864 4341 16904
rect 4299 16855 4341 16864
rect 4300 16770 4340 16855
rect 3627 16568 3669 16577
rect 3627 16528 3628 16568
rect 3668 16528 3669 16568
rect 3627 16519 3669 16528
rect 3628 16409 3668 16519
rect 4588 16409 4628 17200
rect 4875 17191 4917 17200
rect 4684 17072 4724 17081
rect 4684 16997 4724 17032
rect 4779 17072 4821 17081
rect 4779 17032 4780 17072
rect 4820 17032 4821 17072
rect 4779 17023 4821 17032
rect 4876 17072 4916 17191
rect 4876 17023 4916 17032
rect 4972 17072 5012 17081
rect 4683 16988 4725 16997
rect 4683 16948 4684 16988
rect 4724 16948 4725 16988
rect 4683 16939 4725 16948
rect 4684 16493 4724 16939
rect 4780 16938 4820 17023
rect 4972 16913 5012 17032
rect 4971 16904 5013 16913
rect 4971 16864 4972 16904
rect 5012 16864 5013 16904
rect 4971 16855 5013 16864
rect 4683 16484 4725 16493
rect 4683 16444 4684 16484
rect 4724 16444 4725 16484
rect 4683 16435 4725 16444
rect 1420 16400 1460 16409
rect 843 15812 885 15821
rect 843 15772 844 15812
rect 884 15772 885 15812
rect 843 15763 885 15772
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 939 15560 981 15569
rect 939 15520 940 15560
rect 980 15520 981 15560
rect 939 15511 981 15520
rect 1324 15560 1364 15569
rect 1420 15560 1460 16360
rect 2859 16400 2901 16409
rect 2859 16360 2860 16400
rect 2900 16360 2901 16400
rect 2859 16351 2901 16360
rect 3339 16400 3381 16409
rect 3339 16360 3340 16400
rect 3380 16360 3381 16400
rect 3339 16351 3381 16360
rect 3627 16400 3669 16409
rect 3627 16360 3628 16400
rect 3668 16360 3669 16400
rect 3627 16351 3669 16360
rect 4587 16400 4629 16409
rect 4587 16360 4588 16400
rect 4628 16360 4629 16400
rect 4587 16351 4629 16360
rect 1364 15520 1460 15560
rect 2188 15560 2228 15569
rect 1324 15511 1364 15520
rect 940 15426 980 15511
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 1516 14888 1556 14897
rect 652 14552 692 14839
rect 1036 14552 1076 14561
rect 652 14503 692 14512
rect 940 14512 1036 14552
rect 940 14057 980 14512
rect 1036 14503 1076 14512
rect 1035 14132 1077 14141
rect 1035 14092 1036 14132
rect 1076 14092 1077 14132
rect 1035 14083 1077 14092
rect 939 14048 981 14057
rect 939 14008 940 14048
rect 980 14008 981 14048
rect 939 13999 981 14008
rect 1036 14048 1076 14083
rect 1036 13997 1076 14008
rect 1420 14048 1460 14057
rect 1516 14048 1556 14848
rect 1460 14008 1556 14048
rect 2188 14048 2228 15520
rect 2860 14729 2900 16351
rect 3051 16232 3093 16241
rect 3051 16192 3052 16232
rect 3092 16192 3093 16232
rect 3051 16183 3093 16192
rect 3244 16232 3284 16241
rect 3340 16232 3380 16351
rect 3436 16232 3476 16241
rect 3340 16192 3436 16232
rect 3052 16098 3092 16183
rect 3147 16148 3189 16157
rect 3147 16108 3148 16148
rect 3188 16108 3189 16148
rect 3147 16099 3189 16108
rect 3148 16014 3188 16099
rect 3244 15653 3284 16192
rect 3436 16183 3476 16192
rect 3628 16232 3668 16243
rect 3628 16157 3668 16192
rect 3724 16232 3764 16241
rect 4011 16232 4053 16241
rect 3764 16192 3860 16232
rect 3724 16183 3764 16192
rect 3627 16148 3669 16157
rect 3627 16108 3628 16148
rect 3668 16108 3669 16148
rect 3627 16099 3669 16108
rect 3532 16064 3572 16073
rect 3243 15644 3285 15653
rect 3243 15604 3244 15644
rect 3284 15604 3285 15644
rect 3243 15595 3285 15604
rect 3532 15569 3572 16024
rect 3820 15728 3860 16192
rect 4011 16192 4012 16232
rect 4052 16192 4053 16232
rect 4011 16183 4053 16192
rect 4684 16232 4724 16241
rect 4972 16232 5012 16855
rect 4724 16192 4916 16232
rect 4684 16183 4724 16192
rect 4012 15728 4052 16183
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4108 15728 4148 15737
rect 3820 15679 3860 15688
rect 3916 15688 4108 15728
rect 4148 15688 4340 15728
rect 3627 15644 3669 15653
rect 3627 15604 3628 15644
rect 3668 15604 3669 15644
rect 3627 15595 3669 15604
rect 3531 15560 3573 15569
rect 3531 15520 3532 15560
rect 3572 15520 3573 15560
rect 3531 15511 3573 15520
rect 3340 15317 3380 15402
rect 3339 15308 3381 15317
rect 3339 15268 3340 15308
rect 3380 15268 3381 15308
rect 3339 15259 3381 15268
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 2955 14888 2997 14897
rect 2955 14848 2956 14888
rect 2996 14848 2997 14888
rect 2955 14839 2997 14848
rect 3435 14888 3477 14897
rect 3435 14848 3436 14888
rect 3476 14848 3477 14888
rect 3435 14839 3477 14848
rect 2859 14720 2901 14729
rect 2859 14680 2860 14720
rect 2900 14680 2901 14720
rect 2859 14671 2901 14680
rect 2956 14720 2996 14839
rect 3436 14754 3476 14839
rect 2956 14671 2996 14680
rect 3052 14720 3092 14729
rect 2284 14048 2324 14057
rect 2188 14008 2284 14048
rect 1420 13999 1460 14008
rect 2284 13217 2324 14008
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 2283 13208 2325 13217
rect 2283 13168 2284 13208
rect 2324 13168 2325 13208
rect 2283 13159 2325 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 652 12704 692 12713
rect 652 12377 692 12664
rect 2860 12545 2900 14671
rect 3052 13796 3092 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3531 14720 3573 14729
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 3628 14720 3668 15595
rect 3916 15560 3956 15688
rect 4108 15679 4148 15688
rect 3724 15520 3956 15560
rect 4011 15560 4053 15569
rect 4011 15520 4012 15560
rect 4052 15520 4053 15560
rect 3724 14751 3764 15520
rect 4011 15511 4053 15520
rect 4300 15560 4340 15688
rect 4395 15644 4437 15653
rect 4395 15604 4396 15644
rect 4436 15604 4437 15644
rect 4395 15595 4437 15604
rect 4300 15511 4340 15520
rect 4396 15560 4436 15595
rect 4012 15426 4052 15511
rect 3724 14702 3764 14711
rect 3820 15308 3860 15317
rect 4396 15308 4436 15520
rect 4491 15560 4533 15569
rect 4491 15520 4492 15560
rect 4532 15520 4533 15560
rect 4491 15511 4533 15520
rect 4588 15560 4628 15569
rect 4780 15560 4820 15569
rect 4628 15520 4724 15560
rect 4588 15511 4628 15520
rect 3628 14671 3668 14680
rect 3244 14586 3284 14671
rect 3148 14552 3188 14561
rect 3148 14141 3188 14512
rect 3147 14132 3189 14141
rect 3147 14092 3148 14132
rect 3188 14092 3189 14132
rect 3147 14083 3189 14092
rect 3532 14048 3572 14671
rect 3724 14561 3764 14646
rect 3723 14552 3765 14561
rect 3723 14512 3724 14552
rect 3764 14512 3765 14552
rect 3723 14503 3765 14512
rect 3820 14384 3860 15268
rect 4204 15268 4436 15308
rect 4204 14720 4244 15268
rect 4395 15140 4437 15149
rect 4395 15100 4396 15140
rect 4436 15100 4437 15140
rect 4395 15091 4437 15100
rect 4011 14552 4053 14561
rect 4011 14512 4012 14552
rect 4052 14512 4053 14552
rect 4011 14503 4053 14512
rect 3532 13999 3572 14008
rect 3724 14344 3860 14384
rect 3531 13880 3573 13889
rect 3531 13840 3532 13880
rect 3572 13840 3573 13880
rect 3531 13831 3573 13840
rect 2956 13756 3092 13796
rect 2859 12536 2901 12545
rect 2859 12496 2860 12536
rect 2900 12496 2901 12536
rect 2859 12487 2901 12496
rect 2956 12461 2996 13756
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3244 13208 3284 13217
rect 3532 13208 3572 13831
rect 3284 13168 3572 13208
rect 3628 13208 3668 13217
rect 3244 13159 3284 13168
rect 3628 12629 3668 13168
rect 3627 12620 3669 12629
rect 3627 12580 3628 12620
rect 3668 12580 3669 12620
rect 3627 12571 3669 12580
rect 3724 12536 3764 14344
rect 3915 13880 3957 13889
rect 3915 13840 3916 13880
rect 3956 13840 3957 13880
rect 3915 13831 3957 13840
rect 3916 13746 3956 13831
rect 3724 12487 3764 12496
rect 3916 12536 3956 12545
rect 4012 12536 4052 14503
rect 4204 14216 4244 14680
rect 4299 14720 4341 14729
rect 4299 14680 4300 14720
rect 4340 14680 4341 14720
rect 4299 14671 4341 14680
rect 4396 14720 4436 15091
rect 4396 14671 4436 14680
rect 4492 14720 4532 15511
rect 4587 15392 4629 15401
rect 4587 15352 4588 15392
rect 4628 15352 4629 15392
rect 4587 15343 4629 15352
rect 4588 15258 4628 15343
rect 4684 15233 4724 15520
rect 4683 15224 4725 15233
rect 4683 15184 4684 15224
rect 4724 15184 4725 15224
rect 4683 15175 4725 15184
rect 4683 14972 4725 14981
rect 4683 14932 4684 14972
rect 4724 14932 4725 14972
rect 4683 14923 4725 14932
rect 4684 14838 4724 14923
rect 4780 14729 4820 15520
rect 4876 15149 4916 16192
rect 5068 16232 5108 17200
rect 5164 16997 5204 17527
rect 5163 16988 5205 16997
rect 5163 16948 5164 16988
rect 5204 16948 5205 16988
rect 5163 16939 5205 16948
rect 5163 16820 5205 16829
rect 5163 16780 5164 16820
rect 5204 16780 5205 16820
rect 5163 16771 5205 16780
rect 5164 16686 5204 16771
rect 5164 16232 5204 16241
rect 5068 16192 5164 16232
rect 4972 16183 5012 16192
rect 5164 16183 5204 16192
rect 5068 16064 5108 16073
rect 5260 16064 5300 17611
rect 5548 17576 5588 17585
rect 5588 17536 5780 17576
rect 5548 17527 5588 17536
rect 5355 17492 5397 17501
rect 5355 17452 5356 17492
rect 5396 17452 5397 17492
rect 5355 17443 5397 17452
rect 5356 16232 5396 17443
rect 5644 17072 5684 17081
rect 5644 16829 5684 17032
rect 5740 17072 5780 17536
rect 5836 17240 5876 17249
rect 5932 17240 5972 18115
rect 6124 17744 6164 18460
rect 6604 18173 6644 18544
rect 6603 18164 6645 18173
rect 6603 18124 6604 18164
rect 6644 18124 6645 18164
rect 6603 18115 6645 18124
rect 6699 17912 6741 17921
rect 6699 17872 6700 17912
rect 6740 17872 6741 17912
rect 6699 17863 6741 17872
rect 6124 17695 6164 17704
rect 5876 17200 5972 17240
rect 5836 17191 5876 17200
rect 5740 17023 5780 17032
rect 5932 17072 5972 17081
rect 5643 16820 5685 16829
rect 5548 16780 5644 16820
rect 5684 16780 5685 16820
rect 5452 16409 5492 16494
rect 5451 16400 5493 16409
rect 5451 16360 5452 16400
rect 5492 16360 5493 16400
rect 5451 16351 5493 16360
rect 5452 16232 5492 16241
rect 5356 16192 5452 16232
rect 5452 16183 5492 16192
rect 5108 16024 5300 16064
rect 5068 16015 5108 16024
rect 5548 15905 5588 16780
rect 5643 16771 5685 16780
rect 5932 16493 5972 17032
rect 6124 17072 6164 17081
rect 6164 17032 6260 17072
rect 6124 17023 6164 17032
rect 5931 16484 5973 16493
rect 5931 16444 5932 16484
rect 5972 16444 5973 16484
rect 5931 16435 5973 16444
rect 5643 16400 5685 16409
rect 5643 16360 5644 16400
rect 5684 16360 5685 16400
rect 5643 16351 5685 16360
rect 5644 16232 5684 16351
rect 5644 16183 5684 16192
rect 5740 16232 5780 16241
rect 5835 16232 5877 16241
rect 5780 16192 5836 16232
rect 5876 16192 5877 16232
rect 5740 16183 5780 16192
rect 5835 16183 5877 16192
rect 5932 16232 5972 16241
rect 4971 15896 5013 15905
rect 4971 15856 4972 15896
rect 5012 15856 5013 15896
rect 4971 15847 5013 15856
rect 5547 15896 5589 15905
rect 5547 15856 5548 15896
rect 5588 15856 5589 15896
rect 5547 15847 5589 15856
rect 4972 15569 5012 15847
rect 4971 15560 5013 15569
rect 4971 15520 4972 15560
rect 5012 15520 5013 15560
rect 4971 15511 5013 15520
rect 5355 15560 5397 15569
rect 5355 15520 5356 15560
rect 5396 15520 5397 15560
rect 5355 15511 5397 15520
rect 4875 15140 4917 15149
rect 4875 15100 4876 15140
rect 4916 15100 4917 15140
rect 4875 15091 4917 15100
rect 4971 14972 5013 14981
rect 4971 14932 4972 14972
rect 5012 14932 5013 14972
rect 4971 14923 5013 14932
rect 4492 14671 4532 14680
rect 4779 14720 4821 14729
rect 4779 14680 4780 14720
rect 4820 14680 4821 14720
rect 4779 14671 4821 14680
rect 4300 14586 4340 14671
rect 4876 14552 4916 14561
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4780 14216 4820 14225
rect 4204 14176 4780 14216
rect 4780 14167 4820 14176
rect 4588 14048 4628 14057
rect 4204 14008 4588 14048
rect 4204 12704 4244 14008
rect 4588 13999 4628 14008
rect 4491 13208 4533 13217
rect 4491 13168 4492 13208
rect 4532 13168 4533 13208
rect 4491 13159 4533 13168
rect 4492 13074 4532 13159
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4876 12704 4916 14512
rect 4204 12664 4340 12704
rect 4300 12620 4340 12664
rect 4300 12571 4340 12580
rect 4396 12664 4916 12704
rect 3956 12496 4052 12536
rect 4203 12536 4245 12545
rect 4203 12496 4204 12536
rect 4244 12496 4245 12536
rect 3916 12487 3956 12496
rect 4203 12487 4245 12496
rect 4396 12536 4436 12664
rect 4396 12487 4436 12496
rect 4492 12536 4532 12547
rect 4972 12545 5012 14923
rect 5163 14552 5205 14561
rect 5163 14512 5164 14552
rect 5204 14512 5205 14552
rect 5163 14503 5205 14512
rect 2955 12452 2997 12461
rect 2955 12412 2956 12452
rect 2996 12412 2997 12452
rect 2955 12403 2997 12412
rect 3819 12452 3861 12461
rect 3819 12412 3820 12452
rect 3860 12412 3861 12452
rect 3819 12403 3861 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 3820 12318 3860 12403
rect 4204 12402 4244 12487
rect 4492 12461 4532 12496
rect 4683 12536 4725 12545
rect 4683 12496 4684 12536
rect 4724 12496 4725 12536
rect 4683 12487 4725 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 5164 12536 5204 14503
rect 5356 12620 5396 15511
rect 5452 15308 5492 15317
rect 5452 15149 5492 15268
rect 5644 15308 5684 15317
rect 5547 15224 5589 15233
rect 5547 15184 5548 15224
rect 5588 15184 5589 15224
rect 5547 15175 5589 15184
rect 5451 15140 5493 15149
rect 5451 15100 5452 15140
rect 5492 15100 5493 15140
rect 5451 15091 5493 15100
rect 5452 14645 5492 15091
rect 5548 14720 5588 15175
rect 5548 14671 5588 14680
rect 5451 14636 5493 14645
rect 5451 14596 5452 14636
rect 5492 14596 5493 14636
rect 5451 14587 5493 14596
rect 5644 14132 5684 15268
rect 5644 14083 5684 14092
rect 5740 14552 5780 14561
rect 5452 14048 5492 14057
rect 5492 14008 5588 14048
rect 5452 13999 5492 14008
rect 5548 13460 5588 14008
rect 5644 13460 5684 13469
rect 5548 13420 5644 13460
rect 5644 13411 5684 13420
rect 5740 13292 5780 14512
rect 5836 13889 5876 16183
rect 5932 14897 5972 16192
rect 6124 16232 6164 16241
rect 6028 16064 6068 16073
rect 6028 15233 6068 16024
rect 6124 15653 6164 16192
rect 6123 15644 6165 15653
rect 6123 15604 6124 15644
rect 6164 15604 6165 15644
rect 6123 15595 6165 15604
rect 6027 15224 6069 15233
rect 6027 15184 6028 15224
rect 6068 15184 6069 15224
rect 6027 15175 6069 15184
rect 6220 14897 6260 17032
rect 6411 16568 6453 16577
rect 6411 16528 6412 16568
rect 6452 16528 6453 16568
rect 6411 16519 6453 16528
rect 6412 16484 6452 16519
rect 6412 16433 6452 16444
rect 6604 16316 6644 16325
rect 6508 16276 6604 16316
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 6412 16098 6452 16183
rect 6508 16157 6548 16276
rect 6604 16267 6644 16276
rect 6507 16148 6549 16157
rect 6507 16108 6508 16148
rect 6548 16108 6549 16148
rect 6507 16099 6549 16108
rect 6315 15560 6357 15569
rect 6508 15560 6548 15569
rect 6315 15520 6316 15560
rect 6356 15520 6357 15560
rect 6315 15511 6357 15520
rect 6412 15520 6508 15560
rect 6316 15426 6356 15511
rect 6412 15149 6452 15520
rect 6508 15511 6548 15520
rect 6604 15560 6644 15571
rect 6604 15485 6644 15520
rect 6603 15476 6645 15485
rect 6603 15436 6604 15476
rect 6644 15436 6645 15476
rect 6603 15427 6645 15436
rect 6700 15476 6740 17863
rect 6988 17744 7028 18871
rect 7659 18836 7701 18845
rect 7659 18796 7660 18836
rect 7700 18796 7701 18836
rect 7659 18787 7701 18796
rect 7468 18584 7508 18593
rect 7468 18416 7508 18544
rect 7660 18584 7700 18787
rect 7660 18535 7700 18544
rect 7852 18584 7892 19123
rect 7948 18929 7988 19804
rect 7947 18920 7989 18929
rect 7947 18880 7948 18920
rect 7988 18880 7989 18920
rect 7947 18871 7989 18880
rect 7660 18416 7700 18425
rect 7468 18376 7660 18416
rect 7660 18367 7700 18376
rect 6988 17695 7028 17704
rect 7852 17660 7892 18544
rect 7948 18584 7988 18593
rect 8044 18584 8084 21391
rect 8812 20768 8852 20777
rect 8812 20609 8852 20728
rect 9004 20768 9044 20777
rect 9100 20768 9140 23080
rect 9196 23071 9236 23080
rect 9292 23120 9332 23129
rect 9292 22709 9332 23080
rect 9388 23120 9428 23129
rect 9291 22700 9333 22709
rect 9291 22660 9292 22700
rect 9332 22660 9333 22700
rect 9291 22651 9333 22660
rect 9388 22625 9428 23080
rect 9484 23120 9524 23129
rect 9676 23120 9716 23129
rect 9524 23080 9676 23120
rect 9484 23071 9524 23080
rect 9676 23071 9716 23080
rect 9868 23120 9908 23155
rect 9868 23070 9908 23080
rect 9963 23120 10005 23129
rect 9963 23080 9964 23120
rect 10004 23080 10005 23120
rect 9963 23071 10005 23080
rect 11212 23120 11252 25003
rect 11307 23792 11349 23801
rect 11307 23752 11308 23792
rect 11348 23752 11349 23792
rect 11307 23743 11349 23752
rect 11308 23658 11348 23743
rect 11403 23708 11445 23717
rect 11403 23668 11404 23708
rect 11444 23668 11445 23708
rect 11403 23659 11445 23668
rect 11404 23381 11444 23659
rect 11403 23372 11445 23381
rect 11403 23332 11404 23372
rect 11444 23332 11445 23372
rect 11403 23323 11445 23332
rect 11212 23071 11252 23080
rect 11404 23120 11444 23323
rect 11404 23071 11444 23080
rect 9964 22986 10004 23071
rect 10348 22952 10388 22961
rect 10388 22912 10868 22952
rect 10348 22903 10388 22912
rect 9676 22868 9716 22877
rect 9387 22616 9429 22625
rect 9387 22576 9388 22616
rect 9428 22576 9429 22616
rect 9387 22567 9429 22576
rect 9195 22280 9237 22289
rect 9195 22240 9196 22280
rect 9236 22240 9237 22280
rect 9195 22231 9237 22240
rect 9387 22280 9429 22289
rect 9387 22240 9388 22280
rect 9428 22240 9429 22280
rect 9387 22231 9429 22240
rect 9580 22280 9620 22289
rect 9676 22280 9716 22828
rect 10635 22700 10677 22709
rect 10635 22660 10636 22700
rect 10676 22660 10677 22700
rect 10635 22651 10677 22660
rect 9771 22616 9813 22625
rect 9771 22576 9772 22616
rect 9812 22576 9813 22616
rect 9771 22567 9813 22576
rect 9620 22240 9716 22280
rect 9580 22231 9620 22240
rect 9196 21776 9236 22231
rect 9388 22146 9428 22231
rect 9196 21727 9236 21736
rect 9044 20728 9140 20768
rect 9292 20768 9332 20779
rect 8811 20600 8853 20609
rect 8811 20560 8812 20600
rect 8852 20560 8853 20600
rect 8811 20551 8853 20560
rect 9004 20105 9044 20728
rect 9292 20693 9332 20728
rect 9580 20768 9620 20777
rect 9291 20684 9333 20693
rect 9291 20644 9292 20684
rect 9332 20644 9333 20684
rect 9291 20635 9333 20644
rect 9580 20609 9620 20728
rect 9676 20768 9716 20779
rect 9676 20693 9716 20728
rect 9772 20768 9812 22567
rect 10636 22280 10676 22651
rect 10636 22231 10676 22240
rect 10252 22112 10292 22121
rect 10252 21701 10292 22072
rect 10251 21692 10293 21701
rect 10251 21652 10252 21692
rect 10292 21652 10293 21692
rect 10251 21643 10293 21652
rect 10347 21608 10389 21617
rect 10347 21568 10348 21608
rect 10388 21568 10389 21608
rect 10828 21608 10868 22912
rect 11320 22541 11360 22560
rect 11308 22532 11360 22541
rect 11403 22532 11445 22541
rect 11348 22492 11404 22532
rect 11444 22492 11445 22532
rect 11308 22483 11348 22492
rect 11403 22483 11445 22492
rect 10924 22280 10964 22289
rect 10924 21785 10964 22240
rect 11019 22280 11061 22289
rect 11019 22240 11020 22280
rect 11060 22240 11061 22280
rect 11019 22231 11061 22240
rect 11020 22146 11060 22231
rect 10923 21776 10965 21785
rect 10923 21736 10924 21776
rect 10964 21736 10965 21776
rect 10923 21727 10965 21736
rect 11595 21692 11637 21701
rect 11595 21652 11596 21692
rect 11636 21652 11637 21692
rect 11595 21643 11637 21652
rect 11212 21608 11252 21617
rect 10828 21568 11212 21608
rect 10347 21559 10389 21568
rect 11212 21559 11252 21568
rect 10348 21474 10388 21559
rect 11596 21558 11636 21643
rect 11692 21020 11732 25096
rect 11787 24632 11829 24641
rect 11787 24592 11788 24632
rect 11828 24592 11829 24632
rect 11787 24583 11829 24592
rect 11788 24498 11828 24583
rect 11884 22541 11924 28288
rect 12076 28328 12116 28337
rect 11980 28244 12020 28253
rect 11980 27497 12020 28204
rect 11979 27488 12021 27497
rect 11979 27448 11980 27488
rect 12020 27448 12021 27488
rect 11979 27439 12021 27448
rect 11979 27068 12021 27077
rect 11979 27028 11980 27068
rect 12020 27028 12021 27068
rect 11979 27019 12021 27028
rect 11980 26934 12020 27019
rect 12076 26153 12116 28288
rect 12172 27824 12212 28456
rect 12172 27775 12212 27784
rect 12268 28328 12308 28337
rect 12268 27077 12308 28288
rect 12460 28328 12500 28337
rect 12364 28244 12404 28253
rect 12267 27068 12309 27077
rect 12267 27028 12268 27068
rect 12308 27028 12309 27068
rect 12364 27068 12404 28204
rect 12460 27245 12500 28288
rect 12652 28328 12692 32656
rect 12939 32647 12981 32656
rect 12843 31520 12885 31529
rect 12843 31480 12844 31520
rect 12884 31480 12885 31520
rect 12843 31471 12885 31480
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 12844 31352 12884 31471
rect 12844 31303 12884 31312
rect 12940 31352 12980 32647
rect 13132 32192 13172 33076
rect 13132 32143 13172 32152
rect 13228 32864 13268 32873
rect 13228 31529 13268 32824
rect 13420 31613 13460 34336
rect 13516 34327 13556 34336
rect 13612 34301 13652 35251
rect 13804 35216 13844 35227
rect 13804 35141 13844 35176
rect 13803 35132 13845 35141
rect 13803 35092 13804 35132
rect 13844 35092 13845 35132
rect 13803 35083 13845 35092
rect 13707 35048 13749 35057
rect 13707 35008 13708 35048
rect 13748 35008 13749 35048
rect 13707 34999 13749 35008
rect 13611 34292 13653 34301
rect 13611 34252 13612 34292
rect 13652 34252 13653 34292
rect 13611 34243 13653 34252
rect 13611 34040 13653 34049
rect 13611 34000 13612 34040
rect 13652 34000 13653 34040
rect 13611 33991 13653 34000
rect 13515 33116 13557 33125
rect 13515 33076 13516 33116
rect 13556 33076 13557 33116
rect 13515 33067 13557 33076
rect 13516 32864 13556 33067
rect 13516 32815 13556 32824
rect 13612 32864 13652 33991
rect 13708 33704 13748 34999
rect 13804 34376 13844 35083
rect 13900 34460 13940 35848
rect 13996 35839 14036 35848
rect 15340 35888 15380 35897
rect 15436 35888 15476 36436
rect 15380 35848 15476 35888
rect 15724 35888 15764 35897
rect 16300 35888 16340 36520
rect 15764 35848 16340 35888
rect 15340 35839 15380 35848
rect 15724 35839 15764 35848
rect 15148 35720 15188 35729
rect 14476 35344 14708 35384
rect 13995 35300 14037 35309
rect 13995 35260 13996 35300
rect 14036 35260 14037 35300
rect 13995 35251 14037 35260
rect 13996 35166 14036 35251
rect 14092 35216 14132 35225
rect 14092 34889 14132 35176
rect 14283 35216 14325 35225
rect 14283 35176 14284 35216
rect 14324 35176 14325 35216
rect 14283 35167 14325 35176
rect 14380 35216 14420 35227
rect 14284 35082 14324 35167
rect 14380 35141 14420 35176
rect 14476 35216 14516 35344
rect 14476 35167 14516 35176
rect 14571 35216 14613 35225
rect 14571 35176 14572 35216
rect 14612 35176 14613 35216
rect 14571 35167 14613 35176
rect 14379 35132 14421 35141
rect 14379 35092 14380 35132
rect 14420 35092 14421 35132
rect 14379 35083 14421 35092
rect 14572 35082 14612 35167
rect 14668 35132 14708 35344
rect 15148 35216 15188 35680
rect 15436 35216 15476 35225
rect 15148 35176 15436 35216
rect 14668 35092 14900 35132
rect 14764 34964 14804 34973
rect 14091 34880 14133 34889
rect 14091 34840 14092 34880
rect 14132 34840 14133 34880
rect 14091 34831 14133 34840
rect 14667 34880 14709 34889
rect 14764 34880 14804 34924
rect 14860 34889 14900 35092
rect 14667 34840 14668 34880
rect 14708 34840 14804 34880
rect 14859 34880 14901 34889
rect 14859 34840 14860 34880
rect 14900 34840 14901 34880
rect 14667 34831 14709 34840
rect 14859 34831 14901 34840
rect 14379 34796 14421 34805
rect 14379 34756 14380 34796
rect 14420 34756 14421 34796
rect 14379 34747 14421 34756
rect 14188 34544 14228 34553
rect 14092 34504 14188 34544
rect 13900 34420 14036 34460
rect 13804 34327 13844 34336
rect 13899 34292 13941 34301
rect 13899 34252 13900 34292
rect 13940 34252 13941 34292
rect 13899 34243 13941 34252
rect 13900 34158 13940 34243
rect 13996 33713 14036 34420
rect 13804 33704 13844 33713
rect 13708 33664 13804 33704
rect 13804 33655 13844 33664
rect 13995 33704 14037 33713
rect 13995 33664 13996 33704
rect 14036 33664 14037 33704
rect 13995 33655 14037 33664
rect 13804 33125 13844 33210
rect 13803 33116 13845 33125
rect 13803 33076 13804 33116
rect 13844 33076 13845 33116
rect 13803 33067 13845 33076
rect 13612 32815 13652 32824
rect 13803 32864 13845 32873
rect 13803 32824 13804 32864
rect 13844 32824 13845 32864
rect 13803 32815 13845 32824
rect 13804 32730 13844 32815
rect 13995 32696 14037 32705
rect 13995 32656 13996 32696
rect 14036 32656 14037 32696
rect 13995 32647 14037 32656
rect 13996 32562 14036 32647
rect 13803 31940 13845 31949
rect 13803 31900 13804 31940
rect 13844 31900 13845 31940
rect 13803 31891 13845 31900
rect 13419 31604 13461 31613
rect 13419 31564 13420 31604
rect 13460 31564 13461 31604
rect 13419 31555 13461 31564
rect 13227 31520 13269 31529
rect 13227 31480 13228 31520
rect 13268 31480 13269 31520
rect 13227 31471 13269 31480
rect 13707 31520 13749 31529
rect 13707 31480 13708 31520
rect 13748 31480 13749 31520
rect 13707 31471 13749 31480
rect 13035 31436 13077 31445
rect 13035 31396 13036 31436
rect 13076 31396 13077 31436
rect 13035 31387 13077 31396
rect 13323 31436 13365 31445
rect 13323 31396 13324 31436
rect 13364 31396 13365 31436
rect 13323 31387 13365 31396
rect 12940 31303 12980 31312
rect 13036 31352 13076 31387
rect 12748 31218 12788 31303
rect 13036 31025 13076 31312
rect 13228 31352 13268 31361
rect 13035 31016 13077 31025
rect 13035 30976 13036 31016
rect 13076 30976 13077 31016
rect 13035 30967 13077 30976
rect 12940 30848 12980 30857
rect 13228 30848 13268 31312
rect 13324 31302 13364 31387
rect 13611 31352 13653 31361
rect 13611 31312 13612 31352
rect 13652 31312 13653 31352
rect 13611 31303 13653 31312
rect 13612 31218 13652 31303
rect 13516 31184 13556 31193
rect 13420 31144 13516 31184
rect 12980 30808 13268 30848
rect 13323 30848 13365 30857
rect 13323 30808 13324 30848
rect 13364 30808 13365 30848
rect 12940 30799 12980 30808
rect 13323 30799 13365 30808
rect 13132 30680 13172 30689
rect 13132 30437 13172 30640
rect 13324 30680 13364 30799
rect 13324 30631 13364 30640
rect 13131 30428 13173 30437
rect 13131 30388 13132 30428
rect 13172 30388 13173 30428
rect 13131 30379 13173 30388
rect 13228 30428 13268 30437
rect 12844 30008 12884 30017
rect 12844 29849 12884 29968
rect 13131 29924 13173 29933
rect 13131 29884 13132 29924
rect 13172 29884 13173 29924
rect 13131 29875 13173 29884
rect 12843 29840 12885 29849
rect 12843 29800 12844 29840
rect 12884 29800 12885 29840
rect 12843 29791 12885 29800
rect 13132 29840 13172 29875
rect 13132 29789 13172 29800
rect 13228 29681 13268 30388
rect 13420 30269 13460 31144
rect 13516 31135 13556 31144
rect 13611 31016 13653 31025
rect 13611 30976 13612 31016
rect 13652 30976 13653 31016
rect 13611 30967 13653 30976
rect 13515 30764 13557 30773
rect 13515 30724 13516 30764
rect 13556 30724 13557 30764
rect 13515 30715 13557 30724
rect 13516 30680 13556 30715
rect 13516 30629 13556 30640
rect 13612 30680 13652 30967
rect 13515 30344 13557 30353
rect 13515 30304 13516 30344
rect 13556 30304 13557 30344
rect 13515 30295 13557 30304
rect 13419 30260 13461 30269
rect 13419 30220 13420 30260
rect 13460 30220 13461 30260
rect 13419 30211 13461 30220
rect 13323 30176 13365 30185
rect 13323 30136 13324 30176
rect 13364 30136 13365 30176
rect 13323 30127 13365 30136
rect 13324 29840 13364 30127
rect 13420 29840 13460 29849
rect 13324 29800 13420 29840
rect 13420 29791 13460 29800
rect 13516 29840 13556 30295
rect 13612 30269 13652 30640
rect 13611 30260 13653 30269
rect 13611 30220 13612 30260
rect 13652 30220 13653 30260
rect 13611 30211 13653 30220
rect 13227 29672 13269 29681
rect 13516 29672 13556 29800
rect 13227 29632 13228 29672
rect 13268 29632 13269 29672
rect 13227 29623 13269 29632
rect 13324 29632 13556 29672
rect 13324 29336 13364 29632
rect 13324 29287 13364 29296
rect 13708 29000 13748 31471
rect 13804 31352 13844 31891
rect 14092 31772 14132 34504
rect 14188 34495 14228 34504
rect 14380 34376 14420 34747
rect 15436 34637 15476 35176
rect 16300 35216 16340 35227
rect 16300 35141 16340 35176
rect 16299 35132 16341 35141
rect 16299 35092 16300 35132
rect 16340 35092 16341 35132
rect 16299 35083 16341 35092
rect 16107 35048 16149 35057
rect 16107 35008 16108 35048
rect 16148 35008 16149 35048
rect 16107 34999 16149 35008
rect 15628 34964 15668 34973
rect 15435 34628 15477 34637
rect 15435 34588 15436 34628
rect 15476 34588 15477 34628
rect 15435 34579 15477 34588
rect 14955 34544 14997 34553
rect 14955 34504 14956 34544
rect 14996 34504 14997 34544
rect 14955 34495 14997 34504
rect 14380 34327 14420 34336
rect 14476 34376 14516 34385
rect 14668 34376 14708 34385
rect 14516 34336 14668 34376
rect 14476 34327 14516 34336
rect 14668 34327 14708 34336
rect 14764 34376 14804 34385
rect 14764 34217 14804 34336
rect 14956 34376 14996 34495
rect 15628 34385 15668 34924
rect 15819 34880 15861 34889
rect 15819 34840 15820 34880
rect 15860 34840 15861 34880
rect 15819 34831 15861 34840
rect 14956 34327 14996 34336
rect 15148 34376 15188 34385
rect 14859 34292 14901 34301
rect 14859 34252 14860 34292
rect 14900 34252 14901 34292
rect 14859 34243 14901 34252
rect 14763 34208 14805 34217
rect 14763 34168 14764 34208
rect 14804 34168 14805 34208
rect 14763 34159 14805 34168
rect 14860 34158 14900 34243
rect 14188 33704 14228 33713
rect 14380 33704 14420 33713
rect 14228 33664 14380 33704
rect 14188 33655 14228 33664
rect 14380 33655 14420 33664
rect 15052 33704 15092 33713
rect 14859 33452 14901 33461
rect 14859 33412 14860 33452
rect 14900 33412 14901 33452
rect 14859 33403 14901 33412
rect 14668 32864 14708 32873
rect 14284 32824 14668 32864
rect 14284 32360 14324 32824
rect 14284 32311 14324 32320
rect 14379 32108 14421 32117
rect 14379 32068 14380 32108
rect 14420 32068 14421 32108
rect 14379 32059 14421 32068
rect 14092 31732 14324 31772
rect 13804 31303 13844 31312
rect 14092 31520 14132 31529
rect 13899 31268 13941 31277
rect 13899 31228 13900 31268
rect 13940 31228 13941 31268
rect 13899 31219 13941 31228
rect 13900 31134 13940 31219
rect 14092 30857 14132 31480
rect 14091 30848 14133 30857
rect 14091 30808 14092 30848
rect 14132 30808 14133 30848
rect 14091 30799 14133 30808
rect 13804 30689 13844 30774
rect 13803 30680 13845 30689
rect 13803 30640 13804 30680
rect 13844 30640 13845 30680
rect 13803 30631 13845 30640
rect 13996 30680 14036 30689
rect 13804 30512 13844 30521
rect 13996 30512 14036 30640
rect 13844 30472 14036 30512
rect 13804 30463 13844 30472
rect 14187 30428 14229 30437
rect 14187 30388 14188 30428
rect 14228 30388 14229 30428
rect 14187 30379 14229 30388
rect 13516 28960 13748 29000
rect 13804 30008 13844 30017
rect 13419 28496 13461 28505
rect 13419 28456 13420 28496
rect 13460 28456 13461 28496
rect 13419 28447 13461 28456
rect 12747 28412 12789 28421
rect 12747 28372 12748 28412
rect 12788 28372 12789 28412
rect 12747 28363 12789 28372
rect 13323 28412 13365 28421
rect 13323 28372 13324 28412
rect 13364 28372 13365 28412
rect 13323 28363 13365 28372
rect 12652 28279 12692 28288
rect 12748 28328 12788 28363
rect 12748 28277 12788 28288
rect 12940 28328 12980 28337
rect 13131 28328 13173 28337
rect 12980 28288 13076 28328
rect 12940 28279 12980 28288
rect 12844 28160 12884 28169
rect 12844 27665 12884 28120
rect 12652 27656 12692 27665
rect 12652 27413 12692 27616
rect 12843 27656 12885 27665
rect 12843 27616 12844 27656
rect 12884 27616 12885 27656
rect 12843 27607 12885 27616
rect 13036 27656 13076 28288
rect 13131 28288 13132 28328
rect 13172 28288 13173 28328
rect 13131 28279 13173 28288
rect 13132 28194 13172 28279
rect 13132 27656 13172 27665
rect 13036 27616 13132 27656
rect 12651 27404 12693 27413
rect 12651 27364 12652 27404
rect 12692 27364 12693 27404
rect 12651 27355 12693 27364
rect 12459 27236 12501 27245
rect 12459 27196 12460 27236
rect 12500 27196 12501 27236
rect 12459 27187 12501 27196
rect 12364 27028 12596 27068
rect 12267 27019 12309 27028
rect 12459 26900 12501 26909
rect 12459 26860 12460 26900
rect 12500 26860 12501 26900
rect 12459 26851 12501 26860
rect 12171 26816 12213 26825
rect 12171 26776 12172 26816
rect 12212 26776 12213 26816
rect 12171 26767 12213 26776
rect 12268 26816 12308 26825
rect 12172 26682 12212 26767
rect 12268 26312 12308 26776
rect 12364 26816 12404 26825
rect 12364 26396 12404 26776
rect 12460 26816 12500 26851
rect 12460 26765 12500 26776
rect 12556 26573 12596 27028
rect 12555 26564 12597 26573
rect 12555 26524 12556 26564
rect 12596 26524 12597 26564
rect 12555 26515 12597 26524
rect 12652 26489 12692 27355
rect 13036 26825 13076 27616
rect 13132 27607 13172 27616
rect 13324 27656 13364 28363
rect 13324 27607 13364 27616
rect 13420 27656 13460 28447
rect 13420 27607 13460 27616
rect 13132 27404 13172 27413
rect 13172 27364 13364 27404
rect 13132 27355 13172 27364
rect 13227 27236 13269 27245
rect 13227 27196 13228 27236
rect 13268 27196 13269 27236
rect 13227 27187 13269 27196
rect 13035 26816 13077 26825
rect 13035 26776 13036 26816
rect 13076 26776 13077 26816
rect 13035 26767 13077 26776
rect 12843 26732 12885 26741
rect 12843 26692 12844 26732
rect 12884 26692 12885 26732
rect 12843 26683 12885 26692
rect 12651 26480 12693 26489
rect 12651 26440 12652 26480
rect 12692 26440 12693 26480
rect 12651 26431 12693 26440
rect 12364 26356 12500 26396
rect 12268 26272 12404 26312
rect 12075 26144 12117 26153
rect 12075 26104 12076 26144
rect 12116 26104 12117 26144
rect 12075 26095 12117 26104
rect 12268 26144 12308 26153
rect 12268 25565 12308 26104
rect 12267 25556 12309 25565
rect 12267 25516 12268 25556
rect 12308 25516 12309 25556
rect 12267 25507 12309 25516
rect 12364 25220 12404 26272
rect 12171 25136 12213 25145
rect 12171 25096 12172 25136
rect 12212 25096 12213 25136
rect 12171 25087 12213 25096
rect 11979 24968 12021 24977
rect 11979 24928 11980 24968
rect 12020 24928 12021 24968
rect 11979 24919 12021 24928
rect 11883 22532 11925 22541
rect 11883 22492 11884 22532
rect 11924 22492 11925 22532
rect 11883 22483 11925 22492
rect 11980 22280 12020 24919
rect 12172 24632 12212 25087
rect 12364 25061 12404 25180
rect 12363 25052 12405 25061
rect 12363 25012 12364 25052
rect 12404 25012 12405 25052
rect 12363 25003 12405 25012
rect 12460 24977 12500 26356
rect 12556 26144 12596 26153
rect 12556 25985 12596 26104
rect 12651 26144 12693 26153
rect 12844 26144 12884 26683
rect 13132 26144 13172 26153
rect 12651 26104 12652 26144
rect 12692 26104 12693 26144
rect 12651 26095 12693 26104
rect 12748 26104 12844 26144
rect 12652 26010 12692 26095
rect 12555 25976 12597 25985
rect 12555 25936 12556 25976
rect 12596 25936 12597 25976
rect 12555 25927 12597 25936
rect 12459 24968 12501 24977
rect 12459 24928 12460 24968
rect 12500 24928 12501 24968
rect 12459 24919 12501 24928
rect 12364 24760 12692 24800
rect 12268 24632 12308 24641
rect 12172 24592 12268 24632
rect 12075 23288 12117 23297
rect 12075 23248 12076 23288
rect 12116 23248 12117 23288
rect 12075 23239 12117 23248
rect 12076 23154 12116 23239
rect 12172 22709 12212 24592
rect 12268 24583 12308 24592
rect 12267 23624 12309 23633
rect 12267 23584 12268 23624
rect 12308 23584 12309 23624
rect 12267 23575 12309 23584
rect 12268 23120 12308 23575
rect 12364 23381 12404 24760
rect 12652 24716 12692 24760
rect 12652 24667 12692 24676
rect 12748 24641 12788 26104
rect 12844 26095 12884 26104
rect 12940 26104 13132 26144
rect 12843 25976 12885 25985
rect 12843 25936 12844 25976
rect 12884 25936 12885 25976
rect 12843 25927 12885 25936
rect 12844 25842 12884 25927
rect 12940 25472 12980 26104
rect 13132 26095 13172 26104
rect 13036 25901 13076 25986
rect 13035 25892 13077 25901
rect 13035 25852 13036 25892
rect 13076 25852 13077 25892
rect 13035 25843 13077 25852
rect 13035 25724 13077 25733
rect 13035 25684 13036 25724
rect 13076 25684 13077 25724
rect 13035 25675 13077 25684
rect 12844 25432 12980 25472
rect 12556 24632 12596 24641
rect 12460 24044 12500 24053
rect 12556 24044 12596 24592
rect 12747 24632 12789 24641
rect 12747 24592 12748 24632
rect 12788 24592 12789 24632
rect 12747 24583 12789 24592
rect 12500 24004 12596 24044
rect 12460 23995 12500 24004
rect 12459 23876 12501 23885
rect 12459 23836 12460 23876
rect 12500 23836 12501 23876
rect 12459 23827 12501 23836
rect 12363 23372 12405 23381
rect 12363 23332 12364 23372
rect 12404 23332 12405 23372
rect 12363 23323 12405 23332
rect 12268 23071 12308 23080
rect 12364 23120 12404 23129
rect 12460 23120 12500 23827
rect 12556 23801 12596 24004
rect 12844 23969 12884 25432
rect 12940 25304 12980 25315
rect 12940 25229 12980 25264
rect 12939 25220 12981 25229
rect 12939 25180 12940 25220
rect 12980 25180 12981 25220
rect 12939 25171 12981 25180
rect 12939 24380 12981 24389
rect 12939 24340 12940 24380
rect 12980 24340 12981 24380
rect 12939 24331 12981 24340
rect 12940 24246 12980 24331
rect 12843 23960 12885 23969
rect 12843 23920 12844 23960
rect 12884 23920 12885 23960
rect 12843 23911 12885 23920
rect 12555 23792 12597 23801
rect 12555 23752 12556 23792
rect 12596 23752 12597 23792
rect 12555 23743 12597 23752
rect 12652 23792 12692 23801
rect 12652 23297 12692 23752
rect 12939 23792 12981 23801
rect 12939 23752 12940 23792
rect 12980 23752 12981 23792
rect 12939 23743 12981 23752
rect 12940 23658 12980 23743
rect 12747 23624 12789 23633
rect 12747 23584 12748 23624
rect 12788 23584 12789 23624
rect 12747 23575 12789 23584
rect 12748 23490 12788 23575
rect 13036 23540 13076 25675
rect 13131 25556 13173 25565
rect 13131 25516 13132 25556
rect 13172 25516 13173 25556
rect 13131 25507 13173 25516
rect 13132 25422 13172 25507
rect 13132 24632 13172 24641
rect 13132 24389 13172 24592
rect 13228 24632 13268 27187
rect 13324 26146 13364 27364
rect 13516 27068 13556 28960
rect 13804 28505 13844 29968
rect 13899 29924 13941 29933
rect 13899 29884 13900 29924
rect 13940 29884 13941 29924
rect 13899 29875 13941 29884
rect 13900 29168 13940 29875
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 14188 29840 14228 30379
rect 14188 29791 14228 29800
rect 13996 29706 14036 29791
rect 14092 29756 14132 29765
rect 13995 29168 14037 29177
rect 13900 29128 13996 29168
rect 14036 29128 14037 29168
rect 13995 29119 14037 29128
rect 13996 29034 14036 29119
rect 14092 28589 14132 29716
rect 14284 29672 14324 31732
rect 14380 31352 14420 32059
rect 14380 31303 14420 31312
rect 14476 31352 14516 32824
rect 14668 32815 14708 32824
rect 14763 32864 14805 32873
rect 14763 32824 14764 32864
rect 14804 32824 14805 32864
rect 14763 32815 14805 32824
rect 14860 32864 14900 33403
rect 15052 33125 15092 33664
rect 15051 33116 15093 33125
rect 15051 33076 15052 33116
rect 15092 33076 15093 33116
rect 15051 33067 15093 33076
rect 14860 32815 14900 32824
rect 14668 32024 14708 32033
rect 14764 32024 14804 32815
rect 14955 32780 14997 32789
rect 14955 32740 14956 32780
rect 14996 32740 14997 32780
rect 14955 32731 14997 32740
rect 14859 32696 14901 32705
rect 14859 32656 14860 32696
rect 14900 32656 14901 32696
rect 14859 32647 14901 32656
rect 14860 32192 14900 32647
rect 14956 32360 14996 32731
rect 14956 32311 14996 32320
rect 15148 32360 15188 34336
rect 15340 34376 15380 34385
rect 15244 34208 15284 34217
rect 15244 33713 15284 34168
rect 15243 33704 15285 33713
rect 15243 33664 15244 33704
rect 15284 33664 15285 33704
rect 15243 33655 15285 33664
rect 15243 33452 15285 33461
rect 15243 33412 15244 33452
rect 15284 33412 15285 33452
rect 15243 33403 15285 33412
rect 15244 33318 15284 33403
rect 15340 33377 15380 34336
rect 15436 34376 15476 34385
rect 15339 33368 15381 33377
rect 15339 33328 15340 33368
rect 15380 33328 15381 33368
rect 15339 33319 15381 33328
rect 15243 32864 15285 32873
rect 15243 32824 15244 32864
rect 15284 32824 15285 32864
rect 15243 32815 15285 32824
rect 15244 32730 15284 32815
rect 15340 32612 15380 33319
rect 15436 32789 15476 34336
rect 15627 34376 15669 34385
rect 15627 34336 15628 34376
rect 15668 34336 15669 34376
rect 15627 34327 15669 34336
rect 15723 34292 15765 34301
rect 15723 34252 15724 34292
rect 15764 34252 15765 34292
rect 15723 34243 15765 34252
rect 15724 34158 15764 34243
rect 15435 32780 15477 32789
rect 15435 32740 15436 32780
rect 15476 32740 15477 32780
rect 15435 32731 15477 32740
rect 15340 32572 15476 32612
rect 15148 32311 15188 32320
rect 15339 32192 15381 32201
rect 14860 32143 14900 32152
rect 15244 32150 15284 32159
rect 14708 31984 14804 32024
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15339 32143 15381 32152
rect 15436 32192 15476 32572
rect 15820 32360 15860 34831
rect 16108 34376 16148 34999
rect 16396 34964 16436 36688
rect 24459 36560 24501 36569
rect 24459 36520 24460 36560
rect 24500 36520 24501 36560
rect 24459 36511 24501 36520
rect 24940 36560 24980 36569
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 19756 36056 19796 36065
rect 23884 36056 23924 36065
rect 19372 36016 19756 36056
rect 16588 35888 16628 35897
rect 16491 35216 16533 35225
rect 16491 35176 16492 35216
rect 16532 35176 16533 35216
rect 16491 35167 16533 35176
rect 16492 35082 16532 35167
rect 16492 34964 16532 34973
rect 16396 34924 16492 34964
rect 16492 34915 16532 34924
rect 16588 34385 16628 35848
rect 18987 35888 19029 35897
rect 18987 35848 18988 35888
rect 19028 35848 19029 35888
rect 18987 35839 19029 35848
rect 17740 35720 17780 35729
rect 17644 35680 17740 35720
rect 16779 35300 16821 35309
rect 16779 35260 16780 35300
rect 16820 35260 16821 35300
rect 16779 35251 16821 35260
rect 16684 35216 16724 35225
rect 16684 34973 16724 35176
rect 16780 35216 16820 35251
rect 16780 35165 16820 35176
rect 16972 35216 17012 35225
rect 16683 34964 16725 34973
rect 16683 34924 16684 34964
rect 16724 34924 16725 34964
rect 16683 34915 16725 34924
rect 16972 34553 17012 35176
rect 17068 35216 17108 35225
rect 17068 34889 17108 35176
rect 17163 35216 17205 35225
rect 17163 35176 17164 35216
rect 17204 35176 17205 35216
rect 17163 35167 17205 35176
rect 17260 35216 17300 35225
rect 17164 35082 17204 35167
rect 17067 34880 17109 34889
rect 17067 34840 17068 34880
rect 17108 34840 17109 34880
rect 17067 34831 17109 34840
rect 16971 34544 17013 34553
rect 16971 34504 16972 34544
rect 17012 34504 17013 34544
rect 16971 34495 17013 34504
rect 16108 34327 16148 34336
rect 16203 34376 16245 34385
rect 16203 34336 16204 34376
rect 16244 34336 16245 34376
rect 16203 34327 16245 34336
rect 16587 34376 16629 34385
rect 16587 34336 16588 34376
rect 16628 34336 16629 34376
rect 16587 34327 16629 34336
rect 16971 34376 17013 34385
rect 16971 34336 16972 34376
rect 17012 34336 17013 34376
rect 16971 34327 17013 34336
rect 15915 33704 15957 33713
rect 15915 33664 15916 33704
rect 15956 33664 15957 33704
rect 15915 33655 15957 33664
rect 15916 33570 15956 33655
rect 16108 32864 16148 32873
rect 16204 32864 16244 34327
rect 16972 34242 17012 34327
rect 17260 33797 17300 35176
rect 17644 35141 17684 35680
rect 17740 35671 17780 35680
rect 18892 35720 18932 35729
rect 18796 35300 18836 35309
rect 18892 35300 18932 35680
rect 18836 35260 18932 35300
rect 18796 35251 18836 35260
rect 18123 35216 18165 35225
rect 18123 35176 18124 35216
rect 18164 35176 18165 35216
rect 18123 35167 18165 35176
rect 18315 35216 18357 35225
rect 18315 35176 18316 35216
rect 18356 35176 18357 35216
rect 18315 35167 18357 35176
rect 17643 35132 17685 35141
rect 17643 35092 17644 35132
rect 17684 35092 17685 35132
rect 17643 35083 17685 35092
rect 17451 35048 17493 35057
rect 17451 35008 17452 35048
rect 17492 35008 17493 35048
rect 17451 34999 17493 35008
rect 17452 34914 17492 34999
rect 17259 33788 17301 33797
rect 17259 33748 17260 33788
rect 17300 33748 17301 33788
rect 17259 33739 17301 33748
rect 17644 33788 17684 35083
rect 18124 34628 18164 35167
rect 18316 35082 18356 35167
rect 18412 34964 18452 34973
rect 18452 34924 18740 34964
rect 18412 34915 18452 34924
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 18316 34628 18356 34637
rect 18124 34588 18316 34628
rect 18316 34579 18356 34588
rect 18507 34628 18549 34637
rect 18507 34588 18508 34628
rect 18548 34588 18549 34628
rect 18507 34579 18549 34588
rect 17739 34544 17781 34553
rect 17739 34504 17740 34544
rect 17780 34504 17781 34544
rect 17739 34495 17781 34504
rect 17644 33739 17684 33748
rect 17740 33704 17780 34495
rect 18123 34460 18165 34469
rect 18123 34420 18124 34460
rect 18164 34420 18165 34460
rect 18123 34411 18165 34420
rect 18124 34326 18164 34411
rect 17931 33788 17973 33797
rect 17931 33748 17932 33788
rect 17972 33748 17973 33788
rect 17931 33739 17973 33748
rect 17740 33655 17780 33664
rect 17356 33452 17396 33461
rect 17164 33412 17356 33452
rect 16779 32948 16821 32957
rect 16779 32908 16780 32948
rect 16820 32908 16821 32948
rect 16779 32899 16821 32908
rect 15436 32143 15476 32152
rect 15532 32320 15860 32360
rect 16012 32824 16108 32864
rect 16148 32824 16244 32864
rect 14668 31975 14708 31984
rect 15244 31940 15284 32110
rect 15340 32058 15380 32143
rect 15532 31940 15572 32320
rect 15148 31900 15572 31940
rect 15628 32192 15668 32201
rect 14763 31604 14805 31613
rect 14763 31564 14764 31604
rect 14804 31564 14805 31604
rect 14763 31555 14805 31564
rect 14476 31303 14516 31312
rect 14764 31352 14804 31555
rect 14955 31520 14997 31529
rect 14955 31480 14956 31520
rect 14996 31480 14997 31520
rect 14955 31471 14997 31480
rect 14764 31303 14804 31312
rect 14475 30680 14517 30689
rect 14475 30640 14476 30680
rect 14516 30640 14517 30680
rect 14475 30631 14517 30640
rect 14956 30680 14996 31471
rect 14956 30631 14996 30640
rect 14476 29840 14516 30631
rect 14668 30428 14708 30437
rect 14708 30388 14996 30428
rect 14668 30379 14708 30388
rect 14763 30260 14805 30269
rect 14763 30220 14764 30260
rect 14804 30220 14805 30260
rect 14763 30211 14805 30220
rect 14668 29933 14708 29964
rect 14667 29924 14709 29933
rect 14667 29884 14668 29924
rect 14708 29884 14709 29924
rect 14667 29875 14709 29884
rect 14476 29791 14516 29800
rect 14571 29840 14613 29849
rect 14571 29800 14572 29840
rect 14612 29800 14613 29840
rect 14571 29791 14613 29800
rect 14668 29840 14708 29875
rect 14572 29706 14612 29791
rect 14188 29632 14324 29672
rect 13899 28580 13941 28589
rect 13899 28540 13900 28580
rect 13940 28540 13941 28580
rect 13899 28531 13941 28540
rect 14091 28580 14133 28589
rect 14091 28540 14092 28580
rect 14132 28540 14133 28580
rect 14091 28531 14133 28540
rect 13803 28496 13845 28505
rect 13803 28456 13804 28496
rect 13844 28456 13845 28496
rect 13803 28447 13845 28456
rect 13803 28328 13845 28337
rect 13803 28288 13804 28328
rect 13844 28288 13845 28328
rect 13803 28279 13845 28288
rect 13804 28194 13844 28279
rect 13900 27908 13940 28531
rect 14091 28328 14133 28337
rect 14091 28288 14092 28328
rect 14132 28288 14133 28328
rect 14091 28279 14133 28288
rect 14092 28194 14132 28279
rect 13804 27868 13940 27908
rect 14188 27908 14228 29632
rect 14379 29252 14421 29261
rect 14379 29212 14380 29252
rect 14420 29212 14421 29252
rect 14379 29203 14421 29212
rect 14283 29168 14325 29177
rect 14283 29128 14284 29168
rect 14324 29128 14325 29168
rect 14283 29119 14325 29128
rect 14284 29034 14324 29119
rect 14380 29118 14420 29203
rect 14668 29177 14708 29800
rect 14764 29840 14804 30211
rect 14764 29791 14804 29800
rect 14956 29840 14996 30388
rect 15148 30260 15188 31900
rect 15628 31529 15668 32152
rect 15724 32192 15764 32320
rect 15724 32143 15764 32152
rect 15820 32192 15860 32203
rect 15820 32117 15860 32152
rect 15916 32192 15956 32201
rect 15819 32108 15861 32117
rect 15819 32068 15820 32108
rect 15860 32068 15861 32108
rect 15819 32059 15861 32068
rect 15916 32033 15956 32152
rect 15915 32024 15957 32033
rect 15915 31984 15916 32024
rect 15956 31984 15957 32024
rect 15915 31975 15957 31984
rect 15627 31520 15669 31529
rect 15627 31480 15628 31520
rect 15668 31480 15669 31520
rect 15627 31471 15669 31480
rect 16012 31361 16052 32824
rect 16108 32815 16148 32824
rect 16107 32192 16149 32201
rect 16107 32152 16108 32192
rect 16148 32152 16149 32192
rect 16107 32143 16149 32152
rect 16780 32192 16820 32899
rect 16780 32143 16820 32152
rect 15243 31352 15285 31361
rect 15916 31352 15956 31361
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 15820 31312 15916 31352
rect 15244 31218 15284 31303
rect 15052 30220 15188 30260
rect 15052 29849 15092 30220
rect 15820 29933 15860 31312
rect 15916 31303 15956 31312
rect 16011 31352 16053 31361
rect 16011 31312 16012 31352
rect 16052 31312 16053 31352
rect 16108 31352 16148 32143
rect 16587 32024 16629 32033
rect 16587 31984 16588 32024
rect 16628 31984 16629 32024
rect 16587 31975 16629 31984
rect 16491 31436 16533 31445
rect 16491 31396 16492 31436
rect 16532 31396 16533 31436
rect 16491 31387 16533 31396
rect 16204 31352 16244 31361
rect 16108 31312 16204 31352
rect 16011 31303 16053 31312
rect 16204 31303 16244 31312
rect 16492 31352 16532 31387
rect 15916 30680 15956 30689
rect 16012 30680 16052 31303
rect 16492 31301 16532 31312
rect 16588 31352 16628 31975
rect 16972 31940 17012 31949
rect 16779 31688 16821 31697
rect 16779 31648 16780 31688
rect 16820 31648 16821 31688
rect 16779 31639 16821 31648
rect 16683 31520 16725 31529
rect 16683 31480 16684 31520
rect 16724 31480 16725 31520
rect 16683 31471 16725 31480
rect 16780 31520 16820 31639
rect 16780 31471 16820 31480
rect 16684 31352 16724 31471
rect 16780 31352 16820 31361
rect 16684 31312 16780 31352
rect 16588 31303 16628 31312
rect 16780 31303 16820 31312
rect 16972 31352 17012 31900
rect 16972 31303 17012 31312
rect 16108 31184 16148 31193
rect 16108 30773 16148 31144
rect 16107 30764 16149 30773
rect 16107 30724 16108 30764
rect 16148 30724 16149 30764
rect 16107 30715 16149 30724
rect 15956 30640 16052 30680
rect 15916 30631 15956 30640
rect 15819 29924 15861 29933
rect 15819 29884 15820 29924
rect 15860 29884 15861 29924
rect 15819 29875 15861 29884
rect 14956 29791 14996 29800
rect 15051 29840 15093 29849
rect 15340 29840 15380 29849
rect 15051 29800 15052 29840
rect 15092 29800 15093 29840
rect 15051 29791 15093 29800
rect 15244 29800 15340 29840
rect 16012 29840 16052 30640
rect 16299 30596 16341 30605
rect 16299 30556 16300 30596
rect 16340 30556 16341 30596
rect 16299 30547 16341 30556
rect 16107 30428 16149 30437
rect 16107 30388 16108 30428
rect 16148 30388 16149 30428
rect 16107 30379 16149 30388
rect 16108 30294 16148 30379
rect 16204 29840 16244 29849
rect 16012 29800 16204 29840
rect 15051 29672 15093 29681
rect 15051 29632 15052 29672
rect 15092 29632 15093 29672
rect 15051 29623 15093 29632
rect 14667 29168 14709 29177
rect 14667 29128 14668 29168
rect 14708 29128 14709 29168
rect 14667 29119 14709 29128
rect 14668 28916 14708 28925
rect 14475 28328 14517 28337
rect 14475 28288 14476 28328
rect 14516 28288 14517 28328
rect 14475 28279 14517 28288
rect 14188 27868 14324 27908
rect 13612 27656 13652 27667
rect 13612 27581 13652 27616
rect 13707 27656 13749 27665
rect 13707 27616 13708 27656
rect 13748 27616 13749 27656
rect 13707 27607 13749 27616
rect 13804 27652 13844 27868
rect 14151 27665 14191 27750
rect 13900 27656 13940 27665
rect 13804 27616 13900 27652
rect 14150 27656 14192 27665
rect 13804 27612 13940 27616
rect 13900 27607 13940 27612
rect 13996 27627 14036 27636
rect 13611 27572 13653 27581
rect 13611 27532 13612 27572
rect 13652 27532 13653 27572
rect 13611 27523 13653 27532
rect 13708 27522 13748 27607
rect 14150 27616 14151 27656
rect 14191 27616 14192 27656
rect 14150 27607 14192 27616
rect 13899 27488 13941 27497
rect 13996 27488 14036 27587
rect 14284 27488 14324 27868
rect 13899 27448 13900 27488
rect 13940 27448 14036 27488
rect 14092 27448 14324 27488
rect 13899 27439 13941 27448
rect 13612 27404 13652 27413
rect 13652 27364 13844 27404
rect 13612 27355 13652 27364
rect 13804 27320 13844 27364
rect 13804 27280 13940 27320
rect 13516 27019 13556 27028
rect 13900 26909 13940 27280
rect 13899 26900 13941 26909
rect 13899 26860 13900 26900
rect 13940 26860 13941 26900
rect 13899 26851 13941 26860
rect 13708 26816 13748 26825
rect 13324 26137 13398 26146
rect 13324 26104 13358 26137
rect 13358 26088 13398 26097
rect 13516 26144 13556 26153
rect 13323 25472 13365 25481
rect 13323 25432 13324 25472
rect 13364 25432 13365 25472
rect 13323 25423 13365 25432
rect 13324 24800 13364 25423
rect 13516 24893 13556 26104
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13612 26010 13652 26095
rect 13611 25892 13653 25901
rect 13611 25852 13612 25892
rect 13652 25852 13653 25892
rect 13611 25843 13653 25852
rect 13515 24884 13557 24893
rect 13515 24844 13516 24884
rect 13556 24844 13557 24884
rect 13515 24835 13557 24844
rect 13324 24751 13364 24760
rect 13228 24583 13268 24592
rect 13419 24632 13461 24641
rect 13419 24592 13420 24632
rect 13460 24592 13461 24632
rect 13419 24583 13461 24592
rect 13612 24632 13652 25843
rect 13708 25229 13748 26776
rect 14092 26816 14132 27448
rect 14187 27236 14229 27245
rect 14187 27196 14188 27236
rect 14228 27196 14229 27236
rect 14187 27187 14229 27196
rect 14092 26767 14132 26776
rect 14188 26816 14228 27187
rect 14283 27152 14325 27161
rect 14283 27112 14284 27152
rect 14324 27112 14325 27152
rect 14283 27103 14325 27112
rect 14188 26767 14228 26776
rect 14284 26657 14324 27103
rect 14379 27068 14421 27077
rect 14379 27028 14380 27068
rect 14420 27028 14421 27068
rect 14379 27019 14421 27028
rect 14380 26934 14420 27019
rect 14379 26816 14421 26825
rect 14379 26776 14380 26816
rect 14420 26776 14421 26816
rect 14379 26767 14421 26776
rect 14380 26682 14420 26767
rect 13899 26648 13941 26657
rect 13899 26608 13900 26648
rect 13940 26608 13941 26648
rect 13899 26599 13941 26608
rect 14283 26648 14325 26657
rect 14283 26608 14284 26648
rect 14324 26608 14325 26648
rect 14283 26599 14325 26608
rect 13804 26144 13844 26153
rect 13804 25481 13844 26104
rect 13900 26144 13940 26599
rect 14091 26480 14133 26489
rect 14091 26440 14092 26480
rect 14132 26440 14133 26480
rect 14091 26431 14133 26440
rect 13900 26095 13940 26104
rect 13899 25892 13941 25901
rect 13899 25852 13900 25892
rect 13940 25852 13941 25892
rect 13899 25843 13941 25852
rect 13900 25758 13940 25843
rect 13803 25472 13845 25481
rect 13803 25432 13804 25472
rect 13844 25432 13845 25472
rect 13803 25423 13845 25432
rect 13803 25304 13845 25313
rect 13803 25264 13804 25304
rect 13844 25264 13845 25304
rect 13803 25255 13845 25264
rect 13996 25304 14036 25313
rect 13707 25220 13749 25229
rect 13707 25180 13708 25220
rect 13748 25180 13749 25220
rect 13707 25171 13749 25180
rect 13804 25170 13844 25255
rect 13996 24800 14036 25264
rect 14092 25304 14132 26431
rect 14187 26228 14229 26237
rect 14187 26188 14188 26228
rect 14228 26188 14229 26228
rect 14187 26179 14229 26188
rect 14092 25255 14132 25264
rect 14188 25304 14228 26179
rect 14284 26144 14324 26599
rect 14284 26095 14324 26104
rect 14380 26144 14420 26153
rect 14380 25985 14420 26104
rect 14379 25976 14421 25985
rect 14379 25936 14380 25976
rect 14420 25936 14421 25976
rect 14379 25927 14421 25936
rect 14284 25892 14324 25901
rect 14284 25649 14324 25852
rect 14283 25640 14325 25649
rect 14283 25600 14284 25640
rect 14324 25600 14325 25640
rect 14283 25591 14325 25600
rect 14283 25472 14325 25481
rect 14476 25472 14516 28279
rect 14571 28160 14613 28169
rect 14571 28120 14572 28160
rect 14612 28120 14613 28160
rect 14571 28111 14613 28120
rect 14572 28026 14612 28111
rect 14668 27824 14708 28876
rect 14572 27784 14708 27824
rect 14572 26816 14612 27784
rect 14764 27656 14804 27666
rect 14764 27581 14804 27616
rect 14860 27656 14900 27665
rect 14763 27572 14805 27581
rect 14677 27532 14764 27572
rect 14804 27532 14805 27572
rect 14677 27488 14717 27532
rect 14763 27523 14805 27532
rect 14668 27448 14717 27488
rect 14668 27161 14708 27448
rect 14763 27404 14805 27413
rect 14763 27364 14764 27404
rect 14804 27364 14805 27404
rect 14763 27355 14805 27364
rect 14764 27270 14804 27355
rect 14667 27152 14709 27161
rect 14667 27112 14668 27152
rect 14708 27112 14709 27152
rect 14667 27103 14709 27112
rect 14860 27077 14900 27616
rect 14955 27656 14997 27665
rect 14955 27616 14956 27656
rect 14996 27616 14997 27656
rect 14955 27607 14997 27616
rect 15052 27656 15092 29623
rect 15244 29000 15284 29800
rect 15340 29791 15380 29800
rect 16204 29791 16244 29800
rect 16300 29672 16340 30547
rect 16204 29632 16340 29672
rect 15339 29504 15381 29513
rect 15339 29464 15340 29504
rect 15380 29464 15381 29504
rect 15339 29455 15381 29464
rect 15244 28951 15284 28960
rect 15340 27740 15380 29455
rect 16107 29252 16149 29261
rect 16107 29212 16108 29252
rect 16148 29212 16149 29252
rect 16107 29203 16149 29212
rect 15436 29093 15476 29178
rect 16108 29168 16148 29203
rect 16108 29117 16148 29128
rect 15435 29084 15477 29093
rect 15435 29044 15436 29084
rect 15476 29044 15477 29084
rect 15435 29035 15477 29044
rect 16204 29000 16244 29632
rect 16299 29168 16341 29177
rect 16299 29128 16300 29168
rect 16340 29128 16341 29168
rect 16299 29119 16341 29128
rect 16108 28960 16244 29000
rect 15340 27700 15476 27740
rect 15052 27607 15092 27616
rect 15148 27656 15188 27665
rect 14859 27068 14901 27077
rect 14859 27028 14860 27068
rect 14900 27028 14901 27068
rect 14956 27068 14996 27607
rect 15052 27068 15092 27077
rect 14956 27028 15052 27068
rect 14859 27019 14901 27028
rect 15052 27019 15092 27028
rect 14860 26825 14900 26910
rect 14572 26767 14612 26776
rect 14668 26816 14708 26825
rect 14668 26657 14708 26776
rect 14859 26816 14901 26825
rect 15052 26816 15092 26827
rect 14859 26776 14860 26816
rect 14900 26776 14996 26816
rect 14859 26767 14901 26776
rect 14667 26648 14709 26657
rect 14667 26608 14668 26648
rect 14708 26608 14709 26648
rect 14667 26599 14709 26608
rect 14764 26648 14804 26657
rect 14571 26564 14613 26573
rect 14571 26524 14572 26564
rect 14612 26524 14613 26564
rect 14571 26515 14613 26524
rect 14572 26144 14612 26515
rect 14667 26480 14709 26489
rect 14667 26440 14668 26480
rect 14708 26440 14709 26480
rect 14764 26480 14804 26608
rect 14859 26648 14901 26657
rect 14859 26608 14860 26648
rect 14900 26608 14901 26648
rect 14859 26599 14901 26608
rect 14764 26440 14809 26480
rect 14667 26431 14709 26440
rect 14572 26095 14612 26104
rect 14668 26144 14708 26431
rect 14668 26095 14708 26104
rect 14769 26144 14809 26440
rect 14860 26321 14900 26599
rect 14859 26312 14901 26321
rect 14859 26272 14860 26312
rect 14900 26272 14901 26312
rect 14956 26312 14996 26776
rect 15052 26741 15092 26776
rect 15051 26732 15093 26741
rect 15051 26692 15052 26732
rect 15092 26692 15093 26732
rect 15051 26683 15093 26692
rect 15051 26312 15093 26321
rect 14956 26272 15052 26312
rect 15092 26272 15093 26312
rect 14859 26263 14901 26272
rect 15051 26263 15093 26272
rect 15148 26228 15188 27616
rect 15305 27641 15345 27650
rect 15305 27413 15345 27601
rect 15304 27404 15346 27413
rect 15304 27364 15305 27404
rect 15345 27364 15346 27404
rect 15304 27355 15346 27364
rect 15243 27236 15285 27245
rect 15243 27196 15244 27236
rect 15284 27196 15285 27236
rect 15243 27187 15285 27196
rect 15244 26816 15284 27187
rect 15244 26767 15284 26776
rect 15339 26816 15381 26825
rect 15339 26776 15340 26816
rect 15380 26776 15381 26816
rect 15339 26767 15381 26776
rect 15340 26682 15380 26767
rect 15148 26179 15188 26188
rect 15243 26228 15285 26237
rect 15243 26188 15244 26228
rect 15284 26188 15285 26228
rect 15243 26179 15285 26188
rect 15052 26144 15092 26153
rect 14769 26095 14809 26104
rect 14956 26104 15052 26144
rect 14283 25432 14284 25472
rect 14324 25432 14325 25472
rect 14283 25423 14325 25432
rect 14380 25432 14516 25472
rect 14763 25472 14805 25481
rect 14763 25432 14764 25472
rect 14804 25432 14805 25472
rect 14188 25255 14228 25264
rect 14284 25304 14324 25423
rect 14284 25255 14324 25264
rect 14187 24968 14229 24977
rect 14187 24928 14188 24968
rect 14228 24928 14229 24968
rect 14187 24919 14229 24928
rect 13804 24760 14036 24800
rect 13708 24725 13748 24756
rect 13707 24716 13749 24725
rect 13707 24676 13708 24716
rect 13748 24676 13749 24716
rect 13707 24667 13749 24676
rect 13612 24583 13652 24592
rect 13708 24632 13748 24667
rect 13420 24498 13460 24583
rect 13131 24380 13173 24389
rect 13131 24340 13132 24380
rect 13172 24340 13173 24380
rect 13131 24331 13173 24340
rect 13708 24053 13748 24592
rect 13804 24128 13844 24760
rect 13900 24632 13940 24641
rect 14091 24632 14133 24641
rect 13940 24592 14036 24632
rect 13900 24583 13940 24592
rect 13899 24380 13941 24389
rect 13899 24340 13900 24380
rect 13940 24340 13941 24380
rect 13899 24331 13941 24340
rect 13900 24246 13940 24331
rect 13804 24088 13940 24128
rect 13707 24044 13749 24053
rect 13707 24004 13708 24044
rect 13748 24004 13749 24044
rect 13707 23995 13749 24004
rect 13611 23960 13653 23969
rect 13611 23920 13612 23960
rect 13652 23920 13653 23960
rect 13611 23911 13653 23920
rect 13612 23826 13652 23911
rect 13708 23708 13748 23995
rect 12940 23500 13076 23540
rect 13612 23668 13748 23708
rect 12651 23288 12693 23297
rect 12651 23248 12652 23288
rect 12692 23248 12693 23288
rect 12651 23239 12693 23248
rect 12556 23129 12596 23214
rect 12404 23080 12500 23120
rect 12555 23120 12597 23129
rect 12555 23080 12556 23120
rect 12596 23080 12597 23120
rect 12364 23071 12404 23080
rect 12555 23071 12597 23080
rect 12748 23120 12788 23129
rect 12556 22952 12596 22961
rect 12748 22952 12788 23080
rect 12596 22912 12788 22952
rect 12556 22903 12596 22912
rect 12171 22700 12213 22709
rect 12171 22660 12172 22700
rect 12212 22660 12213 22700
rect 12171 22651 12213 22660
rect 12363 22700 12405 22709
rect 12363 22660 12364 22700
rect 12404 22660 12405 22700
rect 12363 22651 12405 22660
rect 12747 22700 12789 22709
rect 12747 22660 12748 22700
rect 12788 22660 12789 22700
rect 12747 22651 12789 22660
rect 12076 22280 12116 22289
rect 11980 22240 12076 22280
rect 12076 22231 12116 22240
rect 11883 21608 11925 21617
rect 11883 21568 11884 21608
rect 11924 21568 11925 21608
rect 11883 21559 11925 21568
rect 11692 20971 11732 20980
rect 11788 21440 11828 21449
rect 9772 20719 9812 20728
rect 9867 20768 9909 20777
rect 9867 20728 9868 20768
rect 9908 20728 9909 20768
rect 9867 20719 9909 20728
rect 10347 20768 10389 20777
rect 10347 20728 10348 20768
rect 10388 20728 10389 20768
rect 10347 20719 10389 20728
rect 10540 20768 10580 20777
rect 9675 20684 9717 20693
rect 9675 20644 9676 20684
rect 9716 20644 9717 20684
rect 9675 20635 9717 20644
rect 9868 20634 9908 20719
rect 10348 20634 10388 20719
rect 10540 20609 10580 20728
rect 10636 20768 10676 20777
rect 9196 20600 9236 20609
rect 9003 20096 9045 20105
rect 9003 20056 9004 20096
rect 9044 20056 9045 20096
rect 9003 20047 9045 20056
rect 9196 19937 9236 20560
rect 9579 20600 9621 20609
rect 9579 20560 9580 20600
rect 9620 20560 9621 20600
rect 9579 20551 9621 20560
rect 10444 20600 10484 20609
rect 9291 20096 9333 20105
rect 9291 20056 9292 20096
rect 9332 20056 9333 20096
rect 9291 20047 9333 20056
rect 10156 20096 10196 20107
rect 9292 19962 9332 20047
rect 10156 20021 10196 20056
rect 10444 20096 10484 20560
rect 10539 20600 10581 20609
rect 10539 20560 10540 20600
rect 10580 20560 10581 20600
rect 10539 20551 10581 20560
rect 10444 20047 10484 20056
rect 10155 20012 10197 20021
rect 10155 19972 10156 20012
rect 10196 19972 10197 20012
rect 10155 19963 10197 19972
rect 9195 19928 9237 19937
rect 9195 19888 9196 19928
rect 9236 19888 9237 19928
rect 9195 19879 9237 19888
rect 10347 19508 10389 19517
rect 10347 19468 10348 19508
rect 10388 19468 10389 19508
rect 10347 19459 10389 19468
rect 10348 19374 10388 19459
rect 8907 19340 8949 19349
rect 8907 19300 8908 19340
rect 8948 19300 8949 19340
rect 8907 19291 8949 19300
rect 8908 19206 8948 19291
rect 10444 19256 10484 19265
rect 8331 19172 8373 19181
rect 8331 19132 8332 19172
rect 8372 19132 8373 19172
rect 8331 19123 8373 19132
rect 7988 18544 8084 18584
rect 7948 18535 7988 18544
rect 7564 17620 7892 17660
rect 6795 17072 6837 17081
rect 6795 17032 6796 17072
rect 6836 17032 6837 17072
rect 6795 17023 6837 17032
rect 6796 16938 6836 17023
rect 6795 16820 6837 16829
rect 6795 16780 6796 16820
rect 6836 16780 6837 16820
rect 6795 16771 6837 16780
rect 6988 16820 7028 16829
rect 6700 15308 6740 15436
rect 6796 15392 6836 16771
rect 6988 16409 7028 16780
rect 6987 16400 7029 16409
rect 6987 16360 6988 16400
rect 7028 16360 7029 16400
rect 6987 16351 7029 16360
rect 6987 16232 7029 16241
rect 7084 16232 7124 16241
rect 6987 16192 6988 16232
rect 7028 16192 7084 16232
rect 6987 16183 7029 16192
rect 7084 16183 7124 16192
rect 7179 16232 7221 16241
rect 7179 16192 7180 16232
rect 7220 16192 7221 16232
rect 7179 16183 7221 16192
rect 7564 16232 7604 17620
rect 8140 17576 8180 17585
rect 7660 17536 8140 17576
rect 7660 17072 7700 17536
rect 8140 17527 8180 17536
rect 7660 17023 7700 17032
rect 7851 17072 7893 17081
rect 7851 17032 7852 17072
rect 7892 17032 7893 17072
rect 7851 17023 7893 17032
rect 7948 17072 7988 17081
rect 7852 16938 7892 17023
rect 7948 16829 7988 17032
rect 8044 17072 8084 17081
rect 7947 16820 7989 16829
rect 7947 16780 7948 16820
rect 7988 16780 7989 16820
rect 7947 16771 7989 16780
rect 8044 16484 8084 17032
rect 8139 17072 8181 17081
rect 8139 17032 8140 17072
rect 8180 17032 8181 17072
rect 8139 17023 8181 17032
rect 8332 17072 8372 19123
rect 10155 18920 10197 18929
rect 10155 18880 10156 18920
rect 10196 18880 10197 18920
rect 10155 18871 10197 18880
rect 8427 18500 8469 18509
rect 8427 18460 8428 18500
rect 8468 18460 8469 18500
rect 8427 18451 8469 18460
rect 8428 17744 8468 18451
rect 9388 18416 9428 18425
rect 8716 17912 8756 17921
rect 8756 17872 8948 17912
rect 8716 17863 8756 17872
rect 8428 17695 8468 17704
rect 8524 17744 8564 17753
rect 8715 17744 8757 17753
rect 8564 17704 8660 17744
rect 8524 17695 8564 17704
rect 8523 17576 8565 17585
rect 8523 17536 8524 17576
rect 8564 17536 8565 17576
rect 8523 17527 8565 17536
rect 8332 17023 8372 17032
rect 8524 17072 8564 17527
rect 8140 16938 8180 17023
rect 8427 16820 8469 16829
rect 8427 16780 8428 16820
rect 8468 16780 8469 16820
rect 8427 16771 8469 16780
rect 8428 16686 8468 16771
rect 8140 16484 8180 16493
rect 8044 16444 8140 16484
rect 8140 16435 8180 16444
rect 8427 16484 8469 16493
rect 8427 16444 8428 16484
rect 8468 16444 8469 16484
rect 8427 16435 8469 16444
rect 8428 16350 8468 16435
rect 7564 16183 7604 16192
rect 7851 16232 7893 16241
rect 7851 16192 7852 16232
rect 7892 16192 7893 16232
rect 7851 16183 7893 16192
rect 7948 16232 7988 16243
rect 8524 16241 8564 17032
rect 7180 16098 7220 16183
rect 7852 15821 7892 16183
rect 7948 16157 7988 16192
rect 8140 16232 8180 16241
rect 7947 16148 7989 16157
rect 7947 16108 7948 16148
rect 7988 16108 7989 16148
rect 7947 16099 7989 16108
rect 7851 15812 7893 15821
rect 7851 15772 7852 15812
rect 7892 15772 7893 15812
rect 7851 15763 7893 15772
rect 7660 15737 7700 15741
rect 7659 15732 7701 15737
rect 7659 15688 7660 15732
rect 7700 15688 7701 15732
rect 7659 15679 7701 15688
rect 7660 15597 7700 15679
rect 8140 15653 8180 16192
rect 8332 16232 8372 16241
rect 8235 15728 8277 15737
rect 8235 15688 8236 15728
rect 8276 15688 8277 15728
rect 8235 15679 8277 15688
rect 7851 15644 7893 15653
rect 7851 15604 7852 15644
rect 7892 15604 7893 15644
rect 7851 15595 7893 15604
rect 8139 15644 8181 15653
rect 8139 15604 8140 15644
rect 8180 15604 8181 15644
rect 8139 15595 8181 15604
rect 7468 15560 7508 15569
rect 6988 15520 7468 15560
rect 6796 15343 6836 15352
rect 6892 15392 6932 15401
rect 6988 15392 7028 15520
rect 7468 15511 7508 15520
rect 7564 15560 7604 15569
rect 6932 15352 7028 15392
rect 6892 15343 6932 15352
rect 6508 15268 6740 15308
rect 7180 15308 7220 15317
rect 6411 15140 6453 15149
rect 6411 15100 6412 15140
rect 6452 15100 6453 15140
rect 6411 15091 6453 15100
rect 5931 14888 5973 14897
rect 5931 14848 5932 14888
rect 5972 14848 5973 14888
rect 5931 14839 5973 14848
rect 6219 14888 6261 14897
rect 6219 14848 6220 14888
rect 6260 14848 6261 14888
rect 6219 14839 6261 14848
rect 6412 14720 6452 14729
rect 6508 14720 6548 15268
rect 6795 15224 6837 15233
rect 6795 15184 6796 15224
rect 6836 15184 6837 15224
rect 6795 15175 6837 15184
rect 6604 14897 6644 14982
rect 6603 14888 6645 14897
rect 6603 14848 6604 14888
rect 6644 14848 6645 14888
rect 6603 14839 6645 14848
rect 6604 14720 6644 14729
rect 6508 14680 6604 14720
rect 6028 14048 6068 14057
rect 6068 14008 6260 14048
rect 6028 13999 6068 14008
rect 5835 13880 5877 13889
rect 5835 13840 5836 13880
rect 5876 13840 5877 13880
rect 5835 13831 5877 13840
rect 6027 13880 6069 13889
rect 6027 13840 6028 13880
rect 6068 13840 6069 13880
rect 6027 13831 6069 13840
rect 5356 12571 5396 12580
rect 5452 13252 5780 13292
rect 5164 12487 5204 12496
rect 5452 12536 5492 13252
rect 5835 13208 5877 13217
rect 5835 13168 5836 13208
rect 5876 13168 5877 13208
rect 5835 13159 5877 13168
rect 5836 13074 5876 13159
rect 5835 12620 5877 12629
rect 5835 12580 5836 12620
rect 5876 12580 5877 12620
rect 5835 12571 5877 12580
rect 5452 12487 5492 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 4491 12452 4533 12461
rect 4491 12412 4492 12452
rect 4532 12412 4533 12452
rect 4491 12403 4533 12412
rect 4684 12368 4724 12487
rect 5740 12402 5780 12487
rect 5836 12486 5876 12571
rect 5931 12536 5973 12545
rect 5931 12496 5932 12536
rect 5972 12496 5973 12536
rect 5931 12487 5973 12496
rect 6028 12536 6068 13831
rect 6028 12487 6068 12496
rect 5932 12402 5972 12487
rect 4684 12319 4724 12328
rect 6220 12368 6260 14008
rect 6412 12629 6452 14680
rect 6604 14671 6644 14680
rect 6700 14720 6740 14729
rect 6796 14720 6836 15175
rect 6891 15140 6933 15149
rect 6891 15100 6892 15140
rect 6932 15100 6933 15140
rect 6891 15091 6933 15100
rect 6740 14680 6836 14720
rect 6892 14720 6932 15091
rect 7083 15056 7125 15065
rect 7083 15016 7084 15056
rect 7124 15016 7125 15056
rect 7083 15007 7125 15016
rect 7084 14972 7124 15007
rect 7084 14921 7124 14932
rect 6700 14671 6740 14680
rect 6892 14671 6932 14680
rect 6892 14048 6932 14057
rect 6892 13469 6932 14008
rect 6507 13460 6549 13469
rect 6507 13420 6508 13460
rect 6548 13420 6549 13460
rect 6507 13411 6549 13420
rect 6891 13460 6933 13469
rect 6891 13420 6892 13460
rect 6932 13420 6933 13460
rect 6891 13411 6933 13420
rect 6508 13326 6548 13411
rect 6795 13208 6837 13217
rect 6795 13168 6796 13208
rect 6836 13168 6837 13208
rect 6795 13159 6837 13168
rect 7180 13208 7220 15268
rect 7564 14225 7604 15520
rect 7852 15560 7892 15595
rect 7852 15509 7892 15520
rect 8140 15560 8180 15595
rect 8236 15594 8276 15679
rect 8332 15569 8372 16192
rect 8523 16232 8565 16241
rect 8523 16192 8524 16232
rect 8564 16192 8565 16232
rect 8523 16183 8565 16192
rect 8620 16064 8660 17704
rect 8715 17704 8716 17744
rect 8756 17704 8757 17744
rect 8715 17695 8757 17704
rect 8908 17744 8948 17872
rect 8908 17695 8948 17704
rect 9292 17744 9332 17753
rect 9388 17744 9428 18376
rect 9332 17704 9428 17744
rect 10156 17744 10196 18871
rect 10444 18845 10484 19216
rect 10443 18836 10485 18845
rect 10443 18796 10444 18836
rect 10484 18796 10485 18836
rect 10443 18787 10485 18796
rect 10540 18752 10580 20551
rect 10636 19517 10676 20728
rect 11499 20768 11541 20777
rect 11499 20728 11500 20768
rect 11540 20728 11541 20768
rect 11499 20719 11541 20728
rect 10827 20684 10869 20693
rect 10827 20644 10828 20684
rect 10868 20644 10869 20684
rect 10827 20635 10869 20644
rect 10828 20550 10868 20635
rect 11500 20634 11540 20719
rect 11788 20273 11828 21400
rect 10827 20264 10869 20273
rect 10827 20224 10828 20264
rect 10868 20224 10869 20264
rect 10827 20215 10869 20224
rect 11787 20264 11829 20273
rect 11787 20224 11788 20264
rect 11828 20224 11829 20264
rect 11787 20215 11829 20224
rect 10828 20096 10868 20215
rect 11307 20180 11349 20189
rect 11307 20140 11308 20180
rect 11348 20140 11349 20180
rect 11307 20131 11349 20140
rect 10828 20047 10868 20056
rect 10635 19508 10677 19517
rect 10635 19468 10636 19508
rect 10676 19468 10677 19508
rect 10635 19459 10677 19468
rect 11308 19349 11348 20131
rect 11692 20096 11732 20105
rect 11884 20096 11924 21559
rect 12076 20768 12116 20777
rect 11732 20056 11924 20096
rect 11980 20684 12020 20693
rect 11692 20047 11732 20056
rect 11980 19424 12020 20644
rect 12076 20105 12116 20728
rect 12364 20768 12404 22651
rect 12748 22532 12788 22651
rect 12748 22483 12788 22492
rect 12940 22373 12980 23500
rect 13612 23381 13652 23668
rect 13804 23624 13844 23633
rect 13708 23584 13804 23624
rect 13611 23372 13653 23381
rect 13611 23332 13612 23372
rect 13652 23332 13653 23372
rect 13611 23323 13653 23332
rect 13612 23204 13652 23213
rect 13708 23204 13748 23584
rect 13804 23575 13844 23584
rect 13803 23372 13845 23381
rect 13803 23332 13804 23372
rect 13844 23332 13845 23372
rect 13803 23323 13845 23332
rect 13652 23164 13748 23204
rect 13612 23155 13652 23164
rect 13515 23120 13557 23129
rect 13515 23080 13516 23120
rect 13556 23080 13557 23120
rect 13515 23071 13557 23080
rect 13420 22868 13460 22877
rect 13036 22828 13420 22868
rect 12939 22364 12981 22373
rect 12939 22324 12940 22364
rect 12980 22324 12981 22364
rect 12939 22315 12981 22324
rect 12940 22280 12980 22315
rect 12940 22230 12980 22240
rect 13036 21692 13076 22828
rect 13420 22819 13460 22828
rect 13419 22448 13461 22457
rect 13419 22408 13420 22448
rect 13460 22408 13461 22448
rect 13419 22399 13461 22408
rect 13227 22364 13269 22373
rect 13227 22324 13228 22364
rect 13268 22324 13269 22364
rect 13227 22315 13269 22324
rect 13036 21643 13076 21652
rect 12939 21440 12981 21449
rect 12939 21400 12940 21440
rect 12980 21400 12981 21440
rect 12939 21391 12981 21400
rect 12940 20777 12980 21391
rect 13228 20852 13268 22315
rect 13420 21608 13460 22399
rect 13516 22280 13556 23071
rect 13611 22700 13653 22709
rect 13611 22660 13612 22700
rect 13652 22660 13653 22700
rect 13611 22651 13653 22660
rect 13516 22231 13556 22240
rect 13612 22280 13652 22651
rect 13612 22231 13652 22240
rect 13708 22280 13748 22289
rect 13708 22121 13748 22240
rect 13804 22280 13844 23323
rect 13804 22231 13844 22240
rect 13707 22112 13749 22121
rect 13707 22072 13708 22112
rect 13748 22072 13749 22112
rect 13707 22063 13749 22072
rect 13420 21559 13460 21568
rect 13900 21449 13940 24088
rect 13996 23717 14036 24592
rect 14091 24592 14092 24632
rect 14132 24592 14133 24632
rect 14091 24583 14133 24592
rect 14188 24632 14228 24919
rect 14380 24884 14420 25432
rect 14763 25423 14805 25432
rect 14475 25304 14517 25313
rect 14475 25264 14476 25304
rect 14516 25264 14517 25304
rect 14475 25255 14517 25264
rect 14668 25304 14708 25313
rect 14476 24968 14516 25255
rect 14572 25145 14612 25227
rect 14571 25136 14613 25145
rect 14571 25092 14572 25136
rect 14612 25092 14613 25136
rect 14571 25087 14613 25092
rect 14572 25083 14612 25087
rect 14476 24928 14612 24968
rect 14380 24844 14516 24884
rect 14380 24725 14420 24748
rect 14379 24716 14421 24725
rect 14379 24676 14380 24716
rect 14420 24676 14421 24716
rect 14379 24667 14421 24676
rect 14380 24653 14420 24667
rect 14092 24498 14132 24583
rect 14188 24305 14228 24592
rect 14284 24632 14324 24641
rect 14380 24604 14420 24613
rect 14187 24296 14229 24305
rect 14187 24256 14188 24296
rect 14228 24256 14229 24296
rect 14187 24247 14229 24256
rect 14187 24128 14229 24137
rect 14187 24088 14188 24128
rect 14228 24088 14229 24128
rect 14187 24079 14229 24088
rect 14091 23876 14133 23885
rect 14091 23836 14092 23876
rect 14132 23836 14133 23876
rect 14091 23827 14133 23836
rect 13995 23708 14037 23717
rect 13995 23668 13996 23708
rect 14036 23668 14037 23708
rect 13995 23659 14037 23668
rect 13995 23120 14037 23129
rect 13995 23080 13996 23120
rect 14036 23080 14037 23120
rect 13995 23071 14037 23080
rect 13996 22986 14036 23071
rect 13995 22448 14037 22457
rect 13995 22408 13996 22448
rect 14036 22408 14037 22448
rect 13995 22399 14037 22408
rect 13996 22314 14036 22399
rect 13899 21440 13941 21449
rect 13899 21400 13900 21440
rect 13940 21400 13941 21440
rect 13899 21391 13941 21400
rect 13228 20803 13268 20812
rect 13995 20852 14037 20861
rect 13995 20812 13996 20852
rect 14036 20812 14037 20852
rect 13995 20803 14037 20812
rect 12364 20719 12404 20728
rect 12939 20768 12981 20777
rect 12939 20728 12940 20768
rect 12980 20728 12981 20768
rect 12939 20719 12981 20728
rect 13996 20768 14036 20803
rect 12075 20096 12117 20105
rect 12075 20056 12076 20096
rect 12116 20056 12117 20096
rect 12075 20047 12117 20056
rect 12940 20096 12980 20719
rect 13996 20717 14036 20728
rect 14092 20180 14132 23827
rect 14188 23633 14228 24079
rect 14284 23969 14324 24592
rect 14476 24548 14516 24844
rect 14380 24508 14516 24548
rect 14283 23960 14325 23969
rect 14283 23920 14284 23960
rect 14324 23920 14325 23960
rect 14283 23911 14325 23920
rect 14187 23624 14229 23633
rect 14187 23584 14188 23624
rect 14228 23584 14229 23624
rect 14187 23575 14229 23584
rect 14283 22280 14325 22289
rect 14283 22240 14284 22280
rect 14324 22240 14325 22280
rect 14283 22231 14325 22240
rect 14284 21617 14324 22231
rect 14283 21608 14325 21617
rect 14283 21568 14284 21608
rect 14324 21568 14325 21608
rect 14283 21559 14325 21568
rect 14284 21474 14324 21559
rect 12940 20047 12980 20056
rect 13996 20140 14132 20180
rect 14380 20180 14420 24508
rect 14475 24380 14517 24389
rect 14475 24340 14476 24380
rect 14516 24340 14517 24380
rect 14475 24331 14517 24340
rect 14476 23792 14516 24331
rect 14476 23743 14516 23752
rect 14572 22280 14612 24928
rect 14668 23969 14708 25264
rect 14764 25304 14804 25423
rect 14764 25255 14804 25264
rect 14859 25304 14901 25313
rect 14859 25264 14860 25304
rect 14900 25264 14901 25304
rect 14859 25255 14901 25264
rect 14860 24884 14900 25255
rect 14956 24968 14996 26104
rect 15052 26095 15092 26104
rect 15244 26144 15284 26179
rect 15051 25976 15093 25985
rect 15051 25936 15052 25976
rect 15092 25936 15093 25976
rect 15051 25927 15093 25936
rect 15052 25556 15092 25927
rect 15052 25507 15092 25516
rect 15244 25313 15284 26104
rect 15436 26144 15476 27700
rect 16012 27665 16052 27750
rect 16011 27656 16053 27665
rect 16011 27616 16012 27656
rect 16052 27616 16053 27656
rect 16011 27607 16053 27616
rect 16011 27404 16053 27413
rect 16011 27364 16012 27404
rect 16052 27364 16053 27404
rect 16011 27355 16053 27364
rect 16012 27270 16052 27355
rect 16108 26564 16148 28960
rect 16300 28496 16340 29119
rect 16300 28447 16340 28456
rect 16588 29000 16628 29009
rect 17164 29000 17204 33412
rect 17356 33403 17396 33412
rect 17259 32948 17301 32957
rect 17259 32908 17260 32948
rect 17300 32908 17301 32948
rect 17259 32899 17301 32908
rect 17260 32814 17300 32899
rect 17644 32873 17684 32882
rect 17684 32833 17876 32864
rect 17644 32824 17876 32833
rect 17452 32780 17492 32789
rect 17492 32740 17780 32780
rect 17452 32731 17492 32740
rect 17644 32192 17684 32201
rect 17644 31697 17684 32152
rect 17643 31688 17685 31697
rect 17643 31648 17644 31688
rect 17684 31648 17685 31688
rect 17643 31639 17685 31648
rect 17740 31520 17780 32740
rect 17644 31480 17780 31520
rect 17356 31352 17396 31361
rect 17396 31312 17492 31352
rect 17356 31303 17396 31312
rect 17452 30512 17492 31312
rect 17452 30463 17492 30472
rect 17355 29924 17397 29933
rect 17355 29884 17356 29924
rect 17396 29884 17397 29924
rect 17355 29875 17397 29884
rect 17356 29790 17396 29875
rect 16588 28253 16628 28960
rect 16972 28960 17204 29000
rect 16587 28244 16629 28253
rect 16587 28204 16588 28244
rect 16628 28204 16629 28244
rect 16587 28195 16629 28204
rect 16204 27656 16244 27665
rect 16204 27245 16244 27616
rect 16299 27656 16341 27665
rect 16299 27616 16300 27656
rect 16340 27616 16341 27656
rect 16299 27607 16341 27616
rect 16300 27522 16340 27607
rect 16491 27572 16533 27581
rect 16491 27532 16492 27572
rect 16532 27532 16533 27572
rect 16491 27523 16533 27532
rect 16203 27236 16245 27245
rect 16203 27196 16204 27236
rect 16244 27196 16245 27236
rect 16203 27187 16245 27196
rect 16492 26741 16532 27523
rect 16779 27236 16821 27245
rect 16779 27196 16780 27236
rect 16820 27196 16821 27236
rect 16779 27187 16821 27196
rect 16780 26816 16820 27187
rect 16780 26767 16820 26776
rect 16972 26816 17012 28960
rect 17068 28244 17108 28253
rect 17068 27245 17108 28204
rect 17547 28244 17589 28253
rect 17547 28204 17548 28244
rect 17588 28204 17589 28244
rect 17547 28195 17589 28204
rect 17452 27656 17492 27665
rect 17452 27497 17492 27616
rect 17451 27488 17493 27497
rect 17451 27448 17452 27488
rect 17492 27448 17493 27488
rect 17451 27439 17493 27448
rect 17067 27236 17109 27245
rect 17067 27196 17068 27236
rect 17108 27196 17109 27236
rect 17067 27187 17109 27196
rect 17355 27236 17397 27245
rect 17355 27196 17356 27236
rect 17396 27196 17397 27236
rect 17355 27187 17397 27196
rect 17164 26816 17204 26825
rect 16972 26767 17012 26776
rect 17068 26776 17164 26816
rect 16491 26732 16533 26741
rect 16491 26692 16492 26732
rect 16532 26692 16533 26732
rect 16491 26683 16533 26692
rect 16876 26732 16916 26741
rect 15820 26524 16148 26564
rect 15627 26312 15669 26321
rect 15627 26272 15628 26312
rect 15668 26272 15669 26312
rect 15627 26263 15669 26272
rect 15436 26095 15476 26104
rect 15628 26144 15668 26263
rect 15436 25892 15476 25901
rect 15436 25565 15476 25852
rect 15435 25556 15477 25565
rect 15435 25516 15436 25556
rect 15476 25516 15477 25556
rect 15435 25507 15477 25516
rect 15243 25304 15285 25313
rect 15243 25264 15244 25304
rect 15284 25264 15285 25304
rect 15243 25255 15285 25264
rect 15243 25136 15285 25145
rect 15243 25096 15244 25136
rect 15284 25096 15285 25136
rect 15243 25087 15285 25096
rect 14956 24928 15092 24968
rect 14860 24844 14996 24884
rect 14859 24716 14901 24725
rect 14859 24676 14860 24716
rect 14900 24676 14901 24716
rect 14859 24667 14901 24676
rect 14764 24632 14804 24641
rect 14667 23960 14709 23969
rect 14667 23920 14668 23960
rect 14708 23920 14709 23960
rect 14667 23911 14709 23920
rect 14764 23885 14804 24592
rect 14860 24632 14900 24667
rect 14860 24581 14900 24592
rect 14956 24632 14996 24844
rect 15052 24800 15092 24928
rect 15052 24760 15188 24800
rect 14956 24583 14996 24592
rect 15051 24632 15093 24641
rect 15051 24592 15052 24632
rect 15092 24592 15093 24632
rect 15051 24583 15093 24592
rect 15052 24498 15092 24583
rect 15148 24380 15188 24760
rect 15244 24725 15284 25087
rect 15628 24800 15668 26104
rect 15820 25304 15860 26524
rect 16011 26396 16053 26405
rect 16011 26356 16012 26396
rect 16052 26356 16053 26396
rect 16011 26347 16053 26356
rect 15915 26312 15957 26321
rect 15915 26272 15916 26312
rect 15956 26272 15957 26312
rect 15915 26263 15957 26272
rect 15916 26144 15956 26263
rect 15916 26095 15956 26104
rect 16012 26144 16052 26347
rect 16012 26095 16052 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16107 26095 16149 26104
rect 16204 26144 16244 26153
rect 16396 26144 16436 26153
rect 16244 26104 16396 26144
rect 16204 26095 16244 26104
rect 16396 26095 16436 26104
rect 16108 25976 16148 26095
rect 16108 25936 16340 25976
rect 16107 25304 16149 25313
rect 15820 25264 16108 25304
rect 16148 25264 16149 25304
rect 16107 25255 16149 25264
rect 16108 25170 16148 25255
rect 16203 24884 16245 24893
rect 16203 24844 16204 24884
rect 16244 24844 16245 24884
rect 16203 24835 16245 24844
rect 16204 24800 16244 24835
rect 15628 24760 15956 24800
rect 15243 24716 15285 24725
rect 15243 24676 15244 24716
rect 15284 24676 15285 24716
rect 15243 24667 15285 24676
rect 14956 24340 15188 24380
rect 15244 24632 15284 24667
rect 15532 24632 15572 24641
rect 14763 23876 14805 23885
rect 14763 23836 14764 23876
rect 14804 23836 14805 23876
rect 14763 23827 14805 23836
rect 14668 23792 14708 23801
rect 14668 23633 14708 23752
rect 14860 23792 14900 23801
rect 14764 23708 14804 23717
rect 14667 23624 14709 23633
rect 14667 23584 14668 23624
rect 14708 23584 14709 23624
rect 14667 23575 14709 23584
rect 14764 23549 14804 23668
rect 14763 23540 14805 23549
rect 14763 23500 14764 23540
rect 14804 23500 14805 23540
rect 14763 23491 14805 23500
rect 14860 23297 14900 23752
rect 14956 23465 14996 24340
rect 15051 24212 15093 24221
rect 15051 24172 15052 24212
rect 15092 24172 15093 24212
rect 15051 24163 15093 24172
rect 15052 23876 15092 24163
rect 15244 24137 15284 24592
rect 15436 24592 15532 24632
rect 15243 24128 15285 24137
rect 15243 24088 15244 24128
rect 15284 24088 15285 24128
rect 15243 24079 15285 24088
rect 15339 24044 15381 24053
rect 15339 24004 15340 24044
rect 15380 24004 15381 24044
rect 15339 23995 15381 24004
rect 15147 23876 15189 23885
rect 15052 23836 15148 23876
rect 15188 23836 15189 23876
rect 15147 23827 15189 23836
rect 15148 23792 15188 23827
rect 15148 23742 15188 23752
rect 15244 23792 15284 23801
rect 15051 23708 15093 23717
rect 15051 23668 15052 23708
rect 15092 23668 15093 23708
rect 15051 23659 15093 23668
rect 15052 23574 15092 23659
rect 15244 23633 15284 23752
rect 15340 23792 15380 23995
rect 15340 23743 15380 23752
rect 15243 23624 15285 23633
rect 15243 23584 15244 23624
rect 15284 23584 15285 23624
rect 15243 23575 15285 23584
rect 14955 23456 14997 23465
rect 14955 23416 14956 23456
rect 14996 23416 14997 23456
rect 14955 23407 14997 23416
rect 15339 23456 15381 23465
rect 15339 23416 15340 23456
rect 15380 23416 15381 23456
rect 15339 23407 15381 23416
rect 14859 23288 14901 23297
rect 14859 23248 14860 23288
rect 14900 23248 14901 23288
rect 14859 23239 14901 23248
rect 15340 23213 15380 23407
rect 15339 23204 15381 23213
rect 15339 23164 15340 23204
rect 15380 23164 15381 23204
rect 15339 23155 15381 23164
rect 14860 23120 14900 23129
rect 14860 22532 14900 23080
rect 14860 22483 14900 22492
rect 15147 22448 15189 22457
rect 15147 22408 15148 22448
rect 15188 22408 15189 22448
rect 15147 22399 15189 22408
rect 14572 22231 14612 22240
rect 15148 21020 15188 22399
rect 15340 21608 15380 23155
rect 15436 22457 15476 24592
rect 15532 24583 15572 24592
rect 15724 24632 15764 24641
rect 15532 24464 15572 24473
rect 15724 24464 15764 24592
rect 15819 24632 15861 24641
rect 15819 24592 15820 24632
rect 15860 24592 15861 24632
rect 15819 24583 15861 24592
rect 15916 24632 15956 24760
rect 16204 24749 16244 24760
rect 15916 24583 15956 24592
rect 16011 24632 16053 24641
rect 16011 24592 16012 24632
rect 16052 24592 16053 24632
rect 16011 24583 16053 24592
rect 16300 24632 16340 25936
rect 16396 25892 16436 25901
rect 16396 24809 16436 25852
rect 16492 25397 16532 26683
rect 16876 26489 16916 26692
rect 16875 26480 16917 26489
rect 16875 26440 16876 26480
rect 16916 26440 16917 26480
rect 16875 26431 16917 26440
rect 16588 26144 16628 26153
rect 16588 25985 16628 26104
rect 16684 26144 16724 26153
rect 16587 25976 16629 25985
rect 16587 25936 16588 25976
rect 16628 25936 16629 25976
rect 16587 25927 16629 25936
rect 16684 25733 16724 26104
rect 16876 25976 16916 25985
rect 17068 25976 17108 26776
rect 17164 26767 17204 26776
rect 17356 26816 17396 27187
rect 17548 26984 17588 28195
rect 17260 26732 17300 26741
rect 17163 26480 17205 26489
rect 17163 26440 17164 26480
rect 17204 26440 17205 26480
rect 17163 26431 17205 26440
rect 17164 26228 17204 26431
rect 17260 26321 17300 26692
rect 17259 26312 17301 26321
rect 17259 26272 17260 26312
rect 17300 26272 17301 26312
rect 17259 26263 17301 26272
rect 17356 26228 17396 26776
rect 17164 26179 17204 26188
rect 17355 26188 17396 26228
rect 17452 26944 17588 26984
rect 17260 26144 17300 26155
rect 17260 26069 17300 26104
rect 17259 26060 17301 26069
rect 17259 26020 17260 26060
rect 17300 26020 17301 26060
rect 17355 26060 17395 26188
rect 17452 26069 17492 26944
rect 17548 26816 17588 26825
rect 17548 26405 17588 26776
rect 17644 26816 17684 31480
rect 17739 31352 17781 31361
rect 17739 31312 17740 31352
rect 17780 31312 17781 31352
rect 17739 31303 17781 31312
rect 17740 29168 17780 31303
rect 17836 30605 17876 32824
rect 17932 32192 17972 33739
rect 18027 33704 18069 33713
rect 18027 33664 18028 33704
rect 18068 33664 18069 33704
rect 18027 33655 18069 33664
rect 18028 33570 18068 33655
rect 18508 33536 18548 34579
rect 18700 34292 18740 34924
rect 18988 34628 19028 35839
rect 19180 35216 19220 35225
rect 19372 35216 19412 36016
rect 19756 36007 19796 36016
rect 23788 36016 23884 36056
rect 19563 35888 19605 35897
rect 19563 35848 19564 35888
rect 19604 35848 19605 35888
rect 19563 35839 19605 35848
rect 21772 35888 21812 35897
rect 19564 35754 19604 35839
rect 21100 35720 21140 35729
rect 20908 35680 21100 35720
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 19220 35176 19412 35216
rect 20044 35216 20084 35225
rect 19180 35167 19220 35176
rect 19275 34880 19317 34889
rect 19275 34840 19276 34880
rect 19316 34840 19317 34880
rect 19275 34831 19317 34840
rect 18604 34252 18740 34292
rect 18796 34588 19028 34628
rect 18604 33704 18644 34252
rect 18796 33872 18836 34588
rect 18987 34376 19029 34385
rect 18987 34327 18988 34376
rect 19028 34327 19029 34376
rect 19276 34376 19316 34831
rect 19371 34544 19413 34553
rect 19371 34504 19372 34544
rect 19412 34504 19413 34544
rect 19371 34495 19413 34504
rect 19372 34418 19412 34495
rect 20044 34385 20084 35176
rect 19372 34369 19412 34378
rect 19468 34376 19508 34385
rect 19276 34327 19316 34336
rect 18891 34208 18933 34217
rect 18891 34168 18892 34208
rect 18932 34168 18933 34208
rect 18891 34159 18933 34168
rect 18796 33823 18836 33832
rect 18699 33788 18741 33797
rect 18699 33748 18700 33788
rect 18740 33748 18741 33788
rect 18699 33739 18741 33748
rect 18604 33655 18644 33664
rect 18700 33704 18740 33739
rect 18700 33653 18740 33664
rect 18892 33704 18932 34159
rect 18988 33788 19028 34311
rect 19179 34208 19221 34217
rect 19468 34208 19508 34336
rect 20043 34376 20085 34385
rect 20043 34336 20044 34376
rect 20084 34336 20085 34376
rect 20043 34327 20085 34336
rect 19179 34168 19180 34208
rect 19220 34168 19221 34208
rect 19179 34159 19221 34168
rect 19372 34168 19508 34208
rect 19180 34074 19220 34159
rect 19372 33797 19412 34168
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 19371 33788 19413 33797
rect 18988 33748 19124 33788
rect 18892 33655 18932 33664
rect 18891 33536 18933 33545
rect 18508 33496 18740 33536
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 18123 33032 18165 33041
rect 18123 32992 18124 33032
rect 18164 32992 18165 33032
rect 18123 32983 18165 32992
rect 18124 32864 18164 32983
rect 18603 32948 18645 32957
rect 18603 32908 18604 32948
rect 18644 32908 18645 32948
rect 18603 32899 18645 32908
rect 18700 32948 18740 33496
rect 18891 33496 18892 33536
rect 18932 33496 18933 33536
rect 18891 33487 18933 33496
rect 18700 32899 18740 32908
rect 18124 32815 18164 32824
rect 18219 32864 18261 32873
rect 18219 32824 18220 32864
rect 18260 32824 18261 32864
rect 18219 32815 18261 32824
rect 18123 32360 18165 32369
rect 18123 32320 18124 32360
rect 18164 32320 18165 32360
rect 18123 32311 18165 32320
rect 18220 32360 18260 32815
rect 18604 32814 18644 32899
rect 18892 32696 18932 33487
rect 19084 32864 19124 33748
rect 19371 33748 19372 33788
rect 19412 33748 19413 33788
rect 19371 33739 19413 33748
rect 19659 33788 19701 33797
rect 19659 33748 19660 33788
rect 19700 33748 19701 33788
rect 19659 33739 19701 33748
rect 19179 33704 19221 33713
rect 19179 33664 19180 33704
rect 19220 33664 19221 33704
rect 19179 33655 19221 33664
rect 19276 33704 19316 33713
rect 19180 33209 19220 33655
rect 19179 33200 19221 33209
rect 19179 33160 19180 33200
rect 19220 33160 19221 33200
rect 19179 33151 19221 33160
rect 19084 32815 19124 32824
rect 19180 32864 19220 33151
rect 19180 32815 19220 32824
rect 18892 32656 19124 32696
rect 18220 32311 18260 32320
rect 19084 32360 19124 32656
rect 19276 32360 19316 33664
rect 19468 33452 19508 33463
rect 19468 33377 19508 33412
rect 19467 33368 19509 33377
rect 19467 33328 19468 33368
rect 19508 33328 19509 33368
rect 19467 33319 19509 33328
rect 19660 33125 19700 33739
rect 20331 33704 20373 33713
rect 20331 33664 20332 33704
rect 20372 33664 20373 33704
rect 20331 33655 20373 33664
rect 20908 33704 20948 35680
rect 21100 35671 21140 35680
rect 21772 35393 21812 35848
rect 21771 35384 21813 35393
rect 21771 35344 21772 35384
rect 21812 35344 21813 35384
rect 21771 35335 21813 35344
rect 21195 35300 21237 35309
rect 21195 35260 21196 35300
rect 21236 35260 21237 35300
rect 21195 35251 21237 35260
rect 23403 35300 23445 35309
rect 23403 35260 23404 35300
rect 23444 35260 23445 35300
rect 23403 35251 23445 35260
rect 21196 34964 21236 35251
rect 22252 35216 22292 35225
rect 21676 35176 22252 35216
rect 21580 34964 21620 34973
rect 21196 34553 21236 34924
rect 21388 34924 21580 34964
rect 21195 34544 21237 34553
rect 21195 34504 21196 34544
rect 21236 34504 21237 34544
rect 21195 34495 21237 34504
rect 21003 34376 21045 34385
rect 21003 34336 21004 34376
rect 21044 34336 21045 34376
rect 21003 34327 21045 34336
rect 21388 34376 21428 34924
rect 21580 34915 21620 34924
rect 21388 34327 21428 34336
rect 20908 33655 20948 33664
rect 20043 33620 20085 33629
rect 20043 33580 20044 33620
rect 20084 33580 20085 33620
rect 20043 33571 20085 33580
rect 19659 33116 19701 33125
rect 19659 33076 19660 33116
rect 19700 33076 19701 33116
rect 19659 33067 19701 33076
rect 19371 33032 19413 33041
rect 19371 32992 19372 33032
rect 19412 32992 19413 33032
rect 19371 32983 19413 32992
rect 19372 32789 19412 32983
rect 19467 32864 19509 32873
rect 19467 32824 19468 32864
rect 19508 32824 19509 32864
rect 19467 32815 19509 32824
rect 19660 32864 19700 33067
rect 19660 32815 19700 32824
rect 19755 32864 19797 32873
rect 19755 32824 19756 32864
rect 19796 32824 19797 32864
rect 19755 32815 19797 32824
rect 20044 32864 20084 33571
rect 20332 33570 20372 33655
rect 20811 33620 20853 33629
rect 20811 33580 20812 33620
rect 20852 33580 20853 33620
rect 20811 33571 20853 33580
rect 20812 33486 20852 33571
rect 20428 33452 20468 33461
rect 20331 33116 20373 33125
rect 20331 33076 20332 33116
rect 20372 33076 20373 33116
rect 20331 33067 20373 33076
rect 20332 32982 20372 33067
rect 20428 32873 20468 33412
rect 20044 32815 20084 32824
rect 20427 32864 20469 32873
rect 20427 32824 20428 32864
rect 20468 32824 20469 32864
rect 20427 32815 20469 32824
rect 19371 32780 19413 32789
rect 19371 32740 19372 32780
rect 19412 32740 19413 32780
rect 19371 32731 19413 32740
rect 19084 32311 19124 32320
rect 19180 32320 19316 32360
rect 17932 32033 17972 32152
rect 18027 32192 18069 32201
rect 18027 32152 18028 32192
rect 18068 32152 18069 32192
rect 18027 32143 18069 32152
rect 18124 32192 18164 32311
rect 18124 32143 18164 32152
rect 18412 32192 18452 32203
rect 18028 32058 18068 32143
rect 18412 32117 18452 32152
rect 18411 32108 18453 32117
rect 18411 32068 18412 32108
rect 18452 32068 18453 32108
rect 18411 32059 18453 32068
rect 17931 32024 17973 32033
rect 17931 31984 17932 32024
rect 17972 31984 17973 32024
rect 17931 31975 17973 31984
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 18219 31352 18261 31361
rect 18219 31312 18220 31352
rect 18260 31312 18261 31352
rect 18219 31303 18261 31312
rect 18220 31218 18260 31303
rect 17835 30596 17877 30605
rect 17835 30556 17836 30596
rect 17876 30556 17877 30596
rect 17835 30547 17877 30556
rect 18988 30428 19028 30437
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 18699 30176 18741 30185
rect 18699 30136 18700 30176
rect 18740 30136 18741 30176
rect 18699 30127 18741 30136
rect 18603 30008 18645 30017
rect 18603 29968 18604 30008
rect 18644 29968 18645 30008
rect 18603 29959 18645 29968
rect 18604 29840 18644 29959
rect 18604 29791 18644 29800
rect 18700 29840 18740 30127
rect 18988 29933 19028 30388
rect 18795 29924 18837 29933
rect 18795 29884 18796 29924
rect 18836 29884 18837 29924
rect 18795 29875 18837 29884
rect 18987 29924 19029 29933
rect 18987 29884 18988 29924
rect 19028 29884 19029 29924
rect 18987 29875 19029 29884
rect 18700 29261 18740 29800
rect 18796 29840 18836 29875
rect 18699 29252 18741 29261
rect 18699 29212 18700 29252
rect 18740 29212 18741 29252
rect 18699 29203 18741 29212
rect 17740 29119 17780 29128
rect 18603 29168 18645 29177
rect 18603 29128 18604 29168
rect 18644 29128 18645 29168
rect 18603 29119 18645 29128
rect 18604 29034 18644 29119
rect 18796 29000 18836 29800
rect 18891 29840 18933 29849
rect 18891 29800 18892 29840
rect 18932 29800 18933 29840
rect 18891 29791 18933 29800
rect 19180 29840 19220 32320
rect 19276 32192 19316 32201
rect 19372 32192 19412 32731
rect 19468 32730 19508 32815
rect 19564 32705 19604 32790
rect 19756 32730 19796 32815
rect 20139 32780 20181 32789
rect 20139 32740 20140 32780
rect 20180 32740 20181 32780
rect 20139 32731 20181 32740
rect 20908 32780 20948 32789
rect 19563 32696 19605 32705
rect 19563 32656 19564 32696
rect 19604 32656 19605 32696
rect 19563 32647 19605 32656
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 20043 32360 20085 32369
rect 20043 32320 20044 32360
rect 20084 32320 20085 32360
rect 20043 32311 20085 32320
rect 20140 32360 20180 32731
rect 20140 32311 20180 32320
rect 19316 32152 19412 32192
rect 19947 32192 19989 32201
rect 19947 32152 19948 32192
rect 19988 32152 19989 32192
rect 19276 32143 19316 32152
rect 19947 32143 19989 32152
rect 19948 32058 19988 32143
rect 19371 32024 19413 32033
rect 19371 31984 19372 32024
rect 19412 31984 19413 32024
rect 19371 31975 19413 31984
rect 19372 31520 19412 31975
rect 19372 31471 19412 31480
rect 19755 31520 19797 31529
rect 19755 31480 19756 31520
rect 19796 31480 19797 31520
rect 19755 31471 19797 31480
rect 19756 31386 19796 31471
rect 19948 31184 19988 31193
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 19659 30680 19701 30689
rect 19659 30640 19660 30680
rect 19700 30640 19701 30680
rect 19659 30631 19701 30640
rect 19948 30680 19988 31144
rect 20044 30689 20084 32311
rect 20331 31520 20373 31529
rect 20812 31520 20852 31529
rect 20331 31480 20332 31520
rect 20372 31480 20373 31520
rect 20331 31471 20373 31480
rect 20620 31480 20812 31520
rect 19948 30631 19988 30640
rect 20043 30680 20085 30689
rect 20043 30640 20044 30680
rect 20084 30640 20085 30680
rect 20043 30631 20085 30640
rect 20332 30680 20372 31471
rect 20620 31352 20660 31480
rect 20812 31471 20852 31480
rect 20620 31303 20660 31312
rect 20812 31352 20852 31361
rect 20908 31352 20948 32740
rect 21004 32192 21044 34327
rect 21291 34208 21333 34217
rect 21291 34168 21292 34208
rect 21332 34168 21333 34208
rect 21291 34159 21333 34168
rect 21099 33704 21141 33713
rect 21099 33664 21100 33704
rect 21140 33664 21141 33704
rect 21099 33655 21141 33664
rect 21196 33704 21236 33713
rect 21100 33570 21140 33655
rect 21196 32369 21236 33664
rect 21292 33704 21332 34159
rect 21676 33872 21716 35176
rect 22252 35167 22292 35176
rect 23404 35166 23444 35251
rect 23788 35216 23828 36016
rect 23884 36007 23924 36016
rect 24460 35888 24500 36511
rect 24460 35839 24500 35848
rect 24844 35888 24884 35897
rect 24940 35888 24980 36520
rect 24884 35848 24980 35888
rect 24844 35839 24884 35848
rect 25612 35561 25652 36688
rect 25708 36728 25748 36856
rect 25708 36679 25748 36688
rect 25900 36728 25940 36737
rect 26092 36728 26132 36737
rect 25940 36688 26092 36728
rect 25900 36679 25940 36688
rect 26092 36679 26132 36688
rect 26188 36728 26228 36737
rect 25899 36560 25941 36569
rect 25899 36520 25900 36560
rect 25940 36520 25941 36560
rect 25899 36511 25941 36520
rect 25900 36426 25940 36511
rect 25995 36476 26037 36485
rect 25995 36436 25996 36476
rect 26036 36436 26037 36476
rect 25995 36427 26037 36436
rect 25708 35888 25748 35897
rect 25748 35848 25940 35888
rect 25708 35839 25748 35848
rect 24075 35552 24117 35561
rect 24075 35512 24076 35552
rect 24116 35512 24117 35552
rect 24075 35503 24117 35512
rect 25611 35552 25653 35561
rect 25611 35512 25612 35552
rect 25652 35512 25653 35552
rect 25611 35503 25653 35512
rect 23788 35167 23828 35176
rect 22444 35048 22484 35057
rect 21772 34376 21812 34385
rect 22444 34376 22484 35008
rect 24076 34628 24116 35503
rect 25803 35468 25845 35477
rect 25803 35428 25804 35468
rect 25844 35428 25845 35468
rect 25803 35419 25845 35428
rect 25611 35384 25653 35393
rect 25611 35344 25612 35384
rect 25652 35344 25653 35384
rect 25611 35335 25653 35344
rect 24652 35216 24692 35225
rect 24076 34579 24116 34588
rect 24556 35176 24652 35216
rect 24556 34385 24596 35176
rect 24652 35167 24692 35176
rect 25419 34460 25461 34469
rect 25419 34420 25420 34460
rect 25460 34420 25461 34460
rect 25419 34411 25461 34420
rect 21812 34336 22484 34376
rect 22635 34376 22677 34385
rect 22635 34336 22636 34376
rect 22676 34336 22677 34376
rect 21772 34327 21812 34336
rect 22635 34327 22677 34336
rect 24172 34376 24212 34385
rect 24364 34376 24404 34385
rect 24212 34336 24364 34376
rect 24172 34327 24212 34336
rect 24364 34327 24404 34336
rect 24555 34376 24597 34385
rect 24555 34336 24556 34376
rect 24596 34336 24597 34376
rect 24555 34327 24597 34336
rect 25036 34376 25076 34385
rect 22636 34242 22676 34327
rect 23787 34208 23829 34217
rect 23787 34168 23788 34208
rect 23828 34168 23829 34208
rect 23787 34159 23829 34168
rect 23788 34074 23828 34159
rect 21772 33872 21812 33881
rect 21676 33832 21772 33872
rect 21772 33823 21812 33832
rect 21292 33655 21332 33664
rect 21388 33704 21428 33713
rect 21580 33704 21620 33715
rect 21428 33664 21524 33704
rect 21388 33655 21428 33664
rect 21484 33461 21524 33664
rect 21580 33629 21620 33664
rect 21676 33704 21716 33713
rect 21579 33620 21621 33629
rect 21579 33580 21580 33620
rect 21620 33580 21621 33620
rect 21579 33571 21621 33580
rect 21676 33461 21716 33664
rect 21867 33704 21909 33713
rect 21867 33664 21868 33704
rect 21908 33664 21909 33704
rect 21867 33655 21909 33664
rect 23595 33704 23637 33713
rect 23595 33664 23596 33704
rect 23636 33664 23637 33704
rect 23595 33655 23637 33664
rect 24171 33704 24213 33713
rect 24171 33664 24172 33704
rect 24212 33664 24213 33704
rect 24171 33655 24213 33664
rect 21868 33570 21908 33655
rect 21483 33452 21525 33461
rect 21483 33412 21484 33452
rect 21524 33412 21525 33452
rect 21483 33403 21525 33412
rect 21675 33452 21717 33461
rect 23500 33452 23540 33461
rect 21675 33412 21676 33452
rect 21716 33412 21717 33452
rect 21675 33403 21717 33412
rect 23308 33412 23500 33452
rect 23211 33200 23253 33209
rect 23211 33160 23212 33200
rect 23252 33160 23253 33200
rect 23211 33151 23253 33160
rect 21387 33032 21429 33041
rect 21387 32992 21388 33032
rect 21428 32992 21429 33032
rect 21387 32983 21429 32992
rect 22155 33032 22197 33041
rect 22155 32992 22156 33032
rect 22196 32992 22197 33032
rect 22155 32983 22197 32992
rect 21388 32898 21428 32983
rect 21195 32360 21237 32369
rect 21195 32320 21196 32360
rect 21236 32320 21237 32360
rect 21195 32311 21237 32320
rect 21292 32192 21332 32201
rect 21004 32152 21292 32192
rect 21292 32143 21332 32152
rect 22156 32192 22196 32983
rect 22539 32696 22581 32705
rect 22539 32656 22540 32696
rect 22580 32656 22581 32696
rect 22539 32647 22581 32656
rect 22540 32276 22580 32647
rect 22540 32227 22580 32236
rect 22156 32143 22196 32152
rect 21291 32024 21333 32033
rect 21291 31984 21292 32024
rect 21332 31984 21333 32024
rect 21291 31975 21333 31984
rect 21004 31352 21044 31361
rect 20908 31312 21004 31352
rect 20332 30631 20372 30640
rect 19660 30546 19700 30631
rect 19467 30008 19509 30017
rect 19467 29968 19468 30008
rect 19508 29968 19509 30008
rect 19467 29959 19509 29968
rect 19468 29874 19508 29959
rect 19220 29800 19316 29840
rect 19180 29791 19220 29800
rect 18892 29706 18932 29791
rect 18988 29168 19028 29177
rect 19180 29168 19220 29177
rect 19028 29128 19180 29168
rect 18988 29119 19028 29128
rect 19180 29119 19220 29128
rect 19276 29000 19316 29800
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 20044 29336 20084 30631
rect 20812 29849 20852 31312
rect 21004 31303 21044 31312
rect 21100 31352 21140 31361
rect 21100 31184 21140 31312
rect 21292 31352 21332 31975
rect 21292 31303 21332 31312
rect 23020 31520 23060 31529
rect 21388 31184 21428 31193
rect 21100 31144 21388 31184
rect 21388 31135 21428 31144
rect 21196 30680 21236 30689
rect 21196 30269 21236 30640
rect 22636 30680 22676 30689
rect 22348 30428 22388 30437
rect 21195 30260 21237 30269
rect 21195 30220 21196 30260
rect 21236 30220 21237 30260
rect 21195 30211 21237 30220
rect 21675 30260 21717 30269
rect 21675 30220 21676 30260
rect 21716 30220 21717 30260
rect 21675 30211 21717 30220
rect 20140 29840 20180 29849
rect 20428 29840 20468 29849
rect 20180 29800 20276 29840
rect 20140 29791 20180 29800
rect 19756 29296 20084 29336
rect 19659 29084 19701 29093
rect 19659 29044 19660 29084
rect 19700 29044 19701 29084
rect 19659 29035 19701 29044
rect 18796 28960 18932 29000
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 17931 28412 17973 28421
rect 17931 28372 17932 28412
rect 17972 28372 17973 28412
rect 17931 28363 17973 28372
rect 17932 28328 17972 28363
rect 17932 28277 17972 28288
rect 18411 28328 18453 28337
rect 18411 28288 18412 28328
rect 18452 28288 18453 28328
rect 18411 28279 18453 28288
rect 18700 28328 18740 28337
rect 18412 27656 18452 28279
rect 18700 28169 18740 28288
rect 18796 28328 18836 28339
rect 18796 28253 18836 28288
rect 18892 28328 18932 28960
rect 19084 28960 19316 29000
rect 18987 28916 19029 28925
rect 18987 28876 18988 28916
rect 19028 28876 19029 28916
rect 18987 28867 19029 28876
rect 18892 28279 18932 28288
rect 18988 28328 19028 28867
rect 18988 28279 19028 28288
rect 18795 28244 18837 28253
rect 18795 28204 18796 28244
rect 18836 28204 18837 28244
rect 18795 28195 18837 28204
rect 18699 28160 18741 28169
rect 18699 28120 18700 28160
rect 18740 28120 18741 28160
rect 18699 28111 18741 28120
rect 19084 28076 19124 28960
rect 19275 28496 19317 28505
rect 19660 28496 19700 29035
rect 19756 28757 19796 29296
rect 20236 29177 20276 29800
rect 19852 29168 19892 29177
rect 19852 29000 19892 29128
rect 20044 29168 20084 29177
rect 20235 29168 20277 29177
rect 20084 29128 20180 29168
rect 20044 29119 20084 29128
rect 20044 29000 20084 29009
rect 19852 28960 20044 29000
rect 20044 28951 20084 28960
rect 20140 28925 20180 29128
rect 20235 29128 20236 29168
rect 20276 29128 20277 29168
rect 20235 29119 20277 29128
rect 20332 29168 20372 29177
rect 20236 29034 20276 29119
rect 20139 28916 20181 28925
rect 20139 28876 20140 28916
rect 20180 28876 20181 28916
rect 20139 28867 20181 28876
rect 20235 28832 20277 28841
rect 20235 28792 20236 28832
rect 20276 28792 20277 28832
rect 20235 28783 20277 28792
rect 19755 28748 19797 28757
rect 19755 28708 19756 28748
rect 19796 28708 19797 28748
rect 19755 28699 19797 28708
rect 19275 28456 19276 28496
rect 19316 28456 19317 28496
rect 19275 28447 19317 28456
rect 19372 28456 19700 28496
rect 19276 28362 19316 28447
rect 19372 28328 19412 28456
rect 19564 28328 19604 28337
rect 19372 28279 19412 28288
rect 19468 28288 19564 28328
rect 19275 28160 19317 28169
rect 19468 28160 19508 28288
rect 19564 28279 19604 28288
rect 19660 28328 19700 28456
rect 19756 28337 19796 28699
rect 20236 28664 20276 28783
rect 20332 28673 20372 29128
rect 20428 28841 20468 29800
rect 20811 29840 20853 29849
rect 20811 29800 20812 29840
rect 20852 29800 20853 29840
rect 20811 29791 20853 29800
rect 21100 29672 21140 29681
rect 20523 29336 20565 29345
rect 20523 29296 20524 29336
rect 20564 29296 20565 29336
rect 20523 29287 20565 29296
rect 20524 29202 20564 29287
rect 21100 29261 21140 29632
rect 21292 29672 21332 29681
rect 21099 29252 21141 29261
rect 21099 29212 21100 29252
rect 21140 29212 21141 29252
rect 21099 29203 21141 29212
rect 21292 29093 21332 29632
rect 21676 29168 21716 30211
rect 22348 30185 22388 30388
rect 22636 30353 22676 30640
rect 23020 30680 23060 31480
rect 23020 30631 23060 30640
rect 22635 30344 22677 30353
rect 22635 30304 22636 30344
rect 22676 30304 22677 30344
rect 22635 30295 22677 30304
rect 22347 30176 22389 30185
rect 22347 30136 22348 30176
rect 22388 30136 22389 30176
rect 22347 30127 22389 30136
rect 23019 30092 23061 30101
rect 23019 30052 23020 30092
rect 23060 30052 23061 30092
rect 23212 30092 23252 33151
rect 23308 32864 23348 33412
rect 23500 33403 23540 33412
rect 23308 32815 23348 32824
rect 23596 32360 23636 33655
rect 24172 33570 24212 33655
rect 24556 33620 24596 34327
rect 25036 34217 25076 34336
rect 25420 34376 25460 34411
rect 25420 34325 25460 34336
rect 25516 34376 25556 34385
rect 25035 34208 25077 34217
rect 25035 34168 25036 34208
rect 25076 34168 25077 34208
rect 25035 34159 25077 34168
rect 25516 34049 25556 34336
rect 25612 34376 25652 35335
rect 25707 35132 25749 35141
rect 25707 35092 25708 35132
rect 25748 35092 25749 35132
rect 25707 35083 25749 35092
rect 25804 35132 25844 35419
rect 25612 34327 25652 34336
rect 25708 34376 25748 35083
rect 25708 34327 25748 34336
rect 25515 34040 25557 34049
rect 25515 34000 25516 34040
rect 25556 34000 25557 34040
rect 25515 33991 25557 34000
rect 25612 33704 25652 33713
rect 25804 33704 25844 35092
rect 25900 34385 25940 35848
rect 25996 35393 26036 36427
rect 25995 35384 26037 35393
rect 25995 35344 25996 35384
rect 26036 35344 26037 35384
rect 25995 35335 26037 35344
rect 25996 35216 26036 35335
rect 25996 35167 26036 35176
rect 26091 35216 26133 35225
rect 26091 35176 26092 35216
rect 26132 35176 26133 35216
rect 26091 35167 26133 35176
rect 26092 35082 26132 35167
rect 25899 34376 25941 34385
rect 25899 34336 25900 34376
rect 25940 34336 25941 34376
rect 25899 34327 25941 34336
rect 25900 34242 25940 34327
rect 25995 34208 26037 34217
rect 25995 34168 25996 34208
rect 26036 34168 26037 34208
rect 25995 34159 26037 34168
rect 25996 33788 26036 34159
rect 26188 34049 26228 36688
rect 26283 36728 26325 36737
rect 26283 36688 26284 36728
rect 26324 36688 26325 36728
rect 26283 36679 26325 36688
rect 26380 36728 26420 36856
rect 26284 36594 26324 36679
rect 26380 35468 26420 36688
rect 26380 35428 26516 35468
rect 26379 35300 26421 35309
rect 26379 35260 26380 35300
rect 26420 35260 26421 35300
rect 26379 35251 26421 35260
rect 26284 35216 26324 35225
rect 26284 34469 26324 35176
rect 26380 35166 26420 35251
rect 26476 35216 26516 35428
rect 26476 35141 26516 35176
rect 26572 35216 26612 37183
rect 27051 36476 27093 36485
rect 27051 36436 27052 36476
rect 27092 36436 27093 36476
rect 27051 36427 27093 36436
rect 27052 36342 27092 36427
rect 27436 35888 27476 37519
rect 27820 37434 27860 37519
rect 27627 37400 27669 37409
rect 27627 37360 27628 37400
rect 27668 37360 27669 37400
rect 27627 37351 27669 37360
rect 30988 37400 31028 37409
rect 27628 37266 27668 37351
rect 27531 37232 27573 37241
rect 27531 37192 27532 37232
rect 27572 37192 27573 37232
rect 27531 37183 27573 37192
rect 30892 37232 30932 37241
rect 27532 37098 27572 37183
rect 27436 35839 27476 35848
rect 27724 36728 27764 36737
rect 27052 35804 27092 35813
rect 27092 35764 27284 35804
rect 27052 35755 27092 35764
rect 26859 35720 26901 35729
rect 26859 35680 26860 35720
rect 26900 35680 26901 35720
rect 26859 35671 26901 35680
rect 26860 35586 26900 35671
rect 27244 35384 27284 35764
rect 27724 35477 27764 36688
rect 28012 36728 28052 36737
rect 28012 35729 28052 36688
rect 28683 36728 28725 36737
rect 28683 36688 28684 36728
rect 28724 36688 28725 36728
rect 28683 36679 28725 36688
rect 28971 36728 29013 36737
rect 28971 36688 28972 36728
rect 29012 36688 29013 36728
rect 28971 36679 29013 36688
rect 30508 36728 30548 36737
rect 28684 36594 28724 36679
rect 28972 36594 29012 36679
rect 29644 36604 30068 36644
rect 29644 36560 29684 36604
rect 29644 36511 29684 36520
rect 29068 36476 29108 36485
rect 29836 36476 29876 36485
rect 29108 36436 29588 36476
rect 29068 36427 29108 36436
rect 29163 36140 29205 36149
rect 29163 36100 29164 36140
rect 29204 36100 29205 36140
rect 29163 36091 29205 36100
rect 29451 36140 29493 36149
rect 29451 36100 29452 36140
rect 29492 36100 29493 36140
rect 29451 36091 29493 36100
rect 28300 35888 28340 35897
rect 28011 35720 28053 35729
rect 28011 35680 28012 35720
rect 28052 35680 28053 35720
rect 28011 35671 28053 35680
rect 27723 35468 27765 35477
rect 27723 35428 27724 35468
rect 27764 35428 27765 35468
rect 27723 35419 27765 35428
rect 27244 35335 27284 35344
rect 26572 35167 26612 35176
rect 26763 35216 26805 35225
rect 26763 35176 26764 35216
rect 26804 35176 26805 35216
rect 26763 35167 26805 35176
rect 26860 35216 26900 35227
rect 26475 35132 26517 35141
rect 26475 35092 26476 35132
rect 26516 35092 26517 35132
rect 26475 35083 26517 35092
rect 26764 35082 26804 35167
rect 26860 35141 26900 35176
rect 27052 35216 27092 35225
rect 27916 35216 27956 35225
rect 27092 35176 27380 35216
rect 27052 35167 27092 35176
rect 26859 35132 26901 35141
rect 26859 35092 26860 35132
rect 26900 35092 26901 35132
rect 26859 35083 26901 35092
rect 27051 35048 27093 35057
rect 27051 35008 27052 35048
rect 27092 35008 27093 35048
rect 27051 34999 27093 35008
rect 27052 34914 27092 34999
rect 26859 34544 26901 34553
rect 26859 34504 26860 34544
rect 26900 34504 26901 34544
rect 26859 34495 26901 34504
rect 26283 34460 26325 34469
rect 26283 34420 26284 34460
rect 26324 34420 26325 34460
rect 26283 34411 26325 34420
rect 26860 34376 26900 34495
rect 26860 34327 26900 34336
rect 27340 34376 27380 35176
rect 27916 35057 27956 35176
rect 27915 35048 27957 35057
rect 27915 35008 27916 35048
rect 27956 35008 27957 35048
rect 27915 34999 27957 35008
rect 28012 34796 28052 35671
rect 28300 35309 28340 35848
rect 28299 35300 28341 35309
rect 28299 35260 28300 35300
rect 28340 35260 28341 35300
rect 28299 35251 28341 35260
rect 28492 35132 28532 35141
rect 28299 35048 28341 35057
rect 28299 35008 28300 35048
rect 28340 35008 28341 35048
rect 28299 34999 28341 35008
rect 28300 34914 28340 34999
rect 28012 34756 28340 34796
rect 27531 34628 27573 34637
rect 27531 34588 27532 34628
rect 27572 34588 27573 34628
rect 27531 34579 27573 34588
rect 28203 34628 28245 34637
rect 28203 34588 28204 34628
rect 28244 34588 28245 34628
rect 28203 34579 28245 34588
rect 27340 34327 27380 34336
rect 27436 34376 27476 34385
rect 26187 34040 26229 34049
rect 26187 34000 26188 34040
rect 26228 34000 26229 34040
rect 26187 33991 26229 34000
rect 26763 34040 26805 34049
rect 26763 34000 26764 34040
rect 26804 34000 26805 34040
rect 26763 33991 26805 34000
rect 25996 33739 26036 33748
rect 25900 33704 25940 33713
rect 25804 33664 25900 33704
rect 25036 33620 25076 33629
rect 24556 33580 25036 33620
rect 23691 33536 23733 33545
rect 23691 33496 23692 33536
rect 23732 33496 23733 33536
rect 23691 33487 23733 33496
rect 24363 33536 24405 33545
rect 24363 33496 24364 33536
rect 24404 33496 24405 33536
rect 24363 33487 24405 33496
rect 23692 32864 23732 33487
rect 23787 33452 23829 33461
rect 23787 33412 23788 33452
rect 23828 33412 23829 33452
rect 23787 33403 23829 33412
rect 23692 32815 23732 32824
rect 23788 32696 23828 33403
rect 24364 33402 24404 33487
rect 24556 32864 24596 33580
rect 25036 33571 25076 33580
rect 25612 33209 25652 33664
rect 25900 33655 25940 33664
rect 25611 33200 25653 33209
rect 26188 33200 26228 33991
rect 26764 33704 26804 33991
rect 26764 33655 26804 33664
rect 27436 33536 27476 34336
rect 27532 34376 27572 34579
rect 27532 34327 27572 34336
rect 27628 34376 27668 34385
rect 27628 33872 27668 34336
rect 27916 34376 27956 34387
rect 27916 34301 27956 34336
rect 28204 34376 28244 34579
rect 28204 34327 28244 34336
rect 28300 34376 28340 34756
rect 28492 34469 28532 35092
rect 28876 35048 28916 35057
rect 28960 35048 29000 35076
rect 28916 35008 29012 35048
rect 28876 34999 28916 35008
rect 28588 34544 28628 34553
rect 28491 34460 28533 34469
rect 28491 34420 28492 34460
rect 28532 34420 28533 34460
rect 28491 34411 28533 34420
rect 28300 34327 28340 34336
rect 27915 34292 27957 34301
rect 27915 34252 27916 34292
rect 27956 34252 27957 34292
rect 27915 34243 27957 34252
rect 26283 33452 26325 33461
rect 26283 33412 26284 33452
rect 26324 33412 26325 33452
rect 26283 33403 26325 33412
rect 26955 33452 26997 33461
rect 26955 33412 26956 33452
rect 26996 33412 26997 33452
rect 26955 33403 26997 33412
rect 26284 33318 26324 33403
rect 25611 33160 25612 33200
rect 25652 33160 25653 33200
rect 25611 33151 25653 33160
rect 25996 33160 26228 33200
rect 25708 32948 25748 32957
rect 24556 32815 24596 32824
rect 25611 32864 25653 32873
rect 25611 32824 25612 32864
rect 25652 32824 25653 32864
rect 25611 32815 25653 32824
rect 23596 32311 23636 32320
rect 23692 32656 23828 32696
rect 23500 32192 23540 32201
rect 23500 31613 23540 32152
rect 23692 32192 23732 32656
rect 23692 32143 23732 32152
rect 23788 32192 23828 32201
rect 24843 32192 24885 32201
rect 23828 32152 24116 32192
rect 23788 32143 23828 32152
rect 23499 31604 23541 31613
rect 23499 31564 23500 31604
rect 23540 31564 23541 31604
rect 23499 31555 23541 31564
rect 24076 31520 24116 32152
rect 24843 32152 24844 32192
rect 24884 32152 24885 32192
rect 24843 32143 24885 32152
rect 25228 32192 25268 32201
rect 24844 32058 24884 32143
rect 25228 31529 25268 32152
rect 24076 31471 24116 31480
rect 24555 31520 24597 31529
rect 24555 31480 24556 31520
rect 24596 31480 24597 31520
rect 24555 31471 24597 31480
rect 25227 31520 25269 31529
rect 25227 31480 25228 31520
rect 25268 31480 25269 31520
rect 25227 31471 25269 31480
rect 24556 31386 24596 31471
rect 24172 31352 24212 31361
rect 24172 31193 24212 31312
rect 25420 31352 25460 31361
rect 24171 31184 24213 31193
rect 24171 31144 24172 31184
rect 24212 31144 24213 31184
rect 24171 31135 24213 31144
rect 24747 31184 24789 31193
rect 24747 31144 24748 31184
rect 24788 31144 24789 31184
rect 24747 31135 24789 31144
rect 24748 31050 24788 31135
rect 25420 30857 25460 31312
rect 25035 30848 25077 30857
rect 25035 30808 25036 30848
rect 25076 30808 25077 30848
rect 25035 30799 25077 30808
rect 25419 30848 25461 30857
rect 25419 30808 25420 30848
rect 25460 30808 25461 30848
rect 25419 30799 25461 30808
rect 25036 30714 25076 30799
rect 23884 30680 23924 30689
rect 23884 30269 23924 30640
rect 24171 30680 24213 30689
rect 24171 30640 24172 30680
rect 24212 30640 24213 30680
rect 24171 30631 24213 30640
rect 25516 30680 25556 30689
rect 23883 30260 23925 30269
rect 23883 30220 23884 30260
rect 23924 30220 23925 30260
rect 23883 30211 23925 30220
rect 23308 30092 23348 30101
rect 23212 30052 23308 30092
rect 23019 30043 23061 30052
rect 23308 30043 23348 30052
rect 24172 30092 24212 30631
rect 25323 30176 25365 30185
rect 25323 30136 25324 30176
rect 25364 30136 25365 30176
rect 25323 30127 25365 30136
rect 24172 30043 24212 30052
rect 24363 30092 24405 30101
rect 24363 30052 24364 30092
rect 24404 30052 24405 30092
rect 24363 30043 24405 30052
rect 22348 30008 22388 30017
rect 21964 29840 22004 29849
rect 21964 29345 22004 29800
rect 21963 29336 22005 29345
rect 21963 29296 21964 29336
rect 22004 29296 22005 29336
rect 21963 29287 22005 29296
rect 22348 29168 22388 29968
rect 23020 29840 23060 30043
rect 23020 29791 23060 29800
rect 23500 29672 23540 29681
rect 22923 29252 22965 29261
rect 22923 29212 22924 29252
rect 22964 29212 22965 29252
rect 22923 29203 22965 29212
rect 22540 29168 22580 29177
rect 22348 29128 22540 29168
rect 21291 29084 21333 29093
rect 21291 29044 21292 29084
rect 21332 29044 21333 29084
rect 21291 29035 21333 29044
rect 20524 28916 20564 28925
rect 20427 28832 20469 28841
rect 20427 28792 20428 28832
rect 20468 28792 20469 28832
rect 20427 28783 20469 28792
rect 20044 28624 20276 28664
rect 20331 28664 20373 28673
rect 20331 28624 20332 28664
rect 20372 28624 20373 28664
rect 20044 28580 20084 28624
rect 20331 28615 20373 28624
rect 20524 28580 20564 28876
rect 20715 28748 20757 28757
rect 20715 28708 20716 28748
rect 20756 28708 20757 28748
rect 20715 28699 20757 28708
rect 20044 28531 20084 28540
rect 20428 28540 20564 28580
rect 19660 28279 19700 28288
rect 19755 28328 19797 28337
rect 19755 28288 19756 28328
rect 19796 28288 19797 28328
rect 19755 28279 19797 28288
rect 19852 28328 19892 28337
rect 20044 28328 20084 28337
rect 19892 28288 20044 28328
rect 19852 28279 19892 28288
rect 20044 28279 20084 28288
rect 20235 28328 20277 28337
rect 20235 28288 20236 28328
rect 20276 28288 20277 28328
rect 20235 28279 20277 28288
rect 20332 28328 20372 28339
rect 19756 28194 19796 28279
rect 20236 28169 20276 28279
rect 20332 28253 20372 28288
rect 20331 28244 20373 28253
rect 20331 28204 20332 28244
rect 20372 28204 20373 28244
rect 20331 28195 20373 28204
rect 19275 28120 19276 28160
rect 19316 28120 19508 28160
rect 20235 28160 20277 28169
rect 20235 28120 20236 28160
rect 20276 28120 20277 28160
rect 19275 28111 19317 28120
rect 20235 28111 20277 28120
rect 19179 28076 19221 28085
rect 19084 28036 19180 28076
rect 19220 28036 19221 28076
rect 19179 28027 19221 28036
rect 18412 27607 18452 27616
rect 19180 27572 19220 28027
rect 19180 27523 19220 27532
rect 18987 27404 19029 27413
rect 19276 27404 19316 28111
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 20428 27824 20468 28540
rect 20523 28328 20565 28337
rect 20523 28288 20524 28328
rect 20564 28288 20565 28328
rect 20523 28279 20565 28288
rect 20620 28328 20660 28337
rect 20524 27992 20564 28279
rect 20620 28160 20660 28288
rect 20716 28328 20756 28699
rect 20716 28279 20756 28288
rect 21100 28328 21140 28337
rect 21003 28244 21045 28253
rect 21003 28204 21004 28244
rect 21044 28204 21045 28244
rect 21003 28195 21045 28204
rect 20715 28160 20757 28169
rect 20620 28120 20716 28160
rect 20756 28120 20757 28160
rect 20715 28111 20757 28120
rect 20812 28160 20852 28169
rect 20852 28120 20948 28160
rect 20812 28111 20852 28120
rect 20524 27952 20756 27992
rect 20044 27784 20468 27824
rect 19851 27740 19893 27749
rect 19851 27700 19852 27740
rect 19892 27700 19893 27740
rect 19851 27691 19893 27700
rect 19563 27656 19605 27665
rect 19563 27616 19564 27656
rect 19604 27616 19605 27656
rect 19563 27607 19605 27616
rect 19564 27488 19604 27607
rect 19852 27606 19892 27691
rect 19948 27656 19988 27665
rect 20044 27656 20084 27784
rect 19988 27616 20084 27656
rect 20236 27656 20276 27665
rect 20524 27656 20564 27665
rect 19948 27607 19988 27616
rect 19564 27439 19604 27448
rect 18987 27364 18988 27404
rect 19028 27364 19029 27404
rect 18987 27355 19029 27364
rect 19180 27364 19316 27404
rect 19371 27404 19413 27413
rect 19371 27364 19372 27404
rect 19412 27364 19413 27404
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 17739 27068 17781 27077
rect 17739 27028 17740 27068
rect 17780 27028 17781 27068
rect 17739 27019 17781 27028
rect 17644 26767 17684 26776
rect 17740 26816 17780 27019
rect 18027 26984 18069 26993
rect 18027 26944 18028 26984
rect 18068 26944 18069 26984
rect 18027 26935 18069 26944
rect 18028 26850 18068 26935
rect 17547 26396 17589 26405
rect 17547 26356 17548 26396
rect 17588 26356 17589 26396
rect 17547 26347 17589 26356
rect 17740 26153 17780 26776
rect 18700 26816 18740 26825
rect 17836 26648 17876 26657
rect 17876 26608 17972 26648
rect 17836 26599 17876 26608
rect 17932 26396 17972 26608
rect 18700 26489 18740 26776
rect 18891 26732 18933 26741
rect 18891 26692 18892 26732
rect 18932 26692 18933 26732
rect 18891 26683 18933 26692
rect 18699 26480 18741 26489
rect 18699 26440 18700 26480
rect 18740 26440 18741 26480
rect 18699 26431 18741 26440
rect 17932 26356 18452 26396
rect 18219 26228 18261 26237
rect 18219 26188 18220 26228
rect 18260 26188 18261 26228
rect 18219 26179 18261 26188
rect 17548 26144 17588 26153
rect 17451 26060 17493 26069
rect 17355 26020 17396 26060
rect 17259 26011 17301 26020
rect 16916 25936 17108 25976
rect 16876 25927 16916 25936
rect 16683 25724 16725 25733
rect 16683 25684 16684 25724
rect 16724 25684 16725 25724
rect 16683 25675 16725 25684
rect 16491 25388 16533 25397
rect 16491 25348 16492 25388
rect 16532 25348 16533 25388
rect 16491 25339 16533 25348
rect 16971 25304 17013 25313
rect 16971 25264 16972 25304
rect 17012 25264 17013 25304
rect 16971 25255 17013 25264
rect 17164 25304 17204 25313
rect 16395 24800 16437 24809
rect 16876 24800 16916 24809
rect 16395 24760 16396 24800
rect 16436 24760 16437 24800
rect 16395 24751 16437 24760
rect 16492 24760 16876 24800
rect 16300 24583 16340 24592
rect 16395 24632 16437 24641
rect 16395 24592 16396 24632
rect 16436 24592 16437 24632
rect 16395 24583 16437 24592
rect 16492 24632 16532 24760
rect 16876 24751 16916 24760
rect 16492 24583 16532 24592
rect 16684 24632 16724 24641
rect 15820 24498 15860 24583
rect 16012 24498 16052 24583
rect 16396 24498 16436 24583
rect 16684 24473 16724 24592
rect 16780 24632 16820 24641
rect 16972 24632 17012 25255
rect 16820 24592 16916 24632
rect 16780 24583 16820 24592
rect 15572 24424 15764 24464
rect 15915 24464 15957 24473
rect 15915 24424 15916 24464
rect 15956 24424 15957 24464
rect 15532 24415 15572 24424
rect 15915 24415 15957 24424
rect 16683 24464 16725 24473
rect 16683 24424 16684 24464
rect 16724 24424 16725 24464
rect 16683 24415 16725 24424
rect 15627 24128 15669 24137
rect 15627 24088 15628 24128
rect 15668 24088 15669 24128
rect 15627 24079 15669 24088
rect 15531 23960 15573 23969
rect 15531 23920 15532 23960
rect 15572 23920 15573 23960
rect 15531 23911 15573 23920
rect 15532 23465 15572 23911
rect 15628 23792 15668 24079
rect 15628 23743 15668 23752
rect 15724 23792 15764 23801
rect 15724 23633 15764 23752
rect 15723 23624 15765 23633
rect 15916 23624 15956 24415
rect 16203 24044 16245 24053
rect 16203 24004 16204 24044
rect 16244 24004 16245 24044
rect 16203 23995 16245 24004
rect 15723 23584 15724 23624
rect 15764 23584 15860 23624
rect 15723 23575 15765 23584
rect 15531 23456 15573 23465
rect 15531 23416 15532 23456
rect 15572 23416 15573 23456
rect 15531 23407 15573 23416
rect 15627 23288 15669 23297
rect 15627 23248 15628 23288
rect 15668 23248 15669 23288
rect 15820 23288 15860 23584
rect 15916 23575 15956 23584
rect 16108 23792 16148 23801
rect 16108 23465 16148 23752
rect 16204 23792 16244 23995
rect 16396 23969 16436 24054
rect 16587 24044 16629 24053
rect 16587 24004 16588 24044
rect 16628 24004 16629 24044
rect 16587 23995 16629 24004
rect 16395 23960 16437 23969
rect 16395 23920 16396 23960
rect 16436 23920 16437 23960
rect 16395 23911 16437 23920
rect 16204 23540 16244 23752
rect 16396 23792 16436 23801
rect 16588 23792 16628 23995
rect 16683 23876 16725 23885
rect 16683 23836 16684 23876
rect 16724 23836 16725 23876
rect 16683 23827 16725 23836
rect 16436 23752 16532 23792
rect 16396 23743 16436 23752
rect 16492 23624 16532 23752
rect 16588 23743 16628 23752
rect 16684 23792 16724 23827
rect 16780 23801 16820 23886
rect 16684 23741 16724 23752
rect 16779 23792 16821 23801
rect 16779 23752 16780 23792
rect 16820 23752 16821 23792
rect 16876 23792 16916 24592
rect 16972 24583 17012 24592
rect 17164 24464 17204 25264
rect 17260 25304 17300 25313
rect 17356 25304 17396 26020
rect 17451 26020 17452 26060
rect 17492 26020 17493 26060
rect 17451 26011 17493 26020
rect 17451 25724 17493 25733
rect 17451 25684 17452 25724
rect 17492 25684 17493 25724
rect 17451 25675 17493 25684
rect 17452 25556 17492 25675
rect 17452 25507 17492 25516
rect 17451 25388 17493 25397
rect 17451 25348 17452 25388
rect 17492 25348 17493 25388
rect 17451 25339 17493 25348
rect 17300 25264 17396 25304
rect 17452 25304 17492 25339
rect 17260 25255 17300 25264
rect 17452 25253 17492 25264
rect 17548 25145 17588 26104
rect 17739 26144 17781 26153
rect 18124 26144 18164 26153
rect 17739 26104 17740 26144
rect 17780 26104 17781 26144
rect 17739 26095 17781 26104
rect 17932 26104 18124 26144
rect 17932 25556 17972 26104
rect 18124 26095 18164 26104
rect 18220 26144 18260 26179
rect 18220 26093 18260 26104
rect 18412 26144 18452 26356
rect 18412 26095 18452 26104
rect 18700 26144 18740 26153
rect 18411 25976 18453 25985
rect 18411 25936 18412 25976
rect 18452 25936 18453 25976
rect 18411 25927 18453 25936
rect 18412 25842 18452 25927
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 17932 25507 17972 25516
rect 17931 25388 17973 25397
rect 17931 25348 17932 25388
rect 17972 25348 18260 25388
rect 17931 25339 17973 25348
rect 17644 25304 17684 25313
rect 17547 25136 17589 25145
rect 17547 25096 17548 25136
rect 17588 25096 17589 25136
rect 17547 25087 17589 25096
rect 17164 24415 17204 24424
rect 17452 24632 17492 24641
rect 17067 23960 17109 23969
rect 17067 23920 17068 23960
rect 17108 23920 17109 23960
rect 17067 23911 17109 23920
rect 17068 23792 17108 23911
rect 16876 23752 17012 23792
rect 16779 23743 16821 23752
rect 16876 23624 16916 23633
rect 16492 23584 16876 23624
rect 16876 23575 16916 23584
rect 16972 23549 17012 23752
rect 17068 23743 17108 23752
rect 17355 23624 17397 23633
rect 17355 23584 17356 23624
rect 17396 23584 17397 23624
rect 17355 23575 17397 23584
rect 16971 23540 17013 23549
rect 16204 23500 16436 23540
rect 16107 23456 16149 23465
rect 16107 23416 16108 23456
rect 16148 23416 16149 23456
rect 16107 23407 16149 23416
rect 16012 23288 16052 23297
rect 15820 23248 16012 23288
rect 16052 23248 16340 23288
rect 15627 23239 15669 23248
rect 16012 23239 16052 23248
rect 15435 22448 15477 22457
rect 15435 22408 15436 22448
rect 15476 22408 15477 22448
rect 15435 22399 15477 22408
rect 15531 22280 15573 22289
rect 15531 22240 15532 22280
rect 15572 22240 15573 22280
rect 15531 22231 15573 22240
rect 15628 22280 15668 23239
rect 15723 23120 15765 23129
rect 15723 23080 15724 23120
rect 15764 23080 15765 23120
rect 15723 23071 15765 23080
rect 16300 23120 16340 23248
rect 16300 23071 16340 23080
rect 15724 22448 15764 23071
rect 15724 22399 15764 22408
rect 16108 22280 16148 22289
rect 15628 22240 16108 22280
rect 15532 22146 15572 22231
rect 15436 21776 15476 21785
rect 15628 21776 15668 22240
rect 16108 22231 16148 22240
rect 16203 22280 16245 22289
rect 16203 22240 16204 22280
rect 16244 22240 16245 22280
rect 16203 22231 16245 22240
rect 15476 21736 15668 21776
rect 15436 21727 15476 21736
rect 15628 21608 15668 21617
rect 15340 21568 15628 21608
rect 15628 21559 15668 21568
rect 15724 21608 15764 21617
rect 15724 21020 15764 21568
rect 15052 20980 15188 21020
rect 15532 20980 15764 21020
rect 14667 20852 14709 20861
rect 14667 20812 14668 20852
rect 14708 20812 14709 20852
rect 14667 20803 14709 20812
rect 14380 20140 14516 20180
rect 12555 20012 12597 20021
rect 12555 19972 12556 20012
rect 12596 19972 12597 20012
rect 12555 19963 12597 19972
rect 11980 19384 12404 19424
rect 11307 19340 11349 19349
rect 11307 19300 11308 19340
rect 11348 19300 11349 19340
rect 11307 19291 11349 19300
rect 10635 19256 10677 19265
rect 10635 19216 10636 19256
rect 10676 19216 10677 19256
rect 10635 19207 10677 19216
rect 10827 19256 10869 19265
rect 10827 19216 10828 19256
rect 10868 19216 10869 19256
rect 10827 19207 10869 19216
rect 11308 19256 11348 19291
rect 10636 19122 10676 19207
rect 10540 18712 10676 18752
rect 10252 18584 10292 18593
rect 10252 17753 10292 18544
rect 10348 18584 10388 18593
rect 9292 17695 9332 17704
rect 10156 17695 10196 17704
rect 10251 17744 10293 17753
rect 10251 17704 10252 17744
rect 10292 17704 10293 17744
rect 10251 17695 10293 17704
rect 8716 17610 8756 17695
rect 10348 17585 10388 18544
rect 10444 18584 10484 18595
rect 10444 18509 10484 18544
rect 10539 18584 10581 18593
rect 10539 18544 10540 18584
rect 10580 18544 10581 18584
rect 10539 18535 10581 18544
rect 10443 18500 10485 18509
rect 10443 18460 10444 18500
rect 10484 18460 10485 18500
rect 10443 18451 10485 18460
rect 10540 18450 10580 18535
rect 10636 18509 10676 18712
rect 10828 18584 10868 19207
rect 11308 19205 11348 19216
rect 11692 19256 11732 19265
rect 11596 18752 11636 18761
rect 11692 18752 11732 19216
rect 11787 19256 11829 19265
rect 11787 19216 11788 19256
rect 11828 19216 11829 19256
rect 11787 19207 11829 19216
rect 11980 19256 12020 19265
rect 11788 19122 11828 19207
rect 11636 18712 11732 18752
rect 11116 18677 11156 18708
rect 11115 18668 11157 18677
rect 11115 18628 11116 18668
rect 11156 18628 11157 18668
rect 11115 18619 11157 18628
rect 10828 18535 10868 18544
rect 11116 18584 11156 18619
rect 11596 18593 11636 18712
rect 11980 18677 12020 19216
rect 12075 19256 12117 19265
rect 12075 19216 12076 19256
rect 12116 19216 12117 19256
rect 12075 19207 12117 19216
rect 12268 19256 12308 19265
rect 12076 19122 12116 19207
rect 12171 19088 12213 19097
rect 12171 19048 12172 19088
rect 12212 19048 12213 19088
rect 12171 19039 12213 19048
rect 12172 18954 12212 19039
rect 12268 18761 12308 19216
rect 12267 18752 12309 18761
rect 12267 18712 12268 18752
rect 12308 18712 12309 18752
rect 12267 18703 12309 18712
rect 11979 18668 12021 18677
rect 11979 18628 11980 18668
rect 12020 18628 12021 18668
rect 11979 18619 12021 18628
rect 11116 18509 11156 18544
rect 11212 18584 11252 18593
rect 10635 18500 10677 18509
rect 10635 18460 10636 18500
rect 10676 18460 10677 18500
rect 10635 18451 10677 18460
rect 11115 18500 11157 18509
rect 11115 18460 11116 18500
rect 11156 18460 11157 18500
rect 11115 18451 11157 18460
rect 11212 18425 11252 18544
rect 11308 18584 11348 18593
rect 11211 18416 11253 18425
rect 11211 18376 11212 18416
rect 11252 18376 11253 18416
rect 11211 18367 11253 18376
rect 10924 18332 10964 18341
rect 10347 17576 10389 17585
rect 10347 17536 10348 17576
rect 10388 17536 10389 17576
rect 10347 17527 10389 17536
rect 9387 17072 9429 17081
rect 9387 17032 9388 17072
rect 9428 17032 9429 17072
rect 9387 17023 9429 17032
rect 9388 16232 9428 17023
rect 9868 16904 9908 16913
rect 9388 16183 9428 16192
rect 9772 16232 9812 16241
rect 9868 16232 9908 16864
rect 9812 16192 9908 16232
rect 10540 16820 10580 16829
rect 9772 16183 9812 16192
rect 8524 16024 8660 16064
rect 8140 15509 8180 15520
rect 8331 15560 8373 15569
rect 8331 15520 8332 15560
rect 8372 15520 8373 15560
rect 8331 15511 8373 15520
rect 8524 15560 8564 16024
rect 10540 15737 10580 16780
rect 10924 16241 10964 18292
rect 11308 18164 11348 18544
rect 11404 18584 11444 18593
rect 11595 18584 11637 18593
rect 11444 18544 11540 18584
rect 11404 18535 11444 18544
rect 11212 18124 11348 18164
rect 11212 17585 11252 18124
rect 11307 17996 11349 18005
rect 11307 17956 11308 17996
rect 11348 17956 11349 17996
rect 11307 17947 11349 17956
rect 11308 17862 11348 17947
rect 11211 17576 11253 17585
rect 11211 17536 11212 17576
rect 11252 17536 11253 17576
rect 11211 17527 11253 17536
rect 11500 17240 11540 18544
rect 11595 18544 11596 18584
rect 11636 18544 11637 18584
rect 11595 18535 11637 18544
rect 11980 18080 12020 18619
rect 12268 18584 12308 18593
rect 12364 18584 12404 19384
rect 12460 19172 12500 19181
rect 12460 18752 12500 19132
rect 12460 18703 12500 18712
rect 12556 18584 12596 19963
rect 13228 19928 13268 19937
rect 12844 19256 12884 19265
rect 13228 19256 13268 19888
rect 12884 19216 13268 19256
rect 13708 19256 13748 19265
rect 13748 19216 13844 19256
rect 12844 19207 12884 19216
rect 13708 19207 13748 19216
rect 13131 19088 13173 19097
rect 13131 19048 13132 19088
rect 13172 19048 13173 19088
rect 13131 19039 13173 19048
rect 12308 18544 12404 18584
rect 12460 18544 12596 18584
rect 13132 18584 13172 19039
rect 13323 18836 13365 18845
rect 13323 18796 13324 18836
rect 13364 18796 13365 18836
rect 13323 18787 13365 18796
rect 13324 18752 13364 18787
rect 13324 18701 13364 18712
rect 11980 18040 12212 18080
rect 11692 17744 11732 17753
rect 11732 17704 12116 17744
rect 11692 17695 11732 17704
rect 11500 17200 11924 17240
rect 11212 17072 11252 17081
rect 11212 16409 11252 17032
rect 11596 17072 11636 17081
rect 11596 16484 11636 17032
rect 11788 16484 11828 16493
rect 11596 16444 11788 16484
rect 11788 16435 11828 16444
rect 11211 16400 11253 16409
rect 11211 16360 11212 16400
rect 11252 16360 11253 16400
rect 11211 16351 11253 16360
rect 11691 16316 11733 16325
rect 11691 16276 11692 16316
rect 11732 16276 11733 16316
rect 11691 16267 11733 16276
rect 10636 16232 10676 16241
rect 8619 15728 8661 15737
rect 10539 15728 10581 15737
rect 8619 15688 8620 15728
rect 8660 15688 8661 15728
rect 8619 15679 8661 15688
rect 9004 15688 9428 15728
rect 7947 15476 7989 15485
rect 7947 15436 7948 15476
rect 7988 15436 7989 15476
rect 7947 15427 7989 15436
rect 7948 15342 7988 15427
rect 8043 15056 8085 15065
rect 8043 15016 8044 15056
rect 8084 15016 8085 15056
rect 8043 15007 8085 15016
rect 7947 14972 7989 14981
rect 7947 14932 7948 14972
rect 7988 14932 7989 14972
rect 7947 14923 7989 14932
rect 7756 14720 7796 14729
rect 7563 14216 7605 14225
rect 7563 14176 7564 14216
rect 7604 14176 7605 14216
rect 7756 14216 7796 14680
rect 7948 14720 7988 14923
rect 7948 14671 7988 14680
rect 8044 14720 8084 15007
rect 8044 14671 8084 14680
rect 8236 14720 8276 14729
rect 8332 14720 8372 15511
rect 8524 15485 8564 15520
rect 8523 15476 8565 15485
rect 8523 15436 8524 15476
rect 8564 15436 8565 15476
rect 8523 15427 8565 15436
rect 8524 15396 8564 15427
rect 8620 15140 8660 15679
rect 8715 15560 8757 15569
rect 8715 15520 8716 15560
rect 8756 15520 8757 15560
rect 8715 15511 8757 15520
rect 8812 15560 8852 15569
rect 9004 15560 9044 15688
rect 8852 15520 9044 15560
rect 9099 15560 9141 15569
rect 9099 15520 9100 15560
rect 9140 15520 9141 15560
rect 8812 15511 8852 15520
rect 9099 15511 9141 15520
rect 9292 15560 9332 15569
rect 8716 15426 8756 15511
rect 9100 15426 9140 15511
rect 8812 15392 8852 15401
rect 8620 15100 8756 15140
rect 8276 14680 8372 14720
rect 8716 14720 8756 15100
rect 8812 14897 8852 15352
rect 9004 15308 9044 15317
rect 8811 14888 8853 14897
rect 8811 14848 8812 14888
rect 8852 14848 8853 14888
rect 8811 14839 8853 14848
rect 8812 14720 8852 14729
rect 8716 14680 8812 14720
rect 8236 14671 8276 14680
rect 8812 14671 8852 14680
rect 8908 14720 8948 14729
rect 9004 14720 9044 15268
rect 9099 14972 9141 14981
rect 9099 14932 9100 14972
rect 9140 14932 9141 14972
rect 9099 14923 9141 14932
rect 9292 14972 9332 15520
rect 9292 14923 9332 14932
rect 9100 14838 9140 14923
rect 8948 14680 9044 14720
rect 9099 14720 9141 14729
rect 9099 14680 9100 14720
rect 9140 14680 9141 14720
rect 8908 14671 8948 14680
rect 9099 14671 9141 14680
rect 9100 14586 9140 14671
rect 8139 14552 8181 14561
rect 8139 14512 8140 14552
rect 8180 14512 8181 14552
rect 8139 14503 8181 14512
rect 8140 14418 8180 14503
rect 8044 14216 8084 14225
rect 7756 14176 8044 14216
rect 7563 14167 7605 14176
rect 8044 14167 8084 14176
rect 8715 14216 8757 14225
rect 8715 14176 8716 14216
rect 8756 14176 8757 14216
rect 8715 14167 8757 14176
rect 8716 14082 8756 14167
rect 9388 14048 9428 15688
rect 10539 15688 10540 15728
rect 10580 15688 10581 15728
rect 10539 15679 10581 15688
rect 9675 15560 9717 15569
rect 9675 15520 9676 15560
rect 9716 15520 9717 15560
rect 9675 15511 9717 15520
rect 10155 15560 10197 15569
rect 10155 15520 10156 15560
rect 10196 15520 10197 15560
rect 10155 15511 10197 15520
rect 10540 15560 10580 15569
rect 10636 15560 10676 16192
rect 10923 16232 10965 16241
rect 10923 16192 10924 16232
rect 10964 16192 10965 16232
rect 10923 16183 10965 16192
rect 11692 15728 11732 16267
rect 11884 16232 11924 17200
rect 12076 16400 12116 17704
rect 12076 16351 12116 16360
rect 12076 16232 12116 16241
rect 11884 16192 12076 16232
rect 12172 16232 12212 18040
rect 12268 18005 12308 18544
rect 12267 17996 12309 18005
rect 12267 17956 12268 17996
rect 12308 17956 12309 17996
rect 12267 17947 12309 17956
rect 12363 17744 12405 17753
rect 12363 17704 12364 17744
rect 12404 17704 12405 17744
rect 12363 17695 12405 17704
rect 12364 17610 12404 17695
rect 12460 17072 12500 18544
rect 13132 18535 13172 18544
rect 12939 18416 12981 18425
rect 12939 18376 12940 18416
rect 12980 18376 12981 18416
rect 12939 18367 12981 18376
rect 12555 17744 12597 17753
rect 12555 17704 12556 17744
rect 12596 17704 12597 17744
rect 12555 17695 12597 17704
rect 12940 17744 12980 18367
rect 13804 17753 13844 19216
rect 13996 18584 14036 20140
rect 14476 20021 14516 20140
rect 14475 20012 14517 20021
rect 14475 19972 14476 20012
rect 14516 19972 14517 20012
rect 14475 19963 14517 19972
rect 13996 18509 14036 18544
rect 13995 18500 14037 18509
rect 13995 18460 13996 18500
rect 14036 18460 14037 18500
rect 13995 18451 14037 18460
rect 14187 18416 14229 18425
rect 14187 18376 14188 18416
rect 14228 18376 14229 18416
rect 14187 18367 14229 18376
rect 14188 18282 14228 18367
rect 12940 17695 12980 17704
rect 13803 17744 13845 17753
rect 13803 17704 13804 17744
rect 13844 17704 13845 17744
rect 13803 17695 13845 17704
rect 14187 17744 14229 17753
rect 14187 17704 14188 17744
rect 14228 17704 14229 17744
rect 14187 17695 14229 17704
rect 12556 17610 12596 17695
rect 12651 17660 12693 17669
rect 12651 17620 12652 17660
rect 12692 17620 12693 17660
rect 12651 17611 12693 17620
rect 13611 17660 13653 17669
rect 13611 17620 13612 17660
rect 13652 17620 13653 17660
rect 13611 17611 13653 17620
rect 12460 17023 12500 17032
rect 12652 17072 12692 17611
rect 12652 17023 12692 17032
rect 13612 17072 13652 17611
rect 13804 17610 13844 17695
rect 14091 17660 14133 17669
rect 14091 17620 14092 17660
rect 14132 17620 14133 17660
rect 14091 17611 14133 17620
rect 13612 17023 13652 17032
rect 12939 16820 12981 16829
rect 12939 16780 12940 16820
rect 12980 16780 12981 16820
rect 12939 16771 12981 16780
rect 12268 16232 12308 16241
rect 12172 16192 12268 16232
rect 12076 16183 12116 16192
rect 12268 16183 12308 16192
rect 12363 16232 12405 16241
rect 12363 16192 12364 16232
rect 12404 16192 12405 16232
rect 12363 16183 12405 16192
rect 12747 16232 12789 16241
rect 12747 16192 12748 16232
rect 12788 16192 12789 16232
rect 12747 16183 12789 16192
rect 12364 16098 12404 16183
rect 11692 15679 11732 15688
rect 10580 15520 10676 15560
rect 9676 15426 9716 15511
rect 9963 14972 10005 14981
rect 9963 14932 9964 14972
rect 10004 14932 10005 14972
rect 9963 14923 10005 14932
rect 9964 14720 10004 14923
rect 10156 14888 10196 15511
rect 10156 14839 10196 14848
rect 9964 14671 10004 14680
rect 9579 14132 9621 14141
rect 9579 14092 9580 14132
rect 9620 14092 9621 14132
rect 9579 14083 9621 14092
rect 8236 13880 8276 13889
rect 8140 13840 8236 13880
rect 7275 13460 7317 13469
rect 7275 13420 7276 13460
rect 7316 13420 7317 13460
rect 7275 13411 7317 13420
rect 7180 13159 7220 13168
rect 6796 13074 6836 13159
rect 6411 12620 6453 12629
rect 6411 12580 6412 12620
rect 6452 12580 6453 12620
rect 6411 12571 6453 12580
rect 7083 12536 7125 12545
rect 7083 12496 7084 12536
rect 7124 12496 7125 12536
rect 7083 12487 7125 12496
rect 7084 12402 7124 12487
rect 6220 12319 6260 12328
rect 6604 12368 6644 12377
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 6027 11696 6069 11705
rect 6027 11656 6028 11696
rect 6068 11656 6069 11696
rect 6027 11647 6069 11656
rect 6412 11696 6452 11705
rect 6604 11696 6644 12328
rect 6987 12368 7029 12377
rect 6987 12328 6988 12368
rect 7028 12328 7029 12368
rect 6987 12319 7029 12328
rect 6988 12234 7028 12319
rect 6452 11656 6644 11696
rect 7276 11696 7316 13411
rect 7564 13208 7604 13217
rect 8140 13208 8180 13840
rect 8236 13831 8276 13840
rect 8716 13796 8756 13805
rect 8427 13292 8469 13301
rect 8427 13252 8428 13292
rect 8468 13252 8469 13292
rect 8427 13243 8469 13252
rect 7604 13168 8180 13208
rect 8428 13208 8468 13243
rect 7564 13159 7604 13168
rect 8428 13157 8468 13168
rect 8332 12536 8372 12547
rect 8332 12461 8372 12496
rect 8619 12536 8661 12545
rect 8619 12496 8620 12536
rect 8660 12496 8661 12536
rect 8619 12487 8661 12496
rect 8331 12452 8373 12461
rect 8331 12412 8332 12452
rect 8372 12412 8373 12452
rect 8331 12403 8373 12412
rect 8620 12402 8660 12487
rect 6412 11647 6452 11656
rect 6028 11562 6068 11647
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 7276 11453 7316 11656
rect 7468 12368 7508 12377
rect 7275 11444 7317 11453
rect 7275 11404 7276 11444
rect 7316 11404 7317 11444
rect 7275 11395 7317 11404
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 652 11192 692 11201
rect 652 10697 692 11152
rect 7468 11033 7508 12328
rect 7660 12284 7700 12293
rect 7660 11705 7700 12244
rect 8043 11948 8085 11957
rect 8043 11908 8044 11948
rect 8084 11908 8085 11948
rect 8043 11899 8085 11908
rect 8427 11948 8469 11957
rect 8427 11908 8428 11948
rect 8468 11908 8469 11948
rect 8427 11899 8469 11908
rect 7659 11696 7701 11705
rect 7659 11656 7660 11696
rect 7700 11656 7701 11696
rect 7659 11647 7701 11656
rect 7467 11024 7509 11033
rect 7467 10984 7468 11024
rect 7508 10984 7509 11024
rect 7467 10975 7509 10984
rect 7275 10772 7317 10781
rect 7275 10732 7276 10772
rect 7316 10732 7317 10772
rect 7275 10723 7317 10732
rect 7851 10772 7893 10781
rect 7851 10732 7852 10772
rect 7892 10732 7893 10772
rect 7851 10723 7893 10732
rect 651 10688 693 10697
rect 651 10648 652 10688
rect 692 10648 693 10688
rect 651 10639 693 10648
rect 7276 10638 7316 10723
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 6028 10352 6068 10361
rect 5547 10100 5589 10109
rect 5547 10060 5548 10100
rect 5588 10060 5589 10100
rect 5547 10051 5589 10060
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 652 9680 692 9689
rect 652 9017 692 9640
rect 5548 9596 5588 10051
rect 5548 9547 5588 9556
rect 5932 9512 5972 9521
rect 6028 9512 6068 10312
rect 6796 10352 6836 10361
rect 6796 9848 6836 10312
rect 7659 10184 7701 10193
rect 7852 10184 7892 10723
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 7756 10144 7852 10184
rect 6987 10100 7029 10109
rect 6987 10060 6988 10100
rect 7028 10060 7029 10100
rect 6987 10051 7029 10060
rect 6988 9966 7028 10051
rect 7660 10050 7700 10135
rect 6796 9808 7124 9848
rect 5972 9472 6068 9512
rect 6796 9512 6836 9521
rect 6836 9472 6932 9512
rect 5932 9463 5972 9472
rect 6796 9463 6836 9472
rect 3916 9344 3956 9353
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 3435 8840 3477 8849
rect 3435 8800 3436 8840
rect 3476 8800 3477 8840
rect 3435 8791 3477 8800
rect 3436 8672 3476 8791
rect 3436 8623 3476 8632
rect 3820 8672 3860 8681
rect 3916 8672 3956 9304
rect 6124 8849 6164 8934
rect 6123 8840 6165 8849
rect 6123 8800 6124 8840
rect 6164 8800 6165 8840
rect 6123 8791 6165 8800
rect 3860 8632 3956 8672
rect 4684 8672 4724 8681
rect 5931 8672 5973 8681
rect 6124 8672 6164 8681
rect 4724 8632 4820 8672
rect 3820 8623 3860 8632
rect 4684 8623 4724 8632
rect 652 8504 692 8513
rect 556 8464 652 8504
rect 556 8177 596 8464
rect 652 8455 692 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 555 8168 597 8177
rect 555 8128 556 8168
rect 596 8128 597 8168
rect 555 8119 597 8128
rect 652 8168 692 8177
rect 652 7337 692 8128
rect 4684 8009 4724 8094
rect 4492 8000 4532 8009
rect 2860 7832 2900 7841
rect 4492 7832 4532 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4684 7832 4724 7841
rect 4492 7792 4684 7832
rect 4780 7832 4820 8632
rect 5931 8632 5932 8672
rect 5972 8632 5973 8672
rect 5931 8623 5973 8632
rect 6028 8632 6124 8672
rect 5932 8538 5972 8623
rect 5260 8212 5588 8252
rect 4875 8084 4917 8093
rect 4875 8044 4876 8084
rect 4916 8044 4917 8084
rect 4875 8035 4917 8044
rect 4876 8000 4916 8035
rect 4876 7949 4916 7960
rect 4972 8000 5012 8009
rect 4972 7841 5012 7960
rect 5163 8000 5205 8009
rect 5163 7960 5164 8000
rect 5204 7960 5205 8000
rect 5163 7951 5205 7960
rect 5260 8000 5300 8212
rect 5452 8093 5492 8124
rect 5451 8084 5493 8093
rect 5451 8044 5452 8084
rect 5492 8044 5493 8084
rect 5451 8035 5493 8044
rect 5260 7951 5300 7960
rect 5356 8000 5396 8009
rect 5164 7866 5204 7951
rect 5356 7841 5396 7960
rect 5452 8000 5492 8035
rect 5548 8000 5588 8212
rect 5644 8168 5684 8177
rect 6028 8168 6068 8632
rect 6124 8623 6164 8632
rect 6219 8672 6261 8681
rect 6219 8632 6220 8672
rect 6260 8632 6261 8672
rect 6219 8623 6261 8632
rect 6316 8672 6356 8681
rect 5684 8128 6068 8168
rect 5644 8119 5684 8128
rect 5740 8000 5780 8009
rect 5548 7960 5740 8000
rect 4971 7832 5013 7841
rect 4780 7792 4916 7832
rect 2379 7748 2421 7757
rect 2379 7708 2380 7748
rect 2420 7708 2421 7748
rect 2379 7699 2421 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 2380 7160 2420 7699
rect 2380 7111 2420 7120
rect 2764 7160 2804 7169
rect 2860 7160 2900 7792
rect 4684 7783 4724 7792
rect 3819 7748 3861 7757
rect 3819 7708 3820 7748
rect 3860 7708 3861 7748
rect 3819 7699 3861 7708
rect 3820 7614 3860 7699
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4779 7496 4821 7505
rect 4779 7456 4780 7496
rect 4820 7456 4821 7496
rect 4779 7447 4821 7456
rect 4780 7412 4820 7447
rect 4780 7361 4820 7372
rect 2804 7120 2900 7160
rect 3627 7160 3669 7169
rect 3627 7120 3628 7160
rect 3668 7120 3669 7160
rect 4876 7160 4916 7792
rect 4971 7792 4972 7832
rect 5012 7792 5013 7832
rect 4971 7783 5013 7792
rect 5355 7832 5397 7841
rect 5355 7792 5356 7832
rect 5396 7792 5397 7832
rect 5355 7783 5397 7792
rect 5163 7496 5205 7505
rect 5163 7456 5164 7496
rect 5204 7456 5205 7496
rect 5163 7447 5205 7456
rect 4971 7160 5013 7169
rect 4876 7120 4972 7160
rect 5012 7120 5013 7160
rect 2764 7111 2804 7120
rect 3627 7111 3669 7120
rect 4971 7111 5013 7120
rect 5164 7160 5204 7447
rect 5452 7421 5492 7960
rect 5451 7412 5493 7421
rect 5451 7372 5452 7412
rect 5492 7372 5493 7412
rect 5451 7363 5493 7372
rect 5164 7111 5204 7120
rect 3628 7026 3668 7111
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 3723 6488 3765 6497
rect 3723 6448 3724 6488
rect 3764 6448 3765 6488
rect 3723 6439 3765 6448
rect 4108 6488 4148 6497
rect 4875 6488 4917 6497
rect 4148 6448 4244 6488
rect 4108 6439 4148 6448
rect 3724 6354 3764 6439
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4204 5816 4244 6448
rect 4875 6448 4876 6488
rect 4916 6448 4917 6488
rect 4875 6439 4917 6448
rect 4972 6488 5012 7111
rect 4684 5825 4724 5910
rect 4876 5900 4916 6439
rect 4876 5851 4916 5860
rect 4204 5767 4244 5776
rect 4683 5816 4725 5825
rect 4683 5776 4684 5816
rect 4724 5776 4725 5816
rect 4683 5767 4725 5776
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 4396 5648 4436 5657
rect 652 5480 692 5599
rect 4396 5489 4436 5608
rect 4587 5648 4629 5657
rect 4587 5608 4588 5648
rect 4628 5608 4629 5648
rect 4587 5599 4629 5608
rect 4684 5648 4724 5657
rect 4588 5514 4628 5599
rect 4684 5489 4724 5608
rect 652 5431 692 5440
rect 4395 5480 4437 5489
rect 4395 5440 4396 5480
rect 4436 5440 4437 5480
rect 4395 5431 4437 5440
rect 4683 5480 4725 5489
rect 4683 5440 4684 5480
rect 4724 5440 4725 5480
rect 4683 5431 4725 5440
rect 4203 5396 4245 5405
rect 4203 5356 4204 5396
rect 4244 5356 4245 5396
rect 4203 5347 4245 5356
rect 652 5144 692 5153
rect 652 4817 692 5104
rect 4204 4976 4244 5347
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4204 4927 4244 4936
rect 4395 4976 4437 4985
rect 4395 4936 4396 4976
rect 4436 4936 4437 4976
rect 4395 4927 4437 4936
rect 4492 4976 4532 4985
rect 4532 4936 4628 4976
rect 4492 4927 4532 4936
rect 4396 4842 4436 4927
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 3820 4808 3860 4817
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 3339 4220 3381 4229
rect 3339 4180 3340 4220
rect 3380 4180 3381 4220
rect 3339 4171 3381 4180
rect 3340 4136 3380 4171
rect 3340 4085 3380 4096
rect 3724 4136 3764 4145
rect 3820 4136 3860 4768
rect 4491 4808 4533 4817
rect 4491 4768 4492 4808
rect 4532 4768 4533 4808
rect 4491 4759 4533 4768
rect 4492 4674 4532 4759
rect 4588 4397 4628 4936
rect 4684 4724 4724 4733
rect 4587 4388 4629 4397
rect 4587 4348 4588 4388
rect 4628 4348 4629 4388
rect 4587 4339 4629 4348
rect 4684 4229 4724 4684
rect 4683 4220 4725 4229
rect 4683 4180 4684 4220
rect 4724 4180 4725 4220
rect 4683 4171 4725 4180
rect 4972 4145 5012 6448
rect 5643 6404 5685 6413
rect 5643 6364 5644 6404
rect 5684 6364 5685 6404
rect 5643 6355 5685 6364
rect 5547 5816 5589 5825
rect 5547 5776 5548 5816
rect 5588 5776 5589 5816
rect 5547 5767 5589 5776
rect 5548 5648 5588 5767
rect 5548 5599 5588 5608
rect 5356 4976 5396 4985
rect 5356 4817 5396 4936
rect 5355 4808 5397 4817
rect 5355 4768 5356 4808
rect 5396 4768 5397 4808
rect 5644 4808 5684 6355
rect 5740 5900 5780 7960
rect 5836 8000 5876 8009
rect 5836 7589 5876 7960
rect 5932 8000 5972 8009
rect 5972 7960 6068 8000
rect 5932 7951 5972 7960
rect 5931 7832 5973 7841
rect 5931 7792 5932 7832
rect 5972 7792 5973 7832
rect 6028 7832 6068 7960
rect 6124 7941 6164 7950
rect 6220 7925 6260 8623
rect 6219 7916 6261 7925
rect 6164 7901 6220 7916
rect 6124 7876 6220 7901
rect 6260 7876 6261 7916
rect 6219 7867 6261 7876
rect 6316 7841 6356 8632
rect 6700 8588 6740 8597
rect 6700 8177 6740 8548
rect 6699 8168 6741 8177
rect 6699 8128 6700 8168
rect 6740 8128 6741 8168
rect 6699 8119 6741 8128
rect 6315 7832 6357 7841
rect 6028 7792 6164 7832
rect 5931 7783 5973 7792
rect 5835 7580 5877 7589
rect 5835 7540 5836 7580
rect 5876 7540 5877 7580
rect 5835 7531 5877 7540
rect 5835 7412 5877 7421
rect 5835 7372 5836 7412
rect 5876 7372 5877 7412
rect 5835 7363 5877 7372
rect 5836 7278 5876 7363
rect 5836 6992 5876 7001
rect 5836 6413 5876 6952
rect 5932 6992 5972 7783
rect 6028 6992 6068 7001
rect 5932 6952 6028 6992
rect 6124 6992 6164 7792
rect 6315 7792 6316 7832
rect 6356 7792 6357 7832
rect 6315 7783 6357 7792
rect 6796 7748 6836 7757
rect 6796 7589 6836 7708
rect 6219 7580 6261 7589
rect 6219 7540 6220 7580
rect 6260 7540 6261 7580
rect 6219 7531 6261 7540
rect 6795 7580 6837 7589
rect 6795 7540 6796 7580
rect 6836 7540 6837 7580
rect 6795 7531 6837 7540
rect 6220 7160 6260 7531
rect 6892 7412 6932 9472
rect 7084 8672 7124 9808
rect 7084 8623 7124 8632
rect 7756 8261 7796 10144
rect 7852 10135 7892 10144
rect 7947 9428 7989 9437
rect 7852 9388 7948 9428
rect 7988 9388 7989 9428
rect 7755 8252 7797 8261
rect 7755 8212 7756 8252
rect 7796 8212 7797 8252
rect 7755 8203 7797 8212
rect 7468 8000 7508 8009
rect 7371 7580 7413 7589
rect 7371 7540 7372 7580
rect 7412 7540 7413 7580
rect 7371 7531 7413 7540
rect 6988 7412 7028 7421
rect 6892 7372 6988 7412
rect 6988 7363 7028 7372
rect 6220 7111 6260 7120
rect 6507 7160 6549 7169
rect 6507 7120 6508 7160
rect 6548 7120 6549 7160
rect 6507 7111 6549 7120
rect 6508 7026 6548 7111
rect 6316 6992 6356 7001
rect 6124 6952 6316 6992
rect 5835 6404 5877 6413
rect 5835 6364 5836 6404
rect 5876 6364 5877 6404
rect 5835 6355 5877 6364
rect 5740 5860 5876 5900
rect 5836 5741 5876 5860
rect 5835 5732 5877 5741
rect 5835 5692 5836 5732
rect 5876 5692 5877 5732
rect 5835 5683 5877 5692
rect 5836 5648 5876 5683
rect 5836 5599 5876 5608
rect 5740 5480 5780 5491
rect 5740 5405 5780 5440
rect 5739 5396 5781 5405
rect 5739 5356 5740 5396
rect 5780 5356 5781 5396
rect 5739 5347 5781 5356
rect 5932 5228 5972 6952
rect 6028 6943 6068 6952
rect 6316 6833 6356 6952
rect 6315 6824 6357 6833
rect 6315 6784 6316 6824
rect 6356 6784 6357 6824
rect 6315 6775 6357 6784
rect 6219 6572 6261 6581
rect 6219 6532 6220 6572
rect 6260 6532 6261 6572
rect 6219 6523 6261 6532
rect 6220 6488 6260 6523
rect 6220 6437 6260 6448
rect 6411 6488 6453 6497
rect 6411 6439 6412 6488
rect 6452 6439 6453 6488
rect 7372 6488 7412 7531
rect 7468 7505 7508 7960
rect 7563 8000 7605 8009
rect 7563 7960 7564 8000
rect 7604 7960 7605 8000
rect 7563 7951 7605 7960
rect 7756 8000 7796 8009
rect 7564 7866 7604 7951
rect 7659 7916 7701 7925
rect 7756 7916 7796 7960
rect 7659 7876 7660 7916
rect 7700 7876 7796 7916
rect 7659 7867 7701 7876
rect 7660 7673 7700 7867
rect 7755 7748 7797 7757
rect 7755 7708 7756 7748
rect 7796 7708 7797 7748
rect 7755 7699 7797 7708
rect 7659 7664 7701 7673
rect 7659 7624 7660 7664
rect 7700 7624 7701 7664
rect 7659 7615 7701 7624
rect 7756 7614 7796 7699
rect 7467 7496 7509 7505
rect 7467 7456 7468 7496
rect 7508 7456 7509 7496
rect 7467 7447 7509 7456
rect 7467 7160 7509 7169
rect 7467 7120 7468 7160
rect 7508 7120 7509 7160
rect 7467 7111 7509 7120
rect 7852 7160 7892 9388
rect 7947 9379 7989 9388
rect 7948 9294 7988 9379
rect 7947 8672 7989 8681
rect 7947 8632 7948 8672
rect 7988 8632 7989 8672
rect 7947 8623 7989 8632
rect 7948 8538 7988 8623
rect 8044 8000 8084 11899
rect 8428 11814 8468 11899
rect 8427 11360 8469 11369
rect 8427 11320 8428 11360
rect 8468 11320 8469 11360
rect 8427 11311 8469 11320
rect 8428 11024 8468 11311
rect 8428 10975 8468 10984
rect 8523 10016 8565 10025
rect 8523 9976 8524 10016
rect 8564 9976 8565 10016
rect 8523 9967 8565 9976
rect 8524 9882 8564 9967
rect 8139 9512 8181 9521
rect 8139 9472 8140 9512
rect 8180 9472 8181 9512
rect 8139 9463 8181 9472
rect 8236 9512 8276 9521
rect 8428 9512 8468 9521
rect 8276 9472 8428 9512
rect 8236 9463 8276 9472
rect 8428 9463 8468 9472
rect 8140 9378 8180 9463
rect 8331 8252 8373 8261
rect 8331 8212 8332 8252
rect 8372 8212 8373 8252
rect 8331 8203 8373 8212
rect 8235 8168 8277 8177
rect 8235 8128 8236 8168
rect 8276 8128 8277 8168
rect 8235 8119 8277 8128
rect 8236 8034 8276 8119
rect 8044 7951 8084 7960
rect 8139 7412 8181 7421
rect 8139 7372 8140 7412
rect 8180 7372 8181 7412
rect 8139 7363 8181 7372
rect 8140 7278 8180 7363
rect 7468 7026 7508 7111
rect 7755 6824 7797 6833
rect 7755 6784 7756 6824
rect 7796 6784 7797 6824
rect 7755 6775 7797 6784
rect 7468 6488 7508 6497
rect 7372 6448 7468 6488
rect 7468 6439 7508 6448
rect 7564 6488 7604 6499
rect 6412 6353 6452 6435
rect 7564 6413 7604 6448
rect 7660 6488 7700 6497
rect 7563 6404 7605 6413
rect 7563 6364 7564 6404
rect 7604 6364 7605 6404
rect 7563 6355 7605 6364
rect 7660 6329 7700 6448
rect 7756 6488 7796 6775
rect 7852 6497 7892 7120
rect 8140 7160 8180 7169
rect 8332 7160 8372 8203
rect 8427 7496 8469 7505
rect 8427 7456 8428 7496
rect 8468 7456 8469 7496
rect 8427 7447 8469 7456
rect 8180 7120 8276 7160
rect 8140 7111 8180 7120
rect 8044 6992 8084 7001
rect 8084 6952 8180 6992
rect 8044 6943 8084 6952
rect 7756 6439 7796 6448
rect 7851 6488 7893 6497
rect 7851 6448 7852 6488
rect 7892 6448 7893 6488
rect 7851 6439 7893 6448
rect 6027 6320 6069 6329
rect 6027 6280 6028 6320
rect 6068 6280 6069 6320
rect 6027 6271 6069 6280
rect 7083 6320 7125 6329
rect 7083 6280 7084 6320
rect 7124 6280 7125 6320
rect 7083 6271 7125 6280
rect 7659 6320 7701 6329
rect 7659 6280 7660 6320
rect 7700 6280 7701 6320
rect 7659 6271 7701 6280
rect 5740 5188 5972 5228
rect 5740 4976 5780 5188
rect 5931 5060 5973 5069
rect 5931 5020 5932 5060
rect 5972 5020 5973 5060
rect 5931 5011 5973 5020
rect 5740 4927 5780 4936
rect 5836 4976 5876 4985
rect 5836 4808 5876 4936
rect 5932 4926 5972 5011
rect 6028 4976 6068 6271
rect 7084 6186 7124 6271
rect 7276 6236 7316 6245
rect 7180 6196 7276 6236
rect 6219 5900 6261 5909
rect 6219 5860 6220 5900
rect 6260 5860 6261 5900
rect 6219 5851 6261 5860
rect 6123 5648 6165 5657
rect 6123 5608 6124 5648
rect 6164 5608 6165 5648
rect 6123 5599 6165 5608
rect 6124 5514 6164 5599
rect 6123 5396 6165 5405
rect 6123 5356 6124 5396
rect 6164 5356 6165 5396
rect 6123 5347 6165 5356
rect 6028 4927 6068 4936
rect 5644 4768 5876 4808
rect 5355 4759 5397 4768
rect 6124 4640 6164 5347
rect 6220 5144 6260 5851
rect 6796 5648 6836 5657
rect 6411 5480 6453 5489
rect 6411 5440 6412 5480
rect 6452 5440 6453 5480
rect 6411 5431 6453 5440
rect 6220 5104 6356 5144
rect 6219 4976 6261 4985
rect 6219 4936 6220 4976
rect 6260 4936 6261 4976
rect 6219 4927 6261 4936
rect 6220 4842 6260 4927
rect 6316 4724 6356 5104
rect 6028 4600 6164 4640
rect 6220 4684 6356 4724
rect 5835 4220 5877 4229
rect 5835 4180 5836 4220
rect 5876 4180 5877 4220
rect 5835 4171 5877 4180
rect 3764 4096 3860 4136
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 3724 4087 3764 4096
rect 4587 4087 4629 4096
rect 4971 4136 5013 4145
rect 4971 4096 4972 4136
rect 5012 4096 5013 4136
rect 4971 4087 5013 4096
rect 5836 4136 5876 4171
rect 4588 4002 4628 4087
rect 5836 4085 5876 4096
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 652 3632 692 3641
rect 652 3137 692 3592
rect 5452 3464 5492 3473
rect 651 3128 693 3137
rect 651 3088 652 3128
rect 692 3088 693 3128
rect 651 3079 693 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 5452 2717 5492 3424
rect 5836 3464 5876 3473
rect 5836 2801 5876 3424
rect 5835 2792 5877 2801
rect 5835 2752 5836 2792
rect 5876 2752 5877 2792
rect 5835 2743 5877 2752
rect 844 2708 884 2717
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 844 1709 884 2668
rect 5451 2708 5493 2717
rect 5451 2668 5452 2708
rect 5492 2668 5493 2708
rect 5451 2659 5493 2668
rect 6028 2624 6068 4600
rect 6124 4229 6164 4248
rect 6123 4220 6165 4229
rect 6220 4220 6260 4684
rect 6123 4180 6124 4220
rect 6164 4180 6260 4220
rect 6123 4171 6165 4180
rect 6220 4136 6260 4180
rect 6315 4220 6357 4229
rect 6315 4180 6316 4220
rect 6356 4180 6357 4220
rect 6315 4171 6357 4180
rect 6220 4087 6260 4096
rect 6316 3968 6356 4171
rect 6220 3928 6356 3968
rect 6123 2708 6165 2717
rect 6123 2668 6124 2708
rect 6164 2668 6165 2708
rect 6123 2659 6165 2668
rect 6028 2575 6068 2584
rect 6124 2574 6164 2659
rect 6220 2624 6260 3928
rect 6220 2575 6260 2584
rect 6412 2624 6452 5431
rect 6796 5069 6836 5608
rect 7180 5648 7220 6196
rect 7276 6187 7316 6196
rect 7371 6236 7413 6245
rect 7371 6196 7372 6236
rect 7412 6196 7413 6236
rect 7371 6187 7413 6196
rect 7947 6236 7989 6245
rect 7947 6196 7948 6236
rect 7988 6196 7989 6236
rect 7947 6187 7989 6196
rect 7180 5489 7220 5608
rect 7276 5648 7316 5657
rect 7372 5648 7412 6187
rect 7316 5608 7412 5648
rect 7564 5776 7892 5816
rect 6988 5480 7028 5489
rect 6795 5060 6837 5069
rect 6795 5020 6796 5060
rect 6836 5020 6837 5060
rect 6795 5011 6837 5020
rect 6892 4976 6932 4985
rect 6699 4136 6741 4145
rect 6892 4136 6932 4936
rect 6988 4229 7028 5440
rect 7179 5480 7221 5489
rect 7179 5440 7180 5480
rect 7220 5440 7221 5480
rect 7179 5431 7221 5440
rect 7276 5312 7316 5608
rect 7467 5480 7509 5489
rect 7467 5440 7468 5480
rect 7508 5440 7509 5480
rect 7467 5431 7509 5440
rect 7084 5272 7316 5312
rect 6987 4220 7029 4229
rect 6987 4180 6988 4220
rect 7028 4180 7029 4220
rect 6987 4171 7029 4180
rect 7084 4145 7124 5272
rect 7179 5060 7221 5069
rect 7179 5020 7180 5060
rect 7220 5020 7221 5060
rect 7179 5011 7221 5020
rect 7180 4976 7220 5011
rect 7180 4925 7220 4936
rect 7276 4976 7316 4985
rect 7276 4388 7316 4936
rect 7180 4348 7316 4388
rect 7372 4976 7412 4985
rect 6699 4096 6700 4136
rect 6740 4096 6741 4136
rect 6699 4087 6741 4096
rect 6796 4096 6932 4136
rect 7083 4136 7125 4145
rect 7083 4096 7084 4136
rect 7124 4096 7125 4136
rect 6507 4052 6549 4061
rect 6507 4012 6508 4052
rect 6548 4012 6549 4052
rect 6507 4003 6549 4012
rect 6412 2575 6452 2584
rect 6508 2624 6548 4003
rect 6700 3464 6740 4087
rect 6700 3415 6740 3424
rect 6700 2876 6740 2885
rect 6796 2876 6836 4096
rect 7083 4087 7125 4096
rect 6892 3968 6932 3977
rect 7180 3968 7220 4348
rect 7372 4313 7412 4936
rect 7468 4976 7508 5431
rect 7371 4304 7413 4313
rect 7371 4264 7372 4304
rect 7412 4264 7413 4304
rect 7371 4255 7413 4264
rect 7276 4145 7316 4230
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 7372 4136 7412 4145
rect 7468 4136 7508 4936
rect 7564 4397 7604 5776
rect 7756 5648 7796 5657
rect 7756 5069 7796 5608
rect 7852 5648 7892 5776
rect 7948 5741 7988 6187
rect 7947 5732 7989 5741
rect 7947 5692 7948 5732
rect 7988 5692 7989 5732
rect 7947 5683 7989 5692
rect 7852 5599 7892 5608
rect 7948 5648 7988 5683
rect 8140 5648 8180 6952
rect 8236 6488 8276 7120
rect 8332 7111 8372 7120
rect 8428 7160 8468 7447
rect 8428 6917 8468 7120
rect 8619 6992 8661 7001
rect 8619 6952 8620 6992
rect 8660 6952 8661 6992
rect 8619 6943 8661 6952
rect 8427 6908 8469 6917
rect 8427 6868 8428 6908
rect 8468 6868 8469 6908
rect 8427 6859 8469 6868
rect 8620 6858 8660 6943
rect 8716 6833 8756 13756
rect 9388 13460 9428 14008
rect 9580 13998 9620 14083
rect 10540 14057 10580 15520
rect 11404 14720 11444 14729
rect 9964 14048 10004 14057
rect 10539 14048 10581 14057
rect 10004 14008 10100 14048
rect 9964 13999 10004 14008
rect 9580 13460 9620 13469
rect 9388 13420 9580 13460
rect 9580 13411 9620 13420
rect 10060 13376 10100 14008
rect 10539 14008 10540 14048
rect 10580 14008 10581 14048
rect 10539 13999 10581 14008
rect 10827 14048 10869 14057
rect 10827 14008 10828 14048
rect 10868 14008 10869 14048
rect 10827 13999 10869 14008
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 10828 13914 10868 13999
rect 10060 13327 10100 13336
rect 11212 13301 11252 13999
rect 11211 13292 11253 13301
rect 11211 13252 11212 13292
rect 11252 13252 11348 13292
rect 11211 13243 11253 13252
rect 8811 13208 8853 13217
rect 8811 13168 8812 13208
rect 8852 13168 8853 13208
rect 8811 13159 8853 13168
rect 8812 12629 8852 13159
rect 11212 13158 11252 13243
rect 8811 12620 8853 12629
rect 8811 12580 8812 12620
rect 8852 12580 8853 12620
rect 8811 12571 8853 12580
rect 9676 12620 9716 12629
rect 8812 11780 8852 12571
rect 9292 12536 9332 12545
rect 9292 11957 9332 12496
rect 9484 12536 9524 12545
rect 9291 11948 9333 11957
rect 9291 11908 9292 11948
rect 9332 11908 9333 11948
rect 9291 11899 9333 11908
rect 8812 11731 8852 11740
rect 9291 11024 9333 11033
rect 9291 10984 9292 11024
rect 9332 10984 9333 11024
rect 9291 10975 9333 10984
rect 9292 10890 9332 10975
rect 9004 10352 9044 10361
rect 9484 10352 9524 12496
rect 9580 12536 9620 12545
rect 9580 12377 9620 12496
rect 9676 12461 9716 12580
rect 9772 12536 9812 12545
rect 10636 12536 10676 12545
rect 9675 12452 9717 12461
rect 9675 12412 9676 12452
rect 9716 12412 9717 12452
rect 9675 12403 9717 12412
rect 9579 12368 9621 12377
rect 9579 12328 9580 12368
rect 9620 12328 9621 12368
rect 9579 12319 9621 12328
rect 8907 8504 8949 8513
rect 8907 8464 8908 8504
rect 8948 8464 8949 8504
rect 8907 8455 8949 8464
rect 8908 8000 8948 8455
rect 8908 7951 8948 7960
rect 8907 7748 8949 7757
rect 8907 7708 8908 7748
rect 8948 7708 8949 7748
rect 8907 7699 8949 7708
rect 8812 7160 8852 7169
rect 8715 6824 8757 6833
rect 8715 6784 8716 6824
rect 8756 6784 8757 6824
rect 8715 6775 8757 6784
rect 8331 6740 8373 6749
rect 8331 6700 8332 6740
rect 8372 6700 8373 6740
rect 8331 6691 8373 6700
rect 8236 6329 8276 6448
rect 8235 6320 8277 6329
rect 8235 6280 8236 6320
rect 8276 6280 8277 6320
rect 8235 6271 8277 6280
rect 8236 5900 8276 5909
rect 8332 5900 8372 6691
rect 8812 6665 8852 7120
rect 8908 7160 8948 7699
rect 9004 7169 9044 10312
rect 9292 10312 9524 10352
rect 9580 11696 9620 11705
rect 9100 9512 9140 9523
rect 9100 9437 9140 9472
rect 9292 9512 9332 10312
rect 9483 10184 9525 10193
rect 9483 10144 9484 10184
rect 9524 10144 9525 10184
rect 9580 10184 9620 11656
rect 9772 11285 9812 12496
rect 10252 12496 10636 12536
rect 9964 12284 10004 12293
rect 9771 11276 9813 11285
rect 9771 11236 9772 11276
rect 9812 11236 9813 11276
rect 9771 11227 9813 11236
rect 9676 11108 9716 11117
rect 9964 11108 10004 12244
rect 10059 11696 10101 11705
rect 10059 11656 10060 11696
rect 10100 11656 10101 11696
rect 10059 11647 10101 11656
rect 10060 11562 10100 11647
rect 9716 11068 10004 11108
rect 9676 11059 9716 11068
rect 10060 11024 10100 11033
rect 10060 10520 10100 10984
rect 9868 10480 10100 10520
rect 10156 11024 10196 11033
rect 9675 10184 9717 10193
rect 9580 10144 9676 10184
rect 9716 10144 9717 10184
rect 9483 10135 9525 10144
rect 9675 10135 9717 10144
rect 9484 9680 9524 10135
rect 9676 10050 9716 10135
rect 9484 9631 9524 9640
rect 9292 9437 9332 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9868 9512 9908 10480
rect 10156 10445 10196 10984
rect 10155 10436 10197 10445
rect 10155 10396 10156 10436
rect 10196 10396 10197 10436
rect 10155 10387 10197 10396
rect 9963 10352 10005 10361
rect 9963 10312 9964 10352
rect 10004 10312 10005 10352
rect 9963 10303 10005 10312
rect 9964 10218 10004 10303
rect 10252 10268 10292 12496
rect 10636 12487 10676 12496
rect 10828 12368 10868 12377
rect 10444 11696 10484 11705
rect 10828 11696 10868 12328
rect 10484 11656 10868 11696
rect 11308 11696 11348 13252
rect 11404 12629 11444 14680
rect 11788 14552 11828 14561
rect 11788 14057 11828 14512
rect 11787 14048 11829 14057
rect 11787 14008 11788 14048
rect 11828 14008 11829 14048
rect 11787 13999 11829 14008
rect 11595 13880 11637 13889
rect 11595 13840 11596 13880
rect 11636 13840 11637 13880
rect 11595 13831 11637 13840
rect 11979 13880 12021 13889
rect 11979 13840 11980 13880
rect 12020 13840 12021 13880
rect 11979 13831 12021 13840
rect 11403 12620 11445 12629
rect 11403 12580 11404 12620
rect 11444 12580 11445 12620
rect 11403 12571 11445 12580
rect 11596 12452 11636 13831
rect 11980 13746 12020 13831
rect 12172 13796 12212 13805
rect 12212 13756 12500 13796
rect 12172 13747 12212 13756
rect 12268 13376 12308 13387
rect 12268 13301 12308 13336
rect 12267 13292 12309 13301
rect 12267 13252 12268 13292
rect 12308 13252 12309 13292
rect 12267 13243 12309 13252
rect 12460 13208 12500 13756
rect 12460 13159 12500 13168
rect 11596 12403 11636 12412
rect 12076 13040 12116 13049
rect 11787 12284 11829 12293
rect 11787 12244 11788 12284
rect 11828 12244 11829 12284
rect 11787 12235 11829 12244
rect 11980 12284 12020 12293
rect 11788 12150 11828 12235
rect 11980 11705 12020 12244
rect 10444 11647 10484 11656
rect 11308 11360 11348 11656
rect 11979 11696 12021 11705
rect 11979 11656 11980 11696
rect 12020 11656 12021 11696
rect 11979 11647 12021 11656
rect 11116 11320 11348 11360
rect 10348 11033 10388 11118
rect 10347 11024 10389 11033
rect 10347 10984 10348 11024
rect 10388 10984 10389 11024
rect 10347 10975 10389 10984
rect 10540 11024 10580 11033
rect 10348 10856 10388 10865
rect 10540 10856 10580 10984
rect 11019 11024 11061 11033
rect 11019 10984 11020 11024
rect 11060 10984 11061 11024
rect 11019 10975 11061 10984
rect 10388 10816 10580 10856
rect 10348 10807 10388 10816
rect 10060 10228 10292 10268
rect 10060 9680 10100 10228
rect 10155 10100 10197 10109
rect 10155 10060 10156 10100
rect 10196 10060 10197 10100
rect 10155 10051 10197 10060
rect 10060 9631 10100 9640
rect 9099 9428 9141 9437
rect 9099 9388 9100 9428
rect 9140 9388 9141 9428
rect 9099 9379 9141 9388
rect 9291 9428 9333 9437
rect 9291 9388 9292 9428
rect 9332 9388 9333 9428
rect 9291 9379 9333 9388
rect 9388 9378 9428 9463
rect 9580 9378 9620 9463
rect 9868 9437 9908 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10156 9512 10196 10051
rect 10347 10016 10389 10025
rect 10347 9976 10348 10016
rect 10388 9976 10389 10016
rect 10347 9967 10389 9976
rect 10156 9463 10196 9472
rect 10348 9512 10388 9967
rect 11020 9680 11060 10975
rect 11116 10184 11156 11320
rect 11691 11276 11733 11285
rect 11691 11236 11692 11276
rect 11732 11236 11733 11276
rect 11691 11227 11733 11236
rect 11308 11152 11540 11192
rect 11211 10772 11253 10781
rect 11211 10732 11212 10772
rect 11252 10732 11253 10772
rect 11211 10723 11253 10732
rect 11212 10638 11252 10723
rect 11308 10520 11348 11152
rect 11116 10135 11156 10144
rect 11212 10480 11348 10520
rect 11404 11024 11444 11033
rect 11212 10016 11252 10480
rect 11307 10352 11349 10361
rect 11307 10312 11308 10352
rect 11348 10312 11349 10352
rect 11307 10303 11349 10312
rect 11020 9631 11060 9640
rect 11116 9976 11252 10016
rect 10348 9463 10388 9472
rect 10443 9512 10485 9521
rect 10443 9472 10444 9512
rect 10484 9472 10485 9512
rect 10443 9463 10485 9472
rect 11116 9512 11156 9976
rect 11308 9848 11348 10303
rect 11404 10109 11444 10984
rect 11500 11024 11540 11152
rect 11500 10975 11540 10984
rect 11596 11024 11636 11033
rect 11499 10856 11541 10865
rect 11499 10816 11500 10856
rect 11540 10816 11541 10856
rect 11499 10807 11541 10816
rect 11403 10100 11445 10109
rect 11403 10060 11404 10100
rect 11444 10060 11445 10100
rect 11403 10051 11445 10060
rect 11308 9808 11444 9848
rect 11307 9680 11349 9689
rect 11307 9640 11308 9680
rect 11348 9640 11349 9680
rect 11307 9631 11349 9640
rect 9867 9428 9909 9437
rect 9867 9388 9868 9428
rect 9908 9388 9909 9428
rect 9867 9379 9909 9388
rect 9868 8933 9908 9379
rect 9964 9378 10004 9463
rect 10444 9378 10484 9463
rect 11116 9437 11156 9472
rect 11211 9512 11253 9521
rect 11211 9472 11212 9512
rect 11252 9472 11253 9512
rect 11211 9463 11253 9472
rect 11308 9512 11348 9631
rect 11308 9463 11348 9472
rect 11115 9428 11157 9437
rect 11115 9388 11116 9428
rect 11156 9388 11157 9428
rect 11115 9379 11157 9388
rect 11019 9260 11061 9269
rect 11019 9220 11020 9260
rect 11060 9220 11061 9260
rect 11019 9211 11061 9220
rect 9867 8924 9909 8933
rect 9867 8884 9868 8924
rect 9908 8884 9909 8924
rect 9867 8875 9909 8884
rect 10347 8924 10389 8933
rect 10347 8884 10348 8924
rect 10388 8884 10389 8924
rect 10347 8875 10389 8884
rect 9484 8672 9524 8681
rect 9100 8504 9140 8513
rect 9484 8504 9524 8632
rect 10348 8672 10388 8875
rect 10635 8840 10677 8849
rect 10635 8800 10636 8840
rect 10676 8800 10677 8840
rect 10635 8791 10677 8800
rect 10348 8623 10388 8632
rect 10444 8672 10484 8681
rect 9140 8464 9524 8504
rect 9100 8455 9140 8464
rect 9387 8252 9429 8261
rect 9387 8212 9388 8252
rect 9428 8212 9429 8252
rect 9387 8203 9429 8212
rect 9292 8168 9332 8177
rect 9100 8000 9140 8009
rect 9100 7421 9140 7960
rect 9195 8000 9237 8009
rect 9195 7960 9196 8000
rect 9236 7960 9237 8000
rect 9195 7951 9237 7960
rect 9196 7866 9236 7951
rect 9195 7748 9237 7757
rect 9195 7708 9196 7748
rect 9236 7708 9237 7748
rect 9195 7699 9237 7708
rect 9099 7412 9141 7421
rect 9099 7372 9100 7412
rect 9140 7372 9141 7412
rect 9099 7363 9141 7372
rect 9196 7328 9236 7699
rect 9292 7412 9332 8128
rect 9388 8000 9428 8203
rect 9484 8168 9524 8464
rect 10156 8504 10196 8513
rect 9484 8128 10100 8168
rect 9388 7951 9428 7960
rect 9484 8000 9524 8009
rect 9484 7832 9524 7960
rect 9639 8000 9679 8128
rect 9639 7951 9679 7960
rect 9964 8000 10004 8009
rect 9868 7832 9908 7841
rect 9484 7792 9868 7832
rect 9868 7783 9908 7792
rect 9867 7664 9909 7673
rect 9867 7624 9868 7664
rect 9908 7624 9909 7664
rect 9867 7615 9909 7624
rect 9292 7372 9716 7412
rect 9196 7288 9337 7328
rect 8908 7111 8948 7120
rect 9003 7160 9045 7169
rect 9003 7120 9004 7160
rect 9044 7120 9045 7160
rect 9003 7111 9045 7120
rect 9100 7160 9140 7169
rect 9100 7001 9140 7120
rect 9196 7160 9236 7169
rect 9099 6992 9141 7001
rect 9099 6952 9100 6992
rect 9140 6952 9141 6992
rect 9099 6943 9141 6952
rect 9196 6824 9236 7120
rect 9297 7160 9337 7288
rect 9297 7111 9337 7120
rect 9676 7160 9716 7372
rect 9676 7111 9716 7120
rect 9772 7160 9812 7169
rect 9292 6992 9332 7001
rect 9580 6992 9620 6997
rect 9332 6988 9620 6992
rect 9332 6952 9580 6988
rect 9292 6943 9332 6952
rect 9580 6939 9620 6948
rect 9387 6824 9429 6833
rect 9196 6784 9332 6824
rect 8427 6656 8469 6665
rect 8427 6616 8428 6656
rect 8468 6616 8469 6656
rect 8427 6607 8469 6616
rect 8716 6656 8756 6665
rect 8428 6522 8468 6607
rect 8523 6488 8565 6497
rect 8523 6448 8524 6488
rect 8564 6448 8565 6488
rect 8523 6439 8565 6448
rect 8524 6354 8564 6439
rect 8276 5860 8372 5900
rect 8236 5851 8276 5860
rect 8236 5648 8276 5657
rect 8140 5608 8236 5648
rect 7948 5597 7988 5608
rect 8236 5599 8276 5608
rect 8427 5648 8469 5657
rect 8427 5608 8428 5648
rect 8468 5608 8469 5648
rect 8427 5599 8469 5608
rect 8524 5648 8564 5657
rect 8716 5648 8756 6616
rect 8811 6656 8853 6665
rect 8811 6616 8812 6656
rect 8852 6616 8853 6656
rect 8811 6607 8853 6616
rect 9292 6581 9332 6784
rect 9387 6784 9388 6824
rect 9428 6784 9429 6824
rect 9387 6775 9429 6784
rect 9291 6572 9333 6581
rect 9291 6532 9292 6572
rect 9332 6532 9333 6572
rect 9291 6523 9333 6532
rect 8908 6488 8948 6497
rect 8908 6329 8948 6448
rect 9003 6488 9045 6497
rect 9003 6448 9004 6488
rect 9044 6448 9045 6488
rect 9003 6439 9045 6448
rect 9196 6488 9236 6497
rect 9004 6354 9044 6439
rect 9196 6329 9236 6448
rect 9292 6488 9332 6523
rect 9292 6437 9332 6448
rect 9388 6404 9428 6775
rect 9772 6749 9812 7120
rect 9771 6740 9813 6749
rect 9771 6700 9772 6740
rect 9812 6700 9813 6740
rect 9771 6691 9813 6700
rect 9868 6665 9908 7615
rect 9964 7589 10004 7960
rect 9963 7580 10005 7589
rect 9963 7540 9964 7580
rect 10004 7540 10005 7580
rect 10060 7580 10100 8128
rect 10156 8000 10196 8464
rect 10156 7951 10196 7960
rect 10444 7757 10484 8632
rect 10636 8672 10676 8791
rect 10636 8623 10676 8632
rect 10731 8672 10773 8681
rect 10731 8632 10732 8672
rect 10772 8632 10773 8672
rect 10731 8623 10773 8632
rect 11020 8672 11060 9211
rect 11020 8623 11060 8632
rect 10539 8504 10581 8513
rect 10539 8464 10540 8504
rect 10580 8464 10581 8504
rect 10539 8455 10581 8464
rect 10540 8370 10580 8455
rect 10251 7748 10293 7757
rect 10251 7708 10252 7748
rect 10292 7708 10293 7748
rect 10251 7699 10293 7708
rect 10443 7748 10485 7757
rect 10443 7708 10444 7748
rect 10484 7708 10485 7748
rect 10443 7699 10485 7708
rect 10252 7614 10292 7699
rect 10732 7673 10772 8623
rect 10731 7664 10773 7673
rect 10731 7624 10732 7664
rect 10772 7624 10773 7664
rect 10731 7615 10773 7624
rect 10347 7580 10389 7589
rect 10060 7540 10196 7580
rect 9963 7531 10005 7540
rect 10060 7328 10100 7337
rect 10060 6833 10100 7288
rect 10156 7160 10196 7540
rect 10347 7540 10348 7580
rect 10388 7540 10389 7580
rect 10347 7531 10389 7540
rect 10635 7580 10677 7589
rect 10635 7540 10636 7580
rect 10676 7540 10677 7580
rect 10635 7531 10677 7540
rect 10252 7160 10292 7169
rect 10156 7120 10252 7160
rect 10252 7111 10292 7120
rect 10348 7160 10388 7531
rect 10059 6824 10101 6833
rect 10059 6784 10060 6824
rect 10100 6784 10101 6824
rect 10059 6775 10101 6784
rect 9963 6740 10005 6749
rect 9963 6700 9964 6740
rect 10004 6700 10005 6740
rect 9963 6691 10005 6700
rect 9483 6656 9525 6665
rect 9483 6616 9484 6656
rect 9524 6616 9525 6656
rect 9483 6607 9525 6616
rect 9867 6656 9909 6665
rect 9867 6616 9868 6656
rect 9908 6616 9909 6656
rect 9867 6607 9909 6616
rect 9484 6497 9524 6607
rect 9771 6572 9813 6581
rect 9771 6532 9772 6572
rect 9812 6532 9813 6572
rect 9771 6523 9813 6532
rect 9964 6572 10004 6691
rect 10348 6665 10388 7120
rect 10540 6992 10580 7001
rect 10444 6952 10540 6992
rect 10060 6656 10100 6665
rect 10347 6656 10389 6665
rect 10100 6616 10292 6656
rect 10060 6607 10100 6616
rect 9964 6523 10004 6532
rect 9483 6488 9525 6497
rect 9483 6448 9484 6488
rect 9524 6448 9525 6488
rect 9483 6439 9525 6448
rect 9772 6488 9812 6523
rect 9388 6355 9428 6364
rect 8907 6320 8949 6329
rect 8907 6280 8908 6320
rect 8948 6280 8949 6320
rect 8907 6271 8949 6280
rect 9195 6320 9237 6329
rect 9195 6280 9196 6320
rect 9236 6280 9237 6320
rect 9195 6271 9237 6280
rect 9484 6320 9524 6439
rect 9772 6437 9812 6448
rect 9868 6488 9908 6497
rect 9868 6329 9908 6448
rect 9484 6271 9524 6280
rect 9867 6320 9909 6329
rect 9867 6280 9868 6320
rect 9908 6280 9909 6320
rect 9867 6271 9909 6280
rect 9580 6236 9620 6245
rect 8564 5608 8756 5648
rect 9388 5648 9428 5657
rect 8524 5599 8564 5608
rect 8428 5514 8468 5599
rect 8044 5480 8084 5489
rect 7852 5440 8044 5480
rect 7755 5060 7797 5069
rect 7755 5020 7756 5060
rect 7796 5020 7797 5060
rect 7755 5011 7797 5020
rect 7852 4976 7892 5440
rect 8044 5431 8084 5440
rect 8716 5480 8756 5489
rect 7852 4927 7892 4936
rect 8716 4976 8756 5440
rect 8716 4927 8756 4936
rect 9100 4976 9140 4985
rect 9140 4936 9236 4976
rect 9100 4927 9140 4936
rect 7660 4724 7700 4733
rect 7563 4388 7605 4397
rect 7563 4348 7564 4388
rect 7604 4348 7605 4388
rect 7563 4339 7605 4348
rect 7564 4254 7604 4339
rect 7412 4096 7508 4136
rect 7372 4087 7412 4096
rect 7276 3968 7316 3977
rect 6932 3928 7276 3968
rect 6892 3919 6932 3928
rect 6740 2836 6836 2876
rect 6700 2827 6740 2836
rect 6891 2792 6933 2801
rect 6891 2752 6892 2792
rect 6932 2752 6933 2792
rect 6891 2743 6933 2752
rect 6892 2658 6932 2743
rect 6508 2575 6548 2584
rect 6700 2624 6740 2633
rect 6700 2540 6740 2584
rect 6988 2540 7028 3928
rect 7276 3919 7316 3928
rect 7660 3809 7700 4684
rect 8524 4724 8564 4733
rect 8564 4684 8660 4724
rect 8524 4675 8564 4684
rect 7851 4304 7893 4313
rect 7851 4264 7852 4304
rect 7892 4264 7893 4304
rect 7851 4255 7893 4264
rect 8140 4304 8180 4313
rect 7852 4136 7892 4255
rect 8140 4145 8180 4264
rect 8523 4304 8565 4313
rect 8523 4264 8524 4304
rect 8564 4264 8565 4304
rect 8523 4255 8565 4264
rect 8139 4136 8181 4145
rect 7892 4096 8084 4136
rect 7852 4087 7892 4096
rect 7659 3800 7701 3809
rect 7659 3760 7660 3800
rect 7700 3760 7701 3800
rect 7659 3751 7701 3760
rect 7947 3800 7989 3809
rect 7947 3760 7948 3800
rect 7988 3760 7989 3800
rect 7947 3751 7989 3760
rect 7851 3380 7893 3389
rect 7851 3340 7852 3380
rect 7892 3340 7893 3380
rect 7851 3331 7893 3340
rect 7852 3246 7892 3331
rect 7948 2624 7988 3751
rect 8044 3632 8084 4096
rect 8139 4096 8140 4136
rect 8180 4096 8181 4136
rect 8139 4087 8181 4096
rect 8044 3583 8084 3592
rect 8235 2792 8277 2801
rect 8235 2752 8236 2792
rect 8276 2752 8277 2792
rect 8235 2743 8277 2752
rect 8044 2633 8084 2718
rect 8043 2624 8085 2633
rect 7948 2584 8044 2624
rect 8084 2584 8085 2624
rect 8043 2575 8085 2584
rect 8140 2624 8180 2633
rect 6700 2500 7028 2540
rect 8140 2465 8180 2584
rect 8236 2624 8276 2743
rect 8428 2633 8468 2718
rect 8524 2708 8564 4255
rect 8524 2659 8564 2668
rect 8236 2575 8276 2584
rect 8427 2624 8469 2633
rect 8427 2584 8428 2624
rect 8468 2584 8469 2624
rect 8427 2575 8469 2584
rect 8620 2624 8660 4684
rect 9196 4304 9236 4936
rect 9388 4313 9428 5608
rect 9580 5153 9620 6196
rect 10060 6236 10100 6245
rect 10060 5741 10100 6196
rect 10059 5732 10101 5741
rect 10059 5692 10060 5732
rect 10100 5692 10101 5732
rect 10059 5683 10101 5692
rect 9676 5480 9716 5489
rect 9579 5144 9621 5153
rect 9579 5104 9580 5144
rect 9620 5104 9621 5144
rect 9579 5095 9621 5104
rect 9676 5069 9716 5440
rect 9675 5060 9717 5069
rect 9675 5020 9676 5060
rect 9716 5020 9717 5060
rect 9675 5011 9717 5020
rect 9963 4976 10005 4985
rect 9963 4936 9964 4976
rect 10004 4936 10005 4976
rect 9963 4927 10005 4936
rect 9964 4842 10004 4927
rect 9196 4255 9236 4264
rect 9387 4304 9429 4313
rect 9387 4264 9388 4304
rect 9428 4264 9429 4304
rect 9387 4255 9429 4264
rect 9676 4145 9716 4230
rect 10252 4145 10292 6616
rect 10347 6616 10348 6656
rect 10388 6616 10389 6656
rect 10347 6607 10389 6616
rect 10348 6488 10388 6497
rect 10348 6329 10388 6448
rect 10347 6320 10389 6329
rect 10347 6280 10348 6320
rect 10388 6280 10389 6320
rect 10347 6271 10389 6280
rect 10444 5657 10484 6952
rect 10540 6943 10580 6952
rect 10539 6488 10581 6497
rect 10539 6448 10540 6488
rect 10580 6448 10581 6488
rect 10539 6439 10581 6448
rect 10636 6488 10676 7531
rect 10732 7244 10772 7615
rect 10732 7195 10772 7204
rect 10923 7160 10965 7169
rect 10923 7120 10924 7160
rect 10964 7120 10965 7160
rect 10923 7111 10965 7120
rect 10540 6354 10580 6439
rect 10636 6245 10676 6448
rect 10924 6488 10964 7111
rect 10924 6439 10964 6448
rect 11116 6320 11156 9379
rect 11212 9378 11252 9463
rect 11404 8840 11444 9808
rect 11500 9680 11540 10807
rect 11596 9680 11636 10984
rect 11692 11024 11732 11227
rect 11692 10975 11732 10984
rect 11884 10856 11924 10865
rect 11884 10184 11924 10816
rect 11980 10184 12020 10193
rect 11884 10144 11980 10184
rect 11980 10135 12020 10144
rect 11787 10100 11829 10109
rect 11787 10060 11788 10100
rect 11828 10060 11829 10100
rect 11787 10051 11829 10060
rect 11596 9640 11732 9680
rect 11500 9631 11540 9640
rect 11596 9512 11636 9523
rect 11692 9521 11732 9640
rect 11596 9437 11636 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 11788 9512 11828 10051
rect 12076 9689 12116 13000
rect 12652 12536 12692 12545
rect 12652 11957 12692 12496
rect 12651 11948 12693 11957
rect 12651 11908 12652 11948
rect 12692 11908 12693 11948
rect 12651 11899 12693 11908
rect 12459 11696 12501 11705
rect 12459 11656 12460 11696
rect 12500 11656 12501 11696
rect 12459 11647 12501 11656
rect 12460 11528 12500 11647
rect 12460 11024 12500 11488
rect 12460 10975 12500 10984
rect 12652 11024 12692 11033
rect 12363 10772 12405 10781
rect 12363 10732 12364 10772
rect 12404 10732 12405 10772
rect 12363 10723 12405 10732
rect 12364 10184 12404 10723
rect 12555 10352 12597 10361
rect 12555 10312 12556 10352
rect 12596 10312 12597 10352
rect 12555 10303 12597 10312
rect 12364 10135 12404 10144
rect 12556 10184 12596 10303
rect 12652 10277 12692 10984
rect 12651 10268 12693 10277
rect 12651 10228 12652 10268
rect 12692 10228 12693 10268
rect 12651 10219 12693 10228
rect 12556 10135 12596 10144
rect 12075 9680 12117 9689
rect 12075 9640 12076 9680
rect 12116 9640 12117 9680
rect 12075 9631 12117 9640
rect 11788 9463 11828 9472
rect 12652 9512 12692 9521
rect 11595 9428 11637 9437
rect 11595 9388 11596 9428
rect 11636 9388 11637 9428
rect 11595 9379 11637 9388
rect 11692 8933 11732 9463
rect 12652 9353 12692 9472
rect 12651 9344 12693 9353
rect 12651 9304 12652 9344
rect 12692 9304 12693 9344
rect 12651 9295 12693 9304
rect 11979 9260 12021 9269
rect 11979 9220 11980 9260
rect 12020 9220 12021 9260
rect 11979 9211 12021 9220
rect 11980 9126 12020 9211
rect 11691 8924 11733 8933
rect 11691 8884 11692 8924
rect 11732 8884 11733 8924
rect 11691 8875 11733 8884
rect 11404 8800 11540 8840
rect 11404 8672 11444 8681
rect 11404 7832 11444 8632
rect 11404 7783 11444 7792
rect 11211 7664 11253 7673
rect 11500 7664 11540 8800
rect 11692 8000 11732 8875
rect 12748 8840 12788 16183
rect 12940 15560 12980 16771
rect 13036 16400 13076 16409
rect 13036 15560 13076 16360
rect 13227 16232 13269 16241
rect 13227 16192 13228 16232
rect 13268 16192 13269 16232
rect 13227 16183 13269 16192
rect 14092 16232 14132 17611
rect 14092 16183 14132 16192
rect 13228 16098 13268 16183
rect 13324 15560 13364 15569
rect 13036 15520 13324 15560
rect 12940 15511 12980 15520
rect 13324 15511 13364 15520
rect 14188 15560 14228 17695
rect 14668 17669 14708 20803
rect 15052 20600 15092 20980
rect 15148 20777 15188 20862
rect 15147 20768 15189 20777
rect 15147 20728 15148 20768
rect 15188 20728 15189 20768
rect 15147 20719 15189 20728
rect 15340 20768 15380 20777
rect 15340 20693 15380 20728
rect 15436 20768 15476 20777
rect 15339 20684 15381 20693
rect 15339 20644 15340 20684
rect 15380 20644 15381 20684
rect 15339 20635 15381 20644
rect 15244 20600 15284 20609
rect 15052 20560 15188 20600
rect 14764 19844 14804 19853
rect 14804 19804 15092 19844
rect 14764 19795 14804 19804
rect 14859 19508 14901 19517
rect 14859 19468 14860 19508
rect 14900 19468 14901 19508
rect 14859 19459 14901 19468
rect 14860 19374 14900 19459
rect 15052 19256 15092 19804
rect 15148 19517 15188 20560
rect 15244 20357 15284 20560
rect 15243 20348 15285 20357
rect 15243 20308 15244 20348
rect 15284 20308 15285 20348
rect 15243 20299 15285 20308
rect 15147 19508 15189 19517
rect 15147 19468 15148 19508
rect 15188 19468 15189 19508
rect 15147 19459 15189 19468
rect 15052 19207 15092 19216
rect 14955 18752 14997 18761
rect 14955 18712 14956 18752
rect 14996 18712 14997 18752
rect 14955 18703 14997 18712
rect 14956 18618 14996 18703
rect 15051 18584 15093 18593
rect 15051 18544 15052 18584
rect 15092 18544 15093 18584
rect 15051 18535 15093 18544
rect 15148 18584 15188 19459
rect 14955 18500 14997 18509
rect 14955 18460 14956 18500
rect 14996 18460 14997 18500
rect 14955 18451 14997 18460
rect 14956 17996 14996 18451
rect 15052 18450 15092 18535
rect 15148 18416 15188 18544
rect 15244 18584 15284 18593
rect 15340 18584 15380 20635
rect 15436 20609 15476 20728
rect 15435 20600 15477 20609
rect 15435 20560 15436 20600
rect 15476 20560 15477 20600
rect 15435 20551 15477 20560
rect 15532 20180 15572 20980
rect 16108 20936 16148 20945
rect 15627 20768 15669 20777
rect 15627 20728 15628 20768
rect 15668 20728 15669 20768
rect 15627 20719 15669 20728
rect 15724 20768 15764 20777
rect 15628 20634 15668 20719
rect 15628 20180 15668 20189
rect 15532 20140 15628 20180
rect 15628 20131 15668 20140
rect 15435 20096 15477 20105
rect 15435 20056 15436 20096
rect 15476 20056 15477 20096
rect 15435 20047 15477 20056
rect 15436 19962 15476 20047
rect 15724 19433 15764 20728
rect 15820 20768 15860 20777
rect 15820 20105 15860 20728
rect 15916 20768 15956 20779
rect 15916 20693 15956 20728
rect 15915 20684 15957 20693
rect 15915 20644 15916 20684
rect 15956 20644 15957 20684
rect 15915 20635 15957 20644
rect 15819 20096 15861 20105
rect 15819 20056 15820 20096
rect 15860 20056 15861 20096
rect 15819 20047 15861 20056
rect 15723 19424 15765 19433
rect 15723 19384 15724 19424
rect 15764 19384 15765 19424
rect 15723 19375 15765 19384
rect 15436 19256 15476 19265
rect 16108 19256 16148 20896
rect 15476 19216 16148 19256
rect 16204 19256 16244 22231
rect 16396 21776 16436 23500
rect 16971 23500 16972 23540
rect 17012 23500 17013 23540
rect 16971 23491 17013 23500
rect 17356 23204 17396 23575
rect 17356 23155 17396 23164
rect 17452 23129 17492 24592
rect 17548 24632 17588 24641
rect 17548 23885 17588 24592
rect 17644 24557 17684 25264
rect 17739 25304 17781 25313
rect 17739 25264 17740 25304
rect 17780 25264 17781 25304
rect 17739 25255 17781 25264
rect 17932 25304 17972 25339
rect 17740 25170 17780 25255
rect 17932 25254 17972 25264
rect 18220 25229 18260 25348
rect 18027 25220 18069 25229
rect 18027 25180 18028 25220
rect 18068 25180 18069 25220
rect 18027 25171 18069 25180
rect 18219 25220 18261 25229
rect 18219 25180 18220 25220
rect 18260 25180 18261 25220
rect 18219 25171 18261 25180
rect 17835 25136 17877 25145
rect 17835 25096 17836 25136
rect 17876 25096 17877 25136
rect 17835 25087 17877 25096
rect 17836 24641 17876 25087
rect 17835 24632 17877 24641
rect 17835 24592 17836 24632
rect 17876 24592 17877 24632
rect 17835 24583 17877 24592
rect 17643 24548 17685 24557
rect 17643 24508 17644 24548
rect 17684 24508 17685 24548
rect 17643 24499 17685 24508
rect 17836 24498 17876 24583
rect 17932 23960 17972 23969
rect 17836 23920 17932 23960
rect 17547 23876 17589 23885
rect 17547 23836 17548 23876
rect 17588 23836 17589 23876
rect 17547 23827 17589 23836
rect 17739 23624 17781 23633
rect 17739 23584 17740 23624
rect 17780 23584 17781 23624
rect 17739 23575 17781 23584
rect 17740 23490 17780 23575
rect 17451 23120 17493 23129
rect 17451 23080 17452 23120
rect 17492 23080 17493 23120
rect 17451 23071 17493 23080
rect 17740 23120 17780 23129
rect 17836 23120 17876 23920
rect 17932 23911 17972 23920
rect 18028 23792 18068 25171
rect 18507 25136 18549 25145
rect 18507 25096 18508 25136
rect 18548 25096 18549 25136
rect 18507 25087 18549 25096
rect 18508 24464 18548 25087
rect 18604 24632 18644 24641
rect 18700 24632 18740 26104
rect 18796 26144 18836 26153
rect 18796 26069 18836 26104
rect 18892 26144 18932 26683
rect 18892 26095 18932 26104
rect 18988 26144 19028 27355
rect 19083 26732 19125 26741
rect 19083 26692 19084 26732
rect 19124 26692 19125 26732
rect 19083 26683 19125 26692
rect 18795 26060 18837 26069
rect 18795 26020 18796 26060
rect 18836 26020 18837 26060
rect 18795 26011 18837 26020
rect 18796 25397 18836 26011
rect 18795 25388 18837 25397
rect 18795 25348 18796 25388
rect 18836 25348 18837 25388
rect 18795 25339 18837 25348
rect 18988 25220 19028 26104
rect 19084 25733 19124 26683
rect 19180 26144 19220 27364
rect 19371 27355 19413 27364
rect 19372 27270 19412 27355
rect 20236 27245 20276 27616
rect 20332 27616 20524 27656
rect 20235 27236 20277 27245
rect 20235 27196 20236 27236
rect 20276 27196 20277 27236
rect 20235 27187 20277 27196
rect 19276 26984 19316 26993
rect 19276 26825 19316 26944
rect 19275 26816 19317 26825
rect 19275 26776 19276 26816
rect 19316 26776 19317 26816
rect 19275 26767 19317 26776
rect 19659 26816 19701 26825
rect 19659 26776 19660 26816
rect 19700 26776 19701 26816
rect 19659 26767 19701 26776
rect 19948 26816 19988 26825
rect 20236 26816 20276 27187
rect 19988 26776 20276 26816
rect 19948 26767 19988 26776
rect 19564 26732 19604 26741
rect 19372 26692 19564 26732
rect 19275 26480 19317 26489
rect 19275 26440 19276 26480
rect 19316 26440 19317 26480
rect 19275 26431 19317 26440
rect 19276 26237 19316 26431
rect 19372 26321 19412 26692
rect 19564 26683 19604 26692
rect 19660 26682 19700 26767
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 19371 26312 19413 26321
rect 19371 26272 19372 26312
rect 19412 26272 19413 26312
rect 19371 26263 19413 26272
rect 19275 26228 19317 26237
rect 19275 26188 19276 26228
rect 19316 26188 19317 26228
rect 19275 26179 19317 26188
rect 19180 26095 19220 26104
rect 19276 26144 19316 26179
rect 19276 26094 19316 26104
rect 19372 26102 19412 26155
rect 20332 26153 20372 27616
rect 20524 27607 20564 27616
rect 20716 27656 20756 27952
rect 20716 27607 20756 27616
rect 20812 27656 20852 27665
rect 20908 27656 20948 28120
rect 21004 28110 21044 28195
rect 21004 27656 21044 27665
rect 20908 27616 21004 27656
rect 20619 27572 20661 27581
rect 20619 27532 20620 27572
rect 20660 27532 20661 27572
rect 20619 27523 20661 27532
rect 20524 27404 20564 27413
rect 20428 26816 20468 26825
rect 20524 26816 20564 27364
rect 20468 26776 20564 26816
rect 20428 26767 20468 26776
rect 20620 26732 20660 27523
rect 20524 26692 20660 26732
rect 19371 26062 19372 26069
rect 19467 26144 19509 26153
rect 19467 26104 19468 26144
rect 19508 26104 19509 26144
rect 19467 26095 19509 26104
rect 19660 26144 19700 26153
rect 19412 26062 19413 26069
rect 19371 26060 19413 26062
rect 19371 26020 19372 26060
rect 19412 26020 19413 26060
rect 19371 26011 19413 26020
rect 19468 26010 19508 26095
rect 19083 25724 19125 25733
rect 19083 25684 19084 25724
rect 19124 25684 19125 25724
rect 19083 25675 19125 25684
rect 19371 25724 19413 25733
rect 19371 25684 19372 25724
rect 19412 25684 19413 25724
rect 19371 25675 19413 25684
rect 19372 25556 19412 25675
rect 19372 25507 19412 25516
rect 19371 25388 19413 25397
rect 19371 25348 19372 25388
rect 19412 25348 19413 25388
rect 19371 25339 19413 25348
rect 18644 24592 18740 24632
rect 18796 25180 19028 25220
rect 19180 25304 19220 25313
rect 18796 24632 18836 25180
rect 19084 25136 19124 25145
rect 18604 24583 18644 24592
rect 18604 24464 18644 24473
rect 18508 24424 18604 24464
rect 18796 24464 18836 24592
rect 18892 25096 19084 25136
rect 18892 24632 18932 25096
rect 19084 25087 19124 25096
rect 19084 24800 19124 24809
rect 19180 24800 19220 25264
rect 19124 24760 19220 24800
rect 19084 24751 19124 24760
rect 19372 24632 19412 25339
rect 19660 25145 19700 26104
rect 20331 26144 20373 26153
rect 20331 26104 20332 26144
rect 20372 26104 20373 26144
rect 20331 26095 20373 26104
rect 20524 26144 20564 26692
rect 20620 26312 20660 26321
rect 20812 26312 20852 27616
rect 21004 27607 21044 27616
rect 21003 27488 21045 27497
rect 21003 27448 21004 27488
rect 21044 27448 21045 27488
rect 21003 27439 21045 27448
rect 21004 27354 21044 27439
rect 21100 27068 21140 28288
rect 21196 27656 21236 27665
rect 21196 27413 21236 27616
rect 21292 27656 21332 27665
rect 21484 27656 21524 27665
rect 21332 27616 21484 27656
rect 21292 27607 21332 27616
rect 21484 27607 21524 27616
rect 21580 27656 21620 27665
rect 21195 27404 21237 27413
rect 21195 27364 21196 27404
rect 21236 27364 21237 27404
rect 21195 27355 21237 27364
rect 21292 27068 21332 27077
rect 21100 27028 21292 27068
rect 21292 27019 21332 27028
rect 20660 26272 20852 26312
rect 21100 26648 21140 26657
rect 20620 26263 20660 26272
rect 21100 26237 21140 26608
rect 20907 26228 20949 26237
rect 20907 26188 20908 26228
rect 20948 26188 20949 26228
rect 20907 26179 20949 26188
rect 21099 26228 21141 26237
rect 21099 26188 21100 26228
rect 21140 26188 21141 26228
rect 21099 26179 21141 26188
rect 20524 26095 20564 26104
rect 20908 26144 20948 26179
rect 20908 26093 20948 26104
rect 20331 25892 20373 25901
rect 20331 25852 20332 25892
rect 20372 25852 20373 25892
rect 20331 25843 20373 25852
rect 20332 25758 20372 25843
rect 20523 25304 20565 25313
rect 20523 25264 20524 25304
rect 20564 25264 20565 25304
rect 20523 25255 20565 25264
rect 21388 25304 21428 25313
rect 20524 25170 20564 25255
rect 19659 25136 19701 25145
rect 19659 25096 19660 25136
rect 19700 25096 19701 25136
rect 19659 25087 19701 25096
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 18892 24583 18932 24592
rect 19276 24592 19412 24632
rect 19564 24760 19988 24800
rect 18796 24424 19124 24464
rect 18604 24415 18644 24424
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 19084 23969 19124 24424
rect 19179 24044 19221 24053
rect 19179 24004 19180 24044
rect 19220 24004 19221 24044
rect 19179 23995 19221 24004
rect 19083 23960 19125 23969
rect 19083 23920 19084 23960
rect 19124 23920 19125 23960
rect 19083 23911 19125 23920
rect 17780 23080 17876 23120
rect 17932 23752 18068 23792
rect 19084 23792 19124 23911
rect 17740 23071 17780 23080
rect 16972 22868 17012 22877
rect 16972 22541 17012 22828
rect 16971 22532 17013 22541
rect 16971 22492 16972 22532
rect 17012 22492 17013 22532
rect 16971 22483 17013 22492
rect 17643 22448 17685 22457
rect 17643 22408 17644 22448
rect 17684 22408 17685 22448
rect 17643 22399 17685 22408
rect 17164 22280 17204 22289
rect 16972 22240 17164 22280
rect 16779 22112 16821 22121
rect 16779 22072 16780 22112
rect 16820 22072 16821 22112
rect 16779 22063 16821 22072
rect 16780 21978 16820 22063
rect 16492 21776 16532 21785
rect 16396 21736 16492 21776
rect 16492 21727 16532 21736
rect 16875 21608 16917 21617
rect 16875 21568 16876 21608
rect 16916 21568 16917 21608
rect 16875 21559 16917 21568
rect 16876 20852 16916 21559
rect 16972 21020 17012 22240
rect 17164 22231 17204 22240
rect 17067 22112 17109 22121
rect 17067 22072 17068 22112
rect 17108 22072 17109 22112
rect 17067 22063 17109 22072
rect 16972 20971 17012 20980
rect 16780 20812 16916 20852
rect 16683 20768 16725 20777
rect 16683 20728 16684 20768
rect 16724 20728 16725 20768
rect 16683 20719 16725 20728
rect 16780 20768 16820 20812
rect 16780 20719 16820 20728
rect 16684 20634 16724 20719
rect 16876 20693 16916 20812
rect 16972 20768 17012 20777
rect 17068 20768 17108 22063
rect 17259 21692 17301 21701
rect 17259 21652 17260 21692
rect 17300 21652 17301 21692
rect 17259 21643 17301 21652
rect 17260 21558 17300 21643
rect 17644 21608 17684 22399
rect 17836 22112 17876 22121
rect 17836 21701 17876 22072
rect 17835 21692 17877 21701
rect 17835 21652 17836 21692
rect 17876 21652 17877 21692
rect 17835 21643 17877 21652
rect 17644 21559 17684 21568
rect 17259 20852 17301 20861
rect 17259 20812 17260 20852
rect 17300 20812 17301 20852
rect 17259 20803 17301 20812
rect 17012 20728 17108 20768
rect 16972 20719 17012 20728
rect 17260 20718 17300 20803
rect 16875 20684 16917 20693
rect 16875 20644 16876 20684
rect 16916 20644 16917 20684
rect 16875 20635 16917 20644
rect 16395 20600 16437 20609
rect 16395 20560 16396 20600
rect 16436 20560 16437 20600
rect 16395 20551 16437 20560
rect 16299 20096 16341 20105
rect 16299 20056 16300 20096
rect 16340 20056 16341 20096
rect 16299 20047 16341 20056
rect 16300 19517 16340 20047
rect 16299 19508 16341 19517
rect 16299 19468 16300 19508
rect 16340 19468 16341 19508
rect 16299 19459 16341 19468
rect 16299 19256 16341 19265
rect 16204 19216 16300 19256
rect 16340 19216 16341 19256
rect 15436 19207 15476 19216
rect 16299 19207 16341 19216
rect 16300 19122 16340 19207
rect 15627 19088 15669 19097
rect 15627 19048 15628 19088
rect 15668 19048 15669 19088
rect 15627 19039 15669 19048
rect 15628 18593 15668 19039
rect 16396 18752 16436 20551
rect 16683 20096 16725 20105
rect 16683 20056 16684 20096
rect 16724 20056 16725 20096
rect 16683 20047 16725 20056
rect 16684 19962 16724 20047
rect 16876 19928 16916 20635
rect 17932 20180 17972 23752
rect 19084 23743 19124 23752
rect 19180 23792 19220 23995
rect 19276 23801 19316 24592
rect 19564 24044 19604 24760
rect 19756 24632 19796 24641
rect 19564 23995 19604 24004
rect 19660 24592 19756 24632
rect 19660 23885 19700 24592
rect 19756 24583 19796 24592
rect 19948 24632 19988 24760
rect 19948 24583 19988 24592
rect 20428 24508 20852 24548
rect 19659 23876 19701 23885
rect 19659 23836 19660 23876
rect 19700 23836 19701 23876
rect 19659 23827 19701 23836
rect 20043 23876 20085 23885
rect 20043 23836 20044 23876
rect 20084 23836 20085 23876
rect 20043 23827 20085 23836
rect 19180 23743 19220 23752
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 19372 23792 19412 23801
rect 19564 23792 19604 23801
rect 19412 23752 19564 23792
rect 19372 23743 19412 23752
rect 19564 23743 19604 23752
rect 19276 23658 19316 23743
rect 19660 23633 19700 23827
rect 19755 23792 19797 23801
rect 19755 23752 19756 23792
rect 19796 23752 19797 23792
rect 19755 23743 19797 23752
rect 19852 23792 19892 23801
rect 20044 23792 20084 23827
rect 19892 23752 19988 23792
rect 19852 23743 19892 23752
rect 19756 23658 19796 23743
rect 19659 23624 19701 23633
rect 19659 23584 19660 23624
rect 19700 23584 19701 23624
rect 19659 23575 19701 23584
rect 19275 23456 19317 23465
rect 19275 23416 19276 23456
rect 19316 23416 19317 23456
rect 19275 23407 19317 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 18604 23120 18644 23129
rect 18644 23080 18740 23120
rect 18604 23071 18644 23080
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 18507 22448 18549 22457
rect 18507 22408 18508 22448
rect 18548 22408 18549 22448
rect 18507 22399 18549 22408
rect 18123 22364 18165 22373
rect 18123 22324 18124 22364
rect 18164 22324 18165 22364
rect 18123 22315 18165 22324
rect 18124 22280 18164 22315
rect 18508 22314 18548 22399
rect 18124 22229 18164 22240
rect 18219 22280 18261 22289
rect 18219 22240 18220 22280
rect 18260 22240 18261 22280
rect 18219 22231 18261 22240
rect 18316 22280 18356 22289
rect 18220 22146 18260 22231
rect 18027 22112 18069 22121
rect 18027 22072 18028 22112
rect 18068 22072 18069 22112
rect 18027 22063 18069 22072
rect 18028 21978 18068 22063
rect 18316 21617 18356 22240
rect 18315 21608 18357 21617
rect 18315 21568 18316 21608
rect 18356 21568 18357 21608
rect 18315 21559 18357 21568
rect 18508 21608 18548 21617
rect 18700 21608 18740 23080
rect 19179 22532 19221 22541
rect 19179 22492 19180 22532
rect 19220 22492 19221 22532
rect 19179 22483 19221 22492
rect 19276 22532 19316 23407
rect 19755 23288 19797 23297
rect 19755 23248 19756 23288
rect 19796 23248 19797 23288
rect 19755 23239 19797 23248
rect 19756 23154 19796 23239
rect 19371 23120 19413 23129
rect 19371 23080 19372 23120
rect 19412 23080 19413 23120
rect 19371 23071 19413 23080
rect 19276 22483 19316 22492
rect 18892 22280 18932 22291
rect 18892 22205 18932 22240
rect 19180 22280 19220 22483
rect 19180 22231 19220 22240
rect 18891 22196 18933 22205
rect 18891 22156 18892 22196
rect 18932 22156 18933 22196
rect 18891 22147 18933 22156
rect 18548 21568 18740 21608
rect 18508 21559 18548 21568
rect 18700 21449 18740 21568
rect 18988 22112 19028 22121
rect 18699 21440 18741 21449
rect 18699 21400 18700 21440
rect 18740 21400 18741 21440
rect 18699 21391 18741 21400
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 18124 20768 18164 20779
rect 18988 20777 19028 22072
rect 19372 21776 19412 23071
rect 19948 23036 19988 23752
rect 20044 23741 20084 23752
rect 20428 23792 20468 24508
rect 20812 24464 20852 24508
rect 20812 24415 20852 24424
rect 21388 24464 21428 25264
rect 21580 24800 21620 27616
rect 21676 26489 21716 29128
rect 22540 29119 22580 29128
rect 22924 29118 22964 29203
rect 23500 29000 23540 29632
rect 23212 28960 23540 29000
rect 22348 28496 22388 28505
rect 21868 27656 21908 27665
rect 21868 27497 21908 27616
rect 22252 27656 22292 27665
rect 22348 27656 22388 28456
rect 22731 28160 22773 28169
rect 22731 28120 22732 28160
rect 22772 28120 22773 28160
rect 22731 28111 22773 28120
rect 22732 28026 22772 28111
rect 22292 27616 22388 27656
rect 23116 27656 23156 27665
rect 22252 27607 22292 27616
rect 21867 27488 21909 27497
rect 21867 27448 21868 27488
rect 21908 27448 21909 27488
rect 21867 27439 21909 27448
rect 22348 26984 22388 26993
rect 21963 26816 22005 26825
rect 21963 26776 21964 26816
rect 22004 26776 22005 26816
rect 21963 26767 22005 26776
rect 21964 26682 22004 26767
rect 21675 26480 21717 26489
rect 21675 26440 21676 26480
rect 21716 26440 21717 26480
rect 21675 26431 21717 26440
rect 22059 26480 22101 26489
rect 22059 26440 22060 26480
rect 22100 26440 22101 26480
rect 22059 26431 22101 26440
rect 22060 26144 22100 26431
rect 22348 26153 22388 26944
rect 23116 26489 23156 27616
rect 23212 27245 23252 28960
rect 23404 28328 23444 28337
rect 23404 27749 23444 28288
rect 24364 28328 24404 30043
rect 25324 29840 25364 30127
rect 25324 29791 25364 29800
rect 25516 29261 25556 30640
rect 25612 30680 25652 32815
rect 25708 32789 25748 32908
rect 25996 32873 26036 33160
rect 26091 33032 26133 33041
rect 26091 32992 26092 33032
rect 26132 32992 26133 33032
rect 26091 32983 26133 32992
rect 25995 32864 26037 32873
rect 25995 32824 25996 32864
rect 26036 32824 26037 32864
rect 25995 32815 26037 32824
rect 26092 32864 26132 32983
rect 26187 32948 26229 32957
rect 26187 32908 26188 32948
rect 26228 32908 26229 32948
rect 26187 32899 26229 32908
rect 26859 32948 26901 32957
rect 26859 32908 26860 32948
rect 26900 32908 26901 32948
rect 26859 32899 26901 32908
rect 26092 32815 26132 32824
rect 26188 32864 26228 32899
rect 25707 32780 25749 32789
rect 25707 32740 25708 32780
rect 25748 32740 25749 32780
rect 25707 32731 25749 32740
rect 25996 32730 26036 32815
rect 26188 32813 26228 32824
rect 26380 32864 26420 32873
rect 26380 32789 26420 32824
rect 26379 32780 26421 32789
rect 26379 32740 26380 32780
rect 26420 32740 26421 32780
rect 26379 32731 26421 32740
rect 25900 32696 25940 32705
rect 25707 31352 25749 31361
rect 25707 31312 25708 31352
rect 25748 31312 25749 31352
rect 25707 31303 25749 31312
rect 25900 31352 25940 32656
rect 26380 32201 26420 32731
rect 25995 32192 26037 32201
rect 25995 32152 25996 32192
rect 26036 32152 26037 32192
rect 25995 32143 26037 32152
rect 26092 32192 26132 32201
rect 25900 31303 25940 31312
rect 25708 30689 25748 31303
rect 25996 31268 26036 32143
rect 26092 31604 26132 32152
rect 26379 32192 26421 32201
rect 26379 32152 26380 32192
rect 26420 32152 26421 32192
rect 26379 32143 26421 32152
rect 26092 31564 26324 31604
rect 25996 31219 26036 31228
rect 26092 31352 26132 31361
rect 26092 31109 26132 31312
rect 26188 31352 26228 31363
rect 26188 31277 26228 31312
rect 26187 31268 26229 31277
rect 26187 31228 26188 31268
rect 26228 31228 26229 31268
rect 26187 31219 26229 31228
rect 26091 31100 26133 31109
rect 26091 31060 26092 31100
rect 26132 31060 26133 31100
rect 26091 31051 26133 31060
rect 25612 30437 25652 30640
rect 25707 30680 25749 30689
rect 25707 30640 25708 30680
rect 25748 30640 25749 30680
rect 25707 30631 25749 30640
rect 25804 30680 25844 30689
rect 25708 30546 25748 30631
rect 25611 30428 25653 30437
rect 25611 30388 25612 30428
rect 25652 30388 25653 30428
rect 25611 30379 25653 30388
rect 25515 29252 25557 29261
rect 25515 29212 25516 29252
rect 25556 29212 25557 29252
rect 25515 29203 25557 29212
rect 25804 29177 25844 30640
rect 25996 30680 26036 30689
rect 25996 30269 26036 30640
rect 25995 30260 26037 30269
rect 25995 30220 25996 30260
rect 26036 30220 26037 30260
rect 25995 30211 26037 30220
rect 26284 30185 26324 31564
rect 26380 31361 26420 31446
rect 26379 31352 26421 31361
rect 26379 31312 26380 31352
rect 26420 31312 26421 31352
rect 26379 31303 26421 31312
rect 26860 31193 26900 32899
rect 26379 31184 26421 31193
rect 26379 31144 26380 31184
rect 26420 31144 26421 31184
rect 26379 31135 26421 31144
rect 26859 31184 26901 31193
rect 26859 31144 26860 31184
rect 26900 31144 26901 31184
rect 26859 31135 26901 31144
rect 26283 30176 26325 30185
rect 26283 30136 26284 30176
rect 26324 30136 26325 30176
rect 26283 30127 26325 30136
rect 26188 29840 26228 29849
rect 25803 29168 25845 29177
rect 25803 29128 25804 29168
rect 25844 29128 25845 29168
rect 25803 29119 25845 29128
rect 25420 29000 25460 29009
rect 26188 29000 26228 29800
rect 26283 29168 26325 29177
rect 26283 29128 26284 29168
rect 26324 29128 26325 29168
rect 26283 29119 26325 29128
rect 26380 29168 26420 31135
rect 26956 31100 26996 33403
rect 27436 33125 27476 33496
rect 27532 33832 27668 33872
rect 27435 33116 27477 33125
rect 27435 33076 27436 33116
rect 27476 33076 27477 33116
rect 27435 33067 27477 33076
rect 27532 32957 27572 33832
rect 27628 33704 27668 33715
rect 27628 33629 27668 33664
rect 27723 33704 27765 33713
rect 27723 33664 27724 33704
rect 27764 33664 27765 33704
rect 27723 33655 27765 33664
rect 27627 33620 27669 33629
rect 27627 33580 27628 33620
rect 27668 33580 27669 33620
rect 27627 33571 27669 33580
rect 27724 33368 27764 33655
rect 27819 33620 27861 33629
rect 27819 33580 27820 33620
rect 27860 33580 27861 33620
rect 27819 33571 27861 33580
rect 27628 33328 27764 33368
rect 27531 32948 27573 32957
rect 27531 32908 27532 32948
rect 27572 32908 27573 32948
rect 27531 32899 27573 32908
rect 27052 32864 27092 32873
rect 27244 32864 27284 32873
rect 27532 32864 27572 32899
rect 27092 32824 27244 32864
rect 27284 32824 27476 32864
rect 27052 32815 27092 32824
rect 27244 32815 27284 32824
rect 27340 32696 27380 32705
rect 27147 32528 27189 32537
rect 27147 32488 27148 32528
rect 27188 32488 27189 32528
rect 27147 32479 27189 32488
rect 27051 31352 27093 31361
rect 27051 31312 27052 31352
rect 27092 31312 27093 31352
rect 27051 31303 27093 31312
rect 27052 31218 27092 31303
rect 26956 31060 27092 31100
rect 26955 30680 26997 30689
rect 26955 30640 26956 30680
rect 26996 30640 26997 30680
rect 26955 30631 26997 30640
rect 26956 30546 26996 30631
rect 26475 30428 26517 30437
rect 26475 30388 26476 30428
rect 26516 30388 26517 30428
rect 26475 30379 26517 30388
rect 26380 29119 26420 29128
rect 26476 29168 26516 30379
rect 26956 30008 26996 30017
rect 26860 29968 26956 30008
rect 26571 29756 26613 29765
rect 26571 29716 26572 29756
rect 26612 29716 26613 29756
rect 26571 29707 26613 29716
rect 26572 29622 26612 29707
rect 26572 29177 26612 29262
rect 26476 29119 26516 29128
rect 26571 29168 26613 29177
rect 26764 29168 26804 29177
rect 26571 29128 26572 29168
rect 26612 29128 26613 29168
rect 26571 29119 26613 29128
rect 26668 29128 26764 29168
rect 26284 29034 26324 29119
rect 25460 28960 26228 29000
rect 25420 28951 25460 28960
rect 26475 28916 26517 28925
rect 26475 28876 26476 28916
rect 26516 28876 26517 28916
rect 26475 28867 26517 28876
rect 24364 28279 24404 28288
rect 25323 28328 25365 28337
rect 25996 28328 26036 28337
rect 25323 28288 25324 28328
rect 25364 28288 25365 28328
rect 25323 28279 25365 28288
rect 25420 28288 25996 28328
rect 25324 28194 25364 28279
rect 23403 27740 23445 27749
rect 23403 27700 23404 27740
rect 23444 27700 23445 27740
rect 23403 27691 23445 27700
rect 24267 27740 24309 27749
rect 24267 27700 24268 27740
rect 24308 27700 24309 27740
rect 24267 27691 24309 27700
rect 24459 27740 24501 27749
rect 24459 27700 24460 27740
rect 24500 27700 24501 27740
rect 24459 27691 24501 27700
rect 24268 27572 24308 27691
rect 24268 27523 24308 27532
rect 23211 27236 23253 27245
rect 23211 27196 23212 27236
rect 23252 27196 23253 27236
rect 23211 27187 23253 27196
rect 23115 26480 23157 26489
rect 23115 26440 23116 26480
rect 23156 26440 23157 26480
rect 23115 26431 23157 26440
rect 22731 26396 22773 26405
rect 22731 26356 22732 26396
rect 22772 26356 22773 26396
rect 22731 26347 22773 26356
rect 21771 25892 21813 25901
rect 21771 25852 21772 25892
rect 21812 25852 21813 25892
rect 21771 25843 21813 25852
rect 21772 25304 21812 25843
rect 22060 25313 22100 26104
rect 22347 26144 22389 26153
rect 22347 26104 22348 26144
rect 22388 26104 22389 26144
rect 22347 26095 22389 26104
rect 22732 25388 22772 26347
rect 22923 26144 22965 26153
rect 22923 26104 22924 26144
rect 22964 26104 22965 26144
rect 22923 26095 22965 26104
rect 22827 26060 22869 26069
rect 22827 26020 22828 26060
rect 22868 26020 22869 26060
rect 22827 26011 22869 26020
rect 22828 25397 22868 26011
rect 22924 26010 22964 26095
rect 22732 25339 22772 25348
rect 22827 25388 22869 25397
rect 22827 25348 22828 25388
rect 22868 25348 22869 25388
rect 22827 25339 22869 25348
rect 21772 25255 21812 25264
rect 22059 25304 22101 25313
rect 22059 25264 22060 25304
rect 22100 25264 22101 25304
rect 22059 25255 22101 25264
rect 21580 24751 21620 24760
rect 22252 24632 22292 24643
rect 22252 24557 22292 24592
rect 22443 24632 22485 24641
rect 22443 24592 22444 24632
rect 22484 24592 22485 24632
rect 22443 24583 22485 24592
rect 22251 24548 22293 24557
rect 22251 24508 22252 24548
rect 22292 24508 22293 24548
rect 22251 24499 22293 24508
rect 21388 24415 21428 24424
rect 20620 24380 20660 24389
rect 20620 23885 20660 24340
rect 22252 24044 22292 24499
rect 22444 24498 22484 24583
rect 22732 24380 22772 24389
rect 22636 24340 22732 24380
rect 22444 24044 22484 24053
rect 22252 24004 22444 24044
rect 22444 23995 22484 24004
rect 20619 23876 20661 23885
rect 20619 23836 20620 23876
rect 20660 23836 20661 23876
rect 20619 23827 20661 23836
rect 20428 23743 20468 23752
rect 21292 23792 21332 23801
rect 20619 23120 20661 23129
rect 20619 23080 20620 23120
rect 20660 23080 20661 23120
rect 20619 23071 20661 23080
rect 19948 22996 20084 23036
rect 19948 22868 19988 22877
rect 19948 22289 19988 22828
rect 20044 22532 20084 22996
rect 20620 22986 20660 23071
rect 20044 22483 20084 22492
rect 19947 22280 19989 22289
rect 19947 22240 19948 22280
rect 19988 22240 19989 22280
rect 19947 22231 19989 22240
rect 19948 22146 19988 22231
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 19660 21776 19700 21785
rect 19372 21736 19660 21776
rect 19660 21727 19700 21736
rect 21196 21608 21236 21617
rect 20235 21440 20277 21449
rect 20235 21400 20236 21440
rect 20276 21400 20277 21440
rect 20235 21391 20277 21400
rect 20236 21104 20276 21391
rect 20140 21064 20276 21104
rect 20140 20779 20180 21064
rect 18124 20693 18164 20728
rect 18987 20768 19029 20777
rect 19276 20768 19316 20777
rect 18987 20728 18988 20768
rect 19028 20728 19029 20768
rect 18987 20719 19029 20728
rect 19084 20728 19276 20768
rect 20140 20730 20180 20739
rect 20811 20768 20853 20777
rect 18123 20684 18165 20693
rect 18123 20644 18124 20684
rect 18164 20644 18165 20684
rect 18123 20635 18165 20644
rect 18892 20684 18932 20693
rect 18892 20273 18932 20644
rect 18891 20264 18933 20273
rect 18891 20224 18892 20264
rect 18932 20224 18933 20264
rect 18891 20215 18933 20224
rect 17932 20140 18068 20180
rect 16876 19879 16916 19888
rect 17451 19508 17493 19517
rect 17451 19468 17452 19508
rect 17492 19468 17493 19508
rect 17451 19459 17493 19468
rect 17452 19374 17492 19459
rect 17931 19424 17973 19433
rect 17931 19384 17932 19424
rect 17972 19384 17973 19424
rect 17931 19375 17973 19384
rect 17644 19256 17684 19265
rect 17644 19097 17684 19216
rect 17932 19256 17972 19375
rect 17932 19207 17972 19216
rect 18028 19097 18068 20140
rect 18891 20012 18933 20021
rect 18891 19972 18892 20012
rect 18932 19972 18933 20012
rect 18891 19963 18933 19972
rect 18508 19928 18548 19937
rect 18548 19888 18740 19928
rect 18508 19879 18548 19888
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 18508 19256 18548 19265
rect 18700 19256 18740 19888
rect 18548 19216 18740 19256
rect 18508 19207 18548 19216
rect 18124 19172 18164 19181
rect 17643 19088 17685 19097
rect 17643 19048 17644 19088
rect 17684 19048 17685 19088
rect 17643 19039 17685 19048
rect 17836 19088 17876 19097
rect 17836 18920 17876 19048
rect 18027 19088 18069 19097
rect 18027 19048 18028 19088
rect 18068 19048 18069 19088
rect 18027 19039 18069 19048
rect 18124 18920 18164 19132
rect 17836 18880 18164 18920
rect 16396 18703 16436 18712
rect 15284 18544 15380 18584
rect 15436 18584 15476 18593
rect 15244 18535 15284 18544
rect 15436 18416 15476 18544
rect 15627 18584 15669 18593
rect 15627 18544 15628 18584
rect 15668 18544 15669 18584
rect 15627 18535 15669 18544
rect 16108 18584 16148 18593
rect 16300 18584 16340 18593
rect 16148 18544 16300 18584
rect 16108 18535 16148 18544
rect 16300 18535 16340 18544
rect 15148 18376 15476 18416
rect 14956 17947 14996 17956
rect 14667 17660 14709 17669
rect 14667 17620 14668 17660
rect 14708 17620 14709 17660
rect 14667 17611 14709 17620
rect 15244 17072 15284 17081
rect 14379 16904 14421 16913
rect 14379 16864 14380 16904
rect 14420 16864 14421 16904
rect 14379 16855 14421 16864
rect 14380 16770 14420 16855
rect 14571 16820 14613 16829
rect 14571 16780 14572 16820
rect 14612 16780 14613 16820
rect 14571 16771 14613 16780
rect 14572 16686 14612 16771
rect 15244 16409 15284 17032
rect 15436 17072 15476 17081
rect 15436 16997 15476 17032
rect 15435 16988 15477 16997
rect 15435 16948 15436 16988
rect 15476 16948 15477 16988
rect 15435 16939 15477 16948
rect 15243 16400 15285 16409
rect 15243 16360 15244 16400
rect 15284 16360 15285 16400
rect 15243 16351 15285 16360
rect 15340 16232 15380 16241
rect 15340 15905 15380 16192
rect 15339 15896 15381 15905
rect 15339 15856 15340 15896
rect 15380 15856 15381 15896
rect 15339 15847 15381 15856
rect 15436 15728 15476 16939
rect 15628 16484 15668 18535
rect 18220 18416 18260 18425
rect 18124 18376 18220 18416
rect 15916 17744 15956 17755
rect 15916 17669 15956 17704
rect 17739 17744 17781 17753
rect 17739 17704 17740 17744
rect 17780 17704 17781 17744
rect 17739 17695 17781 17704
rect 18124 17744 18164 18376
rect 18220 18367 18260 18376
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 18124 17695 18164 17704
rect 15915 17660 15957 17669
rect 15915 17620 15916 17660
rect 15956 17620 15957 17660
rect 15915 17611 15957 17620
rect 16779 17660 16821 17669
rect 16779 17620 16780 17660
rect 16820 17620 16821 17660
rect 16779 17611 16821 17620
rect 16683 17072 16725 17081
rect 15628 16435 15668 16444
rect 16396 17032 16684 17072
rect 16724 17032 16725 17072
rect 15723 16232 15765 16241
rect 15723 16192 15724 16232
rect 15764 16192 15765 16232
rect 15723 16183 15765 16192
rect 14188 15149 14228 15520
rect 15244 15688 15476 15728
rect 14187 15140 14229 15149
rect 14187 15100 14188 15140
rect 14228 15100 14229 15140
rect 14187 15091 14229 15100
rect 15051 14888 15093 14897
rect 15051 14848 15052 14888
rect 15092 14848 15093 14888
rect 15051 14839 15093 14848
rect 13804 14720 13844 14729
rect 13708 14552 13748 14561
rect 13612 14512 13708 14552
rect 13419 14216 13461 14225
rect 13419 14176 13420 14216
rect 13460 14176 13461 14216
rect 13419 14167 13461 14176
rect 13035 14132 13077 14141
rect 13035 14092 13036 14132
rect 13076 14092 13077 14132
rect 13035 14083 13077 14092
rect 12844 14048 12884 14057
rect 12844 13889 12884 14008
rect 13036 13998 13076 14083
rect 13323 14048 13365 14057
rect 13323 14008 13324 14048
rect 13364 14008 13365 14048
rect 13323 13999 13365 14008
rect 12843 13880 12885 13889
rect 12843 13840 12844 13880
rect 12884 13840 12885 13880
rect 12843 13831 12885 13840
rect 13035 13544 13077 13553
rect 13035 13504 13036 13544
rect 13076 13504 13077 13544
rect 13035 13495 13077 13504
rect 13036 13208 13076 13495
rect 13324 13460 13364 13999
rect 13324 13411 13364 13420
rect 13036 13159 13076 13168
rect 13132 13208 13172 13219
rect 13324 13217 13364 13302
rect 13132 13133 13172 13168
rect 13323 13208 13365 13217
rect 13323 13168 13324 13208
rect 13364 13168 13365 13208
rect 13323 13159 13365 13168
rect 13131 13124 13173 13133
rect 13131 13084 13132 13124
rect 13172 13084 13173 13124
rect 13131 13075 13173 13084
rect 13227 13040 13269 13049
rect 13227 13000 13228 13040
rect 13268 13000 13269 13040
rect 13227 12991 13269 13000
rect 13228 12536 13268 12991
rect 13420 12788 13460 14167
rect 13515 14132 13557 14141
rect 13515 14092 13516 14132
rect 13556 14092 13557 14132
rect 13515 14083 13557 14092
rect 12843 11696 12885 11705
rect 12843 11656 12844 11696
rect 12884 11656 12885 11696
rect 12843 11647 12885 11656
rect 12844 11562 12884 11647
rect 13228 10856 13268 12496
rect 13324 12748 13460 12788
rect 13324 12536 13364 12748
rect 13516 12704 13556 14083
rect 13324 12487 13364 12496
rect 13420 12664 13556 12704
rect 13420 12536 13460 12664
rect 13420 12487 13460 12496
rect 13516 12536 13556 12545
rect 13612 12536 13652 14512
rect 13708 14503 13748 14512
rect 13804 14141 13844 14680
rect 13900 14720 13940 14729
rect 13900 14225 13940 14680
rect 13996 14720 14036 14729
rect 14380 14720 14420 14729
rect 14036 14680 14228 14720
rect 13996 14671 14036 14680
rect 13899 14216 13941 14225
rect 13899 14176 13900 14216
rect 13940 14176 13941 14216
rect 13899 14167 13941 14176
rect 13803 14132 13845 14141
rect 13803 14092 13804 14132
rect 13844 14092 13845 14132
rect 13803 14083 13845 14092
rect 13708 14048 13748 14057
rect 14092 14048 14132 14057
rect 13708 12704 13748 14008
rect 13900 14008 14092 14048
rect 13803 13880 13845 13889
rect 13803 13840 13804 13880
rect 13844 13840 13845 13880
rect 13803 13831 13845 13840
rect 13804 13208 13844 13831
rect 13900 13805 13940 14008
rect 14092 13999 14132 14008
rect 14188 14048 14228 14680
rect 13899 13796 13941 13805
rect 13899 13756 13900 13796
rect 13940 13756 13941 13796
rect 13899 13747 13941 13756
rect 13996 13796 14036 13805
rect 14036 13756 14132 13796
rect 13996 13747 14036 13756
rect 13804 13049 13844 13168
rect 13900 13208 13940 13747
rect 13995 13628 14037 13637
rect 13995 13588 13996 13628
rect 14036 13588 14037 13628
rect 13995 13579 14037 13588
rect 13900 13159 13940 13168
rect 13996 13124 14036 13579
rect 14092 13553 14132 13756
rect 14091 13544 14133 13553
rect 14091 13504 14092 13544
rect 14132 13504 14133 13544
rect 14091 13495 14133 13504
rect 14188 13301 14228 14008
rect 14380 13973 14420 14680
rect 14572 14720 14612 14729
rect 14476 14636 14516 14645
rect 14379 13964 14421 13973
rect 14379 13924 14380 13964
rect 14420 13924 14421 13964
rect 14379 13915 14421 13924
rect 14283 13880 14325 13889
rect 14283 13840 14284 13880
rect 14324 13840 14325 13880
rect 14283 13831 14325 13840
rect 14187 13292 14229 13301
rect 14187 13252 14188 13292
rect 14228 13252 14229 13292
rect 14187 13243 14229 13252
rect 14284 13133 14324 13831
rect 14476 13712 14516 14596
rect 14572 13805 14612 14680
rect 15052 14720 15092 14839
rect 15052 14671 15092 14680
rect 15147 14720 15189 14729
rect 15147 14680 15148 14720
rect 15188 14680 15189 14720
rect 15147 14671 15189 14680
rect 15148 14586 15188 14671
rect 14764 14057 14804 14142
rect 14668 14048 14708 14057
rect 14571 13796 14613 13805
rect 14571 13756 14572 13796
rect 14612 13756 14613 13796
rect 14571 13747 14613 13756
rect 14380 13672 14516 13712
rect 14380 13217 14420 13672
rect 14475 13544 14517 13553
rect 14475 13504 14476 13544
rect 14516 13504 14517 13544
rect 14475 13495 14517 13504
rect 14379 13208 14421 13217
rect 14379 13168 14380 13208
rect 14420 13168 14421 13208
rect 14379 13159 14421 13168
rect 14476 13208 14516 13495
rect 14668 13460 14708 14008
rect 14763 14048 14805 14057
rect 14763 14008 14764 14048
rect 14804 14008 14805 14048
rect 14763 13999 14805 14008
rect 14955 14048 14997 14057
rect 14955 14008 14956 14048
rect 14996 14008 14997 14048
rect 14955 13999 14997 14008
rect 15148 14048 15188 14057
rect 14956 13914 14996 13999
rect 15051 13880 15093 13889
rect 15148 13880 15188 14008
rect 15244 13973 15284 15688
rect 15436 15560 15476 15569
rect 15339 14552 15381 14561
rect 15339 14512 15340 14552
rect 15380 14512 15381 14552
rect 15339 14503 15381 14512
rect 15340 14418 15380 14503
rect 15340 14048 15380 14057
rect 15243 13964 15285 13973
rect 15243 13924 15244 13964
rect 15284 13924 15285 13964
rect 15243 13915 15285 13924
rect 15051 13840 15052 13880
rect 15092 13840 15188 13880
rect 15051 13831 15093 13840
rect 14764 13796 14804 13805
rect 14764 13637 14804 13756
rect 14859 13796 14901 13805
rect 15244 13796 15284 13805
rect 14859 13756 14860 13796
rect 14900 13756 14901 13796
rect 14859 13747 14901 13756
rect 15148 13756 15244 13796
rect 14763 13628 14805 13637
rect 14763 13588 14764 13628
rect 14804 13588 14805 13628
rect 14763 13579 14805 13588
rect 14764 13460 14804 13469
rect 14668 13420 14764 13460
rect 14764 13411 14804 13420
rect 14667 13292 14709 13301
rect 14667 13252 14668 13292
rect 14708 13252 14709 13292
rect 14667 13243 14709 13252
rect 14283 13124 14325 13133
rect 13996 13084 14040 13124
rect 13803 13040 13845 13049
rect 13803 13000 13804 13040
rect 13844 13000 13845 13040
rect 13803 12991 13845 13000
rect 14000 12956 14040 13084
rect 14283 13084 14284 13124
rect 14324 13084 14325 13124
rect 14283 13075 14325 13084
rect 14092 13040 14132 13049
rect 14132 13000 14228 13040
rect 14092 12991 14132 13000
rect 13996 12916 14040 12956
rect 13996 12872 14036 12916
rect 13900 12832 14036 12872
rect 14091 12872 14133 12881
rect 14091 12832 14092 12872
rect 14132 12832 14133 12872
rect 13708 12664 13844 12704
rect 13804 12620 13844 12664
rect 13804 12571 13844 12580
rect 13708 12536 13748 12545
rect 13612 12496 13708 12536
rect 13516 11696 13556 12496
rect 13708 12487 13748 12496
rect 13900 12536 13940 12832
rect 14091 12823 14133 12832
rect 13995 12620 14037 12629
rect 13995 12580 13996 12620
rect 14036 12580 14037 12620
rect 13995 12571 14037 12580
rect 13900 12487 13940 12496
rect 13996 12536 14036 12571
rect 13996 12485 14036 12496
rect 14092 12368 14132 12823
rect 14188 12545 14228 13000
rect 14284 13036 14324 13075
rect 14380 13074 14420 13159
rect 14476 13049 14516 13168
rect 14187 12536 14229 12545
rect 14187 12496 14188 12536
rect 14228 12496 14229 12536
rect 14187 12487 14229 12496
rect 13900 12328 14132 12368
rect 14188 12368 14228 12377
rect 14284 12368 14324 12996
rect 14475 13040 14517 13049
rect 14475 13000 14476 13040
rect 14516 13000 14517 13040
rect 14475 12991 14517 13000
rect 14475 12788 14517 12797
rect 14475 12748 14476 12788
rect 14516 12748 14517 12788
rect 14475 12739 14517 12748
rect 14380 12545 14420 12630
rect 14379 12536 14421 12545
rect 14379 12496 14380 12536
rect 14420 12496 14421 12536
rect 14379 12487 14421 12496
rect 14228 12328 14324 12368
rect 14380 12368 14420 12379
rect 13707 11948 13749 11957
rect 13707 11908 13708 11948
rect 13748 11908 13749 11948
rect 13707 11899 13749 11908
rect 13708 11814 13748 11899
rect 13708 11696 13748 11705
rect 13516 11656 13708 11696
rect 13708 11647 13748 11656
rect 13900 11696 13940 12328
rect 14188 12319 14228 12328
rect 14380 12293 14420 12328
rect 14379 12284 14421 12293
rect 14379 12244 14380 12284
rect 14420 12244 14421 12284
rect 14379 12235 14421 12244
rect 14476 12116 14516 12739
rect 14668 12536 14708 13243
rect 14763 12956 14805 12965
rect 14763 12916 14764 12956
rect 14804 12916 14805 12956
rect 14763 12907 14805 12916
rect 14668 12461 14708 12496
rect 14764 12536 14804 12907
rect 14860 12797 14900 13747
rect 14956 13208 14996 13217
rect 14956 12965 14996 13168
rect 15052 13208 15092 13217
rect 14955 12956 14997 12965
rect 14955 12916 14956 12956
rect 14996 12916 14997 12956
rect 14955 12907 14997 12916
rect 14859 12788 14901 12797
rect 14859 12748 14860 12788
rect 14900 12748 14901 12788
rect 14859 12739 14901 12748
rect 14955 12704 14997 12713
rect 14955 12664 14956 12704
rect 14996 12664 14997 12704
rect 14955 12655 14997 12664
rect 14956 12570 14996 12655
rect 15052 12545 15092 13168
rect 15148 12965 15188 13756
rect 15244 13747 15284 13756
rect 15244 13460 15284 13469
rect 15340 13460 15380 14008
rect 15284 13420 15380 13460
rect 15244 13411 15284 13420
rect 15436 13385 15476 15520
rect 15628 15308 15668 15317
rect 15532 15268 15628 15308
rect 15532 14048 15572 15268
rect 15628 15259 15668 15268
rect 15627 14216 15669 14225
rect 15627 14176 15628 14216
rect 15668 14176 15669 14216
rect 15724 14216 15764 16183
rect 16204 16148 16244 16157
rect 16108 16108 16204 16148
rect 16011 15560 16053 15569
rect 16011 15520 16012 15560
rect 16052 15520 16053 15560
rect 16011 15511 16053 15520
rect 15819 15476 15861 15485
rect 15819 15436 15820 15476
rect 15860 15436 15861 15476
rect 15819 15427 15861 15436
rect 15820 14720 15860 15427
rect 16012 14972 16052 15511
rect 16012 14923 16052 14932
rect 15820 14384 15860 14680
rect 15915 14720 15957 14729
rect 15915 14680 15916 14720
rect 15956 14680 15957 14720
rect 15915 14671 15957 14680
rect 15916 14586 15956 14671
rect 15820 14344 15956 14384
rect 15820 14216 15860 14225
rect 15724 14176 15820 14216
rect 15627 14167 15669 14176
rect 15820 14167 15860 14176
rect 15532 13973 15572 14008
rect 15628 14048 15668 14167
rect 15628 13999 15668 14008
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 15531 13964 15573 13973
rect 15531 13924 15532 13964
rect 15572 13924 15573 13964
rect 15531 13915 15573 13924
rect 15435 13376 15477 13385
rect 15435 13336 15436 13376
rect 15476 13336 15477 13376
rect 15435 13327 15477 13336
rect 15244 13217 15284 13302
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15436 13208 15476 13217
rect 15243 13040 15285 13049
rect 15243 13000 15244 13040
rect 15284 13000 15285 13040
rect 15243 12991 15285 13000
rect 15147 12956 15189 12965
rect 15147 12916 15148 12956
rect 15188 12916 15189 12956
rect 15147 12907 15189 12916
rect 15147 12788 15189 12797
rect 15147 12748 15148 12788
rect 15188 12748 15189 12788
rect 15147 12739 15189 12748
rect 14764 12487 14804 12496
rect 14860 12536 14900 12545
rect 14667 12452 14709 12461
rect 14667 12412 14668 12452
rect 14708 12412 14709 12452
rect 14667 12403 14709 12412
rect 14763 12368 14805 12377
rect 14763 12328 14764 12368
rect 14804 12328 14805 12368
rect 14763 12319 14805 12328
rect 14476 12076 14708 12116
rect 13995 11948 14037 11957
rect 13995 11908 13996 11948
rect 14036 11908 14037 11948
rect 13995 11899 14037 11908
rect 13900 11647 13940 11656
rect 13996 11696 14036 11899
rect 13996 11647 14036 11656
rect 14476 11696 14516 11705
rect 13515 11528 13557 11537
rect 13515 11488 13516 11528
rect 13556 11488 13557 11528
rect 13515 11479 13557 11488
rect 13899 11528 13941 11537
rect 13899 11488 13900 11528
rect 13940 11488 13941 11528
rect 13899 11479 13941 11488
rect 13516 11394 13556 11479
rect 13900 11024 13940 11479
rect 13900 10975 13940 10984
rect 13228 10807 13268 10816
rect 13611 10856 13653 10865
rect 13611 10816 13612 10856
rect 13652 10816 13653 10856
rect 14476 10856 14516 11656
rect 14572 11696 14612 11705
rect 14572 11453 14612 11656
rect 14668 11696 14708 12076
rect 14571 11444 14613 11453
rect 14571 11404 14572 11444
rect 14612 11404 14613 11444
rect 14571 11395 14613 11404
rect 14668 11360 14708 11656
rect 14764 11696 14804 12319
rect 14860 11705 14900 12496
rect 15051 12536 15093 12545
rect 15051 12496 15052 12536
rect 15092 12496 15093 12536
rect 15051 12487 15093 12496
rect 14955 12452 14997 12461
rect 14955 12412 14956 12452
rect 14996 12412 14997 12452
rect 14955 12403 14997 12412
rect 14956 11873 14996 12403
rect 15148 12368 15188 12739
rect 15148 12319 15188 12328
rect 15244 12368 15284 12991
rect 15339 12704 15381 12713
rect 15436 12704 15476 13168
rect 15531 13208 15573 13217
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 15628 13208 15668 13217
rect 15532 13074 15572 13159
rect 15628 12881 15668 13168
rect 15724 12965 15764 13999
rect 15819 13880 15861 13889
rect 15819 13840 15820 13880
rect 15860 13840 15861 13880
rect 15819 13831 15861 13840
rect 15723 12956 15765 12965
rect 15723 12916 15724 12956
rect 15764 12916 15765 12956
rect 15723 12907 15765 12916
rect 15627 12872 15669 12881
rect 15627 12832 15628 12872
rect 15668 12832 15669 12872
rect 15627 12823 15669 12832
rect 15723 12704 15765 12713
rect 15339 12664 15340 12704
rect 15380 12664 15476 12704
rect 15628 12664 15724 12704
rect 15764 12664 15765 12704
rect 15339 12655 15381 12664
rect 15628 12620 15668 12664
rect 15723 12655 15765 12664
rect 15436 12580 15668 12620
rect 15339 12536 15381 12545
rect 15339 12496 15340 12536
rect 15380 12496 15381 12536
rect 15339 12487 15381 12496
rect 15436 12536 15476 12580
rect 15723 12536 15765 12545
rect 15340 12452 15380 12487
rect 15340 12401 15380 12412
rect 15244 12319 15284 12328
rect 14955 11864 14997 11873
rect 14955 11824 14956 11864
rect 14996 11824 14997 11864
rect 14955 11815 14997 11824
rect 14764 11647 14804 11656
rect 14859 11696 14901 11705
rect 15244 11696 15284 11705
rect 14859 11656 14860 11696
rect 14900 11656 14901 11696
rect 14859 11647 14901 11656
rect 15148 11656 15244 11696
rect 14860 11360 14900 11647
rect 15148 11369 15188 11656
rect 15244 11647 15284 11656
rect 15339 11696 15381 11705
rect 15339 11656 15340 11696
rect 15380 11656 15381 11696
rect 15339 11647 15381 11656
rect 15340 11562 15380 11647
rect 15243 11528 15285 11537
rect 15243 11488 15244 11528
rect 15284 11488 15285 11528
rect 15243 11479 15285 11488
rect 15147 11360 15189 11369
rect 14668 11320 14900 11360
rect 14860 11024 14900 11320
rect 15052 11320 15148 11360
rect 15188 11320 15189 11360
rect 15052 11117 15092 11320
rect 15147 11311 15189 11320
rect 15051 11108 15093 11117
rect 15244 11108 15284 11479
rect 15339 11360 15381 11369
rect 15339 11320 15340 11360
rect 15380 11320 15381 11360
rect 15339 11311 15381 11320
rect 15051 11068 15052 11108
rect 15092 11068 15093 11108
rect 15051 11059 15093 11068
rect 15148 11068 15284 11108
rect 14860 10975 14900 10984
rect 14956 11024 14996 11033
rect 14956 10856 14996 10984
rect 14476 10816 14996 10856
rect 13611 10807 13653 10816
rect 13515 10436 13557 10445
rect 13515 10396 13516 10436
rect 13556 10396 13557 10436
rect 13515 10387 13557 10396
rect 13516 10302 13556 10387
rect 13228 10184 13268 10193
rect 13420 10184 13460 10193
rect 13268 10144 13420 10184
rect 13228 10135 13268 10144
rect 13420 10135 13460 10144
rect 13324 9680 13364 9689
rect 12844 9640 13324 9680
rect 12844 9512 12884 9640
rect 13324 9631 13364 9640
rect 13419 9680 13461 9689
rect 13419 9640 13420 9680
rect 13460 9640 13461 9680
rect 13419 9631 13461 9640
rect 12844 9463 12884 9472
rect 13036 9512 13076 9521
rect 12843 9344 12885 9353
rect 12843 9304 12844 9344
rect 12884 9304 12885 9344
rect 12843 9295 12885 9304
rect 12844 9210 12884 9295
rect 12748 8800 12884 8840
rect 12267 8672 12309 8681
rect 12267 8632 12268 8672
rect 12308 8632 12309 8672
rect 12267 8623 12309 8632
rect 12747 8672 12789 8681
rect 12747 8632 12748 8672
rect 12788 8632 12789 8672
rect 12747 8623 12789 8632
rect 12268 8538 12308 8623
rect 11788 8000 11828 8009
rect 12652 8000 12692 8009
rect 11692 7960 11788 8000
rect 11788 7951 11828 7960
rect 12556 7960 12652 8000
rect 11211 7624 11212 7664
rect 11252 7624 11253 7664
rect 11211 7615 11253 7624
rect 11404 7624 11540 7664
rect 10924 6280 11156 6320
rect 11212 6320 11252 7615
rect 11404 7169 11444 7624
rect 11308 7160 11348 7169
rect 11308 6917 11348 7120
rect 11403 7160 11445 7169
rect 11403 7120 11404 7160
rect 11444 7120 11445 7160
rect 11403 7111 11445 7120
rect 11788 7160 11828 7169
rect 11595 6992 11637 7001
rect 11595 6952 11596 6992
rect 11636 6952 11637 6992
rect 11595 6943 11637 6952
rect 11307 6908 11349 6917
rect 11307 6868 11308 6908
rect 11348 6868 11349 6908
rect 11307 6859 11349 6868
rect 11596 6858 11636 6943
rect 11788 6749 11828 7120
rect 11883 7160 11925 7169
rect 12364 7160 12404 7169
rect 12556 7160 12596 7960
rect 12652 7951 12692 7960
rect 12748 7169 12788 8623
rect 12844 7589 12884 8800
rect 13036 8168 13076 9472
rect 13132 9512 13172 9521
rect 13132 9353 13172 9472
rect 13420 9512 13460 9631
rect 13420 9437 13460 9472
rect 13515 9512 13557 9521
rect 13515 9472 13516 9512
rect 13556 9472 13557 9512
rect 13515 9463 13557 9472
rect 13612 9512 13652 10807
rect 14668 10184 14708 10193
rect 14091 10016 14133 10025
rect 14091 9976 14092 10016
rect 14132 9976 14133 10016
rect 14091 9967 14133 9976
rect 13899 9680 13941 9689
rect 13899 9640 13900 9680
rect 13940 9640 13941 9680
rect 13899 9631 13941 9640
rect 13803 9596 13845 9605
rect 13803 9556 13804 9596
rect 13844 9556 13845 9596
rect 13803 9547 13845 9556
rect 13612 9463 13652 9472
rect 13419 9428 13461 9437
rect 13419 9388 13420 9428
rect 13460 9388 13461 9428
rect 13419 9379 13461 9388
rect 13131 9344 13173 9353
rect 13420 9348 13460 9379
rect 13131 9304 13132 9344
rect 13172 9304 13173 9344
rect 13131 9295 13173 9304
rect 13132 8177 13172 9295
rect 13516 9092 13556 9463
rect 13804 9462 13844 9547
rect 13900 9512 13940 9631
rect 13900 9260 13940 9472
rect 13995 9512 14037 9521
rect 13995 9472 13996 9512
rect 14036 9472 14037 9512
rect 13995 9463 14037 9472
rect 14092 9512 14132 9967
rect 14668 9689 14708 10144
rect 14956 9689 14996 10816
rect 15051 10100 15093 10109
rect 15148 10100 15188 11068
rect 15243 10940 15285 10949
rect 15243 10900 15244 10940
rect 15284 10900 15285 10940
rect 15243 10891 15285 10900
rect 15244 10806 15284 10891
rect 15051 10060 15052 10100
rect 15092 10060 15188 10100
rect 15051 10051 15093 10060
rect 15340 10016 15380 11311
rect 15436 10949 15476 12496
rect 15532 12494 15572 12503
rect 15723 12496 15724 12536
rect 15764 12496 15765 12536
rect 15723 12487 15765 12496
rect 15532 11780 15572 12454
rect 15724 12402 15764 12487
rect 15820 12368 15860 13831
rect 15916 13385 15956 14344
rect 16108 14057 16148 16108
rect 16204 16099 16244 16108
rect 16300 15560 16340 15571
rect 16300 15485 16340 15520
rect 16299 15476 16341 15485
rect 16299 15436 16300 15476
rect 16340 15436 16341 15476
rect 16299 15427 16341 15436
rect 16396 15149 16436 17032
rect 16683 17023 16725 17032
rect 16684 16938 16724 17023
rect 16492 16409 16532 16494
rect 16491 16400 16533 16409
rect 16491 16360 16492 16400
rect 16532 16360 16533 16400
rect 16491 16351 16533 16360
rect 16491 16232 16533 16241
rect 16491 16192 16492 16232
rect 16532 16192 16533 16232
rect 16491 16183 16533 16192
rect 16683 16232 16725 16241
rect 16683 16192 16684 16232
rect 16724 16192 16725 16232
rect 16683 16183 16725 16192
rect 16492 16098 16532 16183
rect 16684 16098 16724 16183
rect 16780 15905 16820 17611
rect 17740 17610 17780 17695
rect 18892 17669 18932 19963
rect 19084 19928 19124 20728
rect 19276 20719 19316 20728
rect 20811 20728 20812 20768
rect 20852 20728 20853 20768
rect 20811 20719 20853 20728
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 19659 20264 19701 20273
rect 19659 20224 19660 20264
rect 19700 20224 19796 20264
rect 19659 20215 19701 20224
rect 19756 20180 19796 20224
rect 19756 20131 19796 20140
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19372 20096 19412 20107
rect 19276 19962 19316 20047
rect 19372 20021 19412 20056
rect 19468 20096 19508 20105
rect 19371 20012 19413 20021
rect 19371 19972 19372 20012
rect 19412 19972 19413 20012
rect 19371 19963 19413 19972
rect 19468 19937 19508 20056
rect 19564 20096 19604 20105
rect 19084 19879 19124 19888
rect 19467 19928 19509 19937
rect 19467 19888 19468 19928
rect 19508 19888 19509 19928
rect 19467 19879 19509 19888
rect 19275 19424 19317 19433
rect 19275 19384 19276 19424
rect 19316 19384 19317 19424
rect 19275 19375 19317 19384
rect 19276 18752 19316 19375
rect 19564 19349 19604 20056
rect 20428 20096 20468 20105
rect 20428 19928 20468 20056
rect 20620 19928 20660 19937
rect 20428 19888 20620 19928
rect 20620 19879 20660 19888
rect 20812 19508 20852 20719
rect 21099 20600 21141 20609
rect 21099 20560 21100 20600
rect 21140 20560 21141 20600
rect 21099 20551 21141 20560
rect 21100 20322 21140 20551
rect 20907 20096 20949 20105
rect 20907 20056 20908 20096
rect 20948 20056 20949 20096
rect 20907 20047 20949 20056
rect 21004 20096 21044 20105
rect 20908 19962 20948 20047
rect 20812 19459 20852 19468
rect 21004 19424 21044 20056
rect 20908 19384 21044 19424
rect 19563 19340 19605 19349
rect 19563 19300 19564 19340
rect 19604 19300 19605 19340
rect 19563 19291 19605 19300
rect 20715 19340 20757 19349
rect 20715 19300 20716 19340
rect 20756 19300 20757 19340
rect 20715 19291 20757 19300
rect 19371 19256 19413 19265
rect 19371 19216 19372 19256
rect 19412 19216 19413 19256
rect 19371 19207 19413 19216
rect 20716 19256 20756 19291
rect 19372 19122 19412 19207
rect 20716 19205 20756 19216
rect 20811 19256 20853 19265
rect 20811 19216 20812 19256
rect 20852 19216 20853 19256
rect 20811 19207 20853 19216
rect 20524 19088 20564 19097
rect 20812 19088 20852 19207
rect 20564 19048 20852 19088
rect 20524 19039 20564 19048
rect 20908 19004 20948 19384
rect 21003 19256 21045 19265
rect 21003 19216 21004 19256
rect 21044 19216 21045 19256
rect 21003 19207 21045 19216
rect 21004 19122 21044 19207
rect 20812 18964 20948 19004
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 19564 18752 19604 18761
rect 19276 18712 19564 18752
rect 19564 18703 19604 18712
rect 20524 18752 20564 18761
rect 20812 18752 20852 18964
rect 21003 18920 21045 18929
rect 21003 18880 21004 18920
rect 21044 18880 21045 18920
rect 21003 18871 21045 18880
rect 20907 18836 20949 18845
rect 20907 18796 20908 18836
rect 20948 18796 20949 18836
rect 20907 18787 20949 18796
rect 20564 18712 20852 18752
rect 20524 18703 20564 18712
rect 20235 18584 20277 18593
rect 20235 18544 20236 18584
rect 20276 18544 20277 18584
rect 20235 18535 20277 18544
rect 20620 18584 20660 18593
rect 20812 18584 20852 18712
rect 20660 18544 20756 18584
rect 20620 18535 20660 18544
rect 20236 18450 20276 18535
rect 20139 17996 20181 18005
rect 20139 17956 20140 17996
rect 20180 17956 20181 17996
rect 20139 17947 20181 17956
rect 20140 17862 20180 17947
rect 18988 17744 19028 17753
rect 18891 17660 18933 17669
rect 18891 17620 18892 17660
rect 18932 17620 18933 17660
rect 18891 17611 18933 17620
rect 17931 17156 17973 17165
rect 17931 17116 17932 17156
rect 17972 17116 17973 17156
rect 17931 17107 17973 17116
rect 17548 17072 17588 17081
rect 17548 16913 17588 17032
rect 17932 17072 17972 17107
rect 17932 17021 17972 17032
rect 18316 17072 18356 17083
rect 18988 17081 19028 17704
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 19371 17156 19413 17165
rect 19371 17116 19372 17156
rect 19412 17116 19413 17156
rect 19371 17107 19413 17116
rect 18316 16997 18356 17032
rect 18987 17072 19029 17081
rect 18987 17032 18988 17072
rect 19028 17032 19029 17072
rect 18987 17023 19029 17032
rect 19372 17022 19412 17107
rect 20716 17081 20756 18544
rect 20812 18535 20852 18544
rect 20908 18500 20948 18787
rect 21004 18752 21044 18871
rect 21100 18836 21140 20282
rect 21196 20180 21236 21568
rect 21292 21449 21332 23752
rect 22636 23792 22676 24340
rect 22732 24331 22772 24340
rect 22828 23876 22868 25339
rect 23212 24632 23252 27187
rect 24267 27152 24309 27161
rect 24267 27112 24268 27152
rect 24308 27112 24309 27152
rect 24267 27103 24309 27112
rect 24268 26993 24308 27103
rect 24267 26984 24309 26993
rect 24267 26944 24268 26984
rect 24308 26944 24309 26984
rect 24267 26935 24309 26944
rect 24268 26816 24308 26935
rect 24268 26767 24308 26776
rect 24460 26816 24500 27691
rect 24652 27656 24692 27665
rect 24844 27656 24884 27665
rect 24652 27161 24692 27616
rect 24748 27621 24788 27630
rect 24748 27245 24788 27581
rect 24844 27329 24884 27616
rect 25131 27404 25173 27413
rect 25131 27364 25132 27404
rect 25172 27364 25173 27404
rect 25131 27355 25173 27364
rect 24843 27320 24885 27329
rect 24843 27280 24844 27320
rect 24884 27280 24885 27320
rect 24843 27271 24885 27280
rect 25132 27270 25172 27355
rect 24747 27236 24789 27245
rect 24747 27196 24748 27236
rect 24788 27196 24789 27236
rect 24747 27187 24789 27196
rect 24651 27152 24693 27161
rect 24651 27112 24652 27152
rect 24692 27112 24693 27152
rect 24651 27103 24693 27112
rect 24747 27068 24789 27077
rect 24747 27028 24748 27068
rect 24788 27028 24789 27068
rect 24747 27019 24789 27028
rect 24460 26767 24500 26776
rect 24748 26816 24788 27019
rect 24939 26984 24981 26993
rect 24939 26944 24940 26984
rect 24980 26944 24981 26984
rect 24939 26935 24981 26944
rect 23883 26732 23925 26741
rect 23883 26692 23884 26732
rect 23924 26692 23925 26732
rect 23883 26683 23925 26692
rect 24363 26732 24405 26741
rect 24363 26692 24364 26732
rect 24404 26692 24405 26732
rect 24363 26683 24405 26692
rect 23307 26228 23349 26237
rect 23307 26188 23308 26228
rect 23348 26188 23349 26228
rect 23307 26179 23349 26188
rect 23308 26144 23348 26179
rect 23308 26093 23348 26104
rect 23692 26144 23732 26153
rect 23692 25565 23732 26104
rect 23788 26144 23828 26153
rect 23691 25556 23733 25565
rect 23691 25516 23692 25556
rect 23732 25516 23733 25556
rect 23691 25507 23733 25516
rect 23595 25472 23637 25481
rect 23595 25432 23596 25472
rect 23636 25432 23637 25472
rect 23595 25423 23637 25432
rect 23596 25304 23636 25423
rect 23596 25255 23636 25264
rect 23788 24893 23828 26104
rect 23884 26144 23924 26683
rect 24364 26598 24404 26683
rect 24748 26657 24788 26776
rect 24747 26648 24789 26657
rect 24747 26608 24748 26648
rect 24788 26608 24789 26648
rect 24747 26599 24789 26608
rect 24940 26489 24980 26935
rect 24939 26480 24981 26489
rect 24939 26440 24940 26480
rect 24980 26440 24981 26480
rect 24939 26431 24981 26440
rect 25420 26405 25460 28288
rect 25996 28279 26036 28288
rect 26476 28328 26516 28867
rect 26571 28664 26613 28673
rect 26571 28624 26572 28664
rect 26612 28624 26613 28664
rect 26571 28615 26613 28624
rect 26476 28279 26516 28288
rect 26572 28328 26612 28615
rect 26668 28580 26708 29128
rect 26764 29119 26804 29128
rect 26763 28916 26805 28925
rect 26763 28876 26764 28916
rect 26804 28876 26805 28916
rect 26763 28867 26805 28876
rect 26764 28782 26804 28867
rect 26860 28673 26900 29968
rect 26956 29959 26996 29968
rect 26956 29168 26996 29177
rect 26859 28664 26901 28673
rect 26859 28624 26860 28664
rect 26900 28624 26901 28664
rect 26859 28615 26901 28624
rect 26668 28540 26804 28580
rect 26572 28279 26612 28288
rect 26668 28328 26708 28337
rect 26668 28253 26708 28288
rect 26667 28244 26709 28253
rect 26667 28204 26668 28244
rect 26708 28204 26709 28244
rect 26667 28195 26709 28204
rect 26092 28160 26132 28171
rect 26092 28085 26132 28120
rect 26380 28160 26420 28169
rect 26091 28076 26133 28085
rect 26091 28036 26092 28076
rect 26132 28036 26133 28076
rect 26091 28027 26133 28036
rect 26283 28076 26325 28085
rect 26283 28036 26284 28076
rect 26324 28036 26325 28076
rect 26283 28027 26325 28036
rect 26091 27656 26133 27665
rect 26091 27616 26092 27656
rect 26132 27616 26133 27656
rect 26091 27607 26133 27616
rect 26284 27656 26324 28027
rect 26284 27607 26324 27616
rect 25516 27572 25556 27581
rect 24555 26396 24597 26405
rect 24555 26356 24556 26396
rect 24596 26356 24597 26396
rect 24555 26347 24597 26356
rect 25419 26396 25461 26405
rect 25419 26356 25420 26396
rect 25460 26356 25461 26396
rect 25419 26347 25461 26356
rect 23884 26095 23924 26104
rect 23980 26144 24020 26153
rect 24020 26104 24212 26144
rect 23980 26095 24020 26104
rect 23787 24884 23829 24893
rect 23787 24844 23788 24884
rect 23828 24844 23829 24884
rect 23787 24835 23829 24844
rect 23308 24632 23348 24641
rect 23212 24592 23308 24632
rect 23212 24137 23252 24592
rect 23308 24583 23348 24592
rect 23211 24128 23253 24137
rect 23211 24088 23212 24128
rect 23252 24088 23253 24128
rect 23211 24079 23253 24088
rect 24172 24044 24212 26104
rect 24267 26060 24309 26069
rect 24267 26020 24268 26060
rect 24308 26020 24309 26060
rect 24267 26011 24309 26020
rect 24268 25926 24308 26011
rect 24556 25556 24596 26347
rect 25516 26228 25556 27532
rect 26092 27488 26132 27607
rect 26092 27439 26132 27448
rect 26188 26984 26228 26993
rect 25324 26188 25556 26228
rect 25612 26944 26188 26984
rect 25131 26144 25173 26153
rect 25131 26104 25132 26144
rect 25172 26104 25173 26144
rect 25131 26095 25173 26104
rect 25132 26010 25172 26095
rect 24843 25892 24885 25901
rect 24843 25852 24844 25892
rect 24884 25852 24885 25892
rect 24843 25843 24885 25852
rect 24556 24221 24596 25516
rect 24844 25304 24884 25843
rect 24844 25255 24884 25264
rect 25132 25304 25172 25313
rect 25132 24809 25172 25264
rect 25324 25229 25364 26188
rect 25516 25892 25556 25901
rect 25516 25565 25556 25852
rect 25515 25556 25557 25565
rect 25515 25516 25516 25556
rect 25556 25516 25557 25556
rect 25515 25507 25557 25516
rect 25516 25304 25556 25313
rect 25612 25304 25652 26944
rect 26188 26935 26228 26944
rect 25899 26480 25941 26489
rect 25899 26440 25900 26480
rect 25940 26440 25941 26480
rect 25899 26431 25941 26440
rect 25804 26144 25844 26153
rect 25804 25985 25844 26104
rect 25900 26139 25940 26431
rect 26380 26237 26420 28120
rect 26668 26573 26708 28195
rect 26764 27665 26804 28540
rect 26956 28253 26996 29128
rect 27052 29168 27092 31060
rect 27148 30680 27188 32479
rect 27243 32360 27285 32369
rect 27243 32320 27244 32360
rect 27284 32320 27285 32360
rect 27243 32311 27285 32320
rect 27244 32226 27284 32311
rect 27340 31529 27380 32656
rect 27339 31520 27381 31529
rect 27339 31480 27340 31520
rect 27380 31480 27381 31520
rect 27339 31471 27381 31480
rect 27340 31352 27380 31361
rect 27340 31193 27380 31312
rect 27436 31352 27476 32824
rect 27532 32813 27572 32824
rect 27628 32864 27668 33328
rect 27723 33116 27765 33125
rect 27723 33076 27724 33116
rect 27764 33076 27765 33116
rect 27723 33067 27765 33076
rect 27628 32815 27668 32824
rect 27724 32864 27764 33067
rect 27820 32873 27860 33571
rect 27724 32815 27764 32824
rect 27819 32864 27861 32873
rect 27819 32824 27820 32864
rect 27860 32824 27861 32864
rect 27819 32815 27861 32824
rect 27627 32696 27669 32705
rect 27627 32656 27628 32696
rect 27668 32656 27669 32696
rect 27627 32647 27669 32656
rect 27819 32696 27861 32705
rect 27819 32656 27820 32696
rect 27860 32656 27861 32696
rect 27819 32647 27861 32656
rect 27531 32528 27573 32537
rect 27531 32488 27532 32528
rect 27572 32488 27573 32528
rect 27531 32479 27573 32488
rect 27532 32192 27572 32479
rect 27532 32143 27572 32152
rect 27628 32024 27668 32647
rect 27820 32562 27860 32647
rect 27916 32537 27956 34243
rect 28588 34049 28628 34504
rect 28780 34376 28820 34385
rect 28587 34040 28629 34049
rect 28587 34000 28588 34040
rect 28628 34000 28629 34040
rect 28587 33991 28629 34000
rect 28011 33704 28053 33713
rect 28011 33664 28012 33704
rect 28052 33664 28053 33704
rect 28011 33655 28053 33664
rect 28012 33620 28052 33655
rect 28012 33569 28052 33580
rect 28587 33116 28629 33125
rect 28587 33076 28588 33116
rect 28628 33076 28629 33116
rect 28587 33067 28629 33076
rect 28395 33032 28437 33041
rect 28395 32992 28396 33032
rect 28436 32992 28437 33032
rect 28395 32983 28437 32992
rect 28012 32864 28052 32873
rect 27915 32528 27957 32537
rect 27915 32488 27916 32528
rect 27956 32488 27957 32528
rect 27915 32479 27957 32488
rect 28012 32369 28052 32824
rect 28107 32696 28149 32705
rect 28107 32656 28108 32696
rect 28148 32656 28149 32696
rect 28107 32647 28149 32656
rect 28011 32360 28053 32369
rect 28011 32320 28012 32360
rect 28052 32320 28053 32360
rect 28011 32311 28053 32320
rect 27819 32192 27861 32201
rect 27819 32152 27820 32192
rect 27860 32152 27861 32192
rect 27819 32143 27861 32152
rect 27916 32192 27956 32201
rect 28012 32192 28052 32311
rect 27956 32152 28052 32192
rect 27916 32143 27956 32152
rect 27820 32058 27860 32143
rect 27436 31303 27476 31312
rect 27532 31984 27668 32024
rect 27532 31352 27572 31984
rect 27627 31604 27669 31613
rect 27627 31564 27628 31604
rect 27668 31564 27669 31604
rect 27627 31555 27669 31564
rect 27532 31303 27572 31312
rect 27628 31352 27668 31555
rect 27819 31520 27861 31529
rect 27819 31480 27820 31520
rect 27860 31480 27861 31520
rect 27819 31471 27861 31480
rect 28011 31520 28053 31529
rect 28011 31480 28012 31520
rect 28052 31480 28053 31520
rect 28011 31471 28053 31480
rect 27628 31303 27668 31312
rect 27820 31352 27860 31471
rect 27820 31303 27860 31312
rect 27916 31352 27956 31361
rect 27916 31193 27956 31312
rect 28012 31268 28052 31471
rect 28108 31352 28148 32647
rect 28396 32192 28436 32983
rect 28491 32864 28533 32873
rect 28491 32824 28492 32864
rect 28532 32824 28533 32864
rect 28491 32815 28533 32824
rect 28492 32360 28532 32815
rect 28492 32311 28532 32320
rect 28588 32192 28628 33067
rect 28683 33032 28725 33041
rect 28683 32992 28684 33032
rect 28724 32992 28725 33032
rect 28683 32983 28725 32992
rect 28684 32898 28724 32983
rect 28396 32143 28436 32152
rect 28492 32152 28628 32192
rect 28108 31303 28148 31312
rect 28204 31940 28244 31949
rect 28012 31219 28052 31228
rect 27339 31184 27381 31193
rect 27339 31144 27340 31184
rect 27380 31144 27381 31184
rect 27339 31135 27381 31144
rect 27915 31184 27957 31193
rect 27915 31144 27916 31184
rect 27956 31144 27957 31184
rect 27915 31135 27957 31144
rect 27627 30848 27669 30857
rect 27627 30808 27628 30848
rect 27668 30808 27669 30848
rect 27627 30799 27669 30808
rect 27340 30680 27380 30689
rect 27628 30680 27668 30799
rect 27723 30764 27765 30773
rect 27723 30724 27724 30764
rect 27764 30724 27765 30764
rect 27723 30715 27765 30724
rect 27148 30640 27340 30680
rect 27380 30640 27572 30680
rect 27340 30631 27380 30640
rect 27532 30512 27572 30640
rect 27628 30631 27668 30640
rect 27724 30630 27764 30715
rect 27532 30472 27668 30512
rect 27147 30344 27189 30353
rect 27147 30304 27148 30344
rect 27188 30304 27189 30344
rect 27147 30295 27189 30304
rect 27052 29119 27092 29128
rect 27148 29000 27188 30295
rect 27340 29840 27380 29849
rect 27628 29840 27668 30472
rect 27380 29800 27572 29840
rect 27340 29791 27380 29800
rect 27244 29756 27284 29765
rect 27244 29429 27284 29716
rect 27243 29420 27285 29429
rect 27243 29380 27244 29420
rect 27284 29380 27285 29420
rect 27243 29371 27285 29380
rect 27435 29336 27477 29345
rect 27435 29296 27436 29336
rect 27476 29296 27477 29336
rect 27435 29287 27477 29296
rect 27244 29177 27284 29262
rect 27243 29168 27285 29177
rect 27243 29128 27244 29168
rect 27284 29128 27285 29168
rect 27243 29119 27285 29128
rect 27436 29168 27476 29287
rect 27532 29177 27572 29800
rect 27628 29597 27668 29800
rect 28012 30428 28052 30437
rect 28204 30428 28244 31900
rect 28299 31352 28341 31361
rect 28299 31312 28300 31352
rect 28340 31312 28341 31352
rect 28299 31303 28341 31312
rect 28300 31218 28340 31303
rect 28395 31268 28437 31277
rect 28395 31228 28396 31268
rect 28436 31228 28437 31268
rect 28395 31219 28437 31228
rect 28396 31134 28436 31219
rect 28396 30680 28436 30689
rect 28204 30388 28340 30428
rect 27915 29756 27957 29765
rect 27915 29716 27916 29756
rect 27956 29716 27957 29756
rect 27915 29707 27957 29716
rect 27916 29622 27956 29707
rect 27627 29588 27669 29597
rect 27627 29548 27628 29588
rect 27668 29548 27669 29588
rect 27627 29539 27669 29548
rect 27436 29093 27476 29128
rect 27531 29168 27573 29177
rect 27531 29128 27532 29168
rect 27572 29128 27573 29168
rect 27531 29119 27573 29128
rect 27435 29084 27477 29093
rect 27435 29044 27436 29084
rect 27476 29044 27477 29084
rect 27435 29035 27477 29044
rect 27532 29034 27572 29119
rect 27244 29000 27284 29009
rect 27148 28960 27244 29000
rect 27244 28951 27284 28960
rect 27532 28580 27572 28589
rect 27628 28580 27668 29539
rect 27916 29261 27956 29305
rect 27915 29252 27957 29261
rect 27915 29212 27916 29252
rect 27956 29212 27957 29252
rect 27915 29210 27957 29212
rect 27915 29203 27916 29210
rect 27956 29203 27957 29210
rect 27916 29161 27956 29170
rect 27915 29000 27957 29009
rect 27915 28960 27916 29000
rect 27956 28960 27957 29000
rect 28012 29000 28052 30388
rect 28203 29420 28245 29429
rect 28203 29380 28204 29420
rect 28244 29380 28245 29420
rect 28203 29371 28245 29380
rect 28107 29336 28149 29345
rect 28107 29296 28108 29336
rect 28148 29296 28149 29336
rect 28107 29287 28149 29296
rect 28108 29168 28148 29287
rect 28204 29261 28244 29371
rect 28203 29252 28245 29261
rect 28203 29212 28204 29252
rect 28244 29212 28245 29252
rect 28203 29203 28245 29212
rect 28108 29119 28148 29128
rect 28204 29168 28244 29203
rect 28204 29118 28244 29128
rect 28012 28960 28148 29000
rect 27915 28951 27957 28960
rect 27916 28866 27956 28951
rect 27572 28540 27668 28580
rect 27532 28531 27572 28540
rect 27723 28328 27765 28337
rect 27723 28288 27724 28328
rect 27764 28288 27765 28328
rect 27723 28279 27765 28288
rect 26955 28244 26997 28253
rect 26955 28204 26956 28244
rect 26996 28204 26997 28244
rect 26955 28195 26997 28204
rect 27724 28001 27764 28279
rect 27723 27992 27765 28001
rect 27723 27952 27724 27992
rect 27764 27952 27765 27992
rect 27723 27943 27765 27952
rect 26763 27656 26805 27665
rect 26763 27616 26764 27656
rect 26804 27616 26805 27656
rect 26763 27607 26805 27616
rect 27724 27656 27764 27665
rect 26764 27522 26804 27607
rect 27724 27413 27764 27616
rect 28012 27656 28052 27665
rect 28012 27497 28052 27616
rect 28108 27656 28148 28960
rect 28300 28664 28340 30388
rect 28396 30353 28436 30640
rect 28492 30680 28532 32152
rect 28780 32108 28820 34336
rect 28972 32612 29012 35008
rect 29164 34637 29204 36091
rect 29452 36006 29492 36091
rect 29548 35216 29588 36436
rect 29740 36436 29836 36476
rect 29644 35888 29684 35897
rect 29740 35888 29780 36436
rect 29836 36427 29876 36436
rect 29684 35848 29780 35888
rect 30028 35888 30068 36604
rect 29644 35839 29684 35848
rect 30028 35839 30068 35848
rect 30508 35393 30548 36688
rect 30796 36728 30836 36737
rect 30796 36149 30836 36688
rect 30795 36140 30837 36149
rect 30795 36100 30796 36140
rect 30836 36100 30837 36140
rect 30795 36091 30837 36100
rect 30892 36056 30932 37192
rect 30988 36905 31028 37360
rect 31755 37400 31797 37409
rect 32428 37400 32468 37409
rect 31755 37360 31756 37400
rect 31796 37360 31797 37400
rect 31755 37351 31797 37360
rect 32044 37360 32428 37400
rect 31756 37266 31796 37351
rect 30987 36896 31029 36905
rect 30987 36856 30988 36896
rect 31028 36856 31029 36896
rect 30987 36847 31029 36856
rect 31659 36896 31701 36905
rect 31659 36856 31660 36896
rect 31700 36856 31701 36896
rect 31659 36847 31701 36856
rect 31660 36762 31700 36847
rect 32044 36569 32084 37360
rect 32428 37351 32468 37360
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 33292 36821 33332 36906
rect 32715 36812 32757 36821
rect 32715 36772 32716 36812
rect 32756 36772 32757 36812
rect 32715 36763 32757 36772
rect 33291 36812 33333 36821
rect 33291 36772 33292 36812
rect 33332 36772 33333 36812
rect 33291 36763 33333 36772
rect 32332 36728 32372 36737
rect 32620 36728 32660 36737
rect 32140 36688 32332 36728
rect 31371 36560 31413 36569
rect 31371 36520 31372 36560
rect 31412 36520 31413 36560
rect 31371 36511 31413 36520
rect 32043 36560 32085 36569
rect 32043 36520 32044 36560
rect 32084 36520 32085 36560
rect 32043 36511 32085 36520
rect 30892 36016 31124 36056
rect 30892 35888 30932 35897
rect 30603 35720 30645 35729
rect 30603 35680 30604 35720
rect 30644 35680 30645 35720
rect 30603 35671 30645 35680
rect 29739 35384 29781 35393
rect 29739 35344 29740 35384
rect 29780 35344 29781 35384
rect 29739 35335 29781 35344
rect 30507 35384 30549 35393
rect 30507 35344 30508 35384
rect 30548 35344 30549 35384
rect 30507 35335 30549 35344
rect 29740 35300 29780 35335
rect 29740 35249 29780 35260
rect 29548 35167 29588 35176
rect 29644 35216 29684 35225
rect 29644 35057 29684 35176
rect 29835 35216 29877 35225
rect 29835 35176 29836 35216
rect 29876 35176 29877 35216
rect 29835 35167 29877 35176
rect 30411 35216 30453 35225
rect 30411 35176 30412 35216
rect 30452 35176 30453 35216
rect 30411 35167 30453 35176
rect 30508 35216 30548 35225
rect 29836 35082 29876 35167
rect 30123 35132 30165 35141
rect 30123 35092 30124 35132
rect 30164 35092 30165 35132
rect 30123 35083 30165 35092
rect 29260 35048 29300 35057
rect 29643 35048 29685 35057
rect 29300 35008 29588 35048
rect 29260 34999 29300 35008
rect 29163 34628 29205 34637
rect 29163 34588 29164 34628
rect 29204 34588 29205 34628
rect 29163 34579 29205 34588
rect 29452 34208 29492 34217
rect 29452 34049 29492 34168
rect 29451 34040 29493 34049
rect 29451 34000 29452 34040
rect 29492 34000 29493 34040
rect 29451 33991 29493 34000
rect 29067 33956 29109 33965
rect 29067 33916 29068 33956
rect 29108 33916 29109 33956
rect 29067 33907 29109 33916
rect 29068 33545 29108 33907
rect 29164 33704 29204 33713
rect 29548 33704 29588 35008
rect 29643 35008 29644 35048
rect 29684 35008 29685 35048
rect 29643 34999 29685 35008
rect 29835 34460 29877 34469
rect 29835 34420 29836 34460
rect 29876 34420 29877 34460
rect 29835 34411 29877 34420
rect 29836 34376 29876 34411
rect 29836 34325 29876 34336
rect 29932 34376 29972 34385
rect 29932 34217 29972 34336
rect 30028 34376 30068 34385
rect 29931 34208 29973 34217
rect 29931 34168 29932 34208
rect 29972 34168 29973 34208
rect 29931 34159 29973 34168
rect 30028 33965 30068 34336
rect 30124 34376 30164 35083
rect 30412 35082 30452 35167
rect 30220 35048 30260 35057
rect 30260 35008 30356 35048
rect 30220 34999 30260 35008
rect 30219 34544 30261 34553
rect 30219 34504 30220 34544
rect 30260 34504 30261 34544
rect 30219 34495 30261 34504
rect 30124 34327 30164 34336
rect 30027 33956 30069 33965
rect 30027 33916 30028 33956
rect 30068 33916 30069 33956
rect 30027 33907 30069 33916
rect 30028 33704 30068 33713
rect 29204 33664 29492 33704
rect 29548 33664 30028 33704
rect 29164 33655 29204 33664
rect 29067 33536 29109 33545
rect 29067 33496 29068 33536
rect 29108 33496 29109 33536
rect 29067 33487 29109 33496
rect 29163 32948 29205 32957
rect 29163 32908 29164 32948
rect 29204 32908 29205 32948
rect 29163 32899 29205 32908
rect 29067 32864 29109 32873
rect 29067 32824 29068 32864
rect 29108 32824 29109 32864
rect 29067 32815 29109 32824
rect 29164 32864 29204 32899
rect 29356 32873 29396 32958
rect 29068 32730 29108 32815
rect 29164 32813 29204 32824
rect 29355 32864 29397 32873
rect 29355 32824 29356 32864
rect 29396 32824 29397 32864
rect 29355 32815 29397 32824
rect 29260 32696 29300 32705
rect 29300 32656 29396 32696
rect 29260 32647 29300 32656
rect 28972 32572 29108 32612
rect 28588 32068 28820 32108
rect 28588 31529 28628 32068
rect 28684 31940 28724 31949
rect 28724 31900 29012 31940
rect 28684 31891 28724 31900
rect 28587 31520 28629 31529
rect 28587 31480 28588 31520
rect 28628 31480 28629 31520
rect 28587 31471 28629 31480
rect 28780 31520 28820 31529
rect 28587 30848 28629 30857
rect 28587 30808 28588 30848
rect 28628 30808 28629 30848
rect 28587 30799 28629 30808
rect 28492 30631 28532 30640
rect 28588 30680 28628 30799
rect 28588 30631 28628 30640
rect 28684 30680 28724 30689
rect 28491 30428 28533 30437
rect 28491 30388 28492 30428
rect 28532 30388 28533 30428
rect 28491 30379 28533 30388
rect 28395 30344 28437 30353
rect 28395 30304 28396 30344
rect 28436 30304 28437 30344
rect 28395 30295 28437 30304
rect 28395 29168 28437 29177
rect 28395 29128 28396 29168
rect 28436 29128 28437 29168
rect 28395 29119 28437 29128
rect 28492 29168 28532 30379
rect 28492 29119 28532 29128
rect 28588 29840 28628 29849
rect 28396 29034 28436 29119
rect 28588 29093 28628 29800
rect 28684 29345 28724 30640
rect 28780 29849 28820 31480
rect 28972 31352 29012 31900
rect 29068 31352 29108 32572
rect 29356 32192 29396 32656
rect 29356 32143 29396 32152
rect 29356 31352 29396 31361
rect 29068 31312 29356 31352
rect 28972 31303 29012 31312
rect 29356 31303 29396 31312
rect 29068 30428 29108 30437
rect 28876 30388 29068 30428
rect 28779 29840 28821 29849
rect 28779 29800 28780 29840
rect 28820 29800 28821 29840
rect 28779 29791 28821 29800
rect 28876 29840 28916 30388
rect 29068 30379 29108 30388
rect 29163 30344 29205 30353
rect 29163 30304 29164 30344
rect 29204 30304 29205 30344
rect 29163 30295 29205 30304
rect 28876 29791 28916 29800
rect 28683 29336 28725 29345
rect 28683 29296 28684 29336
rect 28724 29296 28725 29336
rect 28683 29287 28725 29296
rect 28971 29336 29013 29345
rect 28971 29296 28972 29336
rect 29012 29296 29013 29336
rect 28971 29287 29013 29296
rect 28684 29177 28724 29287
rect 28683 29168 28725 29177
rect 28683 29128 28684 29168
rect 28724 29128 28725 29168
rect 28683 29119 28725 29128
rect 28587 29084 28629 29093
rect 28587 29044 28588 29084
rect 28628 29044 28629 29084
rect 28587 29035 28629 29044
rect 28972 29000 29012 29287
rect 29068 29168 29108 29177
rect 29164 29168 29204 30295
rect 29452 30269 29492 33664
rect 30028 33655 30068 33664
rect 30220 33116 30260 34495
rect 30316 33293 30356 35008
rect 30508 34889 30548 35176
rect 30604 35216 30644 35671
rect 30892 35309 30932 35848
rect 30891 35300 30933 35309
rect 30891 35260 30892 35300
rect 30932 35260 30933 35300
rect 30891 35251 30933 35260
rect 30604 35167 30644 35176
rect 30700 35216 30740 35225
rect 30507 34880 30549 34889
rect 30507 34840 30508 34880
rect 30548 34840 30549 34880
rect 30507 34831 30549 34840
rect 30411 34040 30453 34049
rect 30411 34000 30412 34040
rect 30452 34000 30453 34040
rect 30411 33991 30453 34000
rect 30412 33788 30452 33991
rect 30412 33739 30452 33748
rect 30411 33620 30453 33629
rect 30411 33580 30412 33620
rect 30452 33580 30453 33620
rect 30411 33571 30453 33580
rect 30315 33284 30357 33293
rect 30315 33244 30316 33284
rect 30356 33244 30357 33284
rect 30315 33235 30357 33244
rect 30220 33067 30260 33076
rect 30315 33116 30357 33125
rect 30315 33076 30316 33116
rect 30356 33076 30357 33116
rect 30315 33067 30357 33076
rect 29547 32864 29589 32873
rect 29547 32824 29548 32864
rect 29588 32824 29589 32864
rect 29547 32815 29589 32824
rect 30219 32864 30261 32873
rect 30219 32824 30220 32864
rect 30260 32824 30261 32864
rect 30219 32815 30261 32824
rect 29548 30857 29588 32815
rect 30028 31940 30068 31949
rect 29547 30848 29589 30857
rect 29547 30808 29548 30848
rect 29588 30808 29589 30848
rect 29547 30799 29589 30808
rect 30028 30689 30068 31900
rect 30220 31352 30260 32815
rect 30220 31303 30260 31312
rect 29740 30680 29780 30689
rect 29451 30260 29493 30269
rect 29451 30220 29452 30260
rect 29492 30220 29493 30260
rect 29451 30211 29493 30220
rect 29259 29840 29301 29849
rect 29259 29800 29260 29840
rect 29300 29800 29301 29840
rect 29259 29791 29301 29800
rect 29260 29706 29300 29791
rect 29740 29345 29780 30640
rect 30027 30680 30069 30689
rect 30027 30640 30028 30680
rect 30068 30640 30069 30680
rect 30027 30631 30069 30640
rect 30316 30521 30356 33067
rect 30315 30512 30357 30521
rect 30315 30472 30316 30512
rect 30356 30472 30357 30512
rect 30315 30463 30357 30472
rect 29931 30428 29973 30437
rect 29931 30388 29932 30428
rect 29972 30388 29973 30428
rect 29931 30379 29973 30388
rect 29932 30294 29972 30379
rect 30412 30344 30452 33571
rect 30508 33032 30548 34831
rect 30700 34469 30740 35176
rect 30892 34973 30932 35251
rect 30988 35216 31028 35225
rect 30891 34964 30933 34973
rect 30891 34924 30892 34964
rect 30932 34924 30933 34964
rect 30891 34915 30933 34924
rect 30699 34460 30741 34469
rect 30699 34420 30700 34460
rect 30740 34420 30741 34460
rect 30699 34411 30741 34420
rect 30988 34301 31028 35176
rect 30987 34292 31029 34301
rect 30987 34252 30988 34292
rect 31028 34252 31029 34292
rect 30987 34243 31029 34252
rect 30699 34208 30741 34217
rect 30699 34168 30700 34208
rect 30740 34168 30741 34208
rect 30699 34159 30741 34168
rect 30796 34208 30836 34217
rect 30603 33704 30645 33713
rect 30603 33664 30604 33704
rect 30644 33664 30645 33704
rect 30603 33655 30645 33664
rect 30604 33570 30644 33655
rect 30700 33125 30740 34159
rect 30699 33116 30741 33125
rect 30699 33076 30700 33116
rect 30740 33076 30741 33116
rect 30699 33067 30741 33076
rect 30508 32992 30644 33032
rect 30508 32864 30548 32873
rect 30508 32285 30548 32824
rect 30507 32276 30549 32285
rect 30507 32236 30508 32276
rect 30548 32236 30549 32276
rect 30507 32227 30549 32236
rect 30220 30304 30452 30344
rect 30508 32192 30548 32227
rect 30123 30260 30165 30269
rect 30123 30220 30124 30260
rect 30164 30220 30165 30260
rect 30123 30211 30165 30220
rect 30124 29840 30164 30211
rect 30124 29791 30164 29800
rect 30123 29588 30165 29597
rect 30123 29548 30124 29588
rect 30164 29548 30165 29588
rect 30123 29539 30165 29548
rect 29739 29336 29781 29345
rect 29739 29296 29740 29336
rect 29780 29296 29781 29336
rect 29739 29287 29781 29296
rect 29931 29252 29973 29261
rect 29931 29212 29932 29252
rect 29972 29212 29973 29252
rect 29931 29203 29973 29212
rect 29108 29128 29204 29168
rect 29260 29168 29300 29179
rect 29068 29119 29108 29128
rect 29260 29093 29300 29128
rect 29356 29168 29396 29177
rect 29836 29168 29876 29177
rect 29396 29128 29836 29168
rect 29356 29119 29396 29128
rect 29836 29119 29876 29128
rect 29932 29168 29972 29203
rect 29932 29117 29972 29128
rect 30124 29168 30164 29539
rect 30124 29119 30164 29128
rect 30220 29168 30260 30304
rect 30315 29336 30357 29345
rect 30315 29296 30316 29336
rect 30356 29296 30357 29336
rect 30315 29287 30357 29296
rect 30220 29119 30260 29128
rect 29259 29084 29301 29093
rect 29259 29044 29260 29084
rect 29300 29044 29301 29084
rect 29259 29035 29301 29044
rect 29068 29000 29108 29009
rect 30316 29000 30356 29287
rect 30411 29168 30453 29177
rect 30411 29128 30412 29168
rect 30452 29128 30453 29168
rect 30411 29119 30453 29128
rect 30412 29034 30452 29119
rect 28972 28960 29068 29000
rect 29068 28951 29108 28960
rect 30220 28960 30356 29000
rect 28300 28624 28724 28664
rect 28492 28328 28532 28337
rect 28492 28169 28532 28288
rect 28587 28328 28629 28337
rect 28587 28288 28588 28328
rect 28628 28288 28629 28328
rect 28684 28328 28724 28624
rect 29643 28496 29685 28505
rect 29643 28456 29644 28496
rect 29684 28456 29685 28496
rect 29643 28447 29685 28456
rect 28875 28412 28917 28421
rect 28875 28372 28876 28412
rect 28916 28372 28917 28412
rect 28875 28363 28917 28372
rect 28780 28328 28820 28337
rect 28684 28288 28780 28328
rect 28587 28279 28629 28288
rect 28780 28279 28820 28288
rect 28876 28328 28916 28363
rect 28588 28194 28628 28279
rect 28876 28277 28916 28288
rect 29068 28328 29108 28337
rect 29108 28288 29204 28328
rect 29068 28279 29108 28288
rect 28971 28244 29013 28253
rect 28971 28204 28972 28244
rect 29012 28204 29013 28244
rect 28971 28195 29013 28204
rect 28108 27607 28148 27616
rect 28300 28160 28340 28169
rect 28011 27488 28053 27497
rect 28011 27448 28012 27488
rect 28052 27448 28053 27488
rect 28011 27439 28053 27448
rect 27147 27404 27189 27413
rect 27147 27364 27148 27404
rect 27188 27364 27189 27404
rect 27147 27355 27189 27364
rect 27723 27404 27765 27413
rect 27723 27364 27724 27404
rect 27764 27364 27765 27404
rect 27723 27355 27765 27364
rect 26667 26564 26709 26573
rect 26667 26524 26668 26564
rect 26708 26524 26709 26564
rect 26667 26515 26709 26524
rect 26379 26228 26421 26237
rect 26379 26188 26380 26228
rect 26420 26188 26421 26228
rect 26379 26179 26421 26188
rect 25900 26090 25940 26099
rect 25995 26144 26037 26153
rect 26956 26144 26996 26153
rect 25995 26104 25996 26144
rect 26036 26104 26037 26144
rect 25995 26095 26037 26104
rect 26860 26104 26956 26144
rect 25996 26010 26036 26095
rect 25803 25976 25845 25985
rect 25803 25936 25804 25976
rect 25844 25936 25845 25976
rect 25803 25927 25845 25936
rect 26283 25892 26325 25901
rect 26283 25852 26284 25892
rect 26324 25852 26325 25892
rect 26283 25843 26325 25852
rect 26284 25758 26324 25843
rect 26860 25481 26900 26104
rect 26956 26095 26996 26104
rect 26955 25892 26997 25901
rect 26955 25852 26956 25892
rect 26996 25852 26997 25892
rect 26955 25843 26997 25852
rect 26859 25472 26901 25481
rect 26859 25432 26860 25472
rect 26900 25432 26901 25472
rect 26859 25423 26901 25432
rect 25556 25264 25652 25304
rect 26379 25304 26421 25313
rect 26379 25264 26380 25304
rect 26420 25264 26421 25304
rect 25516 25255 25556 25264
rect 26379 25255 26421 25264
rect 25323 25220 25365 25229
rect 25323 25180 25324 25220
rect 25364 25180 25365 25220
rect 25323 25171 25365 25180
rect 26380 25170 26420 25255
rect 25131 24800 25173 24809
rect 25131 24760 25132 24800
rect 25172 24760 25173 24800
rect 25131 24751 25173 24760
rect 25803 24800 25845 24809
rect 25803 24760 25804 24800
rect 25844 24760 25845 24800
rect 25803 24751 25845 24760
rect 25804 24666 25844 24751
rect 25708 24632 25748 24641
rect 25612 24592 25708 24632
rect 24555 24212 24597 24221
rect 24555 24172 24556 24212
rect 24596 24172 24597 24212
rect 24555 24163 24597 24172
rect 24172 24004 24980 24044
rect 23404 23960 23444 23969
rect 23444 23920 23732 23960
rect 23404 23911 23444 23920
rect 22636 23743 22676 23752
rect 22732 23836 22868 23876
rect 22732 23792 22772 23836
rect 22924 23801 22964 23886
rect 23308 23801 23348 23832
rect 22732 23717 22772 23752
rect 22923 23792 22965 23801
rect 22923 23752 22924 23792
rect 22964 23752 22965 23792
rect 22923 23743 22965 23752
rect 23307 23792 23349 23801
rect 23307 23752 23308 23792
rect 23348 23752 23349 23792
rect 23307 23743 23349 23752
rect 23404 23792 23444 23803
rect 22731 23708 22773 23717
rect 22731 23668 22732 23708
rect 22772 23668 22773 23708
rect 22731 23659 22773 23668
rect 23308 23708 23348 23743
rect 23404 23717 23444 23752
rect 23499 23792 23541 23801
rect 23499 23752 23500 23792
rect 23540 23752 23541 23792
rect 23499 23743 23541 23752
rect 23692 23792 23732 23920
rect 24652 23801 24692 23886
rect 23692 23743 23732 23752
rect 23883 23792 23925 23801
rect 23883 23752 23884 23792
rect 23924 23752 23925 23792
rect 23883 23743 23925 23752
rect 24075 23792 24117 23801
rect 24075 23752 24076 23792
rect 24116 23752 24117 23792
rect 24075 23743 24117 23752
rect 24651 23792 24693 23801
rect 24651 23752 24652 23792
rect 24692 23752 24693 23792
rect 24651 23743 24693 23752
rect 24844 23792 24884 23803
rect 22732 23628 22772 23659
rect 22924 23624 22964 23633
rect 23116 23624 23156 23633
rect 22964 23584 23060 23624
rect 22924 23575 22964 23584
rect 23020 23120 23060 23584
rect 23116 23288 23156 23584
rect 23212 23624 23252 23635
rect 23212 23549 23252 23584
rect 23211 23540 23253 23549
rect 23211 23500 23212 23540
rect 23252 23500 23253 23540
rect 23211 23491 23253 23500
rect 23116 23248 23252 23288
rect 23116 23120 23156 23129
rect 23020 23080 23116 23120
rect 23116 23071 23156 23080
rect 23212 22532 23252 23248
rect 23308 22952 23348 23668
rect 23403 23708 23445 23717
rect 23403 23668 23404 23708
rect 23444 23668 23445 23708
rect 23403 23659 23445 23668
rect 23500 23658 23540 23743
rect 23788 23708 23828 23717
rect 23403 23540 23445 23549
rect 23403 23500 23404 23540
rect 23444 23500 23445 23540
rect 23403 23491 23445 23500
rect 23404 23127 23444 23491
rect 23404 23078 23444 23087
rect 23692 23120 23732 23129
rect 23404 22952 23444 22961
rect 23692 22952 23732 23080
rect 23788 23120 23828 23668
rect 23884 23658 23924 23743
rect 23788 23071 23828 23080
rect 23883 23120 23925 23129
rect 23883 23080 23884 23120
rect 23924 23080 23925 23120
rect 23883 23071 23925 23080
rect 23980 23120 24020 23129
rect 23884 22986 23924 23071
rect 23308 22912 23351 22952
rect 23311 22793 23351 22912
rect 23444 22912 23732 22952
rect 23404 22903 23444 22912
rect 23307 22784 23351 22793
rect 23307 22744 23308 22784
rect 23348 22744 23351 22784
rect 23595 22784 23637 22793
rect 23595 22744 23596 22784
rect 23636 22744 23637 22784
rect 23307 22735 23349 22744
rect 23595 22735 23637 22744
rect 23020 22492 23252 22532
rect 21676 22448 21716 22457
rect 21580 22408 21676 22448
rect 21580 21608 21620 22408
rect 21676 22399 21716 22408
rect 21580 21559 21620 21568
rect 22444 21608 22484 21617
rect 22444 21449 22484 21568
rect 21291 21440 21333 21449
rect 21291 21400 21292 21440
rect 21332 21400 21333 21440
rect 21291 21391 21333 21400
rect 22443 21440 22485 21449
rect 22443 21400 22444 21440
rect 22484 21400 22485 21440
rect 22443 21391 22485 21400
rect 21291 20852 21333 20861
rect 21291 20812 21292 20852
rect 21332 20812 21333 20852
rect 21291 20803 21333 20812
rect 22155 20852 22197 20861
rect 22155 20812 22156 20852
rect 22196 20812 22197 20852
rect 22155 20803 22197 20812
rect 21292 20718 21332 20803
rect 22156 20768 22196 20803
rect 22156 20717 22196 20728
rect 22347 20768 22389 20777
rect 22347 20728 22348 20768
rect 22388 20728 22389 20768
rect 22347 20719 22389 20728
rect 22444 20768 22484 20777
rect 22348 20634 22388 20719
rect 21483 20600 21525 20609
rect 21483 20560 21484 20600
rect 21524 20560 21525 20600
rect 21483 20551 21525 20560
rect 21675 20600 21717 20609
rect 21675 20560 21676 20600
rect 21716 20560 21717 20600
rect 21675 20551 21717 20560
rect 21484 20466 21524 20551
rect 21484 20180 21524 20189
rect 21196 20140 21484 20180
rect 21484 20131 21524 20140
rect 21676 20096 21716 20551
rect 21676 20047 21716 20056
rect 21772 20264 21812 20273
rect 21772 20021 21812 20224
rect 21964 20264 22004 20273
rect 21867 20180 21909 20189
rect 21867 20140 21868 20180
rect 21908 20140 21909 20180
rect 21867 20131 21909 20140
rect 21771 20012 21813 20021
rect 21771 19972 21772 20012
rect 21812 19972 21813 20012
rect 21771 19963 21813 19972
rect 21868 19769 21908 20131
rect 21964 20105 22004 20224
rect 22059 20180 22101 20189
rect 22059 20140 22060 20180
rect 22100 20140 22196 20180
rect 22059 20131 22101 20140
rect 21963 20096 22005 20105
rect 21963 20056 21964 20096
rect 22004 20056 22005 20096
rect 21963 20047 22005 20056
rect 22156 20096 22196 20140
rect 22444 20105 22484 20728
rect 22540 20768 22580 20777
rect 21964 19937 22004 20047
rect 22156 20045 22196 20056
rect 22252 20096 22292 20105
rect 21963 19928 22005 19937
rect 21963 19888 21964 19928
rect 22004 19888 22005 19928
rect 21963 19879 22005 19888
rect 21867 19760 21909 19769
rect 21867 19720 21868 19760
rect 21908 19720 21909 19760
rect 21867 19711 21909 19720
rect 21676 19088 21716 19097
rect 21100 18796 21332 18836
rect 21004 18712 21140 18752
rect 21003 18584 21045 18593
rect 21003 18544 21004 18584
rect 21044 18544 21045 18584
rect 21003 18535 21045 18544
rect 20908 18451 20948 18460
rect 21004 18416 21044 18535
rect 21100 18500 21140 18712
rect 21195 18584 21237 18593
rect 21195 18544 21196 18584
rect 21236 18544 21237 18584
rect 21195 18535 21237 18544
rect 21100 18451 21140 18460
rect 21004 18367 21044 18376
rect 21196 18248 21236 18535
rect 21004 18208 21236 18248
rect 20811 17744 20853 17753
rect 20811 17704 20812 17744
rect 20852 17704 20853 17744
rect 20811 17695 20853 17704
rect 20812 17610 20852 17695
rect 20811 17240 20853 17249
rect 20811 17200 20812 17240
rect 20852 17200 20853 17240
rect 20811 17191 20853 17200
rect 20812 17106 20852 17191
rect 20044 17072 20084 17081
rect 18315 16988 18357 16997
rect 18315 16948 18316 16988
rect 18356 16948 18357 16988
rect 18315 16939 18357 16948
rect 18795 16988 18837 16997
rect 18795 16948 18796 16988
rect 18836 16948 18837 16988
rect 18795 16939 18837 16948
rect 17547 16904 17589 16913
rect 17547 16864 17548 16904
rect 17588 16864 17589 16904
rect 17547 16855 17589 16864
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 17547 16232 17589 16241
rect 18604 16232 18644 16241
rect 17547 16192 17548 16232
rect 17588 16192 17589 16232
rect 17547 16183 17589 16192
rect 18508 16192 18604 16232
rect 16779 15896 16821 15905
rect 16779 15856 16780 15896
rect 16820 15856 16821 15896
rect 16779 15847 16821 15856
rect 16683 15560 16725 15569
rect 16683 15520 16684 15560
rect 16724 15520 16725 15560
rect 16683 15511 16725 15520
rect 16780 15560 16820 15569
rect 16684 15426 16724 15511
rect 16780 15233 16820 15520
rect 16971 15308 17013 15317
rect 16971 15268 16972 15308
rect 17012 15268 17013 15308
rect 16971 15259 17013 15268
rect 16779 15224 16821 15233
rect 16779 15184 16780 15224
rect 16820 15184 16821 15224
rect 16779 15175 16821 15184
rect 16972 15174 17012 15259
rect 16395 15140 16437 15149
rect 16395 15100 16396 15140
rect 16436 15100 16437 15140
rect 16395 15091 16437 15100
rect 16396 14636 16436 15091
rect 17548 14972 17588 16183
rect 18508 15737 18548 16192
rect 18604 16183 18644 16192
rect 18699 16232 18741 16241
rect 18699 16192 18700 16232
rect 18740 16192 18741 16232
rect 18699 16183 18741 16192
rect 18700 15980 18740 16183
rect 18604 15940 18740 15980
rect 18507 15728 18549 15737
rect 18507 15688 18508 15728
rect 18548 15688 18549 15728
rect 18507 15679 18549 15688
rect 18604 15560 18644 15940
rect 18604 15511 18644 15520
rect 18699 15560 18741 15569
rect 18699 15520 18700 15560
rect 18740 15520 18741 15560
rect 18699 15511 18741 15520
rect 18700 15426 18740 15511
rect 18796 15401 18836 16939
rect 20044 16904 20084 17032
rect 20332 17072 20372 17081
rect 20524 17072 20564 17081
rect 20372 17032 20468 17072
rect 20332 17023 20372 17032
rect 20332 16904 20372 16913
rect 20044 16864 20332 16904
rect 20332 16855 20372 16864
rect 18988 16820 19028 16829
rect 18891 16400 18933 16409
rect 18891 16360 18892 16400
rect 18932 16360 18933 16400
rect 18891 16351 18933 16360
rect 18892 16232 18932 16351
rect 18988 16325 19028 16780
rect 20332 16409 20372 16494
rect 20428 16484 20468 17032
rect 20524 16568 20564 17032
rect 20620 17072 20660 17081
rect 20620 16736 20660 17032
rect 20715 17072 20757 17081
rect 20715 17032 20716 17072
rect 20756 17032 20757 17072
rect 20715 17023 20757 17032
rect 20907 17072 20949 17081
rect 20907 17032 20908 17072
rect 20948 17032 20949 17072
rect 20907 17023 20949 17032
rect 21004 17072 21044 18208
rect 21004 17023 21044 17032
rect 21100 17072 21140 17081
rect 21292 17072 21332 18796
rect 21676 18593 21716 19048
rect 21868 18929 21908 19711
rect 21963 19508 22005 19517
rect 21963 19468 21964 19508
rect 22004 19468 22005 19508
rect 21963 19459 22005 19468
rect 21867 18920 21909 18929
rect 21867 18880 21868 18920
rect 21908 18880 21909 18920
rect 21867 18871 21909 18880
rect 21388 18584 21428 18593
rect 21388 18005 21428 18544
rect 21675 18584 21717 18593
rect 21675 18544 21676 18584
rect 21716 18544 21717 18584
rect 21675 18535 21717 18544
rect 21867 18500 21909 18509
rect 21867 18460 21868 18500
rect 21908 18460 21909 18500
rect 21867 18451 21909 18460
rect 21387 17996 21429 18005
rect 21387 17956 21388 17996
rect 21428 17956 21429 17996
rect 21387 17947 21429 17956
rect 21483 17912 21525 17921
rect 21483 17872 21484 17912
rect 21524 17872 21525 17912
rect 21483 17863 21525 17872
rect 21484 17744 21524 17863
rect 21676 17744 21716 17753
rect 21484 17695 21524 17704
rect 21580 17704 21676 17744
rect 21140 17032 21332 17072
rect 21484 17072 21524 17081
rect 21100 17023 21140 17032
rect 20908 16938 20948 17023
rect 20620 16696 21428 16736
rect 20524 16528 21044 16568
rect 20428 16444 20660 16484
rect 19275 16400 19317 16409
rect 19275 16360 19276 16400
rect 19316 16360 19317 16400
rect 19275 16351 19317 16360
rect 20139 16400 20181 16409
rect 20139 16360 20140 16400
rect 20180 16360 20181 16400
rect 20139 16351 20181 16360
rect 20331 16400 20373 16409
rect 20331 16360 20332 16400
rect 20372 16360 20373 16400
rect 20331 16351 20373 16360
rect 18987 16316 19029 16325
rect 18987 16276 18988 16316
rect 19028 16276 19029 16316
rect 18987 16267 19029 16276
rect 18892 16183 18932 16192
rect 19083 16232 19125 16241
rect 19083 16192 19084 16232
rect 19124 16192 19125 16232
rect 19083 16183 19125 16192
rect 19084 16148 19124 16183
rect 19084 16097 19124 16108
rect 19179 16148 19221 16157
rect 19179 16108 19180 16148
rect 19220 16108 19221 16148
rect 19179 16099 19221 16108
rect 19084 15644 19124 15653
rect 18892 15604 19084 15644
rect 18892 15560 18932 15604
rect 19084 15595 19124 15604
rect 19180 15569 19220 16099
rect 18892 15511 18932 15520
rect 19179 15560 19221 15569
rect 19179 15520 19180 15560
rect 19220 15520 19221 15560
rect 19179 15511 19221 15520
rect 19276 15560 19316 16351
rect 19372 16232 19412 16243
rect 19372 16157 19412 16192
rect 19659 16232 19701 16241
rect 19659 16192 19660 16232
rect 19700 16192 19701 16232
rect 19659 16183 19701 16192
rect 19371 16148 19413 16157
rect 19371 16108 19372 16148
rect 19412 16108 19413 16148
rect 19371 16099 19413 16108
rect 19660 16098 19700 16183
rect 19852 16157 19892 16242
rect 20140 16190 20180 16351
rect 20236 16316 20276 16325
rect 20236 16241 20276 16276
rect 20428 16316 20468 16325
rect 19851 16148 19893 16157
rect 19851 16108 19852 16148
rect 19892 16108 19893 16148
rect 19851 16099 19893 16108
rect 20228 16232 20276 16241
rect 20228 16192 20229 16232
rect 20269 16192 20276 16232
rect 20331 16232 20373 16241
rect 20331 16192 20332 16232
rect 20372 16192 20373 16232
rect 20228 16183 20270 16192
rect 20331 16183 20373 16192
rect 19947 16064 19989 16073
rect 19947 16024 19948 16064
rect 19988 16024 19989 16064
rect 19947 16015 19989 16024
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 19660 15746 19892 15786
rect 19371 15728 19413 15737
rect 19660 15728 19700 15746
rect 19371 15688 19372 15728
rect 19412 15688 19413 15728
rect 19371 15679 19413 15688
rect 19657 15688 19700 15728
rect 19852 15728 19892 15746
rect 19372 15594 19412 15679
rect 19564 15644 19604 15655
rect 19564 15569 19604 15604
rect 19276 15511 19316 15520
rect 19563 15560 19605 15569
rect 19563 15520 19564 15560
rect 19604 15520 19605 15560
rect 19657 15560 19697 15688
rect 19852 15679 19892 15688
rect 19756 15560 19796 15569
rect 19948 15560 19988 16015
rect 20140 15989 20180 16150
rect 20139 15980 20181 15989
rect 20139 15940 20140 15980
rect 20180 15940 20181 15980
rect 20139 15931 20181 15940
rect 20332 15896 20372 16183
rect 20428 16157 20468 16276
rect 20523 16316 20565 16325
rect 20523 16276 20524 16316
rect 20564 16276 20565 16316
rect 20523 16267 20565 16276
rect 20524 16232 20564 16267
rect 20524 16181 20564 16192
rect 20427 16148 20469 16157
rect 20427 16108 20428 16148
rect 20468 16108 20469 16148
rect 20427 16099 20469 16108
rect 20620 15905 20660 16444
rect 20715 16232 20757 16241
rect 20715 16192 20716 16232
rect 20756 16192 20757 16232
rect 20715 16183 20757 16192
rect 20812 16232 20852 16241
rect 20716 16098 20756 16183
rect 20812 16073 20852 16192
rect 20908 16232 20948 16241
rect 20811 16064 20853 16073
rect 20811 16024 20812 16064
rect 20852 16024 20853 16064
rect 20811 16015 20853 16024
rect 20236 15856 20372 15896
rect 20619 15896 20661 15905
rect 20619 15856 20620 15896
rect 20660 15856 20661 15896
rect 20236 15737 20276 15856
rect 20619 15847 20661 15856
rect 20235 15728 20277 15737
rect 20235 15688 20236 15728
rect 20276 15688 20277 15728
rect 20235 15679 20277 15688
rect 20332 15728 20372 15737
rect 20908 15728 20948 16192
rect 21004 16232 21044 16528
rect 21388 16400 21428 16696
rect 21388 16351 21428 16360
rect 21292 16316 21332 16325
rect 21004 16183 21044 16192
rect 21195 16232 21237 16241
rect 21195 16192 21196 16232
rect 21236 16192 21237 16232
rect 21195 16183 21237 16192
rect 21196 16098 21236 16183
rect 21003 15896 21045 15905
rect 21003 15856 21004 15896
rect 21044 15856 21045 15896
rect 21003 15847 21045 15856
rect 20372 15688 20948 15728
rect 20332 15679 20372 15688
rect 21004 15644 21044 15847
rect 21292 15821 21332 16276
rect 21484 16316 21524 17032
rect 21291 15812 21333 15821
rect 21291 15772 21292 15812
rect 21332 15772 21333 15812
rect 21291 15763 21333 15772
rect 21484 15737 21524 16276
rect 21580 16232 21620 17704
rect 21676 17695 21716 17704
rect 21868 17240 21908 18451
rect 21964 17249 22004 19459
rect 22155 19424 22197 19433
rect 22155 19384 22156 19424
rect 22196 19384 22197 19424
rect 22155 19375 22197 19384
rect 22156 19256 22196 19375
rect 22156 19207 22196 19216
rect 22252 18929 22292 20056
rect 22443 20096 22485 20105
rect 22443 20056 22444 20096
rect 22484 20056 22485 20096
rect 22443 20047 22485 20056
rect 22540 19517 22580 20728
rect 22635 20600 22677 20609
rect 22635 20560 22636 20600
rect 22676 20560 22677 20600
rect 22635 20551 22677 20560
rect 22636 20466 22676 20551
rect 23020 20180 23060 22492
rect 23115 22364 23157 22373
rect 23115 22324 23116 22364
rect 23156 22324 23157 22364
rect 23115 22315 23157 22324
rect 23116 22280 23156 22315
rect 23116 22229 23156 22240
rect 23308 22280 23348 22735
rect 23499 22532 23541 22541
rect 23499 22492 23500 22532
rect 23540 22492 23541 22532
rect 23499 22483 23541 22492
rect 23308 22231 23348 22240
rect 23500 22280 23540 22483
rect 23500 22231 23540 22240
rect 23596 22280 23636 22735
rect 23787 22700 23829 22709
rect 23787 22660 23788 22700
rect 23828 22660 23829 22700
rect 23787 22651 23829 22660
rect 23788 22532 23828 22651
rect 23883 22616 23925 22625
rect 23883 22576 23884 22616
rect 23924 22576 23925 22616
rect 23883 22567 23925 22576
rect 23788 22483 23828 22492
rect 23212 22196 23252 22205
rect 23212 22112 23252 22156
rect 23596 22112 23636 22240
rect 23691 22280 23733 22289
rect 23691 22240 23692 22280
rect 23732 22240 23733 22280
rect 23691 22231 23733 22240
rect 23788 22280 23828 22289
rect 23884 22280 23924 22567
rect 23828 22240 23924 22280
rect 23788 22231 23828 22240
rect 23212 22072 23636 22112
rect 23692 21608 23732 22231
rect 23692 21559 23732 21568
rect 23403 21440 23445 21449
rect 23403 21400 23404 21440
rect 23444 21400 23445 21440
rect 23884 21440 23924 22240
rect 23980 22280 24020 23080
rect 24076 22709 24116 23743
rect 24844 23717 24884 23752
rect 24843 23708 24885 23717
rect 24843 23668 24844 23708
rect 24884 23668 24885 23708
rect 24843 23659 24885 23668
rect 24171 23624 24213 23633
rect 24748 23624 24788 23633
rect 24171 23584 24172 23624
rect 24212 23584 24213 23624
rect 24171 23575 24213 23584
rect 24268 23584 24748 23624
rect 24075 22700 24117 22709
rect 24075 22660 24076 22700
rect 24116 22660 24117 22700
rect 24075 22651 24117 22660
rect 23980 22231 24020 22240
rect 24172 22280 24212 23575
rect 24172 22231 24212 22240
rect 24268 22280 24308 23584
rect 24748 23575 24788 23584
rect 24555 23372 24597 23381
rect 24555 23332 24556 23372
rect 24596 23332 24597 23372
rect 24555 23323 24597 23332
rect 24364 23120 24404 23129
rect 24364 22373 24404 23080
rect 24459 23120 24501 23129
rect 24459 23080 24460 23120
rect 24500 23080 24501 23120
rect 24459 23071 24501 23080
rect 24460 22986 24500 23071
rect 24556 22793 24596 23323
rect 24747 23120 24789 23129
rect 24747 23080 24748 23120
rect 24788 23080 24789 23120
rect 24747 23071 24789 23080
rect 24748 23036 24788 23071
rect 24748 22985 24788 22996
rect 24652 22868 24692 22877
rect 24555 22784 24597 22793
rect 24555 22744 24556 22784
rect 24596 22744 24597 22784
rect 24555 22735 24597 22744
rect 24459 22532 24501 22541
rect 24459 22492 24460 22532
rect 24500 22492 24501 22532
rect 24459 22483 24501 22492
rect 24460 22398 24500 22483
rect 24555 22448 24597 22457
rect 24555 22408 24556 22448
rect 24596 22408 24597 22448
rect 24555 22399 24597 22408
rect 24652 22448 24692 22828
rect 24747 22868 24789 22877
rect 24844 22868 24884 23659
rect 24747 22828 24748 22868
rect 24788 22828 24884 22868
rect 24747 22819 24789 22828
rect 24652 22399 24692 22408
rect 24363 22364 24405 22373
rect 24363 22324 24364 22364
rect 24404 22324 24405 22364
rect 24363 22315 24405 22324
rect 24268 22231 24308 22240
rect 24076 22112 24116 22121
rect 24556 22112 24596 22399
rect 24652 22280 24692 22291
rect 24652 22205 24692 22240
rect 24651 22196 24693 22205
rect 24651 22156 24652 22196
rect 24692 22156 24693 22196
rect 24651 22147 24693 22156
rect 24748 22121 24788 22819
rect 24940 22784 24980 24004
rect 25324 23801 25364 23886
rect 25036 23792 25076 23801
rect 25228 23792 25268 23801
rect 25076 23752 25172 23792
rect 25036 23743 25076 23752
rect 25035 23624 25077 23633
rect 25035 23584 25036 23624
rect 25076 23584 25077 23624
rect 25035 23575 25077 23584
rect 25036 23490 25076 23575
rect 25035 23372 25077 23381
rect 25132 23372 25172 23752
rect 25228 23381 25268 23752
rect 25323 23792 25365 23801
rect 25323 23752 25324 23792
rect 25364 23752 25365 23792
rect 25323 23743 25365 23752
rect 25516 23624 25556 23633
rect 25324 23584 25516 23624
rect 25035 23332 25036 23372
rect 25076 23332 25172 23372
rect 25227 23372 25269 23381
rect 25227 23332 25228 23372
rect 25268 23332 25269 23372
rect 25035 23323 25077 23332
rect 25227 23323 25269 23332
rect 25324 23204 25364 23584
rect 25516 23575 25556 23584
rect 25612 23456 25652 24592
rect 25708 24583 25748 24592
rect 25900 24632 25940 24641
rect 25940 24592 26036 24632
rect 25900 24583 25940 24592
rect 25803 24212 25845 24221
rect 25803 24172 25804 24212
rect 25844 24172 25845 24212
rect 25803 24163 25845 24172
rect 25707 23792 25749 23801
rect 25707 23752 25708 23792
rect 25748 23752 25749 23792
rect 25707 23743 25749 23752
rect 25804 23792 25844 24163
rect 25996 23960 26036 24592
rect 25708 23658 25748 23743
rect 25516 23416 25652 23456
rect 25419 23372 25461 23381
rect 25419 23332 25420 23372
rect 25460 23332 25461 23372
rect 25419 23323 25461 23332
rect 25036 23164 25364 23204
rect 25036 23120 25076 23164
rect 25036 23071 25076 23080
rect 25420 23120 25460 23323
rect 25420 23071 25460 23080
rect 25131 23036 25173 23045
rect 25131 22996 25132 23036
rect 25172 22996 25173 23036
rect 25131 22987 25173 22996
rect 25323 23036 25365 23045
rect 25323 22996 25324 23036
rect 25364 22996 25365 23036
rect 25323 22987 25365 22996
rect 25035 22952 25077 22961
rect 25035 22912 25036 22952
rect 25076 22912 25077 22952
rect 25035 22903 25077 22912
rect 24844 22744 24980 22784
rect 24076 21617 24116 22072
rect 24268 22072 24596 22112
rect 24747 22112 24789 22121
rect 24747 22072 24748 22112
rect 24788 22072 24789 22112
rect 24075 21608 24117 21617
rect 24075 21568 24076 21608
rect 24116 21568 24117 21608
rect 24075 21559 24117 21568
rect 24172 21440 24212 21449
rect 23884 21400 24172 21440
rect 23403 21391 23445 21400
rect 24172 21391 24212 21400
rect 22828 20140 23060 20180
rect 22636 19844 22676 19853
rect 22539 19508 22581 19517
rect 22539 19468 22540 19508
rect 22580 19468 22581 19508
rect 22539 19459 22581 19468
rect 22636 19433 22676 19804
rect 22635 19424 22677 19433
rect 22635 19384 22636 19424
rect 22676 19384 22677 19424
rect 22635 19375 22677 19384
rect 22828 19349 22868 20140
rect 23404 20105 23444 21391
rect 24268 21272 24308 22072
rect 24747 22063 24789 22072
rect 24363 21692 24405 21701
rect 24363 21652 24364 21692
rect 24404 21652 24405 21692
rect 24363 21643 24405 21652
rect 24364 21608 24404 21643
rect 24364 21557 24404 21568
rect 24460 21608 24500 21617
rect 24460 21449 24500 21568
rect 24844 21524 24884 22744
rect 25036 22700 25076 22903
rect 24940 22660 25076 22700
rect 24940 22280 24980 22660
rect 25132 22541 25172 22987
rect 25228 22952 25268 22961
rect 25228 22784 25268 22912
rect 25324 22902 25364 22987
rect 25516 22784 25556 23416
rect 25804 23372 25844 23752
rect 25708 23332 25844 23372
rect 25900 23920 26036 23960
rect 26859 23960 26901 23969
rect 26859 23920 26860 23960
rect 26900 23920 26901 23960
rect 25708 23288 25748 23332
rect 25695 23248 25748 23288
rect 25900 23288 25940 23920
rect 26859 23911 26901 23920
rect 26667 23876 26709 23885
rect 26667 23836 26668 23876
rect 26708 23836 26709 23876
rect 26667 23827 26709 23836
rect 25611 23204 25653 23213
rect 25611 23164 25612 23204
rect 25652 23164 25653 23204
rect 25611 23155 25653 23164
rect 25228 22744 25556 22784
rect 25612 23120 25652 23155
rect 25695 23129 25735 23248
rect 25900 23239 25940 23248
rect 25996 23792 26036 23801
rect 25695 23120 25748 23129
rect 25695 23087 25708 23120
rect 25612 22709 25652 23080
rect 25708 23071 25748 23080
rect 25804 23120 25844 23129
rect 25844 23080 25940 23120
rect 25804 23071 25844 23080
rect 25900 22961 25940 23080
rect 25899 22952 25941 22961
rect 25899 22912 25900 22952
rect 25940 22912 25941 22952
rect 25899 22903 25941 22912
rect 25611 22700 25653 22709
rect 25611 22660 25612 22700
rect 25652 22660 25653 22700
rect 25611 22651 25653 22660
rect 25131 22532 25173 22541
rect 25131 22492 25132 22532
rect 25172 22492 25173 22532
rect 25131 22483 25173 22492
rect 25131 22364 25173 22373
rect 25131 22324 25132 22364
rect 25172 22324 25173 22364
rect 25131 22315 25173 22324
rect 24940 22231 24980 22240
rect 25036 22280 25076 22289
rect 25036 22121 25076 22240
rect 25035 22112 25077 22121
rect 25035 22072 25036 22112
rect 25076 22072 25077 22112
rect 25035 22063 25077 22072
rect 25036 21701 25076 22063
rect 25035 21692 25077 21701
rect 25035 21652 25036 21692
rect 25076 21652 25077 21692
rect 25035 21643 25077 21652
rect 24556 21484 24844 21524
rect 24459 21440 24501 21449
rect 24459 21400 24460 21440
rect 24500 21400 24501 21440
rect 24459 21391 24501 21400
rect 24172 21232 24308 21272
rect 23308 20096 23348 20105
rect 22827 19340 22869 19349
rect 22827 19300 22828 19340
rect 22868 19300 22869 19340
rect 22827 19291 22869 19300
rect 22539 19256 22581 19265
rect 22539 19216 22540 19256
rect 22580 19216 22581 19256
rect 22539 19207 22581 19216
rect 22540 19122 22580 19207
rect 23308 18929 23348 20056
rect 23403 20096 23445 20105
rect 23403 20056 23404 20096
rect 23444 20056 23445 20096
rect 23403 20047 23445 20056
rect 24076 20096 24116 20105
rect 24172 20096 24212 21232
rect 24460 20768 24500 20777
rect 24556 20768 24596 21484
rect 24844 21475 24884 21484
rect 25035 21440 25077 21449
rect 25035 21400 25036 21440
rect 25076 21400 25077 21440
rect 25035 21391 25077 21400
rect 25036 21306 25076 21391
rect 25036 20936 25076 20945
rect 25132 20936 25172 22315
rect 25420 22289 25460 22374
rect 25419 22280 25461 22289
rect 25419 22240 25420 22280
rect 25460 22240 25461 22280
rect 25419 22231 25461 22240
rect 25996 22121 26036 23752
rect 26091 23792 26133 23801
rect 26091 23752 26092 23792
rect 26132 23752 26133 23792
rect 26091 23743 26133 23752
rect 26284 23792 26324 23801
rect 26476 23792 26516 23801
rect 26324 23752 26420 23792
rect 26284 23743 26324 23752
rect 26092 23297 26132 23743
rect 26187 23624 26229 23633
rect 26187 23584 26188 23624
rect 26228 23584 26229 23624
rect 26187 23575 26229 23584
rect 26284 23624 26324 23633
rect 26091 23288 26133 23297
rect 26091 23248 26092 23288
rect 26132 23248 26133 23288
rect 26091 23239 26133 23248
rect 26091 23120 26133 23129
rect 26091 23080 26092 23120
rect 26132 23080 26133 23120
rect 26091 23071 26133 23080
rect 26188 23120 26228 23575
rect 26284 23381 26324 23584
rect 26283 23372 26325 23381
rect 26283 23332 26284 23372
rect 26324 23332 26325 23372
rect 26283 23323 26325 23332
rect 26380 23288 26420 23752
rect 26476 23549 26516 23752
rect 26668 23792 26708 23827
rect 26668 23741 26708 23752
rect 26571 23708 26613 23717
rect 26571 23668 26572 23708
rect 26612 23668 26613 23708
rect 26571 23659 26613 23668
rect 26572 23574 26612 23659
rect 26475 23540 26517 23549
rect 26475 23500 26476 23540
rect 26516 23500 26517 23540
rect 26475 23491 26517 23500
rect 26380 23248 26516 23288
rect 26092 22986 26132 23071
rect 26091 22700 26133 22709
rect 26091 22660 26092 22700
rect 26132 22660 26133 22700
rect 26091 22651 26133 22660
rect 26092 22532 26132 22651
rect 26092 22483 26132 22492
rect 26188 22205 26228 23080
rect 26284 23204 26324 23213
rect 26284 23045 26324 23164
rect 26380 23120 26420 23129
rect 26283 23036 26325 23045
rect 26283 22996 26284 23036
rect 26324 22996 26325 23036
rect 26283 22987 26325 22996
rect 26380 22877 26420 23080
rect 26379 22868 26421 22877
rect 26379 22828 26380 22868
rect 26420 22828 26421 22868
rect 26379 22819 26421 22828
rect 26476 22205 26516 23248
rect 26763 23204 26805 23213
rect 26763 23164 26764 23204
rect 26804 23164 26805 23204
rect 26763 23155 26805 23164
rect 26572 23120 26612 23129
rect 26572 22289 26612 23080
rect 26668 23120 26708 23129
rect 26668 22961 26708 23080
rect 26764 23120 26804 23155
rect 26764 23069 26804 23080
rect 26860 23120 26900 23911
rect 26860 23071 26900 23080
rect 26667 22952 26709 22961
rect 26667 22912 26668 22952
rect 26708 22912 26709 22952
rect 26667 22903 26709 22912
rect 26571 22280 26613 22289
rect 26571 22240 26572 22280
rect 26612 22240 26613 22280
rect 26571 22231 26613 22240
rect 26187 22196 26229 22205
rect 26187 22156 26188 22196
rect 26228 22156 26229 22196
rect 26187 22147 26229 22156
rect 26475 22196 26517 22205
rect 26475 22156 26476 22196
rect 26516 22156 26517 22196
rect 26475 22147 26517 22156
rect 25227 22112 25269 22121
rect 25227 22072 25228 22112
rect 25268 22072 25269 22112
rect 25227 22063 25269 22072
rect 25995 22112 26037 22121
rect 25995 22072 25996 22112
rect 26036 22072 26037 22112
rect 25995 22063 26037 22072
rect 26092 22112 26132 22121
rect 25228 21978 25268 22063
rect 25419 22028 25461 22037
rect 25419 21988 25420 22028
rect 25460 21988 25461 22028
rect 25419 21979 25461 21988
rect 25323 21944 25365 21953
rect 25323 21904 25324 21944
rect 25364 21904 25365 21944
rect 25323 21895 25365 21904
rect 25227 21692 25269 21701
rect 25227 21652 25228 21692
rect 25268 21652 25269 21692
rect 25227 21643 25269 21652
rect 25324 21692 25364 21895
rect 25324 21643 25364 21652
rect 25228 21608 25268 21643
rect 25228 21557 25268 21568
rect 25420 21608 25460 21979
rect 25899 21944 25941 21953
rect 25899 21904 25900 21944
rect 25940 21904 25941 21944
rect 25899 21895 25941 21904
rect 25707 21776 25749 21785
rect 25707 21736 25708 21776
rect 25748 21736 25749 21776
rect 25707 21727 25749 21736
rect 25708 21642 25748 21727
rect 25420 21559 25460 21568
rect 25611 21608 25653 21617
rect 25611 21568 25612 21608
rect 25652 21568 25653 21608
rect 25611 21559 25653 21568
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 25803 21559 25845 21568
rect 25612 21474 25652 21559
rect 25707 21524 25749 21533
rect 25707 21484 25708 21524
rect 25748 21484 25749 21524
rect 25707 21475 25749 21484
rect 25515 21440 25557 21449
rect 25515 21400 25516 21440
rect 25556 21400 25557 21440
rect 25515 21391 25557 21400
rect 25076 20896 25172 20936
rect 25036 20887 25076 20896
rect 24500 20728 24596 20768
rect 24460 20719 24500 20728
rect 24844 20140 24980 20180
rect 24116 20056 24212 20096
rect 24268 20096 24308 20105
rect 24844 20096 24884 20140
rect 24308 20056 24788 20096
rect 23404 19256 23444 20047
rect 23500 19928 23540 19937
rect 23500 19265 23540 19888
rect 23404 19207 23444 19216
rect 23499 19256 23541 19265
rect 23499 19216 23500 19256
rect 23540 19216 23541 19256
rect 23499 19207 23541 19216
rect 22251 18920 22293 18929
rect 22251 18880 22252 18920
rect 22292 18880 22293 18920
rect 22251 18871 22293 18880
rect 23307 18920 23349 18929
rect 23307 18880 23308 18920
rect 23348 18880 23349 18920
rect 23307 18871 23349 18880
rect 24076 18761 24116 20056
rect 24268 20047 24308 20056
rect 24172 19844 24212 19853
rect 22060 18752 22100 18761
rect 23307 18752 23349 18761
rect 22100 18712 22580 18752
rect 22060 18703 22100 18712
rect 22251 18584 22293 18593
rect 22251 18544 22252 18584
rect 22292 18544 22293 18584
rect 22251 18535 22293 18544
rect 22252 17837 22292 18535
rect 22347 18500 22389 18509
rect 22347 18460 22348 18500
rect 22388 18460 22389 18500
rect 22347 18451 22389 18460
rect 22540 18500 22580 18712
rect 23307 18712 23308 18752
rect 23348 18712 23349 18752
rect 23307 18703 23349 18712
rect 24075 18752 24117 18761
rect 24075 18712 24076 18752
rect 24116 18712 24117 18752
rect 24075 18703 24117 18712
rect 23116 18668 23156 18677
rect 23020 18628 23116 18668
rect 22348 18366 22388 18451
rect 22444 18416 22484 18425
rect 22347 17996 22389 18005
rect 22347 17956 22348 17996
rect 22388 17956 22389 17996
rect 22347 17947 22389 17956
rect 22251 17828 22293 17837
rect 22251 17788 22252 17828
rect 22292 17788 22293 17828
rect 22251 17779 22293 17788
rect 21868 17191 21908 17200
rect 21963 17240 22005 17249
rect 21963 17200 21964 17240
rect 22004 17200 22005 17240
rect 21963 17191 22005 17200
rect 21867 17072 21909 17081
rect 22348 17072 22388 17947
rect 22444 17753 22484 18376
rect 22540 17996 22580 18460
rect 22636 18584 22676 18593
rect 22636 18425 22676 18544
rect 22635 18416 22677 18425
rect 22635 18376 22636 18416
rect 22676 18376 22677 18416
rect 22635 18367 22677 18376
rect 22540 17956 22676 17996
rect 22539 17828 22581 17837
rect 22539 17788 22540 17828
rect 22580 17788 22581 17828
rect 22539 17779 22581 17788
rect 22443 17744 22485 17753
rect 22443 17704 22444 17744
rect 22484 17704 22485 17744
rect 22443 17695 22485 17704
rect 22540 17744 22580 17779
rect 22540 17693 22580 17704
rect 22636 17081 22676 17956
rect 22923 17744 22965 17753
rect 22923 17704 22924 17744
rect 22964 17704 22965 17744
rect 22923 17695 22965 17704
rect 23020 17744 23060 18628
rect 23116 18619 23156 18628
rect 23308 18593 23348 18703
rect 23212 18584 23252 18593
rect 23187 18544 23212 18584
rect 23187 18542 23252 18544
rect 23116 18535 23252 18542
rect 23307 18584 23349 18593
rect 23307 18544 23308 18584
rect 23348 18544 23349 18584
rect 23307 18535 23349 18544
rect 23404 18584 23444 18593
rect 23499 18584 23541 18593
rect 23444 18544 23500 18584
rect 23540 18544 23541 18584
rect 23404 18535 23444 18544
rect 23499 18535 23541 18544
rect 23596 18584 23636 18593
rect 23116 18502 23227 18535
rect 23116 18080 23156 18502
rect 23308 18450 23348 18535
rect 23499 18164 23541 18173
rect 23499 18124 23500 18164
rect 23540 18124 23541 18164
rect 23499 18115 23541 18124
rect 23116 18040 23348 18080
rect 23020 17695 23060 17704
rect 22924 17610 22964 17695
rect 23116 17669 23156 17754
rect 23211 17744 23253 17753
rect 23211 17704 23212 17744
rect 23252 17704 23253 17744
rect 23211 17695 23253 17704
rect 23115 17660 23157 17669
rect 23115 17620 23116 17660
rect 23156 17620 23157 17660
rect 23115 17611 23157 17620
rect 23212 17610 23252 17695
rect 23115 17492 23157 17501
rect 23115 17452 23116 17492
rect 23156 17452 23157 17492
rect 23115 17443 23157 17452
rect 22540 17072 22580 17081
rect 21867 17032 21868 17072
rect 21908 17032 21909 17072
rect 21867 17023 21909 17032
rect 22060 17032 22540 17072
rect 21675 16820 21717 16829
rect 21675 16780 21676 16820
rect 21716 16780 21717 16820
rect 21675 16771 21717 16780
rect 21676 16686 21716 16771
rect 21771 16400 21813 16409
rect 21771 16360 21772 16400
rect 21812 16360 21813 16400
rect 21771 16351 21813 16360
rect 21580 16073 21620 16192
rect 21579 16064 21621 16073
rect 21579 16024 21580 16064
rect 21620 16024 21621 16064
rect 21579 16015 21621 16024
rect 21772 15989 21812 16351
rect 21771 15980 21813 15989
rect 21771 15940 21772 15980
rect 21812 15940 21813 15980
rect 21868 15980 21908 17023
rect 21964 16409 22004 16494
rect 21963 16400 22005 16409
rect 21963 16360 21964 16400
rect 22004 16360 22005 16400
rect 21963 16351 22005 16360
rect 21964 16232 22004 16241
rect 22060 16232 22100 17032
rect 22540 17023 22580 17032
rect 22635 17072 22677 17081
rect 22635 17032 22636 17072
rect 22676 17032 22677 17072
rect 22635 17023 22677 17032
rect 22004 16192 22100 16232
rect 22156 16400 22196 16409
rect 22156 16232 22196 16360
rect 22443 16316 22485 16325
rect 22443 16276 22444 16316
rect 22484 16276 22485 16316
rect 22443 16267 22485 16276
rect 22347 16232 22389 16241
rect 22156 16192 22348 16232
rect 22388 16192 22389 16232
rect 21964 16183 22004 16192
rect 22347 16183 22389 16192
rect 22444 16232 22484 16267
rect 22348 16098 22388 16183
rect 22444 16181 22484 16192
rect 22636 16232 22676 16241
rect 22636 16157 22676 16192
rect 22828 16232 22868 16243
rect 22828 16157 22868 16192
rect 22923 16232 22965 16241
rect 22923 16192 22924 16232
rect 22964 16192 22965 16232
rect 22923 16183 22965 16192
rect 22635 16148 22677 16157
rect 22635 16108 22636 16148
rect 22676 16108 22677 16148
rect 22635 16099 22677 16108
rect 22827 16148 22869 16157
rect 22827 16108 22828 16148
rect 22868 16108 22869 16148
rect 22827 16099 22869 16108
rect 22636 16097 22676 16099
rect 22924 16098 22964 16183
rect 22539 16064 22581 16073
rect 22539 16024 22540 16064
rect 22580 16024 22581 16064
rect 22539 16015 22581 16024
rect 23116 16064 23156 17443
rect 23308 17240 23348 18040
rect 23404 17744 23444 17753
rect 23404 17501 23444 17704
rect 23500 17744 23540 18115
rect 23596 17837 23636 18544
rect 23692 18584 23732 18593
rect 23692 18005 23732 18544
rect 23788 18584 23828 18593
rect 23788 18089 23828 18544
rect 23883 18584 23925 18593
rect 23883 18544 23884 18584
rect 23924 18544 23925 18584
rect 23883 18535 23925 18544
rect 24075 18584 24117 18593
rect 24075 18544 24076 18584
rect 24116 18544 24117 18584
rect 24075 18535 24117 18544
rect 23787 18080 23829 18089
rect 23787 18040 23788 18080
rect 23828 18040 23829 18080
rect 23787 18031 23829 18040
rect 23691 17996 23733 18005
rect 23691 17956 23692 17996
rect 23732 17956 23733 17996
rect 23691 17947 23733 17956
rect 23884 17912 23924 18535
rect 24076 18450 24116 18535
rect 24172 18173 24212 19804
rect 24556 19256 24596 19265
rect 24556 18593 24596 19216
rect 24748 18752 24788 20056
rect 24844 20047 24884 20056
rect 24843 19928 24885 19937
rect 24843 19888 24844 19928
rect 24884 19888 24885 19928
rect 24843 19879 24885 19888
rect 24844 19794 24884 19879
rect 24940 19349 24980 20140
rect 25036 19853 25076 19938
rect 25035 19844 25077 19853
rect 25035 19804 25036 19844
rect 25076 19804 25077 19844
rect 25035 19795 25077 19804
rect 24939 19340 24981 19349
rect 24939 19300 24940 19340
rect 24980 19300 24981 19340
rect 24939 19291 24981 19300
rect 25132 19004 25172 20896
rect 25420 20189 25460 20199
rect 25227 20180 25269 20189
rect 25227 20140 25228 20180
rect 25268 20140 25269 20180
rect 25227 20131 25269 20140
rect 25419 20180 25461 20189
rect 25419 20140 25420 20180
rect 25460 20140 25461 20180
rect 25419 20131 25461 20140
rect 25228 19937 25268 20131
rect 25420 20104 25460 20131
rect 25420 20055 25460 20064
rect 25227 19928 25269 19937
rect 25227 19888 25228 19928
rect 25268 19888 25269 19928
rect 25227 19879 25269 19888
rect 24748 18703 24788 18712
rect 24844 18964 25172 19004
rect 25324 19844 25364 19853
rect 24555 18584 24597 18593
rect 24555 18544 24556 18584
rect 24596 18544 24597 18584
rect 24555 18535 24597 18544
rect 24748 18332 24788 18341
rect 24460 18292 24748 18332
rect 24171 18164 24213 18173
rect 24171 18124 24172 18164
rect 24212 18124 24213 18164
rect 24171 18115 24213 18124
rect 24364 17996 24404 18005
rect 24172 17956 24364 17996
rect 23788 17872 23924 17912
rect 23979 17912 24021 17921
rect 23979 17872 23980 17912
rect 24020 17872 24021 17912
rect 23595 17828 23637 17837
rect 23595 17788 23596 17828
rect 23636 17788 23637 17828
rect 23595 17779 23637 17788
rect 23500 17695 23540 17704
rect 23691 17744 23733 17753
rect 23691 17704 23692 17744
rect 23732 17704 23733 17744
rect 23691 17695 23733 17704
rect 23595 17660 23637 17669
rect 23595 17620 23596 17660
rect 23636 17620 23637 17660
rect 23595 17611 23637 17620
rect 23499 17576 23541 17585
rect 23499 17536 23500 17576
rect 23540 17536 23541 17576
rect 23499 17527 23541 17536
rect 23403 17492 23445 17501
rect 23403 17452 23404 17492
rect 23444 17452 23445 17492
rect 23403 17443 23445 17452
rect 23404 17240 23444 17249
rect 23308 17200 23404 17240
rect 23404 17191 23444 17200
rect 23500 17072 23540 17527
rect 23596 17526 23636 17611
rect 23692 17610 23732 17695
rect 23500 16997 23540 17032
rect 23596 17072 23636 17081
rect 23499 16988 23541 16997
rect 23499 16948 23500 16988
rect 23540 16948 23541 16988
rect 23499 16939 23541 16948
rect 23212 16820 23252 16829
rect 23252 16780 23444 16820
rect 23212 16771 23252 16780
rect 23211 16232 23253 16241
rect 23211 16192 23212 16232
rect 23252 16192 23253 16232
rect 23211 16183 23253 16192
rect 23404 16232 23444 16780
rect 23596 16325 23636 17032
rect 23692 17072 23732 17081
rect 23595 16316 23637 16325
rect 23595 16276 23596 16316
rect 23636 16276 23637 16316
rect 23595 16267 23637 16276
rect 23404 16183 23444 16192
rect 23116 16015 23156 16024
rect 21868 15940 22388 15980
rect 21771 15931 21813 15940
rect 21676 15759 21716 15768
rect 21483 15728 21525 15737
rect 21483 15688 21484 15728
rect 21524 15688 21525 15728
rect 21771 15728 21813 15737
rect 21716 15719 21772 15728
rect 21676 15688 21772 15719
rect 21812 15688 21813 15728
rect 21483 15679 21525 15688
rect 21771 15679 21813 15688
rect 21004 15595 21044 15604
rect 19657 15520 19700 15560
rect 19563 15511 19605 15520
rect 19371 15476 19413 15485
rect 19371 15436 19372 15476
rect 19412 15436 19413 15476
rect 19371 15427 19413 15436
rect 18795 15392 18837 15401
rect 18795 15352 18796 15392
rect 18836 15352 18837 15392
rect 18795 15343 18837 15352
rect 17835 15308 17877 15317
rect 17835 15268 17836 15308
rect 17876 15268 17877 15308
rect 17835 15259 17877 15268
rect 18892 15308 18932 15317
rect 17643 15056 17685 15065
rect 17643 15016 17644 15056
rect 17684 15016 17685 15056
rect 17643 15007 17685 15016
rect 17548 14923 17588 14932
rect 16875 14720 16917 14729
rect 16875 14680 16876 14720
rect 16916 14680 16917 14720
rect 16875 14671 16917 14680
rect 17164 14720 17204 14729
rect 16107 14048 16149 14057
rect 16107 14008 16108 14048
rect 16148 14008 16149 14048
rect 16107 13999 16149 14008
rect 16396 13889 16436 14596
rect 16876 14141 16916 14671
rect 16971 14552 17013 14561
rect 16971 14512 16972 14552
rect 17012 14512 17013 14552
rect 16971 14503 17013 14512
rect 16875 14132 16917 14141
rect 16875 14092 16876 14132
rect 16916 14092 16917 14132
rect 16875 14083 16917 14092
rect 16876 14048 16916 14083
rect 16876 13998 16916 14008
rect 16395 13880 16437 13889
rect 16395 13840 16396 13880
rect 16436 13840 16437 13880
rect 16395 13831 16437 13840
rect 16299 13796 16341 13805
rect 16299 13756 16300 13796
rect 16340 13756 16341 13796
rect 16299 13747 16341 13756
rect 16300 13662 16340 13747
rect 16299 13460 16341 13469
rect 16299 13420 16300 13460
rect 16340 13420 16341 13460
rect 16299 13411 16341 13420
rect 15915 13376 15957 13385
rect 15915 13336 15916 13376
rect 15956 13336 15957 13376
rect 15915 13327 15957 13336
rect 16300 13326 16340 13411
rect 16012 13208 16052 13217
rect 15915 13040 15957 13049
rect 15915 13000 15916 13040
rect 15956 13000 15957 13040
rect 15915 12991 15957 13000
rect 15916 12536 15956 12991
rect 16012 12797 16052 13168
rect 16108 13208 16148 13217
rect 16108 13049 16148 13168
rect 16299 13208 16341 13217
rect 16299 13168 16300 13208
rect 16340 13168 16341 13208
rect 16299 13159 16341 13168
rect 16972 13208 17012 14503
rect 17067 14048 17109 14057
rect 17067 14008 17068 14048
rect 17108 14008 17109 14048
rect 17067 13999 17109 14008
rect 17068 13469 17108 13999
rect 17067 13460 17109 13469
rect 17067 13420 17068 13460
rect 17108 13420 17109 13460
rect 17067 13411 17109 13420
rect 16972 13159 17012 13168
rect 17068 13208 17108 13411
rect 17164 13376 17204 14680
rect 17259 14720 17301 14729
rect 17259 14680 17260 14720
rect 17300 14680 17301 14720
rect 17259 14671 17301 14680
rect 17548 14720 17588 14729
rect 17260 14057 17300 14671
rect 17355 14552 17397 14561
rect 17355 14512 17356 14552
rect 17396 14512 17397 14552
rect 17355 14503 17397 14512
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17356 14048 17396 14503
rect 17548 14216 17588 14680
rect 17644 14720 17684 15007
rect 17644 14671 17684 14680
rect 17836 14720 17876 15259
rect 18699 15224 18741 15233
rect 18699 15184 18700 15224
rect 18740 15184 18741 15224
rect 18699 15175 18741 15184
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 17931 14888 17973 14897
rect 17931 14848 17932 14888
rect 17972 14848 17973 14888
rect 17931 14839 17973 14848
rect 17836 14671 17876 14680
rect 17932 14720 17972 14839
rect 18033 14720 18073 14729
rect 17835 14300 17877 14309
rect 17835 14260 17836 14300
rect 17876 14260 17877 14300
rect 17835 14251 17877 14260
rect 17548 14176 17684 14216
rect 17356 13999 17396 14008
rect 17452 14048 17492 14057
rect 17260 13914 17300 13999
rect 17164 13336 17396 13376
rect 17068 13159 17108 13168
rect 17259 13208 17301 13217
rect 17259 13168 17260 13208
rect 17300 13168 17301 13208
rect 17259 13159 17301 13168
rect 16300 13074 16340 13159
rect 17163 13124 17205 13133
rect 17163 13084 17164 13124
rect 17204 13084 17205 13124
rect 17163 13075 17205 13084
rect 16107 13040 16149 13049
rect 16107 13000 16108 13040
rect 16148 13000 16149 13040
rect 16107 12991 16149 13000
rect 16491 13040 16533 13049
rect 16491 13000 16492 13040
rect 16532 13000 16533 13040
rect 16491 12991 16533 13000
rect 16011 12788 16053 12797
rect 16011 12748 16012 12788
rect 16052 12748 16053 12788
rect 16011 12739 16053 12748
rect 16203 12704 16245 12713
rect 16203 12664 16204 12704
rect 16244 12664 16245 12704
rect 16203 12655 16245 12664
rect 15916 12487 15956 12496
rect 16012 12536 16052 12545
rect 16204 12536 16244 12655
rect 16396 12536 16436 12545
rect 16052 12496 16148 12536
rect 16012 12487 16052 12496
rect 16108 12368 16148 12496
rect 16204 12487 16244 12496
rect 16300 12496 16396 12536
rect 16204 12368 16244 12377
rect 15820 12328 16052 12368
rect 16108 12328 16204 12368
rect 15723 12284 15765 12293
rect 15723 12244 15724 12284
rect 15764 12244 15765 12284
rect 15723 12235 15765 12244
rect 15724 12150 15764 12235
rect 15532 11705 15572 11740
rect 15723 11780 15765 11789
rect 15723 11740 15724 11780
rect 15764 11740 15765 11780
rect 15723 11731 15765 11740
rect 15531 11696 15573 11705
rect 15531 11656 15532 11696
rect 15572 11656 15573 11696
rect 15531 11647 15573 11656
rect 15724 11696 15764 11731
rect 15532 11616 15572 11647
rect 15724 11645 15764 11656
rect 15916 11696 15956 11705
rect 15820 11612 15860 11621
rect 15820 11528 15860 11572
rect 15724 11488 15860 11528
rect 15627 11360 15669 11369
rect 15627 11320 15628 11360
rect 15668 11320 15669 11360
rect 15627 11311 15669 11320
rect 15435 10940 15477 10949
rect 15435 10900 15436 10940
rect 15476 10900 15477 10940
rect 15435 10891 15477 10900
rect 15628 10940 15668 11311
rect 15724 11033 15764 11488
rect 15916 11117 15956 11656
rect 15915 11108 15957 11117
rect 15915 11068 15916 11108
rect 15956 11068 15957 11108
rect 15915 11059 15957 11068
rect 15723 11024 15765 11033
rect 15723 10984 15724 11024
rect 15764 10984 15765 11024
rect 15723 10975 15765 10984
rect 15148 9976 15380 10016
rect 15436 10772 15476 10781
rect 14667 9680 14709 9689
rect 14667 9640 14668 9680
rect 14708 9640 14709 9680
rect 14667 9631 14709 9640
rect 14955 9680 14997 9689
rect 14955 9640 14956 9680
rect 14996 9640 14997 9680
rect 14955 9631 14997 9640
rect 14092 9463 14132 9472
rect 14284 9512 14324 9521
rect 13996 9378 14036 9463
rect 14284 9353 14324 9472
rect 14380 9512 14420 9521
rect 14572 9512 14612 9521
rect 14283 9344 14325 9353
rect 14283 9304 14284 9344
rect 14324 9304 14325 9344
rect 14283 9295 14325 9304
rect 13900 9220 14132 9260
rect 13516 9052 13748 9092
rect 13708 8933 13748 9052
rect 13707 8924 13749 8933
rect 13707 8884 13708 8924
rect 13748 8884 13749 8924
rect 13707 8875 13749 8884
rect 13420 8756 13460 8767
rect 13420 8681 13460 8716
rect 13419 8672 13461 8681
rect 13419 8632 13420 8672
rect 13460 8632 13461 8672
rect 13419 8623 13461 8632
rect 13612 8504 13652 8513
rect 13516 8464 13612 8504
rect 13036 8119 13076 8128
rect 13131 8168 13173 8177
rect 13131 8128 13132 8168
rect 13172 8128 13173 8168
rect 13131 8119 13173 8128
rect 13132 8000 13172 8009
rect 13516 8000 13556 8464
rect 13612 8455 13652 8464
rect 13612 8168 13652 8177
rect 13708 8168 13748 8875
rect 13652 8128 13748 8168
rect 13612 8119 13652 8128
rect 13172 7960 13556 8000
rect 13996 8000 14036 8009
rect 13132 7951 13172 7960
rect 13035 7916 13077 7925
rect 13035 7876 13036 7916
rect 13076 7876 13077 7916
rect 13035 7867 13077 7876
rect 13803 7916 13845 7925
rect 13803 7876 13804 7916
rect 13844 7876 13845 7916
rect 13803 7867 13845 7876
rect 12843 7580 12885 7589
rect 12843 7540 12844 7580
rect 12884 7540 12885 7580
rect 12843 7531 12885 7540
rect 13036 7412 13076 7867
rect 13804 7782 13844 7867
rect 13996 7589 14036 7960
rect 14092 8000 14132 9220
rect 14283 8672 14325 8681
rect 14283 8632 14284 8672
rect 14324 8632 14325 8672
rect 14283 8623 14325 8632
rect 14284 8538 14324 8623
rect 14283 8420 14325 8429
rect 14283 8380 14284 8420
rect 14324 8380 14325 8420
rect 14283 8371 14325 8380
rect 14092 7951 14132 7960
rect 14188 8000 14228 8011
rect 14188 7925 14228 7960
rect 14284 8000 14324 8371
rect 14284 7951 14324 7960
rect 14187 7916 14229 7925
rect 14187 7876 14188 7916
rect 14228 7876 14229 7916
rect 14187 7867 14229 7876
rect 13995 7580 14037 7589
rect 13995 7540 13996 7580
rect 14036 7540 14037 7580
rect 13995 7531 14037 7540
rect 14380 7496 14420 9472
rect 14476 9472 14572 9512
rect 14476 8168 14516 9472
rect 14572 9463 14612 9472
rect 14764 9512 14804 9521
rect 14667 9428 14709 9437
rect 14667 9388 14668 9428
rect 14708 9388 14709 9428
rect 14667 9379 14709 9388
rect 14571 9260 14613 9269
rect 14571 9220 14572 9260
rect 14612 9220 14613 9260
rect 14571 9211 14613 9220
rect 14572 9126 14612 9211
rect 14668 8672 14708 9379
rect 14764 8849 14804 9472
rect 14860 9512 14900 9523
rect 14860 9437 14900 9472
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 15052 9512 15092 9521
rect 14859 9428 14901 9437
rect 14859 9388 14860 9428
rect 14900 9388 14901 9428
rect 14859 9379 14901 9388
rect 14859 8924 14901 8933
rect 14956 8924 14996 9463
rect 15052 9185 15092 9472
rect 15051 9176 15093 9185
rect 15051 9136 15052 9176
rect 15092 9136 15093 9176
rect 15051 9127 15093 9136
rect 14859 8884 14860 8924
rect 14900 8884 14996 8924
rect 14859 8875 14901 8884
rect 14763 8840 14805 8849
rect 14763 8800 14764 8840
rect 14804 8800 14805 8840
rect 14763 8791 14805 8800
rect 14764 8672 14804 8681
rect 14476 8119 14516 8128
rect 14572 8632 14764 8672
rect 14572 8000 14612 8632
rect 14764 8623 14804 8632
rect 14860 8672 14900 8875
rect 14860 8623 14900 8632
rect 14956 8672 14996 8681
rect 15148 8672 15188 9976
rect 15243 9848 15285 9857
rect 15243 9808 15244 9848
rect 15284 9808 15285 9848
rect 15243 9799 15285 9808
rect 15244 9512 15284 9799
rect 15436 9773 15476 10732
rect 15628 10184 15668 10900
rect 15628 10135 15668 10144
rect 15724 10016 15764 10975
rect 16012 10940 16052 12328
rect 16204 12319 16244 12328
rect 16300 11705 16340 12496
rect 16396 12487 16436 12496
rect 16492 11864 16532 12991
rect 17164 12990 17204 13075
rect 17260 13074 17300 13159
rect 16588 12536 16628 12545
rect 16588 12377 16628 12496
rect 16683 12536 16725 12545
rect 16683 12496 16684 12536
rect 16724 12496 16725 12536
rect 16683 12487 16725 12496
rect 16684 12402 16724 12487
rect 16587 12368 16629 12377
rect 16587 12328 16588 12368
rect 16628 12328 16629 12368
rect 16587 12319 16629 12328
rect 17163 11864 17205 11873
rect 16492 11824 16724 11864
rect 16299 11696 16341 11705
rect 16299 11656 16300 11696
rect 16340 11656 16341 11696
rect 16299 11647 16341 11656
rect 16396 11696 16436 11705
rect 16492 11696 16532 11824
rect 16436 11656 16532 11696
rect 16587 11696 16629 11705
rect 16587 11656 16588 11696
rect 16628 11656 16629 11696
rect 16396 11647 16436 11656
rect 16587 11647 16629 11656
rect 16684 11696 16724 11824
rect 17163 11824 17164 11864
rect 17204 11824 17205 11864
rect 17163 11815 17205 11824
rect 16684 11647 16724 11656
rect 16971 11696 17013 11705
rect 16971 11656 16972 11696
rect 17012 11656 17013 11696
rect 16971 11647 17013 11656
rect 16588 11562 16628 11647
rect 16107 11528 16149 11537
rect 16107 11488 16108 11528
rect 16148 11488 16149 11528
rect 16107 11479 16149 11488
rect 16299 11528 16341 11537
rect 16299 11488 16300 11528
rect 16340 11488 16341 11528
rect 16299 11479 16341 11488
rect 16875 11528 16917 11537
rect 16875 11488 16876 11528
rect 16916 11488 16917 11528
rect 16875 11479 16917 11488
rect 16108 11394 16148 11479
rect 16300 11196 16340 11479
rect 16876 11394 16916 11479
rect 16395 11360 16437 11369
rect 16972 11360 17012 11647
rect 16395 11320 16396 11360
rect 16436 11320 16437 11360
rect 16395 11311 16437 11320
rect 16967 11320 17012 11360
rect 16203 11024 16245 11033
rect 16108 10982 16148 10991
rect 16107 10942 16108 10949
rect 16203 10984 16204 11024
rect 16244 10984 16245 11024
rect 16203 10975 16245 10984
rect 16148 10942 16149 10949
rect 16107 10940 16149 10942
rect 16012 10900 16053 10940
rect 16013 10856 16053 10900
rect 16107 10900 16108 10940
rect 16148 10900 16149 10940
rect 16107 10891 16149 10900
rect 16012 10816 16053 10856
rect 16108 10847 16148 10891
rect 16204 10890 16244 10975
rect 15628 9976 15764 10016
rect 15820 10772 15860 10781
rect 15435 9764 15477 9773
rect 15435 9724 15436 9764
rect 15476 9724 15477 9764
rect 15435 9715 15477 9724
rect 15244 9463 15284 9472
rect 15339 9512 15381 9521
rect 15339 9472 15340 9512
rect 15380 9472 15381 9512
rect 15339 9463 15381 9472
rect 15436 9512 15476 9715
rect 15340 9378 15380 9463
rect 15436 9437 15476 9472
rect 15532 9512 15572 9521
rect 15435 9428 15477 9437
rect 15435 9388 15436 9428
rect 15476 9388 15477 9428
rect 15435 9379 15477 9388
rect 15532 8849 15572 9472
rect 15531 8840 15573 8849
rect 15531 8800 15532 8840
rect 15572 8800 15573 8840
rect 15531 8791 15573 8800
rect 15628 8681 15668 9976
rect 15723 9848 15765 9857
rect 15723 9808 15724 9848
rect 15764 9808 15765 9848
rect 15723 9799 15765 9808
rect 15724 9533 15764 9799
rect 15820 9689 15860 10732
rect 15915 9764 15957 9773
rect 15915 9724 15916 9764
rect 15956 9724 15957 9764
rect 15915 9715 15957 9724
rect 15819 9680 15861 9689
rect 15819 9640 15820 9680
rect 15860 9640 15861 9680
rect 15819 9631 15861 9640
rect 15724 9484 15764 9493
rect 15820 9512 15860 9521
rect 15820 9428 15860 9472
rect 15916 9512 15956 9715
rect 16012 9680 16052 10816
rect 16300 10520 16340 11156
rect 16204 10480 16340 10520
rect 16107 10352 16149 10361
rect 16107 10312 16108 10352
rect 16148 10312 16149 10352
rect 16107 10303 16149 10312
rect 16108 10184 16148 10303
rect 16108 10135 16148 10144
rect 16204 10184 16244 10480
rect 16204 9857 16244 10144
rect 16396 10184 16436 11311
rect 16967 11024 17007 11320
rect 16967 10975 17007 10984
rect 17068 11024 17108 11033
rect 17068 10865 17108 10984
rect 17164 11024 17204 11815
rect 17356 11360 17396 13336
rect 17452 13133 17492 14008
rect 17548 14048 17588 14057
rect 17548 13301 17588 14008
rect 17547 13292 17589 13301
rect 17547 13252 17548 13292
rect 17588 13252 17589 13292
rect 17547 13243 17589 13252
rect 17644 13208 17684 14176
rect 17739 14132 17781 14141
rect 17739 14092 17740 14132
rect 17780 14092 17781 14132
rect 17739 14083 17781 14092
rect 17836 14132 17876 14251
rect 17836 14083 17876 14092
rect 17740 14048 17780 14083
rect 17740 13997 17780 14008
rect 17932 14048 17972 14680
rect 17932 13553 17972 14008
rect 18028 14680 18033 14720
rect 18028 14671 18073 14680
rect 18315 14720 18357 14729
rect 18315 14680 18316 14720
rect 18356 14680 18357 14720
rect 18315 14671 18357 14680
rect 18412 14720 18452 14729
rect 17931 13544 17973 13553
rect 17931 13504 17932 13544
rect 17972 13504 17973 13544
rect 17931 13495 17973 13504
rect 18028 13376 18068 14671
rect 18316 14586 18356 14671
rect 18412 14561 18452 14680
rect 18508 14720 18548 14729
rect 18411 14552 18453 14561
rect 18411 14512 18412 14552
rect 18452 14512 18453 14552
rect 18411 14503 18453 14512
rect 18508 14309 18548 14680
rect 18604 14720 18644 14729
rect 18700 14720 18740 15175
rect 18892 14897 18932 15268
rect 18891 14888 18933 14897
rect 18891 14848 18892 14888
rect 18932 14848 18933 14888
rect 18891 14839 18933 14848
rect 18644 14680 18740 14720
rect 18604 14671 18644 14680
rect 18507 14300 18549 14309
rect 18507 14260 18508 14300
rect 18548 14260 18549 14300
rect 18507 14251 18549 14260
rect 19372 14216 19412 15427
rect 19660 15401 19700 15520
rect 19796 15520 19988 15560
rect 20044 15560 20084 15569
rect 19756 15511 19796 15520
rect 19659 15392 19701 15401
rect 19659 15352 19660 15392
rect 19700 15352 19701 15392
rect 19659 15343 19701 15352
rect 19660 14561 19700 15343
rect 19947 14888 19989 14897
rect 19947 14848 19948 14888
rect 19988 14848 19989 14888
rect 19947 14839 19989 14848
rect 19851 14720 19893 14729
rect 19851 14680 19852 14720
rect 19892 14680 19893 14720
rect 19851 14671 19893 14680
rect 19948 14720 19988 14839
rect 20044 14804 20084 15520
rect 20139 15560 20181 15569
rect 20139 15520 20140 15560
rect 20180 15520 20181 15560
rect 20139 15511 20181 15520
rect 20236 15560 20276 15569
rect 20140 15426 20180 15511
rect 20236 15317 20276 15520
rect 20619 15560 20661 15569
rect 20619 15520 20620 15560
rect 20660 15520 20661 15560
rect 20619 15511 20661 15520
rect 20716 15560 20756 15571
rect 20235 15308 20277 15317
rect 20235 15268 20236 15308
rect 20276 15268 20277 15308
rect 20235 15259 20277 15268
rect 20236 15149 20276 15259
rect 20235 15140 20277 15149
rect 20235 15100 20236 15140
rect 20276 15100 20277 15140
rect 20235 15091 20277 15100
rect 20140 14972 20180 14981
rect 20180 14932 20372 14972
rect 20140 14923 20180 14932
rect 20235 14804 20277 14813
rect 20044 14764 20180 14804
rect 19948 14671 19988 14680
rect 20140 14678 20180 14764
rect 20235 14764 20236 14804
rect 20276 14764 20277 14804
rect 20235 14755 20277 14764
rect 19659 14552 19701 14561
rect 19659 14512 19660 14552
rect 19700 14512 19701 14552
rect 19852 14552 19892 14671
rect 19852 14512 19988 14552
rect 19659 14503 19701 14512
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19948 14225 19988 14512
rect 20140 14393 20180 14638
rect 20139 14384 20181 14393
rect 20139 14344 20140 14384
rect 20180 14344 20181 14384
rect 20139 14335 20181 14344
rect 19852 14216 19892 14225
rect 19947 14216 19989 14225
rect 19372 14176 19796 14216
rect 18987 14132 19029 14141
rect 18987 14092 18988 14132
rect 19028 14092 19029 14132
rect 18987 14083 19029 14092
rect 18796 14048 18836 14057
rect 18796 13889 18836 14008
rect 18891 14048 18933 14057
rect 18891 14008 18892 14048
rect 18932 14008 18933 14048
rect 18891 13999 18933 14008
rect 18988 14048 19028 14083
rect 18892 13914 18932 13999
rect 18988 13997 19028 14008
rect 19084 14048 19124 14057
rect 18795 13880 18837 13889
rect 18795 13840 18796 13880
rect 18836 13840 18837 13880
rect 18795 13831 18837 13840
rect 18987 13796 19029 13805
rect 18987 13756 18988 13796
rect 19028 13756 19029 13796
rect 18987 13747 19029 13756
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 17932 13336 18068 13376
rect 17451 13124 17493 13133
rect 17451 13084 17452 13124
rect 17492 13084 17493 13124
rect 17451 13075 17493 13084
rect 17644 11696 17684 13168
rect 17739 13208 17781 13217
rect 17739 13168 17740 13208
rect 17780 13168 17781 13208
rect 17739 13159 17781 13168
rect 17932 13208 17972 13336
rect 17740 13074 17780 13159
rect 17836 13040 17876 13049
rect 17836 12629 17876 13000
rect 17932 12797 17972 13168
rect 18027 13208 18069 13217
rect 18129 13208 18169 13217
rect 18027 13168 18028 13208
rect 18068 13168 18069 13208
rect 18027 13159 18069 13168
rect 18124 13168 18129 13208
rect 18124 13159 18169 13168
rect 18315 13208 18357 13217
rect 18315 13168 18316 13208
rect 18356 13168 18357 13208
rect 18315 13159 18357 13168
rect 18603 13208 18645 13217
rect 18603 13168 18604 13208
rect 18644 13168 18645 13208
rect 18603 13159 18645 13168
rect 18028 13074 18068 13159
rect 17931 12788 17973 12797
rect 17931 12748 17932 12788
rect 17972 12748 17973 12788
rect 17931 12739 17973 12748
rect 17835 12620 17877 12629
rect 17835 12580 17836 12620
rect 17876 12580 17877 12620
rect 17835 12571 17877 12580
rect 17835 11948 17877 11957
rect 17835 11908 17836 11948
rect 17876 11908 17877 11948
rect 18124 11948 18164 13159
rect 18316 12536 18356 13159
rect 18507 12956 18549 12965
rect 18507 12916 18508 12956
rect 18548 12916 18549 12956
rect 18507 12907 18549 12916
rect 18508 12629 18548 12907
rect 18507 12620 18549 12629
rect 18507 12580 18508 12620
rect 18548 12580 18549 12620
rect 18507 12571 18549 12580
rect 18604 12620 18644 13159
rect 18988 12704 19028 13747
rect 19084 13553 19124 14008
rect 19467 14048 19509 14057
rect 19467 14008 19468 14048
rect 19508 14008 19509 14048
rect 19467 13999 19509 14008
rect 19564 14048 19604 14059
rect 19468 13914 19508 13999
rect 19564 13973 19604 14008
rect 19563 13964 19605 13973
rect 19563 13924 19564 13964
rect 19604 13924 19605 13964
rect 19563 13915 19605 13924
rect 19083 13544 19125 13553
rect 19083 13504 19084 13544
rect 19124 13504 19125 13544
rect 19083 13495 19125 13504
rect 19564 13301 19604 13915
rect 19659 13544 19701 13553
rect 19659 13504 19660 13544
rect 19700 13504 19701 13544
rect 19756 13544 19796 14176
rect 19892 14176 19948 14216
rect 19988 14176 19989 14216
rect 19852 14167 19892 14176
rect 19947 14167 19989 14176
rect 19948 14082 19988 14167
rect 20044 14048 20084 14057
rect 19947 13964 19989 13973
rect 20044 13964 20084 14008
rect 19947 13924 19948 13964
rect 19988 13924 20084 13964
rect 19947 13915 19989 13924
rect 19756 13504 19988 13544
rect 19659 13495 19701 13504
rect 19275 13292 19317 13301
rect 19275 13252 19276 13292
rect 19316 13252 19317 13292
rect 19275 13243 19317 13252
rect 19563 13292 19605 13301
rect 19563 13252 19564 13292
rect 19604 13252 19605 13292
rect 19563 13243 19605 13252
rect 19083 13208 19125 13217
rect 19083 13168 19084 13208
rect 19124 13168 19125 13208
rect 19083 13159 19125 13168
rect 19276 13208 19316 13243
rect 19084 13074 19124 13159
rect 19276 13157 19316 13168
rect 19372 13208 19412 13217
rect 19179 13124 19221 13133
rect 19179 13084 19180 13124
rect 19220 13084 19221 13124
rect 19179 13075 19221 13084
rect 19180 12990 19220 13075
rect 19083 12704 19125 12713
rect 18988 12664 19084 12704
rect 19124 12664 19125 12704
rect 19083 12655 19125 12664
rect 19372 12704 19412 13168
rect 19660 13208 19700 13495
rect 19660 13159 19700 13168
rect 19755 13208 19797 13217
rect 19755 13168 19756 13208
rect 19796 13168 19797 13208
rect 19755 13159 19797 13168
rect 19852 13208 19892 13217
rect 19564 13049 19604 13134
rect 19756 13074 19796 13159
rect 19852 13049 19892 13168
rect 19563 13040 19605 13049
rect 19563 13000 19564 13040
rect 19604 13000 19605 13040
rect 19563 12991 19605 13000
rect 19851 13040 19893 13049
rect 19851 13000 19852 13040
rect 19892 13000 19893 13040
rect 19851 12991 19893 13000
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 19372 12655 19412 12664
rect 19467 12704 19509 12713
rect 19467 12664 19468 12704
rect 19508 12664 19509 12704
rect 19467 12655 19509 12664
rect 18604 12571 18644 12580
rect 18508 12557 18548 12571
rect 18316 12377 18356 12496
rect 18412 12536 18452 12547
rect 18508 12508 18548 12517
rect 18795 12536 18837 12545
rect 18412 12461 18452 12496
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 18795 12487 18837 12496
rect 18988 12536 19028 12547
rect 18411 12452 18453 12461
rect 18411 12412 18412 12452
rect 18452 12412 18453 12452
rect 18411 12403 18453 12412
rect 18796 12402 18836 12487
rect 18988 12461 19028 12496
rect 19084 12536 19124 12545
rect 18987 12452 19029 12461
rect 18987 12412 18988 12452
rect 19028 12412 19029 12452
rect 18987 12403 19029 12412
rect 18315 12368 18357 12377
rect 18315 12328 18316 12368
rect 18356 12328 18357 12368
rect 18315 12319 18357 12328
rect 18795 12284 18837 12293
rect 18795 12244 18796 12284
rect 18836 12244 18837 12284
rect 18795 12235 18837 12244
rect 18796 12150 18836 12235
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 18987 12116 19029 12125
rect 18987 12076 18988 12116
rect 19028 12076 19029 12116
rect 18987 12067 19029 12076
rect 18124 11908 18417 11948
rect 17835 11899 17877 11908
rect 17836 11814 17876 11899
rect 18377 11789 18417 11908
rect 18219 11780 18261 11789
rect 18219 11740 18220 11780
rect 18260 11740 18261 11780
rect 18219 11731 18261 11740
rect 18376 11780 18418 11789
rect 18376 11740 18377 11780
rect 18417 11740 18418 11780
rect 18376 11731 18418 11740
rect 17836 11696 17876 11705
rect 17644 11656 17836 11696
rect 17836 11453 17876 11656
rect 17932 11696 17972 11705
rect 17932 11537 17972 11656
rect 18076 11700 18116 11709
rect 18076 11621 18116 11660
rect 18220 11696 18260 11731
rect 18220 11645 18260 11656
rect 18377 11711 18417 11731
rect 18377 11645 18417 11671
rect 18075 11612 18117 11621
rect 18075 11572 18076 11612
rect 18116 11572 18117 11612
rect 18075 11563 18117 11572
rect 17931 11528 17973 11537
rect 17931 11488 17932 11528
rect 17972 11488 17973 11528
rect 17931 11479 17973 11488
rect 17835 11444 17877 11453
rect 17835 11404 17836 11444
rect 17876 11404 17877 11444
rect 17835 11395 17877 11404
rect 18891 11444 18933 11453
rect 18891 11404 18892 11444
rect 18932 11404 18933 11444
rect 18891 11395 18933 11404
rect 17356 11320 17684 11360
rect 17164 10975 17204 10984
rect 17260 11192 17300 11201
rect 17067 10856 17109 10865
rect 17067 10816 17068 10856
rect 17108 10816 17109 10856
rect 17067 10807 17109 10816
rect 16684 10312 17108 10352
rect 16588 10184 16628 10193
rect 16436 10144 16532 10184
rect 16396 10135 16436 10144
rect 16396 10016 16436 10025
rect 16396 9857 16436 9976
rect 16203 9848 16245 9857
rect 16203 9808 16204 9848
rect 16244 9808 16245 9848
rect 16203 9799 16245 9808
rect 16395 9848 16437 9857
rect 16395 9808 16396 9848
rect 16436 9808 16437 9848
rect 16395 9799 16437 9808
rect 16203 9680 16245 9689
rect 16012 9640 16148 9680
rect 15916 9463 15956 9472
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 15724 9388 15860 9428
rect 15724 8933 15764 9388
rect 16012 9378 16052 9463
rect 15915 9344 15957 9353
rect 15915 9304 15916 9344
rect 15956 9304 15957 9344
rect 16108 9344 16148 9640
rect 16203 9640 16204 9680
rect 16244 9640 16245 9680
rect 16203 9631 16245 9640
rect 16204 9512 16244 9631
rect 16204 9463 16244 9472
rect 16300 9512 16340 9521
rect 16300 9428 16340 9472
rect 16492 9512 16532 10144
rect 16588 9521 16628 10144
rect 16684 10100 16724 10312
rect 16684 10051 16724 10060
rect 16780 10184 16820 10193
rect 16780 9857 16820 10144
rect 16876 10184 16916 10193
rect 16876 10100 16916 10144
rect 17068 10184 17108 10312
rect 17068 10135 17108 10144
rect 16971 10100 17013 10109
rect 16876 10060 16972 10100
rect 17012 10060 17013 10100
rect 16971 10051 17013 10060
rect 16779 9848 16821 9857
rect 16779 9808 16780 9848
rect 16820 9808 16821 9848
rect 16779 9799 16821 9808
rect 16875 9764 16917 9773
rect 16875 9724 16876 9764
rect 16916 9724 16917 9764
rect 16875 9715 16917 9724
rect 16492 9463 16532 9472
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 16300 9388 16436 9428
rect 16108 9304 16244 9344
rect 15915 9295 15957 9304
rect 15819 9260 15861 9269
rect 15819 9220 15820 9260
rect 15860 9220 15861 9260
rect 15819 9211 15861 9220
rect 15723 8924 15765 8933
rect 15723 8884 15724 8924
rect 15764 8884 15765 8924
rect 15723 8875 15765 8884
rect 14996 8632 15188 8672
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 14956 8623 14996 8632
rect 15627 8623 15669 8632
rect 15820 8672 15860 9211
rect 15916 8672 15956 9295
rect 16107 9176 16149 9185
rect 16107 9136 16108 9176
rect 16148 9136 16149 9176
rect 16107 9127 16149 9136
rect 16012 8672 16052 8681
rect 15916 8632 16012 8672
rect 15820 8623 15860 8632
rect 16012 8623 16052 8632
rect 16108 8672 16148 9127
rect 16108 8623 16148 8632
rect 14667 8504 14709 8513
rect 14667 8464 14668 8504
rect 14708 8464 14709 8504
rect 14667 8455 14709 8464
rect 15148 8504 15188 8513
rect 14668 8370 14708 8455
rect 14763 8336 14805 8345
rect 14763 8296 14764 8336
rect 14804 8296 14805 8336
rect 14763 8287 14805 8296
rect 14572 7951 14612 7960
rect 14668 8000 14708 8011
rect 14668 7925 14708 7960
rect 14764 8000 14804 8287
rect 14956 8084 14996 8093
rect 15148 8084 15188 8464
rect 16011 8504 16053 8513
rect 16011 8464 16012 8504
rect 16052 8464 16053 8504
rect 16011 8455 16053 8464
rect 14996 8044 15188 8084
rect 14956 8035 14996 8044
rect 14764 7951 14804 7960
rect 15339 8000 15381 8009
rect 15339 7960 15340 8000
rect 15380 7960 15381 8000
rect 15339 7951 15381 7960
rect 14667 7916 14709 7925
rect 14667 7876 14668 7916
rect 14708 7876 14709 7916
rect 14667 7867 14709 7876
rect 15340 7866 15380 7951
rect 15531 7916 15573 7925
rect 15531 7876 15532 7916
rect 15572 7876 15573 7916
rect 15531 7867 15573 7876
rect 15243 7580 15285 7589
rect 15243 7540 15244 7580
rect 15284 7540 15285 7580
rect 15243 7531 15285 7540
rect 14380 7456 14612 7496
rect 13036 7363 13076 7372
rect 14476 7328 14516 7337
rect 14284 7169 14324 7254
rect 14380 7244 14420 7253
rect 11883 7120 11884 7160
rect 11924 7120 11925 7160
rect 11883 7111 11925 7120
rect 12268 7120 12364 7160
rect 12404 7120 12596 7160
rect 12747 7160 12789 7169
rect 12747 7120 12748 7160
rect 12788 7120 12789 7160
rect 11884 7026 11924 7111
rect 12076 6992 12116 7001
rect 11883 6908 11925 6917
rect 11883 6868 11884 6908
rect 11924 6868 11925 6908
rect 11883 6859 11925 6868
rect 11787 6740 11829 6749
rect 11787 6700 11788 6740
rect 11828 6700 11829 6740
rect 11787 6691 11829 6700
rect 10540 6236 10580 6245
rect 10348 5648 10388 5657
rect 10348 5069 10388 5608
rect 10443 5648 10485 5657
rect 10443 5608 10444 5648
rect 10484 5608 10485 5648
rect 10443 5599 10485 5608
rect 10540 5648 10580 6196
rect 10635 6236 10677 6245
rect 10635 6196 10636 6236
rect 10676 6196 10677 6236
rect 10635 6187 10677 6196
rect 10540 5599 10580 5608
rect 10636 5480 10676 6187
rect 10732 5825 10772 5910
rect 10731 5816 10773 5825
rect 10731 5776 10732 5816
rect 10772 5776 10773 5816
rect 10731 5767 10773 5776
rect 10827 5732 10869 5741
rect 10827 5692 10828 5732
rect 10868 5692 10869 5732
rect 10827 5683 10869 5692
rect 10731 5648 10773 5657
rect 10731 5608 10732 5648
rect 10772 5608 10773 5648
rect 10731 5599 10773 5608
rect 10828 5648 10868 5683
rect 10732 5514 10772 5599
rect 10828 5597 10868 5608
rect 10444 5440 10676 5480
rect 10347 5060 10389 5069
rect 10347 5020 10348 5060
rect 10388 5020 10389 5060
rect 10347 5011 10389 5020
rect 9388 4136 9428 4145
rect 9196 4096 9388 4136
rect 9196 3809 9236 4096
rect 9388 4087 9428 4096
rect 9484 4136 9524 4145
rect 9675 4136 9717 4145
rect 9524 4096 9620 4136
rect 9484 4087 9524 4096
rect 9195 3800 9237 3809
rect 9195 3760 9196 3800
rect 9236 3760 9237 3800
rect 9195 3751 9237 3760
rect 9099 3632 9141 3641
rect 9099 3592 9100 3632
rect 9140 3592 9141 3632
rect 9099 3583 9141 3592
rect 8716 3464 8756 3475
rect 8716 3389 8756 3424
rect 8715 3380 8757 3389
rect 8715 3340 8716 3380
rect 8756 3340 8757 3380
rect 8715 3331 8757 3340
rect 9100 2801 9140 3583
rect 9099 2792 9141 2801
rect 9097 2752 9100 2792
rect 9140 2752 9141 2792
rect 9097 2743 9141 2752
rect 9196 2792 9236 3751
rect 9387 3716 9429 3725
rect 9387 3676 9388 3716
rect 9428 3676 9429 3716
rect 9387 3667 9429 3676
rect 9388 3632 9428 3667
rect 9580 3641 9620 4096
rect 9675 4096 9676 4136
rect 9716 4096 9717 4136
rect 9675 4087 9717 4096
rect 10251 4136 10293 4145
rect 10251 4096 10252 4136
rect 10292 4096 10293 4136
rect 10251 4087 10293 4096
rect 10444 4136 10484 5440
rect 10635 4304 10677 4313
rect 10635 4264 10636 4304
rect 10676 4264 10677 4304
rect 10635 4255 10677 4264
rect 9963 4052 10005 4061
rect 9963 4012 9964 4052
rect 10004 4012 10005 4052
rect 9963 4003 10005 4012
rect 9675 3968 9717 3977
rect 9675 3928 9676 3968
rect 9716 3928 9717 3968
rect 9675 3919 9717 3928
rect 9676 3834 9716 3919
rect 9388 3581 9428 3592
rect 9579 3632 9621 3641
rect 9579 3592 9580 3632
rect 9620 3592 9621 3632
rect 9579 3583 9621 3592
rect 9291 3464 9333 3473
rect 9291 3424 9292 3464
rect 9332 3424 9333 3464
rect 9291 3415 9333 3424
rect 9388 3464 9428 3473
rect 9196 2743 9236 2752
rect 9097 2624 9137 2743
rect 9196 2624 9236 2633
rect 9097 2584 9140 2624
rect 8620 2575 8660 2584
rect 9100 2540 9140 2584
rect 9196 2540 9236 2584
rect 9100 2500 9236 2540
rect 9292 2465 9332 3415
rect 9388 2876 9428 3424
rect 9483 3464 9525 3473
rect 9483 3424 9484 3464
rect 9524 3424 9525 3464
rect 9483 3415 9525 3424
rect 9484 3330 9524 3415
rect 9676 3212 9716 3221
rect 9868 3212 9908 3221
rect 9388 2827 9428 2836
rect 9484 3172 9676 3212
rect 8139 2456 8181 2465
rect 8139 2416 8140 2456
rect 8180 2416 8181 2456
rect 8139 2407 8181 2416
rect 9291 2456 9333 2465
rect 9291 2416 9292 2456
rect 9332 2416 9333 2456
rect 9291 2407 9333 2416
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 9484 1961 9524 3172
rect 9676 3163 9716 3172
rect 9772 3172 9868 3212
rect 9580 2624 9620 2633
rect 9772 2624 9812 3172
rect 9868 3163 9908 3172
rect 9964 3044 10004 4003
rect 9620 2584 9812 2624
rect 9868 3004 10004 3044
rect 9580 2575 9620 2584
rect 9675 2456 9717 2465
rect 9675 2416 9676 2456
rect 9716 2416 9717 2456
rect 9675 2407 9717 2416
rect 9483 1952 9525 1961
rect 9483 1912 9484 1952
rect 9524 1912 9525 1952
rect 9483 1903 9525 1912
rect 9676 1952 9716 2407
rect 9676 1903 9716 1912
rect 9772 1952 9812 1961
rect 9868 1952 9908 3004
rect 9964 2624 10004 2633
rect 9964 2540 10004 2584
rect 9964 2500 10100 2540
rect 9964 1952 10004 1961
rect 9868 1912 9964 1952
rect 843 1700 885 1709
rect 843 1660 844 1700
rect 884 1660 885 1700
rect 843 1651 885 1660
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 9772 1289 9812 1912
rect 9964 1903 10004 1912
rect 9963 1784 10005 1793
rect 9963 1744 9964 1784
rect 10004 1744 10005 1784
rect 10060 1784 10100 2500
rect 10156 1784 10196 1793
rect 10060 1744 10156 1784
rect 9963 1735 10005 1744
rect 10156 1735 10196 1744
rect 9964 1650 10004 1735
rect 9771 1280 9813 1289
rect 9771 1240 9772 1280
rect 9812 1240 9813 1280
rect 9771 1231 9813 1240
rect 10155 1280 10197 1289
rect 10155 1240 10156 1280
rect 10196 1240 10197 1280
rect 10155 1231 10197 1240
rect 10252 1280 10292 4087
rect 10444 3725 10484 4096
rect 10636 4136 10676 4255
rect 10924 4136 10964 6280
rect 11212 6236 11252 6280
rect 11020 6196 11252 6236
rect 11020 4985 11060 6196
rect 11691 6152 11733 6161
rect 11691 6112 11692 6152
rect 11732 6112 11733 6152
rect 11691 6103 11733 6112
rect 11115 6068 11157 6077
rect 11115 6028 11116 6068
rect 11156 6028 11157 6068
rect 11115 6019 11157 6028
rect 11116 5648 11156 6019
rect 11211 5984 11253 5993
rect 11211 5944 11212 5984
rect 11252 5944 11253 5984
rect 11211 5935 11253 5944
rect 11212 5900 11252 5935
rect 11596 5909 11636 5940
rect 11212 5849 11252 5860
rect 11595 5900 11637 5909
rect 11595 5860 11596 5900
rect 11636 5860 11637 5900
rect 11595 5851 11637 5860
rect 11500 5816 11540 5825
rect 11403 5732 11445 5741
rect 11403 5692 11404 5732
rect 11444 5692 11445 5732
rect 11403 5683 11445 5692
rect 11116 5599 11156 5608
rect 11308 5648 11348 5657
rect 11308 5489 11348 5608
rect 11307 5480 11349 5489
rect 11307 5440 11308 5480
rect 11348 5440 11349 5480
rect 11307 5431 11349 5440
rect 11404 5405 11444 5683
rect 11115 5396 11157 5405
rect 11115 5356 11116 5396
rect 11156 5356 11157 5396
rect 11115 5347 11157 5356
rect 11403 5396 11445 5405
rect 11403 5356 11404 5396
rect 11444 5356 11445 5396
rect 11403 5347 11445 5356
rect 11116 5069 11156 5347
rect 11500 5321 11540 5776
rect 11596 5816 11636 5851
rect 11596 5405 11636 5776
rect 11692 5741 11732 6103
rect 11788 5909 11828 6691
rect 11787 5900 11829 5909
rect 11787 5860 11788 5900
rect 11828 5860 11829 5900
rect 11787 5851 11829 5860
rect 11691 5732 11733 5741
rect 11691 5692 11692 5732
rect 11732 5692 11733 5732
rect 11691 5683 11733 5692
rect 11692 5598 11732 5683
rect 11788 5648 11828 5851
rect 11884 5741 11924 6859
rect 12076 6497 12116 6952
rect 12075 6488 12117 6497
rect 12075 6448 12076 6488
rect 12116 6448 12117 6488
rect 12075 6439 12117 6448
rect 12268 6320 12308 7120
rect 12364 7111 12404 7120
rect 12747 7111 12789 7120
rect 13227 7160 13269 7169
rect 13227 7120 13228 7160
rect 13268 7120 13269 7160
rect 13227 7111 13269 7120
rect 13612 7160 13652 7169
rect 14188 7160 14228 7169
rect 12076 6280 12308 6320
rect 12364 6656 12404 6665
rect 11883 5732 11925 5741
rect 11883 5692 11884 5732
rect 11924 5692 11925 5732
rect 11883 5690 11925 5692
rect 11883 5683 11884 5690
rect 11788 5599 11828 5608
rect 11924 5683 11925 5690
rect 11884 5597 11924 5650
rect 11595 5396 11637 5405
rect 11595 5356 11596 5396
rect 11636 5356 11637 5396
rect 11595 5347 11637 5356
rect 11499 5312 11541 5321
rect 11499 5272 11500 5312
rect 11540 5272 11541 5312
rect 11499 5263 11541 5272
rect 11691 5312 11733 5321
rect 11691 5272 11692 5312
rect 11732 5272 11733 5312
rect 11691 5263 11733 5272
rect 11115 5060 11157 5069
rect 11115 5020 11116 5060
rect 11156 5020 11157 5060
rect 11115 5011 11157 5020
rect 11499 5060 11541 5069
rect 11499 5020 11500 5060
rect 11540 5020 11541 5060
rect 11499 5011 11541 5020
rect 11019 4976 11061 4985
rect 11019 4936 11020 4976
rect 11060 4936 11061 4976
rect 11019 4927 11061 4936
rect 11116 4976 11156 5011
rect 11116 4925 11156 4936
rect 11307 4976 11349 4985
rect 11307 4936 11308 4976
rect 11348 4936 11349 4976
rect 11307 4927 11349 4936
rect 11211 4388 11253 4397
rect 11211 4348 11212 4388
rect 11252 4348 11253 4388
rect 11211 4339 11253 4348
rect 11020 4304 11060 4313
rect 11060 4264 11156 4304
rect 11020 4255 11060 4264
rect 11019 4136 11061 4145
rect 10924 4096 11020 4136
rect 11060 4096 11061 4136
rect 10539 4052 10581 4061
rect 10539 4012 10540 4052
rect 10580 4012 10581 4052
rect 10539 4003 10581 4012
rect 10540 3918 10580 4003
rect 10636 3977 10676 4096
rect 11019 4087 11061 4096
rect 10635 3968 10677 3977
rect 10635 3928 10636 3968
rect 10676 3928 10677 3968
rect 10635 3919 10677 3928
rect 10827 3800 10869 3809
rect 10827 3760 10828 3800
rect 10868 3760 10869 3800
rect 10827 3751 10869 3760
rect 10443 3716 10485 3725
rect 10443 3676 10444 3716
rect 10484 3676 10485 3716
rect 10443 3667 10485 3676
rect 10540 3464 10580 3473
rect 10540 1793 10580 3424
rect 10828 2624 10868 3751
rect 11020 3632 11060 4087
rect 11017 3592 11060 3632
rect 11017 3485 11057 3592
rect 11017 3436 11057 3445
rect 11116 3380 11156 4264
rect 11212 4254 11252 4339
rect 11212 3968 11252 3977
rect 11212 3464 11252 3928
rect 11308 3809 11348 4927
rect 11404 4313 11444 4398
rect 11403 4304 11445 4313
rect 11403 4264 11404 4304
rect 11444 4264 11445 4304
rect 11403 4255 11445 4264
rect 11404 4136 11444 4145
rect 11500 4136 11540 5011
rect 11692 4976 11732 5263
rect 11787 5144 11829 5153
rect 11787 5104 11788 5144
rect 11828 5104 11829 5144
rect 11787 5095 11829 5104
rect 11980 5144 12020 5153
rect 11692 4927 11732 4936
rect 11788 4976 11828 5095
rect 11883 5060 11925 5069
rect 11883 5020 11884 5060
rect 11924 5020 11925 5060
rect 11883 5011 11925 5020
rect 11788 4927 11828 4936
rect 11884 4926 11924 5011
rect 11691 4808 11733 4817
rect 11691 4768 11692 4808
rect 11732 4768 11733 4808
rect 11691 4759 11733 4768
rect 11444 4096 11540 4136
rect 11404 4087 11444 4096
rect 11307 3800 11349 3809
rect 11307 3760 11308 3800
rect 11348 3760 11349 3800
rect 11307 3751 11349 3760
rect 11403 3632 11445 3641
rect 11403 3592 11404 3632
rect 11444 3592 11445 3632
rect 11403 3583 11445 3592
rect 11404 3498 11444 3583
rect 11212 3415 11252 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11033 3340 11156 3380
rect 11033 3296 11073 3340
rect 10828 2575 10868 2584
rect 10924 3256 11073 3296
rect 10731 1952 10773 1961
rect 10731 1912 10732 1952
rect 10772 1912 10773 1952
rect 10924 1952 10964 3256
rect 11116 3212 11156 3221
rect 11308 3212 11348 3415
rect 11500 3221 11540 4096
rect 11692 4136 11732 4759
rect 11980 4649 12020 5104
rect 12076 5144 12116 6280
rect 12364 6077 12404 6616
rect 12556 6488 12596 6497
rect 12363 6068 12405 6077
rect 12363 6028 12364 6068
rect 12404 6028 12405 6068
rect 12363 6019 12405 6028
rect 12556 5909 12596 6448
rect 12652 6488 12692 6497
rect 12748 6488 12788 7111
rect 12939 6992 12981 7001
rect 12939 6952 12940 6992
rect 12980 6952 12981 6992
rect 12939 6943 12981 6952
rect 12692 6448 12788 6488
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12652 6439 12692 6448
rect 12843 6439 12885 6448
rect 12940 6488 12980 6943
rect 13132 6656 13172 6665
rect 12940 6439 12980 6448
rect 13036 6572 13076 6581
rect 12844 6354 12884 6439
rect 13036 6077 13076 6532
rect 13035 6068 13077 6077
rect 13035 6028 13036 6068
rect 13076 6028 13077 6068
rect 13035 6019 13077 6028
rect 12555 5900 12597 5909
rect 12555 5860 12556 5900
rect 12596 5860 12597 5900
rect 12555 5851 12597 5860
rect 12268 5741 12308 5772
rect 12267 5732 12309 5741
rect 12267 5692 12268 5732
rect 12308 5692 12309 5732
rect 12267 5683 12309 5692
rect 12171 5648 12213 5657
rect 12171 5608 12172 5648
rect 12212 5608 12213 5648
rect 12171 5599 12213 5608
rect 12268 5648 12308 5683
rect 12172 5514 12212 5599
rect 12076 5095 12116 5104
rect 12268 4976 12308 5608
rect 12747 5564 12789 5573
rect 12747 5524 12748 5564
rect 12788 5524 12789 5564
rect 12747 5515 12789 5524
rect 12459 5480 12501 5489
rect 12459 5440 12460 5480
rect 12500 5440 12501 5480
rect 12459 5431 12501 5440
rect 12460 5346 12500 5431
rect 12748 5430 12788 5515
rect 13132 5489 13172 6616
rect 13228 6656 13268 7111
rect 13612 7001 13652 7120
rect 13900 7120 14188 7160
rect 13131 5480 13173 5489
rect 13131 5440 13132 5480
rect 13172 5440 13173 5480
rect 13131 5431 13173 5440
rect 13228 5144 13268 6616
rect 13516 6992 13556 7001
rect 13516 5993 13556 6952
rect 13611 6992 13653 7001
rect 13804 6992 13844 7001
rect 13611 6952 13612 6992
rect 13652 6952 13653 6992
rect 13611 6943 13653 6952
rect 13708 6952 13804 6992
rect 13611 6656 13653 6665
rect 13611 6616 13612 6656
rect 13652 6616 13653 6656
rect 13611 6607 13653 6616
rect 13515 5984 13557 5993
rect 13515 5944 13516 5984
rect 13556 5944 13557 5984
rect 13515 5935 13557 5944
rect 13612 5816 13652 6607
rect 13708 6488 13748 6952
rect 13804 6943 13844 6952
rect 13803 6824 13845 6833
rect 13803 6784 13804 6824
rect 13844 6784 13845 6824
rect 13803 6775 13845 6784
rect 13708 6439 13748 6448
rect 13804 6488 13844 6775
rect 13804 6439 13844 6448
rect 13803 6320 13845 6329
rect 13803 6280 13804 6320
rect 13844 6280 13845 6320
rect 13803 6271 13845 6280
rect 13612 5776 13748 5816
rect 13708 5732 13748 5776
rect 13708 5683 13748 5692
rect 13419 5648 13461 5657
rect 13419 5608 13420 5648
rect 13460 5608 13461 5648
rect 13419 5599 13461 5608
rect 13612 5648 13652 5659
rect 13420 5514 13460 5599
rect 13612 5573 13652 5608
rect 13804 5648 13844 6271
rect 13804 5599 13844 5608
rect 13900 5816 13940 7120
rect 14188 7111 14228 7120
rect 14283 7160 14325 7169
rect 14283 7120 14284 7160
rect 14324 7120 14325 7160
rect 14283 7111 14325 7120
rect 14284 6992 14324 7001
rect 13996 6952 14284 6992
rect 13996 6488 14036 6952
rect 14284 6943 14324 6952
rect 14188 6656 14228 6665
rect 14228 6616 14324 6656
rect 14188 6607 14228 6616
rect 14284 6572 14324 6616
rect 14284 6532 14325 6572
rect 13996 6439 14036 6448
rect 14092 6488 14132 6497
rect 14092 5900 14132 6448
rect 14192 6488 14234 6497
rect 14192 6448 14193 6488
rect 14233 6448 14234 6488
rect 14192 6439 14234 6448
rect 14193 6354 14233 6439
rect 14285 6404 14325 6532
rect 14380 6497 14420 7204
rect 14476 6665 14516 7288
rect 14572 6749 14612 7456
rect 14764 7160 14804 7169
rect 14571 6740 14613 6749
rect 14571 6700 14572 6740
rect 14612 6700 14708 6740
rect 14571 6691 14613 6700
rect 14475 6656 14517 6665
rect 14475 6616 14476 6656
rect 14516 6616 14517 6656
rect 14475 6607 14517 6616
rect 14379 6488 14421 6497
rect 14379 6448 14380 6488
rect 14420 6448 14421 6488
rect 14379 6439 14421 6448
rect 14284 6364 14325 6404
rect 14284 5984 14324 6364
rect 14380 6320 14420 6439
rect 14668 6329 14708 6700
rect 14572 6320 14612 6329
rect 14380 6280 14572 6320
rect 14572 6271 14612 6280
rect 14667 6320 14709 6329
rect 14667 6280 14668 6320
rect 14708 6280 14709 6320
rect 14667 6271 14709 6280
rect 14764 6161 14804 7120
rect 15051 7160 15093 7169
rect 15051 7120 15052 7160
rect 15092 7120 15093 7160
rect 15051 7111 15093 7120
rect 15052 7026 15092 7111
rect 14956 6992 14996 7001
rect 14860 6952 14956 6992
rect 14860 6488 14900 6952
rect 14956 6943 14996 6952
rect 15051 6740 15093 6749
rect 15051 6691 15052 6740
rect 15092 6691 15093 6740
rect 15052 6605 15092 6674
rect 14860 6439 14900 6448
rect 14956 6488 14996 6497
rect 14763 6152 14805 6161
rect 14763 6112 14764 6152
rect 14804 6112 14805 6152
rect 14763 6103 14805 6112
rect 14284 5944 14516 5984
rect 14092 5860 14324 5900
rect 13900 5776 14132 5816
rect 13611 5564 13653 5573
rect 13611 5524 13612 5564
rect 13652 5524 13653 5564
rect 13611 5515 13653 5524
rect 13803 5144 13845 5153
rect 13228 5104 13748 5144
rect 13132 4985 13172 5070
rect 12076 4936 12308 4976
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 11979 4640 12021 4649
rect 11979 4600 11980 4640
rect 12020 4600 12021 4640
rect 11979 4591 12021 4600
rect 11883 4388 11925 4397
rect 11883 4348 11884 4388
rect 11924 4348 11925 4388
rect 11883 4339 11925 4348
rect 11692 4087 11732 4096
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 11884 4136 11924 4339
rect 11884 4087 11924 4096
rect 11980 4136 12020 4591
rect 11980 4087 12020 4096
rect 11788 4002 11828 4087
rect 12076 3968 12116 4936
rect 12363 4927 12405 4936
rect 12939 4976 12981 4985
rect 12939 4936 12940 4976
rect 12980 4936 12981 4976
rect 12939 4927 12981 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13324 4976 13364 4985
rect 12268 4724 12308 4733
rect 12172 4684 12268 4724
rect 12172 4136 12212 4684
rect 12268 4675 12308 4684
rect 12172 4087 12212 4096
rect 11980 3928 12116 3968
rect 11883 3800 11925 3809
rect 11883 3760 11884 3800
rect 11924 3760 11925 3800
rect 11883 3751 11925 3760
rect 11156 3172 11348 3212
rect 11499 3212 11541 3221
rect 11499 3172 11500 3212
rect 11540 3172 11541 3212
rect 11116 3163 11156 3172
rect 11499 3163 11541 3172
rect 11116 1952 11156 1961
rect 10924 1912 11116 1952
rect 11884 1952 11924 3751
rect 11980 2876 12020 3928
rect 12364 3632 12404 4927
rect 12940 4842 12980 4927
rect 13132 4724 13172 4733
rect 12844 4684 13132 4724
rect 12459 4304 12501 4313
rect 12459 4264 12460 4304
rect 12500 4264 12501 4304
rect 12459 4255 12501 4264
rect 12460 3968 12500 4255
rect 12556 4136 12596 4145
rect 12596 4096 12788 4136
rect 12556 4087 12596 4096
rect 12460 3928 12596 3968
rect 12364 3583 12404 3592
rect 12076 3464 12116 3475
rect 12076 3389 12116 3424
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 12460 3464 12500 3473
rect 12075 3380 12117 3389
rect 12075 3340 12076 3380
rect 12116 3340 12117 3380
rect 12075 3331 12117 3340
rect 12268 3330 12308 3415
rect 12460 3221 12500 3424
rect 12556 3464 12596 3928
rect 12556 3415 12596 3424
rect 12748 3296 12788 4096
rect 12748 3247 12788 3256
rect 12459 3212 12501 3221
rect 12459 3172 12460 3212
rect 12500 3172 12501 3212
rect 12459 3163 12501 3172
rect 11980 2827 12020 2836
rect 12076 2624 12116 2633
rect 11980 1952 12020 1961
rect 11884 1912 11980 1952
rect 10731 1903 10773 1912
rect 11116 1903 11156 1912
rect 11980 1903 12020 1912
rect 10732 1818 10772 1903
rect 10539 1784 10581 1793
rect 10539 1744 10540 1784
rect 10580 1744 10581 1784
rect 10539 1735 10581 1744
rect 11212 1280 11252 1289
rect 10252 1240 11212 1280
rect 10156 1146 10196 1231
rect 10252 1112 10292 1240
rect 11212 1231 11252 1240
rect 10252 1063 10292 1072
rect 11884 1112 11924 1121
rect 12076 1112 12116 2584
rect 12844 2624 12884 4684
rect 13132 4675 13172 4684
rect 13324 4649 13364 4936
rect 13420 4976 13460 4985
rect 13323 4640 13365 4649
rect 13323 4600 13324 4640
rect 13364 4600 13365 4640
rect 13323 4591 13365 4600
rect 13420 4397 13460 4936
rect 13708 4976 13748 5104
rect 13803 5104 13804 5144
rect 13844 5104 13845 5144
rect 13803 5095 13845 5104
rect 13804 5060 13844 5095
rect 13804 5009 13844 5020
rect 13708 4927 13748 4936
rect 13900 4976 13940 5776
rect 14092 5732 14132 5776
rect 14092 5683 14132 5692
rect 13996 5648 14036 5657
rect 13996 5405 14036 5608
rect 14188 5648 14228 5657
rect 14188 5489 14228 5608
rect 14187 5480 14229 5489
rect 14187 5440 14188 5480
rect 14228 5440 14229 5480
rect 14187 5431 14229 5440
rect 13995 5396 14037 5405
rect 13995 5356 13996 5396
rect 14036 5356 14037 5396
rect 13995 5347 14037 5356
rect 13900 4927 13940 4936
rect 13996 4901 14036 5347
rect 14284 5153 14324 5860
rect 14379 5816 14421 5825
rect 14379 5776 14380 5816
rect 14420 5776 14421 5816
rect 14379 5767 14421 5776
rect 14380 5648 14420 5767
rect 14380 5599 14420 5608
rect 14476 5228 14516 5944
rect 14764 5405 14804 6103
rect 14859 5648 14901 5657
rect 14859 5608 14860 5648
rect 14900 5608 14901 5648
rect 14859 5599 14901 5608
rect 14763 5396 14805 5405
rect 14763 5356 14764 5396
rect 14804 5356 14805 5396
rect 14763 5347 14805 5356
rect 14380 5188 14516 5228
rect 14283 5144 14325 5153
rect 14283 5104 14284 5144
rect 14324 5104 14325 5144
rect 14283 5095 14325 5104
rect 14091 4976 14133 4985
rect 14091 4936 14092 4976
rect 14132 4936 14133 4976
rect 14091 4927 14133 4936
rect 14284 4976 14324 4985
rect 13995 4892 14037 4901
rect 13995 4852 13996 4892
rect 14036 4852 14037 4892
rect 13995 4843 14037 4852
rect 14092 4842 14132 4927
rect 14187 4724 14229 4733
rect 14187 4684 14188 4724
rect 14228 4684 14229 4724
rect 14187 4675 14229 4684
rect 14188 4590 14228 4675
rect 13419 4388 13461 4397
rect 13419 4348 13420 4388
rect 13460 4348 13461 4388
rect 13419 4339 13461 4348
rect 13420 4136 13460 4145
rect 13420 3809 13460 4096
rect 14284 3977 14324 4936
rect 14380 4145 14420 5188
rect 14764 5144 14804 5153
rect 14475 5060 14517 5069
rect 14475 5020 14476 5060
rect 14516 5020 14517 5060
rect 14475 5011 14517 5020
rect 14668 5060 14708 5069
rect 14476 4976 14516 5011
rect 14476 4925 14516 4936
rect 14572 4976 14612 4987
rect 14572 4901 14612 4936
rect 14571 4892 14613 4901
rect 14571 4852 14572 4892
rect 14612 4852 14613 4892
rect 14571 4843 14613 4852
rect 14668 4640 14708 5020
rect 14764 4817 14804 5104
rect 14860 5144 14900 5599
rect 14956 5573 14996 6448
rect 15244 6488 15284 7531
rect 15436 7328 15476 7337
rect 15436 6833 15476 7288
rect 15435 6824 15477 6833
rect 15435 6784 15436 6824
rect 15476 6784 15477 6824
rect 15435 6775 15477 6784
rect 15339 6656 15381 6665
rect 15339 6616 15340 6656
rect 15380 6616 15381 6656
rect 15339 6607 15381 6616
rect 15340 6522 15380 6607
rect 15244 6439 15284 6448
rect 15436 6488 15476 6497
rect 15436 5900 15476 6448
rect 15532 6488 15572 7867
rect 15628 7160 15668 7169
rect 15628 6665 15668 7120
rect 15627 6656 15669 6665
rect 15627 6616 15628 6656
rect 15668 6616 15669 6656
rect 15627 6607 15669 6616
rect 15723 6572 15765 6581
rect 15723 6532 15724 6572
rect 15764 6532 15765 6572
rect 15723 6523 15765 6532
rect 15572 6448 15668 6488
rect 15532 6439 15572 6448
rect 15436 5860 15572 5900
rect 15051 5648 15093 5657
rect 15051 5608 15052 5648
rect 15092 5608 15093 5648
rect 15051 5599 15093 5608
rect 15436 5648 15476 5657
rect 14955 5564 14997 5573
rect 14955 5524 14956 5564
rect 14996 5524 14997 5564
rect 14955 5515 14997 5524
rect 14860 5095 14900 5104
rect 14956 5069 14996 5515
rect 15052 5514 15092 5599
rect 15340 5480 15380 5491
rect 15340 5405 15380 5440
rect 15339 5396 15381 5405
rect 15339 5356 15340 5396
rect 15380 5356 15381 5396
rect 15339 5347 15381 5356
rect 14955 5060 14997 5069
rect 14955 5020 14956 5060
rect 14996 5020 14997 5060
rect 14955 5011 14997 5020
rect 15148 4976 15188 4985
rect 15188 4936 15380 4976
rect 15148 4927 15188 4936
rect 14763 4808 14805 4817
rect 14763 4768 14764 4808
rect 14804 4768 14805 4808
rect 14763 4759 14805 4768
rect 15147 4808 15189 4817
rect 15147 4768 15148 4808
rect 15188 4768 15189 4808
rect 15147 4759 15189 4768
rect 14476 4600 14708 4640
rect 14476 4304 14516 4600
rect 14571 4304 14613 4313
rect 14476 4264 14572 4304
rect 14612 4264 14613 4304
rect 14571 4255 14613 4264
rect 14668 4264 15092 4304
rect 14572 4170 14612 4255
rect 14379 4136 14421 4145
rect 14379 4096 14380 4136
rect 14420 4096 14421 4136
rect 14379 4087 14421 4096
rect 14283 3968 14325 3977
rect 14283 3928 14284 3968
rect 14324 3928 14325 3968
rect 14283 3919 14325 3928
rect 13419 3800 13461 3809
rect 13419 3760 13420 3800
rect 13460 3760 13461 3800
rect 13419 3751 13461 3760
rect 14475 3632 14517 3641
rect 14475 3592 14476 3632
rect 14516 3592 14517 3632
rect 14475 3583 14517 3592
rect 14476 3498 14516 3583
rect 14572 3464 14612 3473
rect 14668 3464 14708 4264
rect 14763 4136 14805 4145
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 14860 4136 14900 4145
rect 14764 4002 14804 4087
rect 14860 3884 14900 4096
rect 14764 3844 14900 3884
rect 14956 4136 14996 4145
rect 14764 3557 14804 3844
rect 14859 3716 14901 3725
rect 14859 3676 14860 3716
rect 14900 3676 14901 3716
rect 14859 3667 14901 3676
rect 14763 3548 14805 3557
rect 14763 3508 14764 3548
rect 14804 3508 14805 3548
rect 14763 3499 14805 3508
rect 14612 3424 14708 3464
rect 14860 3464 14900 3667
rect 14956 3632 14996 4096
rect 15052 4136 15092 4264
rect 15052 4087 15092 4096
rect 15052 3632 15092 3641
rect 14956 3592 15052 3632
rect 15052 3583 15092 3592
rect 14956 3464 14996 3473
rect 14860 3424 14956 3464
rect 14572 3415 14612 3424
rect 14956 3415 14996 3424
rect 15148 3464 15188 4759
rect 15243 4304 15285 4313
rect 15243 4264 15244 4304
rect 15284 4264 15285 4304
rect 15243 4255 15285 4264
rect 15244 4136 15284 4255
rect 15244 4087 15284 4096
rect 15148 3415 15188 3424
rect 15244 3464 15284 3475
rect 15244 3389 15284 3424
rect 13131 3380 13173 3389
rect 13131 3340 13132 3380
rect 13172 3340 13173 3380
rect 13131 3331 13173 3340
rect 15243 3380 15285 3389
rect 15243 3340 15244 3380
rect 15284 3340 15285 3380
rect 15243 3331 15285 3340
rect 12844 2575 12884 2584
rect 13132 1952 13172 3331
rect 13324 3296 13364 3305
rect 13228 2624 13268 2633
rect 13324 2624 13364 3256
rect 14764 3212 14804 3221
rect 14092 2633 14132 2718
rect 13268 2584 13364 2624
rect 14091 2624 14133 2633
rect 14091 2584 14092 2624
rect 14132 2584 14133 2624
rect 13228 2575 13268 2584
rect 14091 2575 14133 2584
rect 14764 2540 14804 3172
rect 15244 2876 15284 2885
rect 15340 2876 15380 4936
rect 15436 4817 15476 5608
rect 15532 5489 15572 5860
rect 15628 5825 15668 6448
rect 15724 6438 15764 6523
rect 15627 5816 15669 5825
rect 15627 5776 15628 5816
rect 15668 5776 15669 5816
rect 16012 5816 16052 8455
rect 16204 8000 16244 9304
rect 16396 9092 16436 9388
rect 16491 9344 16533 9353
rect 16491 9304 16492 9344
rect 16532 9304 16533 9344
rect 16491 9295 16533 9304
rect 16492 9210 16532 9295
rect 16300 9052 16436 9092
rect 16300 8924 16340 9052
rect 16300 8875 16340 8884
rect 16587 8840 16629 8849
rect 16587 8800 16588 8840
rect 16628 8800 16629 8840
rect 16587 8791 16629 8800
rect 16779 8840 16821 8849
rect 16779 8800 16780 8840
rect 16820 8800 16821 8840
rect 16779 8791 16821 8800
rect 16299 8672 16341 8681
rect 16299 8632 16300 8672
rect 16340 8632 16341 8672
rect 16299 8623 16341 8632
rect 16300 8538 16340 8623
rect 16204 7951 16244 7960
rect 16491 8000 16533 8009
rect 16491 7960 16492 8000
rect 16532 7960 16533 8000
rect 16491 7951 16533 7960
rect 16492 7328 16532 7951
rect 16492 7279 16532 7288
rect 16300 6992 16340 7001
rect 16107 6824 16149 6833
rect 16107 6784 16108 6824
rect 16148 6784 16149 6824
rect 16107 6775 16149 6784
rect 16108 6488 16148 6775
rect 16300 6581 16340 6952
rect 16299 6572 16341 6581
rect 16299 6532 16300 6572
rect 16340 6532 16341 6572
rect 16299 6523 16341 6532
rect 16108 6439 16148 6448
rect 16299 6320 16341 6329
rect 16299 6280 16300 6320
rect 16340 6280 16341 6320
rect 16299 6271 16341 6280
rect 16012 5776 16148 5816
rect 15627 5767 15669 5776
rect 15723 5732 15765 5741
rect 15723 5692 15724 5732
rect 15764 5692 15765 5732
rect 15723 5683 15765 5692
rect 15725 5665 15765 5683
rect 16012 5648 16052 5657
rect 15725 5598 15765 5625
rect 15916 5608 16012 5648
rect 15531 5480 15573 5489
rect 15820 5480 15860 5489
rect 15531 5440 15532 5480
rect 15572 5440 15573 5480
rect 15531 5431 15573 5440
rect 15724 5440 15820 5480
rect 15531 5060 15573 5069
rect 15531 5020 15532 5060
rect 15572 5020 15573 5060
rect 15531 5011 15573 5020
rect 15435 4808 15477 4817
rect 15435 4768 15436 4808
rect 15476 4768 15477 4808
rect 15435 4759 15477 4768
rect 15435 3464 15477 3473
rect 15435 3424 15436 3464
rect 15476 3424 15477 3464
rect 15435 3415 15477 3424
rect 15436 3053 15476 3415
rect 15532 3380 15572 5011
rect 15724 3809 15764 5440
rect 15820 5431 15860 5440
rect 15819 4808 15861 4817
rect 15819 4768 15820 4808
rect 15860 4768 15861 4808
rect 15819 4759 15861 4768
rect 15820 4674 15860 4759
rect 15916 4136 15956 5608
rect 16012 5599 16052 5608
rect 16108 5228 16148 5776
rect 16300 5648 16340 6271
rect 16395 5816 16437 5825
rect 16395 5776 16396 5816
rect 16436 5776 16437 5816
rect 16395 5767 16437 5776
rect 16300 5599 16340 5608
rect 16203 5480 16245 5489
rect 16396 5480 16436 5767
rect 16203 5440 16204 5480
rect 16244 5440 16245 5480
rect 16203 5431 16245 5440
rect 16300 5440 16436 5480
rect 16204 5346 16244 5431
rect 16108 5188 16244 5228
rect 16107 5060 16149 5069
rect 16107 5020 16108 5060
rect 16148 5020 16149 5060
rect 16107 5011 16149 5020
rect 16011 4976 16053 4985
rect 16011 4936 16012 4976
rect 16052 4936 16053 4976
rect 16011 4927 16053 4936
rect 16108 4976 16148 5011
rect 16012 4842 16052 4927
rect 16108 4925 16148 4936
rect 16108 4145 16148 4230
rect 16107 4136 16149 4145
rect 15916 4096 16052 4136
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 15723 3800 15765 3809
rect 15723 3760 15724 3800
rect 15764 3760 15765 3800
rect 15723 3751 15765 3760
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 15532 3331 15572 3340
rect 15724 3380 15764 3389
rect 15627 3296 15669 3305
rect 15627 3256 15628 3296
rect 15668 3256 15669 3296
rect 15627 3247 15669 3256
rect 15628 3162 15668 3247
rect 15724 3221 15764 3340
rect 15820 3330 15860 3415
rect 15723 3212 15765 3221
rect 15723 3172 15724 3212
rect 15764 3172 15765 3212
rect 15723 3163 15765 3172
rect 15435 3044 15477 3053
rect 15435 3004 15436 3044
rect 15476 3004 15477 3044
rect 15435 2995 15477 3004
rect 15284 2836 15380 2876
rect 15244 2827 15284 2836
rect 15724 2624 15764 3163
rect 15724 2575 15764 2584
rect 15916 2624 15956 3919
rect 16012 2801 16052 4096
rect 16107 4096 16108 4136
rect 16148 4096 16149 4136
rect 16107 4087 16149 4096
rect 16204 3464 16244 5188
rect 16300 4976 16340 5440
rect 16300 4724 16340 4936
rect 16395 4976 16437 4985
rect 16395 4936 16396 4976
rect 16436 4936 16437 4976
rect 16395 4927 16437 4936
rect 16588 4976 16628 8791
rect 16684 8672 16724 8681
rect 16684 8429 16724 8632
rect 16780 8672 16820 8791
rect 16780 8623 16820 8632
rect 16876 8672 16916 9715
rect 16972 9512 17012 9521
rect 17164 9512 17204 9521
rect 17012 9472 17108 9512
rect 16972 9463 17012 9472
rect 16971 9260 17013 9269
rect 16971 9220 16972 9260
rect 17012 9220 17013 9260
rect 16971 9211 17013 9220
rect 16972 9126 17012 9211
rect 16876 8623 16916 8632
rect 16972 8672 17012 8681
rect 17068 8672 17108 9472
rect 17164 9353 17204 9472
rect 17260 9512 17300 11152
rect 17356 11117 17396 11148
rect 17355 11108 17397 11117
rect 17355 11068 17356 11108
rect 17396 11068 17397 11108
rect 17355 11059 17397 11068
rect 17356 11024 17396 11059
rect 17356 10697 17396 10984
rect 17451 11024 17493 11033
rect 17451 10984 17452 11024
rect 17492 10984 17493 11024
rect 17451 10975 17493 10984
rect 17644 11024 17684 11320
rect 17836 11033 17876 11395
rect 17644 10975 17684 10984
rect 17835 11024 17877 11033
rect 17835 10984 17836 11024
rect 17876 10984 17877 11024
rect 17835 10975 17877 10984
rect 18315 11024 18357 11033
rect 18315 10984 18316 11024
rect 18356 10984 18357 11024
rect 18315 10975 18357 10984
rect 18508 11024 18548 11035
rect 17452 10890 17492 10975
rect 17547 10940 17589 10949
rect 17547 10900 17548 10940
rect 17588 10900 17589 10940
rect 17547 10891 17589 10900
rect 17355 10688 17397 10697
rect 17355 10648 17356 10688
rect 17396 10648 17397 10688
rect 17355 10639 17397 10648
rect 17548 10193 17588 10891
rect 18316 10856 18356 10975
rect 18508 10949 18548 10984
rect 18892 11024 18932 11395
rect 18892 10975 18932 10984
rect 18988 11024 19028 12067
rect 19084 12041 19124 12496
rect 19367 12536 19407 12545
rect 19468 12536 19508 12655
rect 19563 12620 19605 12629
rect 19563 12580 19564 12620
rect 19604 12580 19605 12620
rect 19563 12571 19605 12580
rect 19851 12620 19893 12629
rect 19851 12580 19852 12620
rect 19892 12580 19893 12620
rect 19851 12571 19893 12580
rect 19407 12496 19412 12536
rect 19367 12487 19412 12496
rect 19468 12487 19508 12496
rect 19564 12536 19604 12571
rect 19083 12032 19125 12041
rect 19083 11992 19084 12032
rect 19124 11992 19125 12032
rect 19083 11983 19125 11992
rect 19372 11789 19412 12487
rect 19467 12284 19509 12293
rect 19467 12244 19468 12284
rect 19508 12244 19509 12284
rect 19467 12235 19509 12244
rect 19468 11873 19508 12235
rect 19467 11864 19509 11873
rect 19467 11824 19468 11864
rect 19508 11824 19509 11864
rect 19467 11815 19509 11824
rect 19276 11780 19316 11789
rect 18507 10940 18549 10949
rect 18507 10900 18508 10940
rect 18548 10900 18549 10940
rect 18507 10891 18549 10900
rect 18316 10807 18356 10816
rect 18892 10772 18932 10781
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 17547 10184 17589 10193
rect 17547 10144 17548 10184
rect 17588 10144 17589 10184
rect 17547 10135 17589 10144
rect 18316 10184 18356 10193
rect 18356 10144 18740 10184
rect 18316 10135 18356 10144
rect 17260 9463 17300 9472
rect 17548 9512 17588 10135
rect 17740 10100 17780 10109
rect 17932 10100 17972 10109
rect 17780 10060 17932 10100
rect 17740 10051 17780 10060
rect 17932 10051 17972 10060
rect 17548 9463 17588 9472
rect 17163 9344 17205 9353
rect 17163 9304 17164 9344
rect 17204 9304 17205 9344
rect 17163 9295 17205 9304
rect 18700 9344 18740 10144
rect 18892 10109 18932 10732
rect 18891 10100 18933 10109
rect 18891 10060 18892 10100
rect 18932 10060 18933 10100
rect 18891 10051 18933 10060
rect 18988 10025 19028 10984
rect 19084 11740 19276 11780
rect 19084 10781 19124 11740
rect 19276 11731 19316 11740
rect 19371 11780 19413 11789
rect 19371 11740 19372 11780
rect 19412 11740 19413 11780
rect 19371 11731 19413 11740
rect 19179 11612 19221 11621
rect 19179 11572 19180 11612
rect 19220 11572 19221 11612
rect 19179 11563 19221 11572
rect 19180 11024 19220 11563
rect 19275 11528 19317 11537
rect 19275 11488 19276 11528
rect 19316 11488 19317 11528
rect 19275 11479 19317 11488
rect 19180 10975 19220 10984
rect 19276 11024 19316 11479
rect 19372 11033 19412 11731
rect 19564 11705 19604 12496
rect 19756 12536 19796 12547
rect 19756 12461 19796 12496
rect 19852 12536 19892 12571
rect 19755 12452 19797 12461
rect 19755 12412 19756 12452
rect 19796 12412 19797 12452
rect 19755 12403 19797 12412
rect 19852 12284 19892 12496
rect 19660 12244 19892 12284
rect 19563 11696 19605 11705
rect 19563 11656 19564 11696
rect 19604 11656 19605 11696
rect 19563 11647 19605 11656
rect 19660 11696 19700 12244
rect 19755 12032 19797 12041
rect 19755 11992 19756 12032
rect 19796 11992 19892 12032
rect 19755 11983 19797 11992
rect 19755 11864 19797 11873
rect 19755 11824 19756 11864
rect 19796 11824 19797 11864
rect 19755 11815 19797 11824
rect 19660 11537 19700 11656
rect 19756 11696 19796 11815
rect 19756 11647 19796 11656
rect 19659 11528 19701 11537
rect 19659 11488 19660 11528
rect 19700 11488 19701 11528
rect 19659 11479 19701 11488
rect 19852 11528 19892 11992
rect 19948 11873 19988 13504
rect 20139 13208 20181 13217
rect 20139 13168 20140 13208
rect 20180 13168 20181 13208
rect 20139 13159 20181 13168
rect 20140 13082 20180 13159
rect 20140 13033 20180 13042
rect 20139 12956 20181 12965
rect 20139 12916 20140 12956
rect 20180 12916 20181 12956
rect 20236 12956 20276 14755
rect 20332 14720 20372 14932
rect 20332 14671 20372 14680
rect 20620 14720 20660 15511
rect 20716 15485 20756 15520
rect 20812 15560 20852 15569
rect 20715 15476 20757 15485
rect 20715 15436 20716 15476
rect 20756 15436 20757 15476
rect 20715 15427 20757 15436
rect 20812 15149 20852 15520
rect 20908 15560 20948 15569
rect 20811 15140 20853 15149
rect 20620 14671 20660 14680
rect 20716 15100 20812 15140
rect 20852 15100 20853 15140
rect 20523 14552 20565 14561
rect 20523 14512 20524 14552
rect 20564 14512 20565 14552
rect 20523 14503 20565 14512
rect 20524 14418 20564 14503
rect 20619 14468 20661 14477
rect 20619 14428 20620 14468
rect 20660 14428 20661 14468
rect 20619 14419 20661 14428
rect 20428 14057 20468 14142
rect 20524 14132 20564 14141
rect 20427 14048 20469 14057
rect 20427 14008 20428 14048
rect 20468 14008 20469 14048
rect 20427 13999 20469 14008
rect 20427 13880 20469 13889
rect 20427 13840 20428 13880
rect 20468 13840 20469 13880
rect 20427 13831 20469 13840
rect 20331 13208 20373 13217
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 20428 13208 20468 13831
rect 20524 13217 20564 14092
rect 20428 13159 20468 13168
rect 20523 13208 20565 13217
rect 20523 13168 20524 13208
rect 20564 13168 20565 13208
rect 20523 13159 20565 13168
rect 20332 13074 20372 13159
rect 20620 13082 20660 14419
rect 20524 13042 20660 13082
rect 20236 12916 20372 12956
rect 20139 12907 20181 12916
rect 20043 12536 20085 12545
rect 20043 12496 20044 12536
rect 20084 12496 20085 12536
rect 20043 12487 20085 12496
rect 20140 12536 20180 12907
rect 20235 12704 20277 12713
rect 20235 12664 20236 12704
rect 20276 12664 20277 12704
rect 20235 12655 20277 12664
rect 20140 12487 20180 12496
rect 20236 12536 20276 12655
rect 20236 12487 20276 12496
rect 20332 12536 20372 12916
rect 20044 12402 20084 12487
rect 20043 12284 20085 12293
rect 20043 12244 20044 12284
rect 20084 12244 20085 12284
rect 20043 12235 20085 12244
rect 19947 11864 19989 11873
rect 19947 11824 19948 11864
rect 19988 11824 19989 11864
rect 19947 11815 19989 11824
rect 19947 11696 19989 11705
rect 19947 11656 19948 11696
rect 19988 11656 19989 11696
rect 19947 11647 19989 11656
rect 20044 11696 20084 12235
rect 20200 11780 20242 11789
rect 20200 11740 20201 11780
rect 20241 11740 20242 11780
rect 20200 11731 20242 11740
rect 19948 11562 19988 11647
rect 19852 11479 19892 11488
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 19372 11024 19417 11033
rect 19372 10984 19377 11024
rect 19083 10772 19125 10781
rect 19083 10732 19084 10772
rect 19124 10732 19125 10772
rect 19083 10723 19125 10732
rect 19084 10184 19124 10723
rect 19180 10184 19220 10193
rect 19084 10144 19180 10184
rect 18987 10016 19029 10025
rect 18987 9976 18988 10016
rect 19028 9976 19029 10016
rect 18987 9967 19029 9976
rect 18700 9295 18740 9304
rect 17547 9260 17589 9269
rect 18220 9260 18260 9269
rect 17547 9220 17548 9260
rect 17588 9220 17589 9260
rect 17547 9211 17589 9220
rect 18124 9220 18220 9260
rect 17012 8632 17108 8672
rect 17164 8672 17204 8681
rect 16972 8623 17012 8632
rect 16683 8420 16725 8429
rect 16683 8380 16684 8420
rect 16724 8380 16725 8420
rect 16683 8371 16725 8380
rect 17164 8168 17204 8632
rect 17356 8168 17396 8177
rect 17164 8128 17356 8168
rect 17356 8119 17396 8128
rect 17548 8084 17588 9211
rect 18028 8840 18068 8849
rect 17932 8800 18028 8840
rect 17548 8035 17588 8044
rect 17836 8504 17876 8513
rect 16971 8000 17013 8009
rect 16971 7960 16972 8000
rect 17012 7960 17013 8000
rect 16971 7951 17013 7960
rect 16876 6992 16916 7001
rect 16876 6329 16916 6952
rect 16972 6488 17012 7951
rect 17547 7160 17589 7169
rect 17547 7120 17548 7160
rect 17588 7120 17589 7160
rect 17547 7111 17589 7120
rect 17836 7160 17876 8464
rect 17932 8000 17972 8800
rect 18028 8791 18068 8800
rect 17932 7951 17972 7960
rect 17836 7111 17876 7120
rect 18027 7160 18069 7169
rect 18027 7120 18028 7160
rect 18068 7120 18069 7160
rect 18027 7111 18069 7120
rect 17548 7026 17588 7111
rect 17740 6992 17780 7001
rect 17740 6749 17780 6952
rect 17739 6740 17781 6749
rect 17739 6700 17740 6740
rect 17780 6700 17781 6740
rect 17739 6691 17781 6700
rect 16972 6439 17012 6448
rect 16875 6320 16917 6329
rect 16875 6280 16876 6320
rect 16916 6280 16917 6320
rect 18028 6320 18068 7111
rect 18124 6497 18164 9220
rect 18220 9211 18260 9220
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 19180 8009 19220 10144
rect 19276 8429 19316 10984
rect 19377 10975 19417 10984
rect 19851 11024 19893 11033
rect 19851 10984 19852 11024
rect 19892 10984 19893 11024
rect 19851 10975 19893 10984
rect 19852 10890 19892 10975
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 20044 9773 20084 11656
rect 20201 11711 20241 11731
rect 20201 11645 20241 11671
rect 20332 11285 20372 12496
rect 20331 11276 20373 11285
rect 20331 11236 20332 11276
rect 20372 11236 20373 11276
rect 20331 11227 20373 11236
rect 20139 10772 20181 10781
rect 20139 10732 20140 10772
rect 20180 10732 20181 10772
rect 20139 10723 20181 10732
rect 20140 10638 20180 10723
rect 20332 10445 20372 11227
rect 20331 10436 20373 10445
rect 20331 10396 20332 10436
rect 20372 10396 20373 10436
rect 20331 10387 20373 10396
rect 20331 10268 20373 10277
rect 20331 10228 20332 10268
rect 20372 10228 20373 10268
rect 20331 10219 20373 10228
rect 20332 10134 20372 10219
rect 20043 9764 20085 9773
rect 20043 9724 20044 9764
rect 20084 9724 20085 9764
rect 20043 9715 20085 9724
rect 19756 8840 19796 8849
rect 19756 8504 19796 8800
rect 20524 8765 20564 13042
rect 20716 12713 20756 15100
rect 20811 15091 20853 15100
rect 20812 14720 20852 14729
rect 20812 14057 20852 14680
rect 20811 14048 20853 14057
rect 20811 14008 20812 14048
rect 20852 14008 20853 14048
rect 20811 13999 20853 14008
rect 20908 13973 20948 15520
rect 21483 15560 21525 15569
rect 21483 15520 21484 15560
rect 21524 15520 21525 15560
rect 21868 15560 21908 15569
rect 21483 15511 21525 15520
rect 21580 15518 21620 15527
rect 21484 15426 21524 15511
rect 21196 15308 21236 15317
rect 21004 15268 21196 15308
rect 21004 14216 21044 15268
rect 21196 15259 21236 15268
rect 21580 14720 21620 15478
rect 21484 14680 21620 14720
rect 21676 14720 21716 14731
rect 21868 14729 21908 15520
rect 21963 15560 22005 15569
rect 21963 15520 21964 15560
rect 22004 15520 22005 15560
rect 21963 15511 22005 15520
rect 22060 15560 22100 15569
rect 21964 15476 22004 15511
rect 21964 15425 22004 15436
rect 22060 14897 22100 15520
rect 22252 15560 22292 15571
rect 22252 15485 22292 15520
rect 22251 15476 22293 15485
rect 22251 15436 22252 15476
rect 22292 15436 22293 15476
rect 22251 15427 22293 15436
rect 22252 15308 22292 15317
rect 22059 14888 22101 14897
rect 22059 14848 22060 14888
rect 22100 14848 22101 14888
rect 22059 14839 22101 14848
rect 21004 14176 21236 14216
rect 21004 14048 21044 14176
rect 21004 13999 21044 14008
rect 21100 14048 21140 14057
rect 20907 13964 20949 13973
rect 20907 13924 20908 13964
rect 20948 13924 20949 13964
rect 20907 13915 20949 13924
rect 21100 13217 21140 14008
rect 21099 13208 21141 13217
rect 21099 13168 21100 13208
rect 21140 13168 21141 13208
rect 21099 13159 21141 13168
rect 21196 13208 21236 14176
rect 21291 14132 21333 14141
rect 21291 14092 21292 14132
rect 21332 14092 21333 14132
rect 21291 14083 21333 14092
rect 21292 14048 21332 14083
rect 21292 13997 21332 14008
rect 21196 13159 21236 13168
rect 21292 13796 21332 13805
rect 21292 13208 21332 13756
rect 21484 13301 21524 14680
rect 21676 14645 21716 14680
rect 21867 14720 21909 14729
rect 21867 14680 21868 14720
rect 21908 14680 21909 14720
rect 21867 14671 21909 14680
rect 22060 14720 22100 14729
rect 21675 14636 21717 14645
rect 21675 14596 21676 14636
rect 21716 14596 21717 14636
rect 21675 14587 21717 14596
rect 21579 14552 21621 14561
rect 21579 14512 21580 14552
rect 21620 14512 21621 14552
rect 21579 14503 21621 14512
rect 21580 14048 21620 14503
rect 21675 14216 21717 14225
rect 21675 14176 21676 14216
rect 21716 14176 21717 14216
rect 21675 14167 21717 14176
rect 21580 13999 21620 14008
rect 21676 14048 21716 14167
rect 21868 14132 21908 14141
rect 21676 13999 21716 14008
rect 21772 14048 21812 14059
rect 21772 13973 21812 14008
rect 21868 14040 21908 14092
rect 21868 14000 21913 14040
rect 21771 13964 21813 13973
rect 21771 13924 21772 13964
rect 21812 13924 21813 13964
rect 21771 13915 21813 13924
rect 21873 13880 21913 14000
rect 21868 13840 21913 13880
rect 21868 13628 21908 13840
rect 21868 13588 22004 13628
rect 21613 13460 21655 13469
rect 21613 13420 21614 13460
rect 21654 13420 21655 13460
rect 21613 13411 21655 13420
rect 21867 13460 21909 13469
rect 21867 13420 21868 13460
rect 21908 13420 21909 13460
rect 21867 13411 21909 13420
rect 21483 13292 21525 13301
rect 21483 13252 21484 13292
rect 21524 13252 21525 13292
rect 21483 13243 21525 13252
rect 21614 13223 21654 13411
rect 21614 13174 21654 13183
rect 21772 13208 21812 13217
rect 21292 13159 21332 13168
rect 21100 13074 21140 13159
rect 21388 13040 21428 13049
rect 21292 13000 21388 13040
rect 20715 12704 20757 12713
rect 20715 12664 20716 12704
rect 20756 12664 20757 12704
rect 20715 12655 20757 12664
rect 20620 12536 20660 12545
rect 20620 12125 20660 12496
rect 20716 12536 20756 12655
rect 21195 12620 21237 12629
rect 21195 12580 21196 12620
rect 21236 12580 21237 12620
rect 21195 12571 21237 12580
rect 20716 12487 20756 12496
rect 20811 12536 20853 12545
rect 20811 12496 20812 12536
rect 20852 12496 20853 12536
rect 20811 12487 20853 12496
rect 20908 12536 20948 12545
rect 21100 12536 21140 12545
rect 20948 12496 21100 12536
rect 20908 12487 20948 12496
rect 21100 12487 21140 12496
rect 20812 12402 20852 12487
rect 21196 12486 21236 12571
rect 21292 12536 21332 13000
rect 21388 12991 21428 13000
rect 21483 13040 21525 13049
rect 21483 13000 21484 13040
rect 21524 13000 21525 13040
rect 21483 12991 21525 13000
rect 21675 13040 21717 13049
rect 21675 13000 21676 13040
rect 21716 13000 21717 13040
rect 21675 12991 21717 13000
rect 21484 12788 21524 12991
rect 21676 12906 21716 12991
rect 21292 12487 21332 12496
rect 21388 12748 21524 12788
rect 21388 12536 21428 12748
rect 21579 12620 21621 12629
rect 21579 12580 21580 12620
rect 21620 12580 21621 12620
rect 21579 12571 21621 12580
rect 21388 12487 21428 12496
rect 21580 12536 21620 12571
rect 21580 12485 21620 12496
rect 20619 12116 20661 12125
rect 20619 12076 20620 12116
rect 20660 12076 20661 12116
rect 20619 12067 20661 12076
rect 20620 11285 20660 12067
rect 21196 11864 21236 11873
rect 21772 11864 21812 13168
rect 21868 13208 21908 13411
rect 21868 12797 21908 13168
rect 21867 12788 21909 12797
rect 21867 12748 21868 12788
rect 21908 12748 21909 12788
rect 21867 12739 21909 12748
rect 21196 11360 21236 11824
rect 21484 11824 21812 11864
rect 21484 11360 21524 11824
rect 21771 11696 21813 11705
rect 21771 11656 21772 11696
rect 21812 11656 21813 11696
rect 21771 11647 21813 11656
rect 21772 11562 21812 11647
rect 21100 11320 21236 11360
rect 21388 11320 21524 11360
rect 20619 11276 20661 11285
rect 20619 11236 20620 11276
rect 20660 11236 20661 11276
rect 20619 11227 20661 11236
rect 20812 11024 20852 11033
rect 20715 10772 20757 10781
rect 20715 10732 20716 10772
rect 20756 10732 20757 10772
rect 20715 10723 20757 10732
rect 20716 10184 20756 10723
rect 20812 10193 20852 10984
rect 21004 10772 21044 10781
rect 20716 10135 20756 10144
rect 20811 10184 20853 10193
rect 20811 10144 20812 10184
rect 20852 10144 20853 10184
rect 20811 10135 20853 10144
rect 20907 10100 20949 10109
rect 20907 10060 20908 10100
rect 20948 10060 20949 10100
rect 20907 10051 20949 10060
rect 20908 9344 20948 10051
rect 21004 9512 21044 10732
rect 21100 10184 21140 11320
rect 21388 10697 21428 11320
rect 21676 11024 21716 11033
rect 21484 10984 21676 11024
rect 21387 10688 21429 10697
rect 21387 10648 21388 10688
rect 21428 10648 21429 10688
rect 21387 10639 21429 10648
rect 21100 10135 21140 10144
rect 21388 10109 21428 10639
rect 21484 10277 21524 10984
rect 21676 10975 21716 10984
rect 21868 11024 21908 11033
rect 21964 11024 22004 13588
rect 22060 13469 22100 14680
rect 22252 14225 22292 15268
rect 22251 14216 22293 14225
rect 22251 14176 22252 14216
rect 22292 14176 22293 14216
rect 22251 14167 22293 14176
rect 22155 14048 22197 14057
rect 22155 14008 22156 14048
rect 22196 14008 22197 14048
rect 22155 13999 22197 14008
rect 22059 13460 22101 13469
rect 22059 13420 22060 13460
rect 22100 13420 22101 13460
rect 22059 13411 22101 13420
rect 22059 13292 22101 13301
rect 22059 13252 22060 13292
rect 22100 13252 22101 13292
rect 22059 13243 22101 13252
rect 22060 13208 22100 13243
rect 22060 13157 22100 13168
rect 22156 13208 22196 13999
rect 22156 13159 22196 13168
rect 22348 12956 22388 15940
rect 22540 15930 22580 16015
rect 22827 15812 22869 15821
rect 22827 15772 22828 15812
rect 22868 15772 22869 15812
rect 22827 15763 22869 15772
rect 22731 15644 22773 15653
rect 22731 15604 22732 15644
rect 22772 15604 22773 15644
rect 22731 15595 22773 15604
rect 22444 15560 22484 15569
rect 22444 15401 22484 15520
rect 22539 15560 22581 15569
rect 22539 15520 22540 15560
rect 22580 15520 22581 15560
rect 22539 15511 22581 15520
rect 22732 15560 22772 15595
rect 22540 15426 22580 15511
rect 22732 15509 22772 15520
rect 22828 15476 22868 15763
rect 23019 15728 23061 15737
rect 23019 15688 23020 15728
rect 23060 15688 23061 15728
rect 23019 15679 23061 15688
rect 22923 15560 22965 15569
rect 22923 15520 22924 15560
rect 22964 15520 22965 15560
rect 22923 15511 22965 15520
rect 22828 15427 22868 15436
rect 22443 15392 22485 15401
rect 22443 15352 22444 15392
rect 22484 15352 22485 15392
rect 22443 15343 22485 15352
rect 22924 15392 22964 15511
rect 22924 15343 22964 15352
rect 23020 15476 23060 15679
rect 23020 15224 23060 15436
rect 22924 15184 23060 15224
rect 23116 15560 23156 15569
rect 22924 14720 22964 15184
rect 22924 14671 22964 14680
rect 23019 14636 23061 14645
rect 23019 14596 23020 14636
rect 23060 14596 23061 14636
rect 23019 14587 23061 14596
rect 23020 14057 23060 14587
rect 23019 14048 23061 14057
rect 23019 14008 23020 14048
rect 23060 14008 23061 14048
rect 23019 13999 23061 14008
rect 23020 13914 23060 13999
rect 22540 13796 22580 13805
rect 22443 13208 22485 13217
rect 22443 13168 22444 13208
rect 22484 13168 22485 13208
rect 22443 13159 22485 13168
rect 22444 13074 22484 13159
rect 22348 12916 22484 12956
rect 22252 12284 22292 12293
rect 22252 11705 22292 12244
rect 22156 11696 22196 11705
rect 22156 11360 22196 11656
rect 22251 11696 22293 11705
rect 22251 11656 22252 11696
rect 22292 11656 22293 11696
rect 22251 11647 22293 11656
rect 22156 11320 22388 11360
rect 22155 11108 22197 11117
rect 22155 11068 22156 11108
rect 22196 11068 22197 11108
rect 22155 11059 22197 11068
rect 21908 10984 22004 11024
rect 22059 11024 22101 11033
rect 22059 10984 22060 11024
rect 22100 10984 22101 11024
rect 21868 10975 21908 10984
rect 22059 10975 22101 10984
rect 22156 11024 22196 11059
rect 22060 10890 22100 10975
rect 22156 10973 22196 10984
rect 22348 10856 22388 11320
rect 22348 10807 22388 10816
rect 21867 10772 21909 10781
rect 21867 10732 21868 10772
rect 21908 10732 21909 10772
rect 21867 10723 21909 10732
rect 21868 10638 21908 10723
rect 22444 10604 22484 12916
rect 22540 12713 22580 13756
rect 22828 13208 22868 13217
rect 22868 13168 22964 13208
rect 22828 13159 22868 13168
rect 22539 12704 22581 12713
rect 22539 12664 22540 12704
rect 22580 12664 22581 12704
rect 22539 12655 22581 12664
rect 22540 11117 22580 12655
rect 22924 12368 22964 13168
rect 22924 12319 22964 12328
rect 23019 11696 23061 11705
rect 23019 11656 23020 11696
rect 23060 11656 23061 11696
rect 23019 11647 23061 11656
rect 22539 11108 22581 11117
rect 22539 11068 22540 11108
rect 22580 11068 22581 11108
rect 22539 11059 22581 11068
rect 21964 10564 22484 10604
rect 21964 10352 22004 10564
rect 22059 10436 22101 10445
rect 22059 10396 22060 10436
rect 22100 10396 22101 10436
rect 22059 10387 22101 10396
rect 21868 10312 22004 10352
rect 21483 10268 21525 10277
rect 21483 10228 21484 10268
rect 21524 10228 21525 10268
rect 21483 10219 21525 10228
rect 21387 10100 21429 10109
rect 21387 10060 21388 10100
rect 21428 10060 21429 10100
rect 21387 10051 21429 10060
rect 21100 9512 21140 9521
rect 21004 9472 21100 9512
rect 21100 9463 21140 9472
rect 21484 9512 21524 10219
rect 21484 9463 21524 9472
rect 21676 9512 21716 9521
rect 20908 9295 20948 9304
rect 21676 8933 21716 9472
rect 21675 8924 21717 8933
rect 21675 8884 21676 8924
rect 21716 8884 21717 8924
rect 21675 8875 21717 8884
rect 20523 8756 20565 8765
rect 20523 8716 20524 8756
rect 20564 8716 20565 8756
rect 20523 8707 20565 8716
rect 20331 8672 20373 8681
rect 20331 8632 20332 8672
rect 20372 8632 20373 8672
rect 20331 8623 20373 8632
rect 19372 8464 19796 8504
rect 19275 8420 19317 8429
rect 19275 8380 19276 8420
rect 19316 8380 19317 8420
rect 19275 8371 19317 8380
rect 18795 8000 18837 8009
rect 18795 7960 18796 8000
rect 18836 7960 18837 8000
rect 18795 7951 18837 7960
rect 19179 8000 19221 8009
rect 19179 7960 19180 8000
rect 19220 7960 19221 8000
rect 19179 7951 19221 7960
rect 18796 7866 18836 7951
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 19372 7160 19412 8464
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 20236 8000 20276 8009
rect 20332 8000 20372 8623
rect 20524 8009 20564 8707
rect 21004 8672 21044 8681
rect 20620 8504 20660 8513
rect 20620 8345 20660 8464
rect 20619 8336 20661 8345
rect 20619 8296 20620 8336
rect 20660 8296 20661 8336
rect 20619 8287 20661 8296
rect 20908 8168 20948 8177
rect 21004 8168 21044 8632
rect 20948 8128 21044 8168
rect 20908 8119 20948 8128
rect 19948 7960 20236 8000
rect 20276 7960 20372 8000
rect 20523 8000 20565 8009
rect 20523 7960 20524 8000
rect 20564 7960 20565 8000
rect 19948 7916 19988 7960
rect 20236 7951 20276 7960
rect 20523 7951 20565 7960
rect 21195 8000 21237 8009
rect 21195 7960 21196 8000
rect 21236 7960 21237 8000
rect 21195 7951 21237 7960
rect 21484 8000 21524 8009
rect 21676 8000 21716 8009
rect 21524 7960 21620 8000
rect 21484 7951 21524 7960
rect 19948 7867 19988 7876
rect 21196 7866 21236 7951
rect 21483 7748 21525 7757
rect 21483 7708 21484 7748
rect 21524 7708 21525 7748
rect 21483 7699 21525 7708
rect 21484 7614 21524 7699
rect 19372 7111 19412 7120
rect 20236 7160 20276 7169
rect 20276 7120 20468 7160
rect 20236 7111 20276 7120
rect 18988 7026 19028 7111
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 18123 6488 18165 6497
rect 18123 6448 18124 6488
rect 18164 6448 18165 6488
rect 18123 6439 18165 6448
rect 19371 6488 19413 6497
rect 19371 6448 19372 6488
rect 19412 6448 19413 6488
rect 19371 6439 19413 6448
rect 19563 6488 19605 6497
rect 19563 6448 19564 6488
rect 19604 6448 19605 6488
rect 19563 6439 19605 6448
rect 18412 6329 18452 6414
rect 18796 6404 18836 6413
rect 18124 6320 18164 6329
rect 18028 6280 18124 6320
rect 16875 6271 16917 6280
rect 18124 6271 18164 6280
rect 18411 6320 18453 6329
rect 18411 6280 18412 6320
rect 18452 6280 18453 6320
rect 18411 6271 18453 6280
rect 18123 6152 18165 6161
rect 18123 6112 18124 6152
rect 18164 6112 18165 6152
rect 18123 6103 18165 6112
rect 18124 5900 18164 6103
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18124 5860 18356 5900
rect 17452 5816 17492 5825
rect 17356 5776 17452 5816
rect 16588 4927 16628 4936
rect 16780 4976 16820 4985
rect 16396 4842 16436 4927
rect 16588 4808 16628 4817
rect 16780 4808 16820 4936
rect 16628 4768 16820 4808
rect 16588 4759 16628 4768
rect 16300 4684 16436 4724
rect 16299 4136 16341 4145
rect 16299 4096 16300 4136
rect 16340 4096 16341 4136
rect 16299 4087 16341 4096
rect 16300 3632 16340 4087
rect 16396 3632 16436 4684
rect 17356 4136 17396 5776
rect 17452 5767 17492 5776
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 17931 5599 17973 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18316 5648 18356 5860
rect 18316 5599 18356 5608
rect 17932 5514 17972 5599
rect 17739 5060 17781 5069
rect 17739 5020 17740 5060
rect 17780 5020 17781 5060
rect 17739 5011 17781 5020
rect 17740 4926 17780 5011
rect 17356 4087 17396 4096
rect 17452 4724 17492 4733
rect 16972 4052 17012 4061
rect 16780 3968 16820 3977
rect 16972 3968 17012 4012
rect 17452 3968 17492 4684
rect 18027 4724 18069 4733
rect 18027 4684 18028 4724
rect 18068 4684 18069 4724
rect 18027 4675 18069 4684
rect 16972 3928 17492 3968
rect 16396 3592 16532 3632
rect 16300 3583 16340 3592
rect 16204 3415 16244 3424
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 16299 3415 16341 3424
rect 16396 3464 16436 3473
rect 16107 3044 16149 3053
rect 16107 3004 16108 3044
rect 16148 3004 16149 3044
rect 16107 2995 16149 3004
rect 16011 2792 16053 2801
rect 16011 2752 16012 2792
rect 16052 2752 16053 2792
rect 16011 2743 16053 2752
rect 15916 2575 15956 2584
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 16108 2624 16148 2995
rect 16203 2792 16245 2801
rect 16203 2752 16204 2792
rect 16244 2752 16245 2792
rect 16203 2743 16245 2752
rect 16108 2575 16148 2584
rect 14764 2500 15092 2540
rect 15052 2036 15092 2500
rect 15052 1987 15092 1996
rect 13132 1903 13172 1912
rect 15436 1952 15476 1961
rect 16012 1952 16052 2575
rect 16204 2540 16244 2743
rect 16300 2717 16340 3415
rect 16396 3389 16436 3424
rect 16492 3464 16532 3592
rect 16587 3548 16629 3557
rect 16587 3508 16588 3548
rect 16628 3508 16629 3548
rect 16587 3499 16629 3508
rect 16780 3548 16820 3928
rect 16780 3499 16820 3508
rect 16492 3415 16532 3424
rect 16395 3380 16437 3389
rect 16395 3340 16396 3380
rect 16436 3340 16437 3380
rect 16395 3331 16437 3340
rect 16396 2885 16436 3331
rect 16491 3128 16533 3137
rect 16491 3088 16492 3128
rect 16532 3088 16533 3128
rect 16491 3079 16533 3088
rect 16395 2876 16437 2885
rect 16395 2836 16396 2876
rect 16436 2836 16437 2876
rect 16395 2827 16437 2836
rect 16299 2708 16341 2717
rect 16299 2668 16300 2708
rect 16340 2668 16341 2708
rect 16299 2659 16341 2668
rect 16300 2624 16340 2659
rect 16300 2574 16340 2584
rect 16492 2624 16532 3079
rect 16492 2575 16532 2584
rect 16204 2491 16244 2500
rect 16588 2540 16628 3499
rect 17164 3464 17204 3473
rect 18028 3464 18068 4675
rect 18124 4136 18164 5599
rect 18412 4976 18452 4985
rect 18412 4817 18452 4936
rect 18411 4808 18453 4817
rect 18411 4768 18412 4808
rect 18452 4768 18453 4808
rect 18411 4759 18453 4768
rect 18796 4724 18836 6364
rect 19179 5648 19221 5657
rect 19179 5608 19180 5648
rect 19220 5608 19221 5648
rect 19179 5599 19221 5608
rect 19180 5514 19220 5599
rect 19372 4976 19412 6439
rect 19564 6354 19604 6439
rect 20236 6236 20276 6245
rect 20236 5657 20276 6196
rect 20235 5648 20277 5657
rect 20235 5608 20236 5648
rect 20276 5608 20277 5648
rect 20235 5599 20277 5608
rect 20332 5648 20372 5657
rect 20332 5405 20372 5608
rect 20331 5396 20373 5405
rect 20331 5356 20332 5396
rect 20372 5356 20373 5396
rect 20331 5347 20373 5356
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 19468 4976 19508 4985
rect 19372 4936 19468 4976
rect 19468 4927 19508 4936
rect 19948 4976 19988 4985
rect 19371 4808 19413 4817
rect 19371 4768 19372 4808
rect 19412 4768 19413 4808
rect 19371 4759 19413 4768
rect 18891 4724 18933 4733
rect 18796 4684 18892 4724
rect 18932 4684 18933 4724
rect 18891 4675 18933 4684
rect 18892 4590 18932 4675
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 19372 4388 19412 4759
rect 19372 4339 19412 4348
rect 19756 4145 19796 4230
rect 18220 4136 18260 4145
rect 18124 4096 18220 4136
rect 18220 4087 18260 4096
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 19564 3977 19604 4062
rect 19851 4052 19893 4061
rect 19851 4012 19852 4052
rect 19892 4012 19893 4052
rect 19851 4003 19893 4012
rect 19563 3968 19605 3977
rect 19563 3928 19564 3968
rect 19604 3928 19605 3968
rect 19563 3919 19605 3928
rect 19852 3968 19892 4003
rect 19852 3917 19892 3928
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 19948 3716 19988 4936
rect 20428 4733 20468 7120
rect 21387 6992 21429 7001
rect 21387 6952 21388 6992
rect 21428 6952 21429 6992
rect 21387 6943 21429 6952
rect 21388 6858 21428 6943
rect 21580 6497 21620 7960
rect 21716 7960 21812 8000
rect 21676 7951 21716 7960
rect 21772 7001 21812 7960
rect 21771 6992 21813 7001
rect 21771 6952 21772 6992
rect 21812 6952 21813 6992
rect 21771 6943 21813 6952
rect 21868 6572 21908 10312
rect 21963 10184 22005 10193
rect 21963 10144 21964 10184
rect 22004 10144 22005 10184
rect 21963 10135 22005 10144
rect 21964 10050 22004 10135
rect 22060 8672 22100 10387
rect 23020 10193 23060 11647
rect 23116 11285 23156 15520
rect 23212 14141 23252 16183
rect 23596 15728 23636 16267
rect 23692 16241 23732 17032
rect 23691 16232 23733 16241
rect 23691 16192 23692 16232
rect 23732 16192 23733 16232
rect 23691 16183 23733 16192
rect 23691 15980 23733 15989
rect 23691 15940 23692 15980
rect 23732 15940 23733 15980
rect 23691 15931 23733 15940
rect 23596 15679 23636 15688
rect 23692 15560 23732 15931
rect 23788 15728 23828 17872
rect 23979 17863 24021 17872
rect 23884 17744 23924 17753
rect 23884 17408 23924 17704
rect 23980 17660 24020 17863
rect 23980 17611 24020 17620
rect 24076 17744 24116 17753
rect 24076 17585 24116 17704
rect 24172 17744 24212 17956
rect 24364 17947 24404 17956
rect 24267 17828 24309 17837
rect 24267 17788 24268 17828
rect 24308 17788 24309 17828
rect 24267 17779 24309 17788
rect 24172 17695 24212 17704
rect 24075 17576 24117 17585
rect 24075 17536 24076 17576
rect 24116 17536 24117 17576
rect 24075 17527 24117 17536
rect 23884 17368 24212 17408
rect 24075 17240 24117 17249
rect 24075 17200 24076 17240
rect 24116 17200 24117 17240
rect 24075 17191 24117 17200
rect 24172 17240 24212 17368
rect 24172 17191 24212 17200
rect 23883 17072 23925 17081
rect 23883 17032 23884 17072
rect 23924 17032 23925 17072
rect 23883 17023 23925 17032
rect 23980 17072 24020 17081
rect 23884 16938 23924 17023
rect 23980 16997 24020 17032
rect 24076 17072 24116 17191
rect 24268 17072 24308 17779
rect 24364 17744 24404 17755
rect 24364 17669 24404 17704
rect 24460 17744 24500 18292
rect 24748 18283 24788 18292
rect 24844 18164 24884 18964
rect 25324 18920 25364 19804
rect 25516 19601 25556 21391
rect 25708 20852 25748 21475
rect 25804 21474 25844 21559
rect 25708 20180 25748 20812
rect 25612 20140 25748 20180
rect 25515 19592 25557 19601
rect 25515 19552 25516 19592
rect 25556 19552 25557 19592
rect 25515 19543 25557 19552
rect 25612 19424 25652 20140
rect 25804 20096 25844 20105
rect 25708 20056 25804 20096
rect 25708 19937 25748 20056
rect 25804 20047 25844 20056
rect 25707 19928 25749 19937
rect 25707 19888 25708 19928
rect 25748 19888 25749 19928
rect 25707 19879 25749 19888
rect 25132 18880 25364 18920
rect 25516 19384 25652 19424
rect 25132 18584 25172 18880
rect 25516 18593 25556 19384
rect 25612 19256 25652 19265
rect 25708 19256 25748 19879
rect 25652 19216 25748 19256
rect 25804 19256 25844 19265
rect 25900 19256 25940 21895
rect 26092 21608 26132 22072
rect 26572 22112 26612 22121
rect 26572 21617 26612 22072
rect 26092 21559 26132 21568
rect 26571 21608 26613 21617
rect 26571 21568 26572 21608
rect 26612 21568 26613 21608
rect 26571 21559 26613 21568
rect 26379 21440 26421 21449
rect 26379 21400 26380 21440
rect 26420 21400 26421 21440
rect 26379 21391 26421 21400
rect 26091 20348 26133 20357
rect 26091 20308 26092 20348
rect 26132 20308 26133 20348
rect 26091 20299 26133 20308
rect 26092 20096 26132 20299
rect 26283 20264 26325 20273
rect 26283 20224 26284 20264
rect 26324 20224 26325 20264
rect 26283 20215 26325 20224
rect 26284 20096 26324 20215
rect 26380 20189 26420 21391
rect 26572 20768 26612 20777
rect 26956 20768 26996 25843
rect 27148 23960 27188 27355
rect 27916 27068 27956 27077
rect 28012 27068 28052 27439
rect 27956 27028 28052 27068
rect 27916 27019 27956 27028
rect 27340 26816 27380 26825
rect 27340 26573 27380 26776
rect 28300 26732 28340 28120
rect 28491 28160 28533 28169
rect 28491 28120 28492 28160
rect 28532 28120 28533 28160
rect 28491 28111 28533 28120
rect 28683 28160 28725 28169
rect 28683 28120 28684 28160
rect 28724 28120 28725 28160
rect 28683 28111 28725 28120
rect 28684 28001 28724 28111
rect 28972 28110 29012 28195
rect 28683 27992 28725 28001
rect 28683 27952 28684 27992
rect 28724 27952 28725 27992
rect 28683 27943 28725 27952
rect 28491 27656 28533 27665
rect 28491 27616 28492 27656
rect 28532 27616 28533 27656
rect 28491 27607 28533 27616
rect 29067 27656 29109 27665
rect 29067 27616 29068 27656
rect 29108 27616 29109 27656
rect 29067 27607 29109 27616
rect 29164 27656 29204 28288
rect 29259 27656 29301 27665
rect 29164 27616 29260 27656
rect 29300 27616 29301 27656
rect 28492 27522 28532 27607
rect 28587 27572 28629 27581
rect 28587 27532 28588 27572
rect 28628 27532 28629 27572
rect 28587 27523 28629 27532
rect 28588 27438 28628 27523
rect 29068 27522 29108 27607
rect 28683 27488 28725 27497
rect 28683 27448 28684 27488
rect 28724 27448 28725 27488
rect 28683 27439 28725 27448
rect 28491 27404 28533 27413
rect 28491 27364 28492 27404
rect 28532 27364 28533 27404
rect 28491 27355 28533 27364
rect 28012 26692 28340 26732
rect 27339 26564 27381 26573
rect 27339 26524 27340 26564
rect 27380 26524 27381 26564
rect 27339 26515 27381 26524
rect 27627 26228 27669 26237
rect 27627 26188 27628 26228
rect 27668 26188 27669 26228
rect 27627 26179 27669 26188
rect 27532 26144 27572 26153
rect 27243 25892 27285 25901
rect 27243 25852 27244 25892
rect 27284 25852 27285 25892
rect 27243 25843 27285 25852
rect 27244 25758 27284 25843
rect 27532 25817 27572 26104
rect 27628 26139 27668 26179
rect 27628 26090 27668 26099
rect 27723 26144 27765 26153
rect 27723 26104 27724 26144
rect 27764 26104 27765 26144
rect 27723 26095 27765 26104
rect 27724 26010 27764 26095
rect 27531 25808 27573 25817
rect 27531 25768 27532 25808
rect 27572 25768 27573 25808
rect 27531 25759 27573 25768
rect 27531 25472 27573 25481
rect 27531 25432 27532 25472
rect 27572 25432 27573 25472
rect 27531 25423 27573 25432
rect 27532 25338 27572 25423
rect 27916 25304 27956 25313
rect 27628 25264 27916 25304
rect 27628 24464 27668 25264
rect 27916 25255 27956 25264
rect 27915 24632 27957 24641
rect 27915 24592 27916 24632
rect 27956 24592 27957 24632
rect 27915 24583 27957 24592
rect 28012 24632 28052 26692
rect 28395 26480 28437 26489
rect 28395 26440 28396 26480
rect 28436 26440 28437 26480
rect 28395 26431 28437 26440
rect 28299 26144 28341 26153
rect 28299 26104 28300 26144
rect 28340 26104 28341 26144
rect 28299 26095 28341 26104
rect 28396 26144 28436 26431
rect 28204 25472 28244 25481
rect 28107 24884 28149 24893
rect 28107 24835 28108 24884
rect 28148 24835 28149 24884
rect 28108 24749 28148 24818
rect 28012 24583 28052 24592
rect 27916 24498 27956 24583
rect 27628 24415 27668 24424
rect 27052 23920 27188 23960
rect 27052 23120 27092 23920
rect 27243 23876 27285 23885
rect 27243 23836 27244 23876
rect 27284 23836 27285 23876
rect 27243 23827 27285 23836
rect 27531 23876 27573 23885
rect 27531 23836 27532 23876
rect 27572 23836 27573 23876
rect 27531 23827 27573 23836
rect 27723 23876 27765 23885
rect 27723 23836 27724 23876
rect 27764 23836 27765 23876
rect 27723 23827 27765 23836
rect 27148 23792 27188 23803
rect 27148 23717 27188 23752
rect 27244 23792 27284 23827
rect 27244 23741 27284 23752
rect 27436 23792 27476 23801
rect 27147 23708 27189 23717
rect 27147 23668 27148 23708
rect 27188 23668 27189 23708
rect 27147 23659 27189 23668
rect 27339 23624 27381 23633
rect 27339 23584 27340 23624
rect 27380 23584 27381 23624
rect 27339 23575 27381 23584
rect 27340 23490 27380 23575
rect 27243 23372 27285 23381
rect 27243 23332 27244 23372
rect 27284 23332 27285 23372
rect 27243 23323 27285 23332
rect 27244 23120 27284 23323
rect 27436 23297 27476 23752
rect 27532 23465 27572 23827
rect 27627 23792 27669 23801
rect 27627 23752 27628 23792
rect 27668 23752 27669 23792
rect 27627 23743 27669 23752
rect 27628 23658 27668 23743
rect 27724 23742 27764 23827
rect 27820 23792 27860 23801
rect 27915 23792 27957 23801
rect 27860 23752 27916 23792
rect 27956 23752 27957 23792
rect 27820 23743 27860 23752
rect 27915 23743 27957 23752
rect 28108 23792 28148 23801
rect 27723 23624 27765 23633
rect 27723 23584 27724 23624
rect 27764 23584 27765 23624
rect 27723 23575 27765 23584
rect 27531 23456 27573 23465
rect 27531 23416 27532 23456
rect 27572 23416 27573 23456
rect 27531 23407 27573 23416
rect 27435 23288 27477 23297
rect 27435 23248 27436 23288
rect 27476 23248 27477 23288
rect 27435 23239 27477 23248
rect 27092 23080 27188 23120
rect 27052 23071 27092 23080
rect 27052 22877 27092 22962
rect 27051 22868 27093 22877
rect 27051 22828 27052 22868
rect 27092 22828 27093 22868
rect 27051 22819 27093 22828
rect 27051 22196 27093 22205
rect 27051 22156 27052 22196
rect 27092 22156 27093 22196
rect 27051 22147 27093 22156
rect 26612 20728 26956 20768
rect 26572 20719 26612 20728
rect 26956 20719 26996 20728
rect 27052 21608 27092 22147
rect 27052 20600 27092 21568
rect 26860 20560 27092 20600
rect 26668 20273 26708 20275
rect 26667 20264 26709 20273
rect 26667 20224 26668 20264
rect 26708 20224 26709 20264
rect 26667 20215 26709 20224
rect 26379 20180 26421 20189
rect 26379 20140 26380 20180
rect 26420 20140 26421 20180
rect 26379 20131 26421 20140
rect 26668 20180 26708 20215
rect 26860 20180 26900 20560
rect 27148 20357 27188 23080
rect 27244 23071 27284 23080
rect 27340 23120 27380 23129
rect 27243 22280 27285 22289
rect 27243 22240 27244 22280
rect 27284 22240 27285 22280
rect 27243 22231 27285 22240
rect 27244 22146 27284 22231
rect 27340 21776 27380 23080
rect 27724 23120 27764 23575
rect 27819 23456 27861 23465
rect 27819 23416 27820 23456
rect 27860 23416 27861 23456
rect 27819 23407 27861 23416
rect 27724 22793 27764 23080
rect 27820 23120 27860 23407
rect 27820 23071 27860 23080
rect 27723 22784 27765 22793
rect 27723 22744 27724 22784
rect 27764 22744 27765 22784
rect 27723 22735 27765 22744
rect 27531 22616 27573 22625
rect 27531 22576 27532 22616
rect 27572 22576 27573 22616
rect 27531 22567 27573 22576
rect 27436 22280 27476 22289
rect 27436 21785 27476 22240
rect 27340 21727 27380 21736
rect 27435 21776 27477 21785
rect 27435 21736 27436 21776
rect 27476 21736 27477 21776
rect 27435 21727 27477 21736
rect 27532 21608 27572 22567
rect 27916 22205 27956 23743
rect 28012 23624 28052 23633
rect 28012 23036 28052 23584
rect 28108 23213 28148 23752
rect 28204 23717 28244 25432
rect 28300 24800 28340 26095
rect 28396 26069 28436 26104
rect 28395 26060 28437 26069
rect 28395 26020 28396 26060
rect 28436 26020 28437 26060
rect 28395 26011 28437 26020
rect 28396 24800 28436 24809
rect 28300 24760 28396 24800
rect 28396 24751 28436 24760
rect 28300 24632 28340 24641
rect 28300 24137 28340 24592
rect 28492 24632 28532 27355
rect 28684 26732 28724 27439
rect 29164 27413 29204 27616
rect 29259 27607 29301 27616
rect 29547 27656 29589 27665
rect 29547 27611 29548 27656
rect 29588 27611 29589 27656
rect 29547 27607 29589 27611
rect 29548 27521 29588 27607
rect 29163 27404 29205 27413
rect 29163 27364 29164 27404
rect 29204 27364 29205 27404
rect 29163 27355 29205 27364
rect 29644 27320 29684 28447
rect 29739 27740 29781 27749
rect 29739 27700 29740 27740
rect 29780 27700 29781 27740
rect 29739 27691 29781 27700
rect 29740 27606 29780 27691
rect 29644 27280 29780 27320
rect 28779 27068 28821 27077
rect 28779 27028 28780 27068
rect 28820 27028 28821 27068
rect 28779 27019 28821 27028
rect 28588 26692 28724 26732
rect 28780 26816 28820 27019
rect 29643 26984 29685 26993
rect 29643 26944 29644 26984
rect 29684 26944 29685 26984
rect 29643 26935 29685 26944
rect 28588 24800 28628 26692
rect 28588 24760 28724 24800
rect 28492 24583 28532 24592
rect 28587 24632 28629 24641
rect 28587 24592 28588 24632
rect 28628 24592 28629 24632
rect 28587 24583 28629 24592
rect 28588 24498 28628 24583
rect 28684 24380 28724 24760
rect 28588 24340 28724 24380
rect 28299 24128 28341 24137
rect 28299 24088 28300 24128
rect 28340 24088 28341 24128
rect 28299 24079 28341 24088
rect 28492 23801 28532 23886
rect 28491 23792 28533 23801
rect 28491 23752 28492 23792
rect 28532 23752 28533 23792
rect 28491 23743 28533 23752
rect 28588 23792 28628 24340
rect 28780 23960 28820 26776
rect 28971 26816 29013 26825
rect 28971 26776 28972 26816
rect 29012 26776 29013 26816
rect 28971 26767 29013 26776
rect 29068 26816 29108 26825
rect 29452 26816 29492 26825
rect 29108 26776 29300 26816
rect 29068 26767 29108 26776
rect 28972 26682 29012 26767
rect 28876 26648 28916 26657
rect 28876 24893 28916 26608
rect 29067 26564 29109 26573
rect 29067 26524 29068 26564
rect 29108 26524 29109 26564
rect 29067 26515 29109 26524
rect 29068 25976 29108 26515
rect 29260 26312 29300 26776
rect 29452 26489 29492 26776
rect 29547 26816 29589 26825
rect 29547 26776 29548 26816
rect 29588 26776 29589 26816
rect 29547 26767 29589 26776
rect 29644 26816 29684 26935
rect 29644 26767 29684 26776
rect 29548 26682 29588 26767
rect 29451 26480 29493 26489
rect 29451 26440 29452 26480
rect 29492 26440 29493 26480
rect 29451 26431 29493 26440
rect 29740 26321 29780 27280
rect 30028 26648 30068 26657
rect 29644 26312 29684 26321
rect 29260 26272 29644 26312
rect 29644 26263 29684 26272
rect 29739 26312 29781 26321
rect 29739 26272 29740 26312
rect 29780 26272 29781 26312
rect 29739 26263 29781 26272
rect 29068 25927 29108 25936
rect 29356 26144 29396 26153
rect 29356 25481 29396 26104
rect 29548 26144 29588 26153
rect 29548 25565 29588 26104
rect 29740 26144 29780 26263
rect 29740 26095 29780 26104
rect 29835 26144 29877 26153
rect 29835 26104 29836 26144
rect 29876 26104 29877 26144
rect 29835 26095 29877 26104
rect 29836 26010 29876 26095
rect 29547 25556 29589 25565
rect 29547 25516 29548 25556
rect 29588 25516 29589 25556
rect 29547 25507 29589 25516
rect 29355 25472 29397 25481
rect 29355 25432 29356 25472
rect 29396 25432 29397 25472
rect 29355 25423 29397 25432
rect 29836 25472 29876 25481
rect 28875 24884 28917 24893
rect 28875 24844 28876 24884
rect 28916 24844 28917 24884
rect 28875 24835 28917 24844
rect 29356 24632 29396 24641
rect 29356 24044 29396 24592
rect 29740 24632 29780 24641
rect 29836 24632 29876 25432
rect 29780 24592 29876 24632
rect 29740 24583 29780 24592
rect 29452 24044 29492 24053
rect 29356 24004 29452 24044
rect 29452 23995 29492 24004
rect 28875 23960 28917 23969
rect 30028 23960 30068 26608
rect 30220 25481 30260 28960
rect 30412 28916 30452 28925
rect 30412 28337 30452 28876
rect 30411 28328 30453 28337
rect 30411 28288 30412 28328
rect 30452 28288 30453 28328
rect 30411 28279 30453 28288
rect 30508 28160 30548 32152
rect 30604 30941 30644 32992
rect 30796 32957 30836 34168
rect 30891 33452 30933 33461
rect 30891 33412 30892 33452
rect 30932 33412 30933 33452
rect 30891 33403 30933 33412
rect 30795 32948 30837 32957
rect 30700 32908 30796 32948
rect 30836 32908 30837 32948
rect 30603 30932 30645 30941
rect 30603 30892 30604 30932
rect 30644 30892 30645 30932
rect 30603 30883 30645 30892
rect 30603 30764 30645 30773
rect 30603 30724 30604 30764
rect 30644 30724 30645 30764
rect 30603 30715 30645 30724
rect 30604 30680 30644 30715
rect 30700 30680 30740 32908
rect 30795 32899 30837 32908
rect 30892 32864 30932 33403
rect 30892 32815 30932 32824
rect 30796 32696 30836 32705
rect 30796 32024 30836 32656
rect 30988 32612 31028 34243
rect 31084 33629 31124 36016
rect 31372 35300 31412 36511
rect 31372 35251 31412 35260
rect 31468 36476 31508 36485
rect 31276 35216 31316 35225
rect 31276 35057 31316 35176
rect 31468 35141 31508 36436
rect 32044 36140 32084 36149
rect 32140 36140 32180 36688
rect 32332 36679 32372 36688
rect 32428 36688 32620 36728
rect 32084 36100 32180 36140
rect 32236 36140 32276 36149
rect 32428 36140 32468 36688
rect 32620 36679 32660 36688
rect 32276 36100 32468 36140
rect 32044 36091 32084 36100
rect 32236 36091 32276 36100
rect 32236 35888 32276 35897
rect 32043 35720 32085 35729
rect 32043 35680 32044 35720
rect 32084 35680 32085 35720
rect 32043 35671 32085 35680
rect 32044 35586 32084 35671
rect 32236 35225 32276 35848
rect 32428 35888 32468 35897
rect 31948 35216 31988 35225
rect 31467 35132 31509 35141
rect 31467 35092 31468 35132
rect 31508 35092 31509 35132
rect 31467 35083 31509 35092
rect 31275 35048 31317 35057
rect 31275 35008 31276 35048
rect 31316 35008 31317 35048
rect 31275 34999 31317 35008
rect 31660 34964 31700 34973
rect 31660 34721 31700 34924
rect 31659 34712 31701 34721
rect 31659 34672 31660 34712
rect 31700 34672 31701 34712
rect 31659 34663 31701 34672
rect 31755 34628 31797 34637
rect 31755 34588 31756 34628
rect 31796 34588 31797 34628
rect 31755 34579 31797 34588
rect 31275 34460 31317 34469
rect 31275 34420 31276 34460
rect 31316 34420 31317 34460
rect 31275 34411 31317 34420
rect 31276 34376 31316 34411
rect 31660 34376 31700 34385
rect 31276 34325 31316 34336
rect 31564 34336 31660 34376
rect 31083 33620 31125 33629
rect 31083 33580 31084 33620
rect 31124 33580 31125 33620
rect 31083 33571 31125 33580
rect 31275 33452 31317 33461
rect 31468 33452 31508 33461
rect 31275 33412 31276 33452
rect 31316 33412 31317 33452
rect 31275 33403 31317 33412
rect 31372 33412 31468 33452
rect 31276 33318 31316 33403
rect 31084 32864 31124 32873
rect 31372 32864 31412 33412
rect 31468 33403 31508 33412
rect 31467 33284 31509 33293
rect 31467 33244 31468 33284
rect 31508 33244 31509 33284
rect 31467 33235 31509 33244
rect 31124 32824 31412 32864
rect 31468 32864 31508 33235
rect 31084 32815 31124 32824
rect 31468 32815 31508 32824
rect 30892 32572 31028 32612
rect 30892 32192 30932 32572
rect 30892 32143 30932 32152
rect 31180 32192 31220 32201
rect 31180 32024 31220 32152
rect 30796 31984 31220 32024
rect 31180 31361 31220 31984
rect 31276 32192 31316 32201
rect 31179 31352 31221 31361
rect 31179 31312 31180 31352
rect 31220 31312 31221 31352
rect 31179 31303 31221 31312
rect 30891 31184 30933 31193
rect 30891 31144 30892 31184
rect 30932 31144 30933 31184
rect 30891 31135 30933 31144
rect 30796 30680 30836 30689
rect 30700 30640 30796 30680
rect 30604 30629 30644 30640
rect 30796 30631 30836 30640
rect 30892 30680 30932 31135
rect 31276 31025 31316 32152
rect 31564 32108 31604 34336
rect 31660 34327 31700 34336
rect 31756 34376 31796 34579
rect 31948 34553 31988 35176
rect 32235 35216 32277 35225
rect 32235 35176 32236 35216
rect 32276 35176 32277 35216
rect 32235 35167 32277 35176
rect 32235 34964 32277 34973
rect 32235 34924 32236 34964
rect 32276 34924 32372 34964
rect 32235 34915 32277 34924
rect 32236 34830 32276 34915
rect 32139 34712 32181 34721
rect 32139 34672 32140 34712
rect 32180 34672 32181 34712
rect 32139 34663 32181 34672
rect 31947 34544 31989 34553
rect 31947 34504 31948 34544
rect 31988 34504 31989 34544
rect 31947 34495 31989 34504
rect 31756 34327 31796 34336
rect 31948 34376 31988 34385
rect 31852 34208 31892 34217
rect 31755 33956 31797 33965
rect 31755 33916 31756 33956
rect 31796 33916 31797 33956
rect 31755 33907 31797 33916
rect 31756 32192 31796 33907
rect 31852 33713 31892 34168
rect 31851 33704 31893 33713
rect 31851 33664 31852 33704
rect 31892 33664 31893 33704
rect 31851 33655 31893 33664
rect 31852 32360 31892 32369
rect 31948 32360 31988 34336
rect 32140 33872 32180 34663
rect 32236 34385 32276 34470
rect 32235 34376 32277 34385
rect 32235 34336 32236 34376
rect 32276 34336 32277 34376
rect 32235 34327 32277 34336
rect 32140 33832 32276 33872
rect 32139 33704 32181 33713
rect 32139 33664 32140 33704
rect 32180 33664 32181 33704
rect 32139 33655 32181 33664
rect 32140 33570 32180 33655
rect 31892 32320 31988 32360
rect 31852 32311 31892 32320
rect 31948 32192 31988 32201
rect 31756 32152 31948 32192
rect 31468 32068 31604 32108
rect 31371 31184 31413 31193
rect 31371 31144 31372 31184
rect 31412 31144 31413 31184
rect 31371 31135 31413 31144
rect 31372 31050 31412 31135
rect 31275 31016 31317 31025
rect 31275 30976 31276 31016
rect 31316 30976 31317 31016
rect 31275 30967 31317 30976
rect 30987 30932 31029 30941
rect 30987 30892 30988 30932
rect 31028 30892 31029 30932
rect 30987 30883 31029 30892
rect 30892 30631 30932 30640
rect 30988 30680 31028 30883
rect 31083 30848 31125 30857
rect 31083 30808 31084 30848
rect 31124 30808 31125 30848
rect 31083 30799 31125 30808
rect 31276 30848 31316 30857
rect 31468 30848 31508 32068
rect 31564 31940 31604 31949
rect 31604 31900 31892 31940
rect 31564 31891 31604 31900
rect 31564 31352 31604 31361
rect 31564 31193 31604 31312
rect 31563 31184 31605 31193
rect 31755 31184 31797 31193
rect 31563 31144 31564 31184
rect 31604 31144 31605 31184
rect 31563 31135 31605 31144
rect 31660 31144 31756 31184
rect 31796 31144 31797 31184
rect 31563 31016 31605 31025
rect 31563 30976 31564 31016
rect 31604 30976 31605 31016
rect 31563 30967 31605 30976
rect 31316 30808 31508 30848
rect 31564 30848 31604 30967
rect 31276 30799 31316 30808
rect 31564 30799 31604 30808
rect 31084 30714 31124 30799
rect 31179 30764 31221 30773
rect 31179 30724 31180 30764
rect 31220 30724 31221 30764
rect 31179 30715 31221 30724
rect 30891 30512 30933 30521
rect 30891 30472 30892 30512
rect 30932 30472 30933 30512
rect 30891 30463 30933 30472
rect 30699 29336 30741 29345
rect 30699 29296 30700 29336
rect 30740 29296 30741 29336
rect 30699 29287 30741 29296
rect 30603 29168 30645 29177
rect 30603 29128 30604 29168
rect 30644 29128 30645 29168
rect 30603 29119 30645 29128
rect 30700 29168 30740 29287
rect 30700 29119 30740 29128
rect 30796 29168 30836 29177
rect 30604 29034 30644 29119
rect 30699 29000 30741 29009
rect 30699 28960 30700 29000
rect 30740 28960 30741 29000
rect 30699 28951 30741 28960
rect 30603 28916 30645 28925
rect 30603 28876 30604 28916
rect 30644 28876 30645 28916
rect 30603 28867 30645 28876
rect 30604 28328 30644 28867
rect 30604 28279 30644 28288
rect 30700 28328 30740 28951
rect 30796 28505 30836 29128
rect 30892 29168 30932 30463
rect 30988 30008 31028 30640
rect 31180 30092 31220 30715
rect 31372 30680 31412 30689
rect 31372 30521 31412 30640
rect 31660 30680 31700 31144
rect 31755 31135 31797 31144
rect 31660 30631 31700 30640
rect 31371 30512 31413 30521
rect 31371 30472 31372 30512
rect 31412 30472 31413 30512
rect 31371 30463 31413 30472
rect 31276 30092 31316 30101
rect 31180 30052 31276 30092
rect 31276 30043 31316 30052
rect 30988 29968 31220 30008
rect 30987 29840 31029 29849
rect 30987 29800 30988 29840
rect 31028 29800 31029 29840
rect 30987 29791 31029 29800
rect 30892 29119 30932 29128
rect 30988 29009 31028 29791
rect 31083 29168 31125 29177
rect 31083 29128 31084 29168
rect 31124 29128 31125 29168
rect 31083 29119 31125 29128
rect 31084 29034 31124 29119
rect 30987 29000 31029 29009
rect 30987 28960 30988 29000
rect 31028 28960 31029 29000
rect 30987 28951 31029 28960
rect 31083 28580 31125 28589
rect 31083 28540 31084 28580
rect 31124 28540 31125 28580
rect 31083 28531 31125 28540
rect 30795 28496 30837 28505
rect 30795 28456 30796 28496
rect 30836 28456 30837 28496
rect 30795 28447 30837 28456
rect 31084 28446 31124 28531
rect 30700 28279 30740 28288
rect 30796 28328 30836 28337
rect 30508 28120 30644 28160
rect 30316 27784 30548 27824
rect 30316 27077 30356 27784
rect 30411 27656 30453 27665
rect 30411 27616 30412 27656
rect 30452 27616 30453 27656
rect 30411 27607 30453 27616
rect 30508 27656 30548 27784
rect 30508 27607 30548 27616
rect 30315 27068 30357 27077
rect 30315 27028 30316 27068
rect 30356 27028 30357 27068
rect 30315 27019 30357 27028
rect 30315 26900 30357 26909
rect 30315 26860 30316 26900
rect 30356 26860 30357 26900
rect 30315 26851 30357 26860
rect 30412 26851 30452 27607
rect 30316 26816 30356 26851
rect 30412 26802 30452 26811
rect 30508 27404 30548 27413
rect 30508 26816 30548 27364
rect 30316 26765 30356 26776
rect 30508 26767 30548 26776
rect 30604 26648 30644 28120
rect 30796 27824 30836 28288
rect 30891 28328 30933 28337
rect 30891 28288 30892 28328
rect 30932 28288 30933 28328
rect 30891 28279 30933 28288
rect 30892 28194 30932 28279
rect 31180 27917 31220 29968
rect 31468 29840 31508 29849
rect 31371 28496 31413 28505
rect 31371 28456 31372 28496
rect 31412 28456 31413 28496
rect 31371 28447 31413 28456
rect 31179 27908 31221 27917
rect 31179 27868 31180 27908
rect 31220 27868 31221 27908
rect 31179 27859 31221 27868
rect 31275 27824 31317 27833
rect 30796 27784 30932 27824
rect 30700 27749 30740 27780
rect 30699 27740 30741 27749
rect 30699 27700 30700 27740
rect 30740 27700 30741 27740
rect 30699 27691 30741 27700
rect 30700 27656 30740 27691
rect 30700 27077 30740 27616
rect 30796 27656 30836 27665
rect 30796 27329 30836 27616
rect 30795 27320 30837 27329
rect 30795 27280 30796 27320
rect 30836 27280 30837 27320
rect 30795 27271 30837 27280
rect 30699 27068 30741 27077
rect 30699 27028 30700 27068
rect 30740 27028 30741 27068
rect 30699 27019 30741 27028
rect 30892 26984 30932 27784
rect 31275 27784 31276 27824
rect 31316 27784 31317 27824
rect 31275 27775 31317 27784
rect 30987 27740 31029 27749
rect 30987 27700 30988 27740
rect 31028 27700 31029 27740
rect 30987 27691 31029 27700
rect 30988 27656 31028 27691
rect 30988 27605 31028 27616
rect 31180 27656 31220 27665
rect 31180 27488 31220 27616
rect 31276 27656 31316 27775
rect 31276 27607 31316 27616
rect 31275 27488 31317 27497
rect 31180 27448 31276 27488
rect 31316 27448 31317 27488
rect 31275 27439 31317 27448
rect 30988 27404 31028 27413
rect 30988 27320 31028 27364
rect 30988 27280 31220 27320
rect 30987 27068 31029 27077
rect 30987 27028 30988 27068
rect 31028 27028 31029 27068
rect 30987 27019 31029 27028
rect 30796 26944 30932 26984
rect 30699 26816 30741 26825
rect 30699 26776 30700 26816
rect 30740 26776 30741 26816
rect 30699 26767 30741 26776
rect 30700 26657 30740 26767
rect 30508 26608 30644 26648
rect 30699 26648 30741 26657
rect 30699 26608 30700 26648
rect 30740 26608 30741 26648
rect 30219 25472 30261 25481
rect 30219 25432 30220 25472
rect 30260 25432 30261 25472
rect 30219 25423 30261 25432
rect 28780 23920 28876 23960
rect 28916 23920 28917 23960
rect 28875 23911 28917 23920
rect 29932 23920 30068 23960
rect 28203 23708 28245 23717
rect 28203 23668 28204 23708
rect 28244 23668 28245 23708
rect 28203 23659 28245 23668
rect 28300 23624 28340 23633
rect 28340 23584 28532 23624
rect 28300 23575 28340 23584
rect 28299 23288 28341 23297
rect 28299 23248 28300 23288
rect 28340 23248 28341 23288
rect 28299 23239 28341 23248
rect 28107 23204 28149 23213
rect 28107 23164 28108 23204
rect 28148 23164 28149 23204
rect 28107 23155 28149 23164
rect 28300 23120 28340 23239
rect 28300 23071 28340 23080
rect 28492 23120 28532 23584
rect 28588 23465 28628 23752
rect 28684 23792 28724 23801
rect 28587 23456 28629 23465
rect 28587 23416 28588 23456
rect 28628 23416 28629 23456
rect 28587 23407 28629 23416
rect 28492 23071 28532 23080
rect 28588 23120 28628 23129
rect 28107 23036 28149 23045
rect 28012 22996 28108 23036
rect 28148 22996 28149 23036
rect 28107 22987 28149 22996
rect 28108 22902 28148 22987
rect 28588 22877 28628 23080
rect 28684 23045 28724 23752
rect 28779 23792 28821 23801
rect 28779 23752 28780 23792
rect 28820 23752 28821 23792
rect 28779 23743 28821 23752
rect 28780 23658 28820 23743
rect 28779 23288 28821 23297
rect 28779 23248 28780 23288
rect 28820 23248 28821 23288
rect 28779 23239 28821 23248
rect 28780 23154 28820 23239
rect 28683 23036 28725 23045
rect 28683 22996 28684 23036
rect 28724 22996 28725 23036
rect 28683 22987 28725 22996
rect 28876 22961 28916 23911
rect 28971 23876 29013 23885
rect 29163 23876 29205 23885
rect 28971 23836 28972 23876
rect 29012 23836 29108 23876
rect 28971 23827 29013 23836
rect 29068 23792 29108 23836
rect 29163 23836 29164 23876
rect 29204 23836 29205 23876
rect 29163 23827 29205 23836
rect 29068 23743 29108 23752
rect 29164 23792 29204 23827
rect 29452 23801 29492 23886
rect 29164 23741 29204 23752
rect 29260 23792 29300 23801
rect 28971 23624 29013 23633
rect 28971 23584 28972 23624
rect 29012 23584 29013 23624
rect 28971 23575 29013 23584
rect 28972 23490 29012 23575
rect 29260 23465 29300 23752
rect 29451 23792 29493 23801
rect 29644 23792 29684 23801
rect 29451 23752 29452 23792
rect 29492 23752 29493 23792
rect 29451 23743 29493 23752
rect 29548 23752 29644 23792
rect 29451 23624 29493 23633
rect 29548 23624 29588 23752
rect 29644 23743 29684 23752
rect 29740 23792 29780 23801
rect 29451 23584 29452 23624
rect 29492 23584 29588 23624
rect 29451 23575 29493 23584
rect 29259 23456 29301 23465
rect 29259 23416 29260 23456
rect 29300 23416 29301 23456
rect 29259 23407 29301 23416
rect 29451 23456 29493 23465
rect 29451 23416 29452 23456
rect 29492 23416 29493 23456
rect 29451 23407 29493 23416
rect 29067 23372 29109 23381
rect 29067 23332 29068 23372
rect 29108 23332 29109 23372
rect 29067 23323 29109 23332
rect 29068 23288 29108 23323
rect 29068 23237 29108 23248
rect 29163 23204 29205 23213
rect 29163 23164 29164 23204
rect 29204 23164 29205 23204
rect 29163 23155 29205 23164
rect 28971 23120 29013 23129
rect 28971 23080 28972 23120
rect 29012 23080 29013 23120
rect 28971 23071 29013 23080
rect 29164 23120 29204 23155
rect 28972 22986 29012 23071
rect 29164 23069 29204 23080
rect 29452 23120 29492 23407
rect 29740 23297 29780 23752
rect 29739 23288 29781 23297
rect 29739 23248 29740 23288
rect 29780 23248 29781 23288
rect 29739 23239 29781 23248
rect 29547 23204 29589 23213
rect 29547 23164 29548 23204
rect 29588 23164 29589 23204
rect 29547 23155 29589 23164
rect 29452 23071 29492 23080
rect 29548 23070 29588 23155
rect 29644 23120 29684 23129
rect 29932 23120 29972 23920
rect 29684 23080 29972 23120
rect 30123 23120 30165 23129
rect 30123 23080 30124 23120
rect 30164 23080 30165 23120
rect 28875 22952 28917 22961
rect 28875 22912 28876 22952
rect 28916 22912 28917 22952
rect 28875 22903 28917 22912
rect 28587 22868 28629 22877
rect 28587 22828 28588 22868
rect 28628 22828 28724 22868
rect 28587 22819 28629 22828
rect 28588 22373 28628 22404
rect 28587 22364 28629 22373
rect 28587 22324 28588 22364
rect 28628 22324 28629 22364
rect 28587 22315 28629 22324
rect 28588 22280 28628 22315
rect 27915 22196 27957 22205
rect 27915 22156 27916 22196
rect 27956 22156 27957 22196
rect 27915 22147 27957 22156
rect 28108 22112 28148 22121
rect 28108 21692 28148 22072
rect 28588 21953 28628 22240
rect 28684 22280 28724 22828
rect 29163 22364 29205 22373
rect 29163 22324 29164 22364
rect 29204 22324 29205 22364
rect 29163 22315 29205 22324
rect 28684 22231 28724 22240
rect 28780 22280 28820 22291
rect 28780 22205 28820 22240
rect 28875 22280 28917 22289
rect 28875 22240 28876 22280
rect 28916 22240 28917 22280
rect 28875 22231 28917 22240
rect 28779 22196 28821 22205
rect 28779 22156 28780 22196
rect 28820 22156 28821 22196
rect 28779 22147 28821 22156
rect 28876 22146 28916 22231
rect 29164 22230 29204 22315
rect 29644 22280 29684 23080
rect 30123 23071 30165 23080
rect 30411 23120 30453 23129
rect 30411 23080 30412 23120
rect 30452 23080 30453 23120
rect 30411 23071 30453 23080
rect 30124 23036 30164 23071
rect 30124 22985 30164 22996
rect 30412 22986 30452 23071
rect 29931 22952 29973 22961
rect 29931 22912 29932 22952
rect 29972 22912 29973 22952
rect 29931 22903 29973 22912
rect 29932 22818 29972 22903
rect 29932 22280 29972 22289
rect 30412 22280 30452 22289
rect 29644 22240 29932 22280
rect 29932 22231 29972 22240
rect 30316 22240 30412 22280
rect 29451 22112 29493 22121
rect 29451 22072 29452 22112
rect 29492 22072 29493 22112
rect 29451 22063 29493 22072
rect 28587 21944 28629 21953
rect 28587 21904 28588 21944
rect 28628 21904 28629 21944
rect 28587 21895 28629 21904
rect 28204 21692 28244 21701
rect 28108 21652 28204 21692
rect 28204 21643 28244 21652
rect 27532 21449 27572 21568
rect 27627 21608 27669 21617
rect 28588 21608 28628 21617
rect 27627 21568 27628 21608
rect 27668 21568 27669 21608
rect 27627 21559 27669 21568
rect 28300 21568 28588 21608
rect 27628 21474 27668 21559
rect 28300 21524 28340 21568
rect 28588 21559 28628 21568
rect 29452 21608 29492 22063
rect 29452 21559 29492 21568
rect 28012 21484 28340 21524
rect 27531 21440 27573 21449
rect 27531 21400 27532 21440
rect 27572 21400 27573 21440
rect 27531 21391 27573 21400
rect 28012 21440 28052 21484
rect 28012 21391 28052 21400
rect 27628 20936 27668 20945
rect 29068 20936 29108 20945
rect 27147 20348 27189 20357
rect 27147 20308 27148 20348
rect 27188 20308 27189 20348
rect 27147 20299 27189 20308
rect 26668 20131 26708 20140
rect 26764 20140 26900 20180
rect 26092 19937 26132 20056
rect 26188 20056 26284 20096
rect 26091 19928 26133 19937
rect 26091 19888 26092 19928
rect 26132 19888 26133 19928
rect 26091 19879 26133 19888
rect 26188 19760 26228 20056
rect 26284 20047 26324 20056
rect 26380 20021 26420 20131
rect 26572 20096 26612 20105
rect 26476 20056 26572 20096
rect 26379 20012 26421 20021
rect 26379 19972 26380 20012
rect 26420 19972 26421 20012
rect 26379 19963 26421 19972
rect 26092 19720 26228 19760
rect 26284 19928 26324 19937
rect 25995 19592 26037 19601
rect 25995 19552 25996 19592
rect 26036 19552 26037 19592
rect 25995 19543 26037 19552
rect 25844 19216 25940 19256
rect 25612 18929 25652 19216
rect 25804 19172 25844 19216
rect 25804 19132 25845 19172
rect 25805 19088 25845 19132
rect 25804 19048 25845 19088
rect 25900 19088 25940 19097
rect 25611 18920 25653 18929
rect 25611 18880 25612 18920
rect 25652 18880 25653 18920
rect 25611 18871 25653 18880
rect 25804 18836 25844 19048
rect 25900 19013 25940 19048
rect 25898 19004 25940 19013
rect 25898 18964 25899 19004
rect 25939 18964 25940 19004
rect 25898 18955 25940 18964
rect 25804 18796 25940 18836
rect 24748 18124 24884 18164
rect 24940 18544 25132 18584
rect 24460 17695 24500 17704
rect 24555 17744 24597 17753
rect 24555 17704 24556 17744
rect 24596 17704 24597 17744
rect 24555 17695 24597 17704
rect 24652 17744 24692 17753
rect 24363 17660 24405 17669
rect 24363 17620 24364 17660
rect 24404 17620 24405 17660
rect 24363 17611 24405 17620
rect 24459 17492 24501 17501
rect 24459 17452 24460 17492
rect 24500 17452 24501 17492
rect 24459 17443 24501 17452
rect 24364 17072 24404 17081
rect 24268 17032 24364 17072
rect 23979 16988 24021 16997
rect 23979 16948 23980 16988
rect 24020 16948 24021 16988
rect 23979 16939 24021 16948
rect 23980 16493 24020 16939
rect 23979 16484 24021 16493
rect 23979 16444 23980 16484
rect 24020 16444 24021 16484
rect 23979 16435 24021 16444
rect 24076 16316 24116 17032
rect 24364 17023 24404 17032
rect 24460 17072 24500 17443
rect 24556 17240 24596 17695
rect 24652 17501 24692 17704
rect 24748 17744 24788 18124
rect 24940 18080 24980 18544
rect 25132 18535 25172 18544
rect 25515 18584 25557 18593
rect 25515 18544 25516 18584
rect 25556 18544 25652 18584
rect 25515 18535 25557 18544
rect 25035 18416 25077 18425
rect 25035 18376 25036 18416
rect 25076 18376 25077 18416
rect 25035 18367 25077 18376
rect 24905 18040 24980 18080
rect 24905 17759 24945 18040
rect 24905 17710 24945 17719
rect 24651 17492 24693 17501
rect 24651 17452 24652 17492
rect 24692 17452 24693 17492
rect 24651 17443 24693 17452
rect 24652 17240 24692 17249
rect 24556 17200 24652 17240
rect 24652 17191 24692 17200
rect 24460 17023 24500 17032
rect 24556 17072 24596 17081
rect 24171 16736 24213 16745
rect 24171 16696 24172 16736
rect 24212 16696 24213 16736
rect 24171 16687 24213 16696
rect 23980 16276 24116 16316
rect 23884 15728 23924 15737
rect 23788 15688 23884 15728
rect 23788 15560 23828 15569
rect 23692 15520 23788 15560
rect 23307 15476 23349 15485
rect 23307 15436 23308 15476
rect 23348 15436 23349 15476
rect 23307 15427 23349 15436
rect 23308 14720 23348 15427
rect 23788 15233 23828 15520
rect 23787 15224 23829 15233
rect 23787 15184 23788 15224
rect 23828 15184 23829 15224
rect 23787 15175 23829 15184
rect 23308 14671 23348 14680
rect 23211 14132 23253 14141
rect 23211 14092 23212 14132
rect 23252 14092 23253 14132
rect 23211 14083 23253 14092
rect 23692 13208 23732 13217
rect 23692 11705 23732 13168
rect 23691 11696 23733 11705
rect 23691 11656 23692 11696
rect 23732 11656 23733 11696
rect 23691 11647 23733 11656
rect 23884 11360 23924 15688
rect 23980 14981 24020 16276
rect 24172 15821 24212 16687
rect 24556 16316 24596 17032
rect 24748 16409 24788 17704
rect 24939 17492 24981 17501
rect 24939 17452 24940 17492
rect 24980 17452 24981 17492
rect 24939 17443 24981 17452
rect 24940 16577 24980 17443
rect 24939 16568 24981 16577
rect 24939 16528 24940 16568
rect 24980 16528 24981 16568
rect 24939 16519 24981 16528
rect 24747 16400 24789 16409
rect 24747 16360 24748 16400
rect 24788 16360 24789 16400
rect 24747 16351 24789 16360
rect 24460 16276 24596 16316
rect 24267 16232 24309 16241
rect 24267 16192 24268 16232
rect 24308 16192 24309 16232
rect 24267 16183 24309 16192
rect 24364 16232 24404 16241
rect 24171 15812 24213 15821
rect 24171 15772 24172 15812
rect 24212 15772 24213 15812
rect 24171 15763 24213 15772
rect 24076 15560 24116 15569
rect 24172 15560 24212 15763
rect 24116 15520 24212 15560
rect 24268 15560 24308 16183
rect 24364 15989 24404 16192
rect 24363 15980 24405 15989
rect 24363 15940 24364 15980
rect 24404 15940 24405 15980
rect 24363 15931 24405 15940
rect 24460 15905 24500 16276
rect 24748 16232 24788 16351
rect 24748 16183 24788 16192
rect 24555 16148 24597 16157
rect 24555 16108 24556 16148
rect 24596 16108 24597 16148
rect 24555 16099 24597 16108
rect 24556 16014 24596 16099
rect 24844 16064 24884 16073
rect 24747 15980 24789 15989
rect 24844 15980 24884 16024
rect 24747 15940 24748 15980
rect 24788 15940 24884 15980
rect 24747 15931 24789 15940
rect 24459 15896 24501 15905
rect 24940 15896 24980 16519
rect 25036 16241 25076 18367
rect 25419 17576 25461 17585
rect 25419 17536 25420 17576
rect 25460 17536 25461 17576
rect 25419 17527 25461 17536
rect 25420 17240 25460 17527
rect 25515 17408 25557 17417
rect 25515 17368 25516 17408
rect 25556 17368 25557 17408
rect 25515 17359 25557 17368
rect 25420 17191 25460 17200
rect 25227 17072 25269 17081
rect 25132 17032 25228 17072
rect 25268 17032 25269 17072
rect 25035 16232 25077 16241
rect 25035 16192 25036 16232
rect 25076 16192 25077 16232
rect 25035 16183 25077 16192
rect 25035 15980 25077 15989
rect 25035 15940 25036 15980
rect 25076 15940 25077 15980
rect 25035 15931 25077 15940
rect 24459 15856 24460 15896
rect 24500 15856 24501 15896
rect 24459 15847 24501 15856
rect 24844 15856 24980 15896
rect 24844 15737 24884 15856
rect 24843 15728 24885 15737
rect 24843 15688 24844 15728
rect 24884 15688 24885 15728
rect 24843 15679 24885 15688
rect 24076 15511 24116 15520
rect 24268 15511 24308 15520
rect 24748 15560 24788 15569
rect 24748 15485 24788 15520
rect 24459 15476 24501 15485
rect 24459 15436 24460 15476
rect 24500 15436 24501 15476
rect 24459 15427 24501 15436
rect 24747 15476 24789 15485
rect 24747 15436 24748 15476
rect 24788 15436 24789 15476
rect 24747 15427 24789 15436
rect 24844 15476 24884 15679
rect 24939 15560 24981 15569
rect 24939 15520 24940 15560
rect 24980 15520 24981 15560
rect 24939 15511 24981 15520
rect 24844 15427 24884 15436
rect 24171 15392 24213 15401
rect 24171 15352 24172 15392
rect 24212 15352 24213 15392
rect 24171 15343 24213 15352
rect 24172 15258 24212 15343
rect 24267 15140 24309 15149
rect 24267 15100 24268 15140
rect 24308 15100 24309 15140
rect 24267 15091 24309 15100
rect 23979 14972 24021 14981
rect 23979 14932 23980 14972
rect 24020 14932 24021 14972
rect 23979 14923 24021 14932
rect 24268 14720 24308 15091
rect 24268 14671 24308 14680
rect 24364 11696 24404 11705
rect 24172 11528 24212 11537
rect 24364 11528 24404 11656
rect 24212 11488 24404 11528
rect 24172 11479 24212 11488
rect 23596 11320 23924 11360
rect 23115 11276 23157 11285
rect 23115 11236 23116 11276
rect 23156 11236 23157 11276
rect 23115 11227 23157 11236
rect 23308 10940 23348 10949
rect 23116 10352 23156 10361
rect 23308 10352 23348 10900
rect 23156 10312 23348 10352
rect 23116 10303 23156 10312
rect 23019 10184 23061 10193
rect 23019 10144 23020 10184
rect 23060 10144 23061 10184
rect 23019 10135 23061 10144
rect 23308 10184 23348 10312
rect 23500 10772 23540 10781
rect 23403 10268 23445 10277
rect 23403 10228 23404 10268
rect 23444 10228 23445 10268
rect 23403 10219 23445 10228
rect 23308 10135 23348 10144
rect 22443 10100 22485 10109
rect 22443 10060 22444 10100
rect 22484 10060 22485 10100
rect 22443 10051 22485 10060
rect 22444 9512 22484 10051
rect 23404 9521 23444 10219
rect 22444 9463 22484 9472
rect 23403 9512 23445 9521
rect 23403 9472 23404 9512
rect 23444 9472 23445 9512
rect 23403 9463 23445 9472
rect 22827 9428 22869 9437
rect 22827 9388 22828 9428
rect 22868 9388 22869 9428
rect 22827 9379 22869 9388
rect 22828 9294 22868 9379
rect 23404 9344 23444 9463
rect 23404 9295 23444 9304
rect 22540 9260 22580 9269
rect 22540 9101 22580 9220
rect 22539 9092 22581 9101
rect 22539 9052 22540 9092
rect 22580 9052 22581 9092
rect 22539 9043 22581 9052
rect 23500 8924 23540 10732
rect 23020 8884 23540 8924
rect 22731 8756 22773 8765
rect 22731 8716 22732 8756
rect 22772 8716 22773 8756
rect 22731 8707 22773 8716
rect 22060 8009 22100 8632
rect 22348 8672 22388 8681
rect 22388 8632 22676 8672
rect 22348 8623 22388 8632
rect 22252 8504 22292 8513
rect 22059 8000 22101 8009
rect 22059 7960 22060 8000
rect 22100 7960 22101 8000
rect 22059 7951 22101 7960
rect 22060 7412 22100 7951
rect 22252 7589 22292 8464
rect 22539 8000 22581 8009
rect 22539 7960 22540 8000
rect 22580 7960 22581 8000
rect 22539 7951 22581 7960
rect 22636 8000 22676 8632
rect 22540 7866 22580 7951
rect 22348 7748 22388 7757
rect 22251 7580 22293 7589
rect 22251 7540 22252 7580
rect 22292 7540 22293 7580
rect 22251 7531 22293 7540
rect 22060 7363 22100 7372
rect 22251 7412 22293 7421
rect 22251 7372 22252 7412
rect 22292 7372 22293 7412
rect 22251 7363 22293 7372
rect 22155 7328 22197 7337
rect 22155 7288 22156 7328
rect 22196 7288 22197 7328
rect 22155 7279 22197 7288
rect 22156 6656 22196 7279
rect 22156 6607 22196 6616
rect 21908 6532 22100 6572
rect 21868 6523 21908 6532
rect 21004 6488 21044 6497
rect 20908 5648 20948 5657
rect 20620 5608 20908 5648
rect 20620 5144 20660 5608
rect 20908 5599 20948 5608
rect 20620 5095 20660 5104
rect 20812 5060 20852 5069
rect 21004 5060 21044 6448
rect 21579 6488 21621 6497
rect 21579 6448 21580 6488
rect 21620 6448 21621 6488
rect 21579 6439 21621 6448
rect 20852 5020 21044 5060
rect 21292 5648 21332 5657
rect 20812 5011 20852 5020
rect 20427 4724 20469 4733
rect 20427 4684 20428 4724
rect 20468 4684 20469 4724
rect 20427 4675 20469 4684
rect 20043 4136 20085 4145
rect 20043 4096 20044 4136
rect 20084 4096 20085 4136
rect 20043 4087 20085 4096
rect 20715 4136 20757 4145
rect 20715 4096 20716 4136
rect 20756 4096 20757 4136
rect 20715 4087 20757 4096
rect 20908 4136 20948 4145
rect 21292 4136 21332 5608
rect 21867 5648 21909 5657
rect 21867 5608 21868 5648
rect 21908 5608 21909 5648
rect 21867 5599 21909 5608
rect 21483 5396 21525 5405
rect 21483 5356 21484 5396
rect 21524 5356 21525 5396
rect 21483 5347 21525 5356
rect 21484 4976 21524 5347
rect 21484 4927 21524 4936
rect 21483 4808 21525 4817
rect 21483 4768 21484 4808
rect 21524 4768 21525 4808
rect 21483 4759 21525 4768
rect 20948 4096 21236 4136
rect 20908 4087 20948 4096
rect 20044 4002 20084 4087
rect 20331 4052 20373 4061
rect 20331 4012 20332 4052
rect 20372 4012 20373 4052
rect 20331 4003 20373 4012
rect 19948 3676 20084 3716
rect 17204 3424 17300 3464
rect 17164 3415 17204 3424
rect 16683 3296 16725 3305
rect 16683 3256 16684 3296
rect 16724 3256 16725 3296
rect 16683 3247 16725 3256
rect 16684 2624 16724 3247
rect 16875 2876 16917 2885
rect 16875 2836 16876 2876
rect 16916 2836 16917 2876
rect 16875 2827 16917 2836
rect 16876 2742 16916 2827
rect 17260 2792 17300 3424
rect 17260 2743 17300 2752
rect 18028 2717 18068 3424
rect 19756 3464 19796 3473
rect 19796 3424 19988 3464
rect 19756 3415 19796 3424
rect 19180 3212 19220 3221
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 16971 2708 17013 2717
rect 16971 2668 16972 2708
rect 17012 2668 17013 2708
rect 16971 2659 17013 2668
rect 17835 2708 17877 2717
rect 17835 2668 17836 2708
rect 17876 2668 17877 2708
rect 17835 2659 17877 2668
rect 18027 2708 18069 2717
rect 18027 2668 18028 2708
rect 18068 2668 18069 2708
rect 18027 2659 18069 2668
rect 16684 2575 16724 2584
rect 16972 2624 17012 2659
rect 16972 2573 17012 2584
rect 17836 2540 17876 2659
rect 18700 2633 18740 2718
rect 19180 2633 19220 3172
rect 19948 2708 19988 3424
rect 19948 2659 19988 2668
rect 18699 2624 18741 2633
rect 18699 2584 18700 2624
rect 18740 2584 18741 2624
rect 18699 2575 18741 2584
rect 19179 2624 19221 2633
rect 19179 2584 19180 2624
rect 19220 2584 19221 2624
rect 19179 2575 19221 2584
rect 18028 2540 18068 2549
rect 17836 2500 18028 2540
rect 16588 2491 16628 2500
rect 18028 2491 18068 2500
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 20044 2129 20084 3676
rect 20235 3212 20277 3221
rect 20235 3172 20236 3212
rect 20276 3172 20277 3212
rect 20235 3163 20277 3172
rect 20236 2624 20276 3163
rect 20236 2575 20276 2584
rect 20332 2624 20372 4003
rect 20716 4002 20756 4087
rect 20715 3884 20757 3893
rect 20715 3844 20716 3884
rect 20756 3844 20757 3884
rect 20715 3835 20757 3844
rect 20428 3464 20468 3473
rect 20620 3464 20660 3473
rect 20468 3424 20620 3464
rect 20428 3415 20468 3424
rect 20620 3415 20660 3424
rect 20332 2575 20372 2584
rect 20716 2624 20756 3835
rect 21003 3800 21045 3809
rect 21003 3760 21004 3800
rect 21044 3760 21045 3800
rect 21003 3751 21045 3760
rect 21004 3464 21044 3751
rect 21004 3415 21044 3424
rect 21196 3296 21236 4096
rect 21292 3809 21332 4096
rect 21291 3800 21333 3809
rect 21291 3760 21292 3800
rect 21332 3760 21333 3800
rect 21291 3751 21333 3760
rect 21196 3256 21428 3296
rect 21388 2876 21428 3256
rect 21388 2827 21428 2836
rect 21484 2708 21524 4759
rect 21676 4724 21716 4733
rect 21676 4145 21716 4684
rect 21675 4136 21717 4145
rect 21675 4096 21676 4136
rect 21716 4096 21717 4136
rect 21675 4087 21717 4096
rect 20716 2575 20756 2584
rect 21292 2668 21524 2708
rect 21868 3464 21908 5599
rect 22060 5396 22100 6532
rect 22252 6488 22292 7363
rect 22348 7160 22388 7708
rect 22636 7169 22676 7960
rect 22444 7160 22484 7169
rect 22348 7120 22444 7160
rect 22444 7111 22484 7120
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 22252 6329 22292 6448
rect 22443 6488 22485 6497
rect 22443 6448 22444 6488
rect 22484 6448 22485 6488
rect 22443 6439 22485 6448
rect 22444 6354 22484 6439
rect 22251 6320 22293 6329
rect 22251 6280 22252 6320
rect 22292 6280 22293 6320
rect 22636 6320 22676 7111
rect 22732 6581 22772 8707
rect 22923 8504 22965 8513
rect 22923 8464 22924 8504
rect 22964 8464 22965 8504
rect 22923 8455 22965 8464
rect 22924 8370 22964 8455
rect 23020 8429 23060 8884
rect 23403 8756 23445 8765
rect 23596 8756 23636 11320
rect 24171 11276 24213 11285
rect 24171 11236 24172 11276
rect 24212 11236 24213 11276
rect 24171 11227 24213 11236
rect 23692 11024 23732 11033
rect 23692 10277 23732 10984
rect 23787 11024 23829 11033
rect 24172 11024 24212 11227
rect 24364 11117 24404 11488
rect 24363 11108 24405 11117
rect 24363 11068 24364 11108
rect 24404 11068 24405 11108
rect 24363 11059 24405 11068
rect 23787 10984 23788 11024
rect 23828 10984 23829 11024
rect 23787 10975 23829 10984
rect 24076 10984 24172 11024
rect 23788 10890 23828 10975
rect 23691 10268 23733 10277
rect 23691 10228 23692 10268
rect 23732 10228 23733 10268
rect 23691 10219 23733 10228
rect 23980 10100 24020 10109
rect 23692 10060 23980 10100
rect 23692 9512 23732 10060
rect 23980 10051 24020 10060
rect 24076 9680 24116 10984
rect 24172 10975 24212 10984
rect 24460 10940 24500 15427
rect 24748 15425 24788 15427
rect 24940 15392 24980 15511
rect 24940 15343 24980 15352
rect 25036 15476 25076 15931
rect 25132 15653 25172 17032
rect 25227 17023 25269 17032
rect 25324 17072 25364 17081
rect 25228 16938 25268 17023
rect 25324 16661 25364 17032
rect 25516 17072 25556 17359
rect 25516 17023 25556 17032
rect 25612 16745 25652 18544
rect 25803 18500 25845 18509
rect 25803 18460 25804 18500
rect 25844 18460 25845 18500
rect 25803 18451 25845 18460
rect 25707 18416 25749 18425
rect 25707 18376 25708 18416
rect 25748 18376 25749 18416
rect 25707 18367 25749 18376
rect 25708 18282 25748 18367
rect 25707 17576 25749 17585
rect 25707 17536 25708 17576
rect 25748 17536 25749 17576
rect 25707 17527 25749 17536
rect 25611 16736 25653 16745
rect 25611 16696 25612 16736
rect 25652 16696 25653 16736
rect 25611 16687 25653 16696
rect 25323 16652 25365 16661
rect 25323 16612 25324 16652
rect 25364 16612 25365 16652
rect 25323 16603 25365 16612
rect 25324 16064 25364 16603
rect 25419 16484 25461 16493
rect 25419 16444 25420 16484
rect 25460 16444 25461 16484
rect 25419 16435 25461 16444
rect 25228 16024 25364 16064
rect 25131 15644 25173 15653
rect 25131 15604 25132 15644
rect 25172 15604 25173 15644
rect 25131 15595 25173 15604
rect 25132 15560 25172 15595
rect 25132 15510 25172 15520
rect 24747 14972 24789 14981
rect 24747 14932 24748 14972
rect 24788 14932 24789 14972
rect 24747 14923 24789 14932
rect 24748 14720 24788 14923
rect 25036 14720 25076 15436
rect 24748 14671 24788 14680
rect 24940 14680 25076 14720
rect 24843 13292 24885 13301
rect 24843 13252 24844 13292
rect 24884 13252 24885 13292
rect 24843 13243 24885 13252
rect 24844 13158 24884 13243
rect 24748 12536 24788 12545
rect 24748 12377 24788 12496
rect 24747 12368 24789 12377
rect 24747 12328 24748 12368
rect 24788 12328 24789 12368
rect 24747 12319 24789 12328
rect 24747 11024 24789 11033
rect 24747 10984 24748 11024
rect 24788 10984 24789 11024
rect 24747 10975 24789 10984
rect 24364 10900 24500 10940
rect 24364 10193 24404 10900
rect 24460 10772 24500 10781
rect 24363 10184 24405 10193
rect 24363 10144 24364 10184
rect 24404 10144 24405 10184
rect 24363 10135 24405 10144
rect 24460 10184 24500 10732
rect 24652 10184 24692 10193
rect 24460 10135 24500 10144
rect 24556 10144 24652 10184
rect 24172 10016 24212 10025
rect 24556 10016 24596 10144
rect 24652 10135 24692 10144
rect 24748 10184 24788 10975
rect 24940 10352 24980 14680
rect 25132 14552 25172 14561
rect 25132 13973 25172 14512
rect 25131 13964 25173 13973
rect 25131 13924 25132 13964
rect 25172 13924 25173 13964
rect 25131 13915 25173 13924
rect 25036 11528 25076 11537
rect 25036 11024 25076 11488
rect 25131 11108 25173 11117
rect 25131 11068 25132 11108
rect 25172 11068 25173 11108
rect 25131 11059 25173 11068
rect 25036 10975 25076 10984
rect 24940 10312 25076 10352
rect 24748 10135 24788 10144
rect 24940 10184 24980 10193
rect 24843 10100 24885 10109
rect 24940 10100 24980 10144
rect 24843 10060 24844 10100
rect 24884 10060 24885 10100
rect 24843 10051 24885 10060
rect 24938 10060 24980 10100
rect 24212 9976 24596 10016
rect 24172 9967 24212 9976
rect 23692 9463 23732 9472
rect 23980 9640 24116 9680
rect 23980 8849 24020 9640
rect 24076 9512 24116 9521
rect 23979 8840 24021 8849
rect 23979 8800 23980 8840
rect 24020 8800 24021 8840
rect 23979 8791 24021 8800
rect 23403 8716 23404 8756
rect 23444 8716 23445 8756
rect 23403 8707 23445 8716
rect 23500 8716 23636 8756
rect 23116 8672 23156 8681
rect 23019 8420 23061 8429
rect 23019 8380 23020 8420
rect 23060 8380 23061 8420
rect 23019 8371 23061 8380
rect 22828 8168 22868 8177
rect 22828 6992 22868 8128
rect 23020 7925 23060 8371
rect 23116 8009 23156 8632
rect 23212 8672 23252 8681
rect 23115 8000 23157 8009
rect 23115 7960 23116 8000
rect 23156 7960 23157 8000
rect 23115 7951 23157 7960
rect 23212 8000 23252 8632
rect 23404 8672 23444 8707
rect 23404 8621 23444 8632
rect 23500 8672 23540 8716
rect 23884 8672 23924 8681
rect 23500 8252 23540 8632
rect 23596 8632 23884 8672
rect 23596 8513 23636 8632
rect 23884 8623 23924 8632
rect 23980 8672 24020 8681
rect 23595 8504 23637 8513
rect 23595 8464 23596 8504
rect 23636 8464 23637 8504
rect 23595 8455 23637 8464
rect 23692 8504 23732 8513
rect 23980 8504 24020 8632
rect 24076 8597 24116 9472
rect 24171 9512 24213 9521
rect 24171 9472 24172 9512
rect 24212 9472 24213 9512
rect 24171 9463 24213 9472
rect 24268 9512 24308 9976
rect 24844 9966 24884 10051
rect 24938 10016 24978 10060
rect 24938 9976 24980 10016
rect 24843 9596 24885 9605
rect 24843 9556 24844 9596
rect 24884 9556 24885 9596
rect 24843 9547 24885 9556
rect 24268 9463 24308 9472
rect 24364 9512 24404 9521
rect 24556 9512 24596 9521
rect 24404 9472 24556 9512
rect 24364 9463 24404 9472
rect 24556 9463 24596 9472
rect 24652 9512 24692 9521
rect 24172 9378 24212 9463
rect 24555 9344 24597 9353
rect 24555 9304 24556 9344
rect 24596 9304 24597 9344
rect 24555 9295 24597 9304
rect 24171 9008 24213 9017
rect 24171 8968 24172 9008
rect 24212 8968 24213 9008
rect 24171 8959 24213 8968
rect 24172 8924 24212 8959
rect 24172 8873 24212 8884
rect 24172 8672 24212 8681
rect 24075 8588 24117 8597
rect 24075 8548 24076 8588
rect 24116 8548 24117 8588
rect 24075 8539 24117 8548
rect 23732 8464 24020 8504
rect 23692 8455 23732 8464
rect 23500 8212 23636 8252
rect 23403 8168 23445 8177
rect 23403 8128 23404 8168
rect 23444 8128 23445 8168
rect 23403 8119 23445 8128
rect 23404 8034 23444 8119
rect 23019 7916 23061 7925
rect 23019 7876 23020 7916
rect 23060 7876 23061 7916
rect 23019 7867 23061 7876
rect 23019 7748 23061 7757
rect 23019 7708 23020 7748
rect 23060 7708 23061 7748
rect 23019 7699 23061 7708
rect 22923 7580 22965 7589
rect 22923 7540 22924 7580
rect 22964 7540 22965 7580
rect 22923 7531 22965 7540
rect 22924 7160 22964 7531
rect 22924 7111 22964 7120
rect 23020 7160 23060 7699
rect 23212 7589 23252 7960
rect 23500 8000 23540 8011
rect 23500 7925 23540 7960
rect 23307 7916 23349 7925
rect 23307 7876 23308 7916
rect 23348 7876 23349 7916
rect 23307 7867 23349 7876
rect 23499 7916 23541 7925
rect 23499 7876 23500 7916
rect 23540 7876 23541 7916
rect 23499 7867 23541 7876
rect 23211 7580 23253 7589
rect 23211 7540 23212 7580
rect 23252 7540 23253 7580
rect 23211 7531 23253 7540
rect 23020 7111 23060 7120
rect 23212 7160 23252 7169
rect 23212 6992 23252 7120
rect 23308 7160 23348 7867
rect 23464 7328 23506 7337
rect 23464 7288 23465 7328
rect 23505 7288 23506 7328
rect 23464 7279 23506 7288
rect 23465 7175 23505 7279
rect 23465 7126 23505 7135
rect 23308 7111 23348 7120
rect 22828 6952 23252 6992
rect 23307 6992 23349 7001
rect 23307 6952 23308 6992
rect 23348 6952 23349 6992
rect 23307 6943 23349 6952
rect 23404 6992 23444 7001
rect 23115 6740 23157 6749
rect 23115 6700 23116 6740
rect 23156 6700 23157 6740
rect 23115 6691 23157 6700
rect 23116 6656 23156 6691
rect 23116 6605 23156 6616
rect 22731 6572 22773 6581
rect 22731 6532 22732 6572
rect 22772 6532 22773 6572
rect 22731 6523 22773 6532
rect 23211 6488 23253 6497
rect 23211 6448 23212 6488
rect 23252 6448 23253 6488
rect 23211 6439 23253 6448
rect 22923 6320 22965 6329
rect 22636 6280 22772 6320
rect 22251 6271 22293 6280
rect 22155 5648 22197 5657
rect 22155 5608 22156 5648
rect 22196 5608 22197 5648
rect 22155 5599 22197 5608
rect 22156 5514 22196 5599
rect 22060 5356 22196 5396
rect 22156 5202 22196 5356
rect 21963 4976 22005 4985
rect 21963 4936 21964 4976
rect 22004 4936 22005 4976
rect 21963 4927 22005 4936
rect 22060 4976 22100 4985
rect 21964 4842 22004 4927
rect 22060 4817 22100 4936
rect 22156 4901 22196 5162
rect 22732 5069 22772 6280
rect 22923 6280 22924 6320
rect 22964 6280 22965 6320
rect 22923 6271 22965 6280
rect 22347 5060 22389 5069
rect 22347 5020 22348 5060
rect 22388 5020 22389 5060
rect 22347 5011 22389 5020
rect 22731 5060 22773 5069
rect 22731 5020 22732 5060
rect 22772 5020 22773 5060
rect 22731 5011 22773 5020
rect 22348 4976 22388 5011
rect 22348 4925 22388 4936
rect 22155 4892 22197 4901
rect 22155 4852 22156 4892
rect 22196 4852 22292 4892
rect 22155 4843 22197 4852
rect 22059 4808 22101 4817
rect 22059 4768 22060 4808
rect 22100 4768 22101 4808
rect 22059 4759 22101 4768
rect 22155 4724 22197 4733
rect 22155 4684 22156 4724
rect 22196 4684 22197 4724
rect 22155 4675 22197 4684
rect 22156 4145 22196 4675
rect 22155 4136 22197 4145
rect 22155 4096 22156 4136
rect 22196 4096 22197 4136
rect 22155 4087 22197 4096
rect 22156 4002 22196 4087
rect 22059 3800 22101 3809
rect 22059 3760 22060 3800
rect 22100 3760 22101 3800
rect 22059 3751 22101 3760
rect 20043 2120 20085 2129
rect 20043 2080 20044 2120
rect 20084 2080 20085 2120
rect 20043 2071 20085 2080
rect 20811 2120 20853 2129
rect 20811 2080 20812 2120
rect 20852 2080 20853 2120
rect 20811 2071 20853 2080
rect 20812 1986 20852 2071
rect 16300 1952 16340 1961
rect 16012 1912 16300 1952
rect 15436 1280 15476 1912
rect 16300 1903 16340 1912
rect 21003 1952 21045 1961
rect 21003 1912 21004 1952
rect 21044 1912 21045 1952
rect 21003 1903 21045 1912
rect 21292 1952 21332 2668
rect 21868 2633 21908 3424
rect 22060 2885 22100 3751
rect 22059 2876 22101 2885
rect 22059 2836 22060 2876
rect 22100 2836 22101 2876
rect 22059 2827 22101 2836
rect 21963 2708 22005 2717
rect 21963 2668 21964 2708
rect 22004 2668 22005 2708
rect 21963 2659 22005 2668
rect 21867 2624 21909 2633
rect 21867 2584 21868 2624
rect 21908 2584 21909 2624
rect 21867 2575 21909 2584
rect 21964 2574 22004 2659
rect 22060 2120 22100 2827
rect 22060 2071 22100 2080
rect 22252 1961 22292 4852
rect 22924 3464 22964 6271
rect 23212 5900 23252 6439
rect 23308 6404 23348 6943
rect 23404 6833 23444 6952
rect 23499 6992 23541 7001
rect 23499 6952 23500 6992
rect 23540 6952 23541 6992
rect 23499 6943 23541 6952
rect 23403 6824 23445 6833
rect 23403 6784 23404 6824
rect 23444 6784 23445 6824
rect 23403 6775 23445 6784
rect 23500 6656 23540 6943
rect 23500 6607 23540 6616
rect 23596 6497 23636 8212
rect 24172 8177 24212 8632
rect 24171 8168 24213 8177
rect 24171 8128 24172 8168
rect 24212 8128 24213 8168
rect 24171 8119 24213 8128
rect 24076 8000 24116 8009
rect 23788 7991 23828 8000
rect 23691 7916 23733 7925
rect 23788 7916 23828 7951
rect 23691 7876 23692 7916
rect 23732 7876 23828 7916
rect 23980 7960 24076 8000
rect 23691 7867 23733 7876
rect 23692 7160 23732 7867
rect 23883 7580 23925 7589
rect 23883 7540 23884 7580
rect 23924 7540 23925 7580
rect 23883 7531 23925 7540
rect 23788 7169 23828 7254
rect 23692 7111 23732 7120
rect 23787 7160 23829 7169
rect 23787 7120 23788 7160
rect 23828 7120 23829 7160
rect 23787 7111 23829 7120
rect 23884 7085 23924 7531
rect 23980 7169 24020 7960
rect 24076 7951 24116 7960
rect 24171 8000 24213 8009
rect 24171 7960 24172 8000
rect 24212 7960 24213 8000
rect 24171 7951 24213 7960
rect 24076 7748 24116 7757
rect 23979 7160 24021 7169
rect 23979 7120 23980 7160
rect 24020 7120 24021 7160
rect 24076 7160 24116 7708
rect 24172 7412 24212 7951
rect 24172 7363 24212 7372
rect 24556 7253 24596 9295
rect 24652 9017 24692 9472
rect 24748 9512 24788 9521
rect 24748 9260 24788 9472
rect 24844 9462 24884 9547
rect 24940 9353 24980 9976
rect 24939 9344 24981 9353
rect 24939 9304 24940 9344
rect 24980 9304 24981 9344
rect 24939 9295 24981 9304
rect 24748 9220 24884 9260
rect 24651 9008 24693 9017
rect 24651 8968 24652 9008
rect 24692 8968 24693 9008
rect 24651 8959 24693 8968
rect 24844 8882 24884 9220
rect 24651 8840 24693 8849
rect 24651 8800 24652 8840
rect 24692 8800 24693 8840
rect 25036 8849 25076 10312
rect 25132 10268 25172 11059
rect 25132 10219 25172 10228
rect 25228 9512 25268 16024
rect 25323 15560 25365 15569
rect 25323 15520 25324 15560
rect 25364 15520 25365 15560
rect 25323 15511 25365 15520
rect 25420 15560 25460 16435
rect 25611 16400 25653 16409
rect 25611 16360 25612 16400
rect 25652 16360 25653 16400
rect 25611 16351 25653 16360
rect 25612 15728 25652 16351
rect 25612 15679 25652 15688
rect 25420 15511 25460 15520
rect 25612 15560 25652 15569
rect 25324 15426 25364 15511
rect 25612 15401 25652 15520
rect 25708 15485 25748 17527
rect 25707 15476 25749 15485
rect 25707 15436 25708 15476
rect 25748 15436 25749 15476
rect 25707 15427 25749 15436
rect 25611 15392 25653 15401
rect 25611 15352 25612 15392
rect 25652 15352 25653 15392
rect 25611 15343 25653 15352
rect 25611 15056 25653 15065
rect 25611 15016 25612 15056
rect 25652 15016 25653 15056
rect 25611 15007 25653 15016
rect 25612 14720 25652 15007
rect 25612 14671 25652 14680
rect 25804 14216 25844 18451
rect 25900 17585 25940 18796
rect 25996 18164 26036 19543
rect 26092 19256 26132 19720
rect 26092 19207 26132 19216
rect 25996 18124 26228 18164
rect 26091 17996 26133 18005
rect 26091 17956 26092 17996
rect 26132 17956 26133 17996
rect 26091 17947 26133 17956
rect 25995 17912 26037 17921
rect 25995 17872 25996 17912
rect 26036 17872 26037 17912
rect 25995 17863 26037 17872
rect 25899 17576 25941 17585
rect 25899 17536 25900 17576
rect 25940 17536 25941 17576
rect 25899 17527 25941 17536
rect 25899 17408 25941 17417
rect 25899 17368 25900 17408
rect 25940 17368 25941 17408
rect 25899 17359 25941 17368
rect 25900 15644 25940 17359
rect 25900 15595 25940 15604
rect 25996 15560 26036 17863
rect 26092 17862 26132 17947
rect 26092 17744 26132 17753
rect 26092 16232 26132 17704
rect 26188 17669 26228 18124
rect 26284 17921 26324 19888
rect 26476 19853 26516 20056
rect 26572 20047 26612 20056
rect 26764 20096 26804 20140
rect 26475 19844 26517 19853
rect 26475 19804 26476 19844
rect 26516 19804 26517 19844
rect 26475 19795 26517 19804
rect 26476 18416 26516 19795
rect 26764 19769 26804 20056
rect 26955 20096 26997 20105
rect 26955 20056 26956 20096
rect 26996 20056 26997 20096
rect 26955 20047 26997 20056
rect 26956 19962 26996 20047
rect 26763 19760 26805 19769
rect 26763 19720 26764 19760
rect 26804 19720 26805 19760
rect 26763 19711 26805 19720
rect 26667 19256 26709 19265
rect 26667 19216 26668 19256
rect 26708 19216 26709 19256
rect 26667 19207 26709 19216
rect 26668 19122 26708 19207
rect 27147 19088 27189 19097
rect 27147 19048 27148 19088
rect 27188 19048 27189 19088
rect 27147 19039 27189 19048
rect 27148 18954 27188 19039
rect 26763 18920 26805 18929
rect 26763 18880 26764 18920
rect 26804 18880 26805 18920
rect 26763 18871 26805 18880
rect 26668 18761 26708 18846
rect 26667 18752 26709 18761
rect 26667 18712 26668 18752
rect 26708 18712 26709 18752
rect 26667 18703 26709 18712
rect 26667 18584 26709 18593
rect 26667 18544 26668 18584
rect 26708 18544 26709 18584
rect 26667 18535 26709 18544
rect 26764 18584 26804 18871
rect 26764 18535 26804 18544
rect 27148 18584 27188 18593
rect 27532 18584 27572 18593
rect 26571 18500 26613 18509
rect 26571 18460 26572 18500
rect 26612 18460 26613 18500
rect 26571 18451 26613 18460
rect 26476 18367 26516 18376
rect 26572 18366 26612 18451
rect 26668 18450 26708 18535
rect 27148 18005 27188 18544
rect 27244 18544 27532 18584
rect 27147 17996 27189 18005
rect 27147 17956 27148 17996
rect 27188 17956 27189 17996
rect 27147 17947 27189 17956
rect 26283 17912 26325 17921
rect 27244 17912 27284 18544
rect 27532 18535 27572 18544
rect 27628 17912 27668 20896
rect 28972 20896 29068 20936
rect 27915 20096 27957 20105
rect 27915 20056 27916 20096
rect 27956 20056 27957 20096
rect 27915 20047 27957 20056
rect 28588 20096 28628 20105
rect 27916 19962 27956 20047
rect 28011 20012 28053 20021
rect 28011 19972 28012 20012
rect 28052 19972 28053 20012
rect 28011 19963 28053 19972
rect 28012 19256 28052 19963
rect 28395 19928 28437 19937
rect 28395 19888 28396 19928
rect 28436 19888 28437 19928
rect 28395 19879 28437 19888
rect 28396 19794 28436 19879
rect 28299 19760 28341 19769
rect 28299 19720 28300 19760
rect 28340 19720 28341 19760
rect 28299 19711 28341 19720
rect 28012 19207 28052 19216
rect 28108 19256 28148 19265
rect 26283 17872 26284 17912
rect 26324 17872 26612 17912
rect 26283 17863 26325 17872
rect 26284 17744 26324 17753
rect 26572 17744 26612 17872
rect 27244 17863 27284 17872
rect 27436 17872 27668 17912
rect 27820 19088 27860 19097
rect 26324 17704 26420 17744
rect 26284 17695 26324 17704
rect 26187 17660 26229 17669
rect 26187 17620 26188 17660
rect 26228 17620 26229 17660
rect 26187 17611 26229 17620
rect 26283 17492 26325 17501
rect 26283 17452 26284 17492
rect 26324 17452 26325 17492
rect 26283 17443 26325 17452
rect 26284 16736 26324 17443
rect 26380 17240 26420 17704
rect 26572 17695 26612 17704
rect 27436 17744 27476 17872
rect 26763 17660 26805 17669
rect 26763 17620 26764 17660
rect 26804 17620 26805 17660
rect 26763 17611 26805 17620
rect 26475 17576 26517 17585
rect 26475 17536 26476 17576
rect 26516 17536 26517 17576
rect 26475 17527 26517 17536
rect 26476 17442 26516 17527
rect 26764 17526 26804 17611
rect 27243 17576 27285 17585
rect 27243 17536 27244 17576
rect 27284 17536 27285 17576
rect 27243 17527 27285 17536
rect 26667 17324 26709 17333
rect 26667 17284 26668 17324
rect 26708 17284 26709 17324
rect 26667 17275 26709 17284
rect 27051 17324 27093 17333
rect 27051 17284 27052 17324
rect 27092 17284 27093 17324
rect 27051 17275 27093 17284
rect 26572 17240 26612 17249
rect 26380 17200 26572 17240
rect 26572 17191 26612 17200
rect 26476 17072 26516 17081
rect 26284 16696 26420 16736
rect 26380 16493 26420 16696
rect 26379 16484 26421 16493
rect 26379 16444 26380 16484
rect 26420 16444 26421 16484
rect 26379 16435 26421 16444
rect 26188 16232 26228 16241
rect 26092 16192 26188 16232
rect 26188 16183 26228 16192
rect 26284 16232 26324 16241
rect 26092 15560 26132 15569
rect 25996 15520 26092 15560
rect 25899 15476 25941 15485
rect 25899 15436 25900 15476
rect 25940 15436 25941 15476
rect 25899 15427 25941 15436
rect 25900 14813 25940 15427
rect 25899 14804 25941 14813
rect 25899 14764 25900 14804
rect 25940 14764 25941 14804
rect 25899 14755 25941 14764
rect 25996 14720 26036 15520
rect 26092 15511 26132 15520
rect 26284 15065 26324 16192
rect 26380 16232 26420 16435
rect 26476 16409 26516 17032
rect 26668 17072 26708 17275
rect 26668 17023 26708 17032
rect 26764 17072 26804 17081
rect 26571 16652 26613 16661
rect 26571 16612 26572 16652
rect 26612 16612 26613 16652
rect 26571 16603 26613 16612
rect 26475 16400 26517 16409
rect 26475 16360 26476 16400
rect 26516 16360 26517 16400
rect 26475 16351 26517 16360
rect 26380 16183 26420 16192
rect 26476 16232 26516 16241
rect 26572 16232 26612 16603
rect 26668 16484 26708 16493
rect 26764 16484 26804 17032
rect 26955 16820 26997 16829
rect 26955 16780 26956 16820
rect 26996 16780 26997 16820
rect 26955 16771 26997 16780
rect 26708 16444 26804 16484
rect 26668 16435 26708 16444
rect 26668 16325 26708 16356
rect 26667 16316 26709 16325
rect 26667 16276 26668 16316
rect 26708 16276 26709 16316
rect 26667 16267 26709 16276
rect 26516 16192 26612 16232
rect 26668 16232 26708 16267
rect 26476 16183 26516 16192
rect 26668 15737 26708 16192
rect 26860 16232 26900 16241
rect 26860 16073 26900 16192
rect 26956 16232 26996 16771
rect 27052 16241 27092 17275
rect 27147 17240 27189 17249
rect 27147 17200 27148 17240
rect 27188 17200 27189 17240
rect 27147 17191 27189 17200
rect 27148 16829 27188 17191
rect 27244 17072 27284 17527
rect 27244 16997 27284 17032
rect 27340 17072 27380 17081
rect 27436 17072 27476 17704
rect 27628 17744 27668 17753
rect 27532 17660 27572 17669
rect 27532 17072 27572 17620
rect 27628 17585 27668 17704
rect 27627 17576 27669 17585
rect 27627 17536 27628 17576
rect 27668 17536 27669 17576
rect 27627 17527 27669 17536
rect 27724 17333 27764 17393
rect 27723 17324 27765 17333
rect 27723 17275 27724 17324
rect 27764 17275 27765 17324
rect 27724 17249 27764 17258
rect 27820 17156 27860 19048
rect 28108 19013 28148 19216
rect 28204 19256 28244 19265
rect 28107 19004 28149 19013
rect 28107 18964 28108 19004
rect 28148 18964 28149 19004
rect 28107 18955 28149 18964
rect 28204 18929 28244 19216
rect 28300 19256 28340 19711
rect 28300 19207 28340 19216
rect 28588 18929 28628 20056
rect 28972 20096 29012 20896
rect 29068 20887 29108 20896
rect 30316 20105 30356 22240
rect 30412 22231 30452 22240
rect 30508 20180 30548 26608
rect 30699 26599 30741 26608
rect 30603 25892 30645 25901
rect 30603 25852 30604 25892
rect 30644 25852 30645 25892
rect 30603 25843 30645 25852
rect 30604 25758 30644 25843
rect 30603 25304 30645 25313
rect 30603 25264 30604 25304
rect 30644 25264 30645 25304
rect 30603 25255 30645 25264
rect 30604 24641 30644 25255
rect 30603 24632 30645 24641
rect 30603 24592 30604 24632
rect 30644 24592 30645 24632
rect 30603 24583 30645 24592
rect 30604 22532 30644 24583
rect 30700 23381 30740 26599
rect 30796 25565 30836 26944
rect 30988 26909 31028 27019
rect 30987 26900 31029 26909
rect 30987 26860 30988 26900
rect 31028 26860 31029 26900
rect 30987 26851 31029 26860
rect 31084 26825 31124 26910
rect 30891 26816 30933 26825
rect 30891 26776 30892 26816
rect 30932 26776 30933 26816
rect 30891 26767 30933 26776
rect 31083 26816 31125 26825
rect 31083 26776 31084 26816
rect 31124 26776 31125 26816
rect 31083 26767 31125 26776
rect 31180 26816 31220 27280
rect 31372 27245 31412 28447
rect 31468 28337 31508 29800
rect 31659 29840 31701 29849
rect 31659 29800 31660 29840
rect 31700 29800 31701 29840
rect 31659 29791 31701 29800
rect 31756 29840 31796 29849
rect 31660 29706 31700 29791
rect 31564 29672 31604 29681
rect 31564 29177 31604 29632
rect 31756 29345 31796 29800
rect 31755 29336 31797 29345
rect 31755 29296 31756 29336
rect 31796 29296 31797 29336
rect 31755 29287 31797 29296
rect 31563 29168 31605 29177
rect 31563 29128 31564 29168
rect 31604 29128 31605 29168
rect 31563 29119 31605 29128
rect 31756 29093 31796 29178
rect 31755 29084 31797 29093
rect 31755 29044 31756 29084
rect 31796 29044 31797 29084
rect 31755 29035 31797 29044
rect 31852 28748 31892 31900
rect 31948 31529 31988 32152
rect 32043 32192 32085 32201
rect 32043 32152 32044 32192
rect 32084 32152 32085 32192
rect 32043 32143 32085 32152
rect 32140 32192 32180 32203
rect 32044 32058 32084 32143
rect 32140 32117 32180 32152
rect 32139 32108 32181 32117
rect 32139 32068 32140 32108
rect 32180 32068 32181 32108
rect 32139 32059 32181 32068
rect 32236 31940 32276 33832
rect 32332 32873 32372 34924
rect 32428 34385 32468 35848
rect 32524 35888 32564 35897
rect 32524 35309 32564 35848
rect 32716 35888 32756 36763
rect 36076 36728 36116 36737
rect 40012 36728 40052 36737
rect 32716 35839 32756 35848
rect 33100 36604 33428 36644
rect 33100 35888 33140 36604
rect 33388 36560 33428 36604
rect 33484 36560 33524 36569
rect 33388 36520 33484 36560
rect 33484 36511 33524 36520
rect 35595 36560 35637 36569
rect 35595 36520 35596 36560
rect 35636 36520 35637 36560
rect 35595 36511 35637 36520
rect 35404 36476 35444 36485
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 33100 35839 33140 35848
rect 33964 35888 34004 35897
rect 32523 35300 32565 35309
rect 32523 35260 32524 35300
rect 32564 35260 32565 35300
rect 32523 35251 32565 35260
rect 33195 35300 33237 35309
rect 33195 35260 33196 35300
rect 33236 35260 33237 35300
rect 33195 35251 33237 35260
rect 32907 35216 32949 35225
rect 32907 35176 32908 35216
rect 32948 35176 32949 35216
rect 32907 35167 32949 35176
rect 33100 35216 33140 35227
rect 32908 35082 32948 35167
rect 33100 35141 33140 35176
rect 33196 35166 33236 35251
rect 33964 35225 34004 35848
rect 35211 35888 35253 35897
rect 35211 35848 35212 35888
rect 35252 35848 35253 35888
rect 35211 35839 35253 35848
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 34731 35384 34773 35393
rect 34731 35344 34732 35384
rect 34772 35344 34773 35384
rect 34731 35335 34773 35344
rect 34635 35300 34677 35309
rect 34635 35260 34636 35300
rect 34676 35260 34677 35300
rect 34635 35251 34677 35260
rect 33963 35216 34005 35225
rect 33963 35176 33964 35216
rect 34004 35176 34005 35216
rect 33963 35167 34005 35176
rect 34252 35216 34292 35225
rect 33099 35132 33141 35141
rect 33099 35092 33100 35132
rect 33140 35092 33141 35132
rect 33099 35083 33141 35092
rect 33868 34964 33908 34973
rect 33908 34924 34004 34964
rect 33868 34915 33908 34924
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 32523 34628 32565 34637
rect 32523 34588 32524 34628
rect 32564 34588 32565 34628
rect 32523 34579 32565 34588
rect 32427 34376 32469 34385
rect 32427 34336 32428 34376
rect 32468 34336 32469 34376
rect 32427 34327 32469 34336
rect 32428 33788 32468 34327
rect 32428 33739 32468 33748
rect 32331 32864 32373 32873
rect 32331 32824 32332 32864
rect 32372 32824 32373 32864
rect 32331 32815 32373 32824
rect 32332 32730 32372 32815
rect 32524 32528 32564 34579
rect 33388 34504 33908 34544
rect 33196 34376 33236 34385
rect 33196 34049 33236 34336
rect 33388 34376 33428 34504
rect 33388 34327 33428 34336
rect 33771 34376 33813 34385
rect 33771 34336 33772 34376
rect 33812 34336 33813 34376
rect 33771 34327 33813 34336
rect 33772 34242 33812 34327
rect 33195 34040 33237 34049
rect 33195 34000 33196 34040
rect 33236 34000 33237 34040
rect 33195 33991 33237 34000
rect 33771 34040 33813 34049
rect 33771 34000 33772 34040
rect 33812 34000 33813 34040
rect 33771 33991 33813 34000
rect 33196 33704 33236 33713
rect 32332 32488 32564 32528
rect 33004 33664 33196 33704
rect 32332 32192 32372 32488
rect 32427 32360 32469 32369
rect 32427 32320 32428 32360
rect 32468 32320 32469 32360
rect 32427 32311 32469 32320
rect 32332 32117 32372 32152
rect 32428 32192 32468 32311
rect 32428 32143 32468 32152
rect 32524 32192 32564 32201
rect 32331 32108 32373 32117
rect 32331 32068 32332 32108
rect 32372 32068 32373 32108
rect 32331 32059 32373 32068
rect 32332 32028 32372 32059
rect 32524 32024 32564 32152
rect 32620 32192 32660 32201
rect 32660 32152 32948 32192
rect 32620 32143 32660 32152
rect 32140 31900 32276 31940
rect 32428 31984 32564 32024
rect 31947 31520 31989 31529
rect 31947 31480 31948 31520
rect 31988 31480 31989 31520
rect 31947 31471 31989 31480
rect 31948 30596 31988 30605
rect 31948 30269 31988 30556
rect 31947 30260 31989 30269
rect 31947 30220 31948 30260
rect 31988 30220 31989 30260
rect 31947 30211 31989 30220
rect 31947 29840 31989 29849
rect 31947 29800 31948 29840
rect 31988 29800 31989 29840
rect 31947 29791 31989 29800
rect 31948 29706 31988 29791
rect 31947 29168 31989 29177
rect 31947 29128 31948 29168
rect 31988 29128 31989 29168
rect 31947 29119 31989 29128
rect 31948 29034 31988 29119
rect 31564 28708 31892 28748
rect 31467 28328 31509 28337
rect 31467 28288 31468 28328
rect 31508 28288 31509 28328
rect 31467 28279 31509 28288
rect 31468 27656 31508 27665
rect 31468 27497 31508 27616
rect 31564 27656 31604 28708
rect 32140 27833 32180 31900
rect 32428 31529 32468 31984
rect 32812 31940 32852 31949
rect 32524 31900 32812 31940
rect 32427 31520 32469 31529
rect 32427 31480 32428 31520
rect 32468 31480 32469 31520
rect 32427 31471 32469 31480
rect 32524 31352 32564 31900
rect 32812 31891 32852 31900
rect 32908 31529 32948 32152
rect 32907 31520 32949 31529
rect 32907 31480 32908 31520
rect 32948 31480 32949 31520
rect 32907 31471 32949 31480
rect 32524 31303 32564 31312
rect 32236 31193 32276 31278
rect 32235 31184 32277 31193
rect 32235 31144 32236 31184
rect 32276 31144 32277 31184
rect 32235 31135 32277 31144
rect 32428 31184 32468 31193
rect 32428 30848 32468 31144
rect 32332 30808 32468 30848
rect 32235 30260 32277 30269
rect 32235 30220 32236 30260
rect 32276 30220 32277 30260
rect 32235 30211 32277 30220
rect 32236 28328 32276 30211
rect 32332 29429 32372 30808
rect 32427 30680 32469 30689
rect 32427 30640 32428 30680
rect 32468 30640 32469 30680
rect 32427 30631 32469 30640
rect 32428 30546 32468 30631
rect 33004 30596 33044 33664
rect 33196 33655 33236 33664
rect 33676 33704 33716 33715
rect 33676 33629 33716 33664
rect 33772 33704 33812 33991
rect 33868 33872 33908 34504
rect 33964 34208 34004 34924
rect 34252 34889 34292 35176
rect 34539 35216 34581 35225
rect 34539 35176 34540 35216
rect 34580 35176 34581 35216
rect 34539 35167 34581 35176
rect 34347 35132 34389 35141
rect 34347 35092 34348 35132
rect 34388 35092 34389 35132
rect 34347 35083 34389 35092
rect 34251 34880 34293 34889
rect 34251 34840 34252 34880
rect 34292 34840 34293 34880
rect 34251 34831 34293 34840
rect 33964 34168 34100 34208
rect 34060 34040 34100 34168
rect 34348 34049 34388 35083
rect 34540 34376 34580 35167
rect 34636 35166 34676 35251
rect 34732 35216 34772 35335
rect 34732 35167 34772 35176
rect 35115 35048 35157 35057
rect 35115 35008 35116 35048
rect 35156 35008 35157 35048
rect 35115 34999 35157 35008
rect 35116 34914 35156 34999
rect 34636 34376 34676 34385
rect 34540 34336 34636 34376
rect 34636 34327 34676 34336
rect 35019 34376 35061 34385
rect 35019 34336 35020 34376
rect 35060 34336 35061 34376
rect 35019 34327 35061 34336
rect 34347 34040 34389 34049
rect 34060 34000 34292 34040
rect 33868 33823 33908 33832
rect 33772 33655 33812 33664
rect 33964 33704 34004 33713
rect 34156 33704 34196 33713
rect 34004 33664 34156 33704
rect 33964 33655 34004 33664
rect 34156 33655 34196 33664
rect 34252 33704 34292 34000
rect 34347 34000 34348 34040
rect 34388 34000 34389 34040
rect 34347 33991 34389 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 34348 33872 34388 33991
rect 34348 33832 34484 33872
rect 34252 33629 34292 33664
rect 34347 33704 34389 33713
rect 34347 33664 34348 33704
rect 34388 33664 34389 33704
rect 34347 33655 34389 33664
rect 34444 33704 34484 33832
rect 34444 33655 34484 33664
rect 33675 33620 33717 33629
rect 33675 33580 33676 33620
rect 33716 33580 33717 33620
rect 33675 33571 33717 33580
rect 33867 33620 33909 33629
rect 33867 33580 33868 33620
rect 33908 33580 33909 33620
rect 33867 33571 33909 33580
rect 34251 33620 34293 33629
rect 34251 33580 34252 33620
rect 34292 33580 34293 33620
rect 34251 33571 34293 33580
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 33484 32696 33524 32705
rect 33484 32201 33524 32656
rect 33772 32696 33812 32705
rect 33676 32276 33716 32285
rect 33772 32276 33812 32656
rect 33716 32236 33812 32276
rect 33676 32227 33716 32236
rect 33483 32192 33525 32201
rect 33483 32152 33484 32192
rect 33524 32152 33525 32192
rect 33483 32143 33525 32152
rect 33195 32108 33237 32117
rect 33195 32068 33196 32108
rect 33236 32068 33237 32108
rect 33195 32059 33237 32068
rect 33196 31604 33236 32059
rect 33484 32058 33524 32143
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 33196 31564 33428 31604
rect 32908 30556 33044 30596
rect 33100 31520 33140 31529
rect 32716 30428 32756 30437
rect 32716 30269 32756 30388
rect 32715 30260 32757 30269
rect 32715 30220 32716 30260
rect 32756 30220 32757 30260
rect 32715 30211 32757 30220
rect 32908 29840 32948 30556
rect 33003 30428 33045 30437
rect 33003 30388 33004 30428
rect 33044 30388 33045 30428
rect 33003 30379 33045 30388
rect 32331 29420 32373 29429
rect 32331 29380 32332 29420
rect 32372 29380 32373 29420
rect 32331 29371 32373 29380
rect 32908 29261 32948 29800
rect 32907 29252 32949 29261
rect 32907 29212 32908 29252
rect 32948 29212 32949 29252
rect 32907 29203 32949 29212
rect 32620 29168 32660 29177
rect 33004 29168 33044 30379
rect 33100 29849 33140 31480
rect 33291 31352 33333 31361
rect 33291 31312 33292 31352
rect 33332 31312 33333 31352
rect 33291 31303 33333 31312
rect 33388 31352 33428 31564
rect 33579 31520 33621 31529
rect 33579 31480 33580 31520
rect 33620 31480 33621 31520
rect 33579 31471 33621 31480
rect 33483 31436 33525 31445
rect 33483 31396 33484 31436
rect 33524 31396 33525 31436
rect 33483 31387 33525 31396
rect 33388 31303 33428 31312
rect 33292 31218 33332 31303
rect 33484 31268 33524 31387
rect 33580 31352 33620 31471
rect 33580 31303 33620 31312
rect 33868 31352 33908 33571
rect 34348 33570 34388 33655
rect 34636 33536 34676 33545
rect 35020 33536 35060 34327
rect 35212 34133 35252 35839
rect 35404 35393 35444 36436
rect 35596 36140 35636 36511
rect 35636 36100 35924 36140
rect 35596 36091 35636 36100
rect 35403 35384 35445 35393
rect 35403 35344 35404 35384
rect 35444 35344 35445 35384
rect 35403 35335 35445 35344
rect 35307 35300 35349 35309
rect 35307 35260 35308 35300
rect 35348 35260 35349 35300
rect 35307 35251 35349 35260
rect 35308 35216 35348 35251
rect 35788 35225 35828 35310
rect 35308 35165 35348 35176
rect 35403 35216 35445 35225
rect 35596 35216 35636 35225
rect 35403 35176 35404 35216
rect 35444 35176 35445 35216
rect 35403 35167 35445 35176
rect 35500 35176 35596 35216
rect 35404 35082 35444 35167
rect 35211 34124 35253 34133
rect 35211 34084 35212 34124
rect 35252 34084 35253 34124
rect 35211 34075 35253 34084
rect 35500 33965 35540 35176
rect 35596 35167 35636 35176
rect 35787 35216 35829 35225
rect 35787 35176 35788 35216
rect 35828 35176 35829 35216
rect 35787 35167 35829 35176
rect 35884 35216 35924 36100
rect 36076 35897 36116 36688
rect 39724 36688 40012 36728
rect 39148 36604 39476 36644
rect 36459 36560 36501 36569
rect 36459 36520 36460 36560
rect 36500 36520 36501 36560
rect 36459 36511 36501 36520
rect 37611 36560 37653 36569
rect 37611 36520 37612 36560
rect 37652 36520 37653 36560
rect 37611 36511 37653 36520
rect 39148 36560 39188 36604
rect 39148 36511 39188 36520
rect 36460 36426 36500 36511
rect 36075 35888 36117 35897
rect 36075 35848 36076 35888
rect 36116 35848 36117 35888
rect 36075 35839 36117 35848
rect 36748 35888 36788 35897
rect 37612 35888 37652 36511
rect 39340 36476 39380 36485
rect 39244 36436 39340 36476
rect 36788 35848 37076 35888
rect 36748 35839 36788 35848
rect 35980 35225 36020 35310
rect 36075 35300 36117 35309
rect 36075 35260 36076 35300
rect 36116 35260 36117 35300
rect 36075 35251 36117 35260
rect 35884 35167 35924 35176
rect 35979 35216 36021 35225
rect 35979 35176 35980 35216
rect 36020 35176 36021 35216
rect 35979 35167 36021 35176
rect 36076 35166 36116 35251
rect 36459 35216 36501 35225
rect 36459 35176 36460 35216
rect 36500 35176 36501 35216
rect 36459 35167 36501 35176
rect 36940 35216 36980 35227
rect 36363 35048 36405 35057
rect 36363 35008 36364 35048
rect 36404 35008 36405 35048
rect 36363 34999 36405 35008
rect 35596 34964 35636 34973
rect 36268 34964 36308 34973
rect 35636 34924 36020 34964
rect 35596 34915 35636 34924
rect 35980 34376 36020 34924
rect 35980 34327 36020 34336
rect 35787 34208 35829 34217
rect 35787 34168 35788 34208
rect 35828 34168 35829 34208
rect 35787 34159 35829 34168
rect 35788 34074 35828 34159
rect 35499 33956 35541 33965
rect 35499 33916 35500 33956
rect 35540 33916 35541 33956
rect 35499 33907 35541 33916
rect 34676 33496 35060 33536
rect 34636 33487 34676 33496
rect 36268 33116 36308 34924
rect 36364 34376 36404 34999
rect 36364 34327 36404 34336
rect 36363 33956 36405 33965
rect 36363 33916 36364 33956
rect 36404 33916 36405 33956
rect 36363 33907 36405 33916
rect 36364 33872 36404 33907
rect 36460 33881 36500 35167
rect 36940 35141 36980 35176
rect 36939 35132 36981 35141
rect 36939 35092 36940 35132
rect 36980 35092 36981 35132
rect 37036 35132 37076 35848
rect 37612 35839 37652 35848
rect 37996 35888 38036 35897
rect 38188 35888 38228 35897
rect 38860 35888 38900 35897
rect 38036 35848 38188 35888
rect 37996 35839 38036 35848
rect 38188 35839 38228 35848
rect 38476 35848 38860 35888
rect 37611 35384 37653 35393
rect 37611 35344 37612 35384
rect 37652 35344 37653 35384
rect 37611 35335 37653 35344
rect 38476 35384 38516 35848
rect 38860 35839 38900 35848
rect 39052 35888 39092 35897
rect 39244 35888 39284 36436
rect 39340 36427 39380 36436
rect 39092 35848 39284 35888
rect 39436 35888 39476 36604
rect 39052 35839 39092 35848
rect 39436 35839 39476 35848
rect 39147 35468 39189 35477
rect 39147 35428 39148 35468
rect 39188 35428 39189 35468
rect 39147 35419 39189 35428
rect 38476 35335 38516 35344
rect 37612 35250 37652 35335
rect 38283 35300 38325 35309
rect 38667 35300 38709 35309
rect 38283 35260 38284 35300
rect 38324 35260 38420 35300
rect 38283 35251 38325 35260
rect 38091 35216 38133 35225
rect 38091 35176 38092 35216
rect 38132 35176 38133 35216
rect 38091 35167 38133 35176
rect 38380 35216 38420 35260
rect 38667 35260 38668 35300
rect 38708 35260 38709 35300
rect 38667 35251 38709 35260
rect 39051 35300 39093 35309
rect 39051 35260 39052 35300
rect 39092 35260 39093 35300
rect 39051 35251 39093 35260
rect 38380 35167 38420 35176
rect 38572 35216 38612 35225
rect 37228 35132 37268 35141
rect 37036 35092 37228 35132
rect 36939 35083 36981 35092
rect 36940 34301 36980 35083
rect 37228 34376 37268 35092
rect 38092 35082 38132 35167
rect 38475 34544 38517 34553
rect 38475 34504 38476 34544
rect 38516 34504 38517 34544
rect 38475 34495 38517 34504
rect 37611 34460 37653 34469
rect 37611 34420 37612 34460
rect 37652 34420 37653 34460
rect 37611 34411 37653 34420
rect 36939 34292 36981 34301
rect 36939 34252 36940 34292
rect 36980 34252 36981 34292
rect 36939 34243 36981 34252
rect 36843 34208 36885 34217
rect 36843 34168 36844 34208
rect 36884 34168 36885 34208
rect 36843 34159 36885 34168
rect 36364 33821 36404 33832
rect 36459 33872 36501 33881
rect 36459 33832 36460 33872
rect 36500 33832 36501 33872
rect 36459 33823 36501 33832
rect 36460 33704 36500 33823
rect 36460 33655 36500 33664
rect 36556 33704 36596 33713
rect 36556 33545 36596 33664
rect 36651 33704 36693 33713
rect 36651 33664 36652 33704
rect 36692 33664 36693 33704
rect 36651 33655 36693 33664
rect 36844 33704 36884 34159
rect 36884 33664 37076 33704
rect 36844 33655 36884 33664
rect 36652 33570 36692 33655
rect 36555 33536 36597 33545
rect 36555 33496 36556 33536
rect 36596 33496 36597 33536
rect 36555 33487 36597 33496
rect 36172 33076 36308 33116
rect 34636 33032 34676 33041
rect 34348 32992 34636 33032
rect 34060 32192 34100 32201
rect 34348 32192 34388 32992
rect 34636 32983 34676 32992
rect 34100 32152 34388 32192
rect 34444 32864 34484 32873
rect 34060 32143 34100 32152
rect 34444 31529 34484 32824
rect 36076 32864 36116 32873
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 36076 32369 36116 32824
rect 36075 32360 36117 32369
rect 36075 32320 36076 32360
rect 36116 32320 36117 32360
rect 36075 32311 36117 32320
rect 36076 32226 36116 32311
rect 34923 32192 34965 32201
rect 34923 32152 34924 32192
rect 34964 32152 34965 32192
rect 34923 32143 34965 32152
rect 34924 32058 34964 32143
rect 34443 31520 34485 31529
rect 34156 31480 34388 31520
rect 33484 31219 33524 31228
rect 33868 31193 33908 31312
rect 33963 31352 34005 31361
rect 33963 31312 33964 31352
rect 34004 31312 34005 31352
rect 33963 31303 34005 31312
rect 34060 31352 34100 31361
rect 34156 31352 34196 31480
rect 34100 31312 34196 31352
rect 34252 31352 34292 31361
rect 33964 31218 34004 31303
rect 33772 31184 33812 31193
rect 33580 30428 33620 30437
rect 33196 30388 33580 30428
rect 33099 29840 33141 29849
rect 33099 29800 33100 29840
rect 33140 29800 33141 29840
rect 33099 29791 33141 29800
rect 33196 29840 33236 30388
rect 33580 30379 33620 30388
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 33772 30092 33812 31144
rect 33867 31184 33909 31193
rect 33867 31144 33868 31184
rect 33908 31144 33909 31184
rect 33867 31135 33909 31144
rect 33867 30680 33909 30689
rect 33867 30640 33868 30680
rect 33908 30640 33909 30680
rect 33867 30631 33909 30640
rect 33196 29791 33236 29800
rect 33484 30052 33812 30092
rect 33196 29345 33236 29430
rect 33195 29336 33237 29345
rect 33195 29296 33196 29336
rect 33236 29296 33237 29336
rect 33195 29287 33237 29296
rect 33292 29168 33332 29177
rect 33004 29128 33292 29168
rect 32620 28589 32660 29128
rect 33292 29119 33332 29128
rect 33484 29168 33524 30052
rect 33579 29840 33621 29849
rect 33579 29800 33580 29840
rect 33620 29800 33621 29840
rect 33579 29791 33621 29800
rect 33580 29706 33620 29791
rect 33580 29336 33620 29345
rect 33868 29336 33908 30631
rect 34060 30101 34100 31312
rect 34252 31025 34292 31312
rect 34348 31352 34388 31480
rect 34443 31480 34444 31520
rect 34484 31480 34485 31520
rect 34443 31471 34485 31480
rect 34540 31520 34580 31529
rect 34580 31480 35060 31520
rect 34540 31471 34580 31480
rect 34540 31352 34580 31361
rect 34348 31303 34388 31312
rect 34444 31312 34540 31352
rect 34251 31016 34293 31025
rect 34251 30976 34252 31016
rect 34292 30976 34293 31016
rect 34251 30967 34293 30976
rect 34444 30689 34484 31312
rect 34540 31303 34580 31312
rect 35020 31352 35060 31480
rect 35020 31303 35060 31312
rect 35115 31352 35157 31361
rect 35404 31352 35444 31361
rect 35115 31312 35116 31352
rect 35156 31312 35157 31352
rect 35115 31303 35157 31312
rect 35308 31312 35404 31352
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 34251 30680 34293 30689
rect 34251 30640 34252 30680
rect 34292 30640 34293 30680
rect 34251 30631 34293 30640
rect 34443 30680 34485 30689
rect 34443 30640 34444 30680
rect 34484 30640 34485 30680
rect 34443 30631 34485 30640
rect 35116 30680 35156 31303
rect 35308 30932 35348 31312
rect 35404 31303 35444 31312
rect 35403 31184 35445 31193
rect 35403 31144 35404 31184
rect 35444 31144 35445 31184
rect 35403 31135 35445 31144
rect 34252 30546 34292 30631
rect 34347 30596 34389 30605
rect 34347 30556 34348 30596
rect 34388 30556 34389 30596
rect 34347 30547 34389 30556
rect 34059 30092 34101 30101
rect 34059 30052 34060 30092
rect 34100 30052 34101 30092
rect 34059 30043 34101 30052
rect 33620 29296 33908 29336
rect 33580 29287 33620 29296
rect 33963 29252 34005 29261
rect 33963 29212 33964 29252
rect 34004 29212 34005 29252
rect 33963 29203 34005 29212
rect 33484 29119 33524 29128
rect 33676 29168 33716 29179
rect 33676 29093 33716 29128
rect 33771 29168 33813 29177
rect 33771 29128 33772 29168
rect 33812 29128 33813 29168
rect 33771 29119 33813 29128
rect 33964 29168 34004 29203
rect 33675 29084 33717 29093
rect 33675 29044 33676 29084
rect 33716 29044 33717 29084
rect 33675 29035 33717 29044
rect 33772 29034 33812 29119
rect 33964 29117 34004 29128
rect 34251 29168 34293 29177
rect 34251 29128 34252 29168
rect 34292 29128 34293 29168
rect 34251 29119 34293 29128
rect 33004 29000 33044 29009
rect 32427 28580 32469 28589
rect 32427 28540 32428 28580
rect 32468 28540 32469 28580
rect 32427 28531 32469 28540
rect 32619 28580 32661 28589
rect 32619 28540 32620 28580
rect 32660 28540 32661 28580
rect 32619 28531 32661 28540
rect 32236 28279 32276 28288
rect 32139 27824 32181 27833
rect 32139 27784 32140 27824
rect 32180 27784 32181 27824
rect 32139 27775 32181 27784
rect 32151 27669 32191 27678
rect 31564 27607 31604 27616
rect 31660 27656 31700 27665
rect 31467 27488 31509 27497
rect 31467 27448 31468 27488
rect 31508 27448 31509 27488
rect 31467 27439 31509 27448
rect 31371 27236 31413 27245
rect 31180 26767 31220 26776
rect 31276 27196 31372 27236
rect 31412 27196 31413 27236
rect 30892 26682 30932 26767
rect 30988 26648 31028 26657
rect 31028 26608 31124 26648
rect 30988 26599 31028 26608
rect 30892 26144 30932 26153
rect 31084 26144 31124 26608
rect 31179 26396 31221 26405
rect 31179 26356 31180 26396
rect 31220 26356 31221 26396
rect 31179 26347 31221 26356
rect 30892 25649 30932 26104
rect 30988 26109 31028 26118
rect 31084 26095 31124 26104
rect 30988 25985 31028 26069
rect 30987 25976 31029 25985
rect 30987 25936 30988 25976
rect 31028 25936 31029 25976
rect 30987 25927 31029 25936
rect 30891 25640 30933 25649
rect 30891 25600 30892 25640
rect 30932 25600 30933 25640
rect 30891 25591 30933 25600
rect 30795 25556 30837 25565
rect 30795 25516 30796 25556
rect 30836 25516 30837 25556
rect 30795 25507 30837 25516
rect 31180 25304 31220 26347
rect 31276 25976 31316 27196
rect 31371 27187 31413 27196
rect 31372 27068 31412 27077
rect 31660 27068 31700 27616
rect 31755 27656 31797 27665
rect 31948 27656 31988 27665
rect 31755 27616 31756 27656
rect 31796 27616 31797 27656
rect 31755 27607 31797 27616
rect 31852 27616 31948 27656
rect 32191 27629 32372 27656
rect 32151 27616 32372 27629
rect 31756 27522 31796 27607
rect 31412 27028 31700 27068
rect 31755 27068 31797 27077
rect 31755 27028 31756 27068
rect 31796 27028 31797 27068
rect 31372 27019 31412 27028
rect 31755 27019 31797 27028
rect 31852 27068 31892 27616
rect 31948 27607 31988 27616
rect 32044 27488 32084 27497
rect 31947 27448 32044 27488
rect 31947 27404 31987 27448
rect 32044 27439 32084 27448
rect 31947 27364 31988 27404
rect 31852 27019 31892 27028
rect 31372 26909 31412 26940
rect 31371 26900 31413 26909
rect 31371 26860 31372 26900
rect 31412 26860 31413 26900
rect 31371 26851 31413 26860
rect 31372 26816 31412 26851
rect 31372 26153 31412 26776
rect 31564 26816 31604 26825
rect 31564 26489 31604 26776
rect 31660 26816 31700 26825
rect 31756 26816 31796 27019
rect 31948 26825 31988 27364
rect 32139 26900 32181 26909
rect 32139 26860 32140 26900
rect 32180 26860 32181 26900
rect 32139 26851 32181 26860
rect 31700 26776 31796 26816
rect 31947 26816 31989 26825
rect 31947 26776 31948 26816
rect 31988 26776 31989 26816
rect 31660 26767 31700 26776
rect 31947 26767 31989 26776
rect 32140 26816 32180 26851
rect 32140 26765 32180 26776
rect 32235 26816 32277 26825
rect 32235 26776 32236 26816
rect 32276 26776 32277 26816
rect 32235 26767 32277 26776
rect 32236 26682 32276 26767
rect 31563 26480 31605 26489
rect 31563 26440 31564 26480
rect 31604 26440 31605 26480
rect 31563 26431 31605 26440
rect 31755 26480 31797 26489
rect 31755 26440 31756 26480
rect 31796 26440 31797 26480
rect 31755 26431 31797 26440
rect 31756 26312 31796 26431
rect 32332 26321 32372 27616
rect 32428 26909 32468 28531
rect 33004 28328 33044 28960
rect 33099 29000 33141 29009
rect 33099 28960 33100 29000
rect 33140 28960 33236 29000
rect 33099 28951 33141 28960
rect 33100 28328 33140 28337
rect 33004 28288 33100 28328
rect 33196 28328 33236 28960
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 34252 28580 34292 29119
rect 34252 28531 34292 28540
rect 33484 28328 33524 28337
rect 33196 28288 33484 28328
rect 33100 28279 33140 28288
rect 33484 28279 33524 28288
rect 34348 28328 34388 30547
rect 34444 30437 34484 30522
rect 34443 30428 34485 30437
rect 34443 30388 34444 30428
rect 34484 30388 34485 30428
rect 34443 30379 34485 30388
rect 35116 30269 35156 30640
rect 35212 30892 35348 30932
rect 35212 30512 35252 30892
rect 35308 30689 35348 30774
rect 35307 30680 35349 30689
rect 35307 30640 35308 30680
rect 35348 30640 35349 30680
rect 35307 30631 35349 30640
rect 35404 30680 35444 31135
rect 35404 30631 35444 30640
rect 35500 30680 35540 30691
rect 35500 30605 35540 30640
rect 35596 30680 35636 30689
rect 35636 30640 35732 30680
rect 35596 30631 35636 30640
rect 35499 30596 35541 30605
rect 35499 30556 35500 30596
rect 35540 30556 35541 30596
rect 35499 30547 35541 30556
rect 35212 30472 35444 30512
rect 35115 30260 35157 30269
rect 35115 30220 35116 30260
rect 35156 30220 35157 30260
rect 35115 30211 35157 30220
rect 34443 30176 34485 30185
rect 34443 30136 34444 30176
rect 34484 30136 34485 30176
rect 34443 30127 34485 30136
rect 34444 29840 34484 30127
rect 34444 29791 34484 29800
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 34828 29168 34868 29177
rect 34828 29000 34868 29128
rect 34348 28279 34388 28288
rect 34444 28960 34868 29000
rect 35404 29000 35444 30472
rect 35595 30260 35637 30269
rect 35595 30220 35596 30260
rect 35636 30220 35637 30260
rect 35595 30211 35637 30220
rect 35596 30092 35636 30211
rect 35692 30101 35732 30640
rect 35979 30596 36021 30605
rect 35979 30556 35980 30596
rect 36020 30556 36021 30596
rect 35979 30547 36021 30556
rect 35980 30462 36020 30547
rect 36172 30521 36212 33076
rect 36940 33032 36980 33041
rect 36267 32948 36309 32957
rect 36267 32908 36268 32948
rect 36308 32908 36309 32948
rect 36267 32899 36309 32908
rect 36268 32201 36308 32899
rect 36748 32696 36788 32705
rect 36267 32192 36309 32201
rect 36267 32152 36268 32192
rect 36308 32152 36309 32192
rect 36267 32143 36309 32152
rect 36652 32192 36692 32201
rect 36748 32192 36788 32656
rect 36692 32152 36788 32192
rect 36652 32143 36692 32152
rect 36268 31352 36308 32143
rect 36268 31303 36308 31312
rect 36556 31940 36596 31949
rect 36171 30512 36213 30521
rect 36171 30472 36172 30512
rect 36212 30472 36213 30512
rect 36171 30463 36213 30472
rect 35883 30260 35925 30269
rect 35883 30220 35884 30260
rect 35924 30220 35925 30260
rect 35883 30211 35925 30220
rect 35596 30043 35636 30052
rect 35691 30092 35733 30101
rect 35691 30052 35692 30092
rect 35732 30052 35733 30092
rect 35691 30043 35733 30052
rect 35596 29093 35636 29095
rect 35595 29084 35637 29093
rect 35692 29084 35732 30043
rect 35787 29252 35829 29261
rect 35787 29212 35788 29252
rect 35828 29212 35829 29252
rect 35787 29203 35829 29212
rect 35595 29044 35596 29084
rect 35636 29044 35732 29084
rect 35788 29084 35828 29203
rect 35595 29035 35637 29044
rect 35788 29035 35828 29044
rect 34444 27824 34484 28960
rect 35404 28951 35444 28960
rect 35596 29000 35636 29035
rect 35596 28951 35636 28960
rect 35884 28832 35924 30211
rect 36268 30101 36308 30186
rect 36267 30092 36309 30101
rect 36267 30052 36268 30092
rect 36308 30052 36309 30092
rect 36267 30043 36309 30052
rect 35979 29924 36021 29933
rect 35979 29884 35980 29924
rect 36020 29884 36021 29924
rect 35979 29875 36021 29884
rect 35980 29840 36020 29875
rect 36268 29849 36308 29934
rect 36556 29933 36596 31900
rect 36651 30680 36693 30689
rect 36651 30640 36652 30680
rect 36692 30640 36693 30680
rect 36651 30631 36693 30640
rect 36652 30546 36692 30631
rect 36555 29924 36597 29933
rect 36555 29884 36556 29924
rect 36596 29884 36597 29924
rect 36555 29875 36597 29884
rect 35980 29789 36020 29800
rect 36076 29840 36116 29849
rect 35979 29672 36021 29681
rect 35979 29632 35980 29672
rect 36020 29632 36021 29672
rect 35979 29623 36021 29632
rect 35980 29252 36020 29623
rect 35980 29203 36020 29212
rect 36076 29093 36116 29800
rect 36267 29840 36309 29849
rect 36267 29800 36268 29840
rect 36308 29800 36309 29840
rect 36267 29791 36309 29800
rect 36459 29672 36501 29681
rect 36459 29632 36460 29672
rect 36500 29632 36501 29672
rect 36459 29623 36501 29632
rect 36460 29538 36500 29623
rect 36364 29168 36404 29177
rect 36075 29084 36117 29093
rect 36075 29044 36076 29084
rect 36116 29044 36117 29084
rect 36075 29035 36117 29044
rect 36364 29000 36404 29128
rect 36364 28960 36500 29000
rect 35884 28792 36212 28832
rect 35308 28496 35348 28505
rect 35211 28244 35253 28253
rect 35211 28204 35212 28244
rect 35252 28204 35253 28244
rect 35211 28195 35253 28204
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 34444 27784 34580 27824
rect 32811 27656 32853 27665
rect 32811 27616 32812 27656
rect 32852 27616 32853 27656
rect 32811 27607 32853 27616
rect 33291 27656 33333 27665
rect 33291 27616 33292 27656
rect 33332 27616 33333 27656
rect 33291 27607 33333 27616
rect 33963 27656 34005 27665
rect 33963 27616 33964 27656
rect 34004 27616 34005 27656
rect 33963 27607 34005 27616
rect 34156 27656 34196 27665
rect 32523 27236 32565 27245
rect 32523 27196 32524 27236
rect 32564 27196 32565 27236
rect 32523 27187 32565 27196
rect 32427 26900 32469 26909
rect 32427 26860 32428 26900
rect 32468 26860 32469 26900
rect 32427 26851 32469 26860
rect 32524 26816 32564 27187
rect 32812 27068 32852 27607
rect 33292 27522 33332 27607
rect 33099 27488 33141 27497
rect 33099 27448 33100 27488
rect 33140 27448 33141 27488
rect 33099 27439 33141 27448
rect 33100 27354 33140 27439
rect 33964 27404 34004 27607
rect 33772 27364 33964 27404
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 32812 26825 32852 27028
rect 32524 26741 32564 26776
rect 32811 26816 32853 26825
rect 32811 26776 32812 26816
rect 32852 26776 32853 26816
rect 32811 26767 32853 26776
rect 32523 26732 32565 26741
rect 32523 26692 32524 26732
rect 32564 26692 32565 26732
rect 32523 26683 32565 26692
rect 32524 26652 32564 26683
rect 31756 26263 31796 26272
rect 32331 26312 32373 26321
rect 32331 26272 32332 26312
rect 32372 26272 32373 26312
rect 32331 26263 32373 26272
rect 31371 26144 31413 26153
rect 32140 26144 32180 26153
rect 31371 26104 31372 26144
rect 31412 26104 31413 26144
rect 31371 26095 31413 26104
rect 31756 26104 32140 26144
rect 31276 25936 31508 25976
rect 31275 25556 31317 25565
rect 31275 25516 31276 25556
rect 31316 25516 31317 25556
rect 31275 25507 31317 25516
rect 31180 25229 31220 25264
rect 31179 25220 31221 25229
rect 31179 25180 31180 25220
rect 31220 25180 31221 25220
rect 31179 25171 31221 25180
rect 31180 25140 31220 25171
rect 30795 23792 30837 23801
rect 30795 23752 30796 23792
rect 30836 23752 30837 23792
rect 30795 23743 30837 23752
rect 31084 23792 31124 23801
rect 30796 23658 30836 23743
rect 30892 23624 30932 23633
rect 31084 23624 31124 23752
rect 30932 23584 31124 23624
rect 30892 23575 30932 23584
rect 30699 23372 30741 23381
rect 30699 23332 30700 23372
rect 30740 23332 30741 23372
rect 30699 23323 30741 23332
rect 30891 23372 30933 23381
rect 30891 23332 30892 23372
rect 30932 23332 30933 23372
rect 30891 23323 30933 23332
rect 30892 23288 30932 23323
rect 30892 23237 30932 23248
rect 31084 23129 31124 23584
rect 31180 23792 31220 23801
rect 31180 23213 31220 23752
rect 31276 23792 31316 25507
rect 31468 23801 31508 25936
rect 31659 25556 31701 25565
rect 31659 25516 31660 25556
rect 31700 25516 31701 25556
rect 31659 25507 31701 25516
rect 31660 25422 31700 25507
rect 31756 24800 31796 26104
rect 32140 26095 32180 26104
rect 32332 25817 32372 26263
rect 33676 26144 33716 26153
rect 33772 26144 33812 27364
rect 33964 27355 34004 27364
rect 33867 27236 33909 27245
rect 33867 27196 33868 27236
rect 33908 27196 33909 27236
rect 33867 27187 33909 27196
rect 33716 26104 33812 26144
rect 33868 26159 33908 27187
rect 33964 26816 34004 26825
rect 33964 26312 34004 26776
rect 33964 26272 34100 26312
rect 33868 26110 33908 26119
rect 33964 26144 34004 26153
rect 33676 26095 33716 26104
rect 33964 26060 34004 26104
rect 33877 26020 34004 26060
rect 33580 25901 33620 25986
rect 33877 25976 33917 26020
rect 34060 25976 34100 26272
rect 34156 26144 34196 27616
rect 34156 26095 34196 26104
rect 34252 27656 34292 27665
rect 33868 25936 33917 25976
rect 33964 25936 34100 25976
rect 34155 25976 34197 25985
rect 34155 25936 34156 25976
rect 34196 25936 34197 25976
rect 32715 25892 32757 25901
rect 32715 25852 32716 25892
rect 32756 25852 32757 25892
rect 32715 25843 32757 25852
rect 33579 25892 33621 25901
rect 33579 25852 33580 25892
rect 33620 25852 33621 25892
rect 33579 25843 33621 25852
rect 32331 25808 32373 25817
rect 32331 25768 32332 25808
rect 32372 25768 32373 25808
rect 32331 25759 32373 25768
rect 32523 25472 32565 25481
rect 32523 25432 32524 25472
rect 32564 25432 32565 25472
rect 32523 25423 32565 25432
rect 32524 25338 32564 25423
rect 32716 25304 32756 25843
rect 33868 25733 33908 25936
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 33867 25724 33909 25733
rect 33867 25684 33868 25724
rect 33908 25684 33909 25724
rect 33867 25675 33909 25684
rect 32811 25472 32853 25481
rect 32811 25432 32812 25472
rect 32852 25432 32853 25472
rect 32811 25423 32853 25432
rect 33004 25472 33044 25481
rect 33044 25432 33908 25472
rect 33004 25423 33044 25432
rect 32716 25255 32756 25264
rect 32812 25304 32852 25423
rect 32812 25255 32852 25264
rect 33003 25304 33045 25313
rect 33003 25264 33004 25304
rect 33044 25264 33045 25304
rect 33003 25255 33045 25264
rect 33868 25304 33908 25432
rect 33868 25255 33908 25264
rect 32427 25220 32469 25229
rect 32427 25180 32428 25220
rect 32468 25180 32469 25220
rect 32427 25171 32469 25180
rect 31756 24751 31796 24760
rect 32428 23960 32468 25171
rect 33004 25170 33044 25255
rect 33291 25220 33333 25229
rect 33291 25180 33292 25220
rect 33332 25180 33333 25220
rect 33291 25171 33333 25180
rect 33196 25136 33236 25145
rect 33100 25096 33196 25136
rect 33100 24884 33140 25096
rect 33196 25087 33236 25096
rect 32812 24844 33140 24884
rect 32812 24716 32852 24844
rect 32812 24667 32852 24676
rect 33196 24632 33236 24641
rect 33292 24632 33332 25171
rect 33964 24641 34004 25936
rect 34155 25927 34197 25936
rect 34156 25842 34196 25927
rect 34252 25724 34292 27616
rect 34347 27656 34389 27665
rect 34347 27616 34348 27656
rect 34388 27616 34389 27656
rect 34347 27607 34389 27616
rect 34444 27656 34484 27665
rect 34348 27522 34388 27607
rect 34444 26825 34484 27616
rect 34443 26816 34485 26825
rect 34348 26776 34444 26816
rect 34484 26776 34485 26816
rect 34348 25733 34388 26776
rect 34443 26767 34485 26776
rect 34540 26648 34580 27784
rect 35212 27665 35252 28195
rect 35019 27656 35061 27665
rect 35019 27616 35020 27656
rect 35060 27616 35061 27656
rect 35019 27607 35061 27616
rect 35211 27656 35253 27665
rect 35211 27616 35212 27656
rect 35252 27616 35253 27656
rect 35211 27607 35253 27616
rect 34827 27488 34869 27497
rect 34827 27448 34828 27488
rect 34868 27448 34869 27488
rect 34827 27439 34869 27448
rect 34828 26816 34868 27439
rect 34828 26767 34868 26776
rect 34444 26608 34580 26648
rect 34156 25684 34292 25724
rect 34347 25724 34389 25733
rect 34347 25684 34348 25724
rect 34388 25684 34389 25724
rect 34059 25304 34101 25313
rect 34059 25264 34060 25304
rect 34100 25264 34101 25304
rect 34059 25255 34101 25264
rect 34156 25304 34196 25684
rect 34347 25675 34389 25684
rect 34348 25481 34388 25675
rect 34347 25472 34389 25481
rect 34347 25432 34348 25472
rect 34388 25432 34389 25472
rect 34347 25423 34389 25432
rect 34060 25170 34100 25255
rect 34156 25229 34196 25264
rect 34251 25304 34293 25313
rect 34251 25264 34252 25304
rect 34292 25264 34293 25304
rect 34251 25255 34293 25264
rect 34348 25304 34388 25423
rect 34155 25220 34197 25229
rect 34155 25180 34156 25220
rect 34196 25180 34197 25220
rect 34155 25171 34197 25180
rect 34156 25140 34196 25171
rect 34252 25170 34292 25255
rect 34348 25229 34388 25264
rect 34347 25220 34389 25229
rect 34347 25180 34348 25220
rect 34388 25180 34389 25220
rect 34347 25171 34389 25180
rect 34155 25052 34197 25061
rect 34348 25052 34388 25171
rect 34155 25012 34156 25052
rect 34196 25012 34197 25052
rect 34155 25003 34197 25012
rect 34252 25012 34388 25052
rect 33236 24592 33332 24632
rect 33963 24632 34005 24641
rect 34060 24632 34100 24641
rect 33963 24592 33964 24632
rect 34004 24592 34060 24632
rect 33196 24583 33236 24592
rect 33963 24583 34005 24592
rect 34060 24583 34100 24592
rect 33964 24498 34004 24583
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 32428 23911 32468 23920
rect 31179 23204 31221 23213
rect 31179 23164 31180 23204
rect 31220 23164 31221 23204
rect 31179 23155 31221 23164
rect 30795 23120 30837 23129
rect 30795 23080 30796 23120
rect 30836 23080 30837 23120
rect 30795 23071 30837 23080
rect 31083 23120 31125 23129
rect 31083 23080 31084 23120
rect 31124 23080 31125 23120
rect 31083 23071 31125 23080
rect 30700 22532 30740 22541
rect 30604 22492 30700 22532
rect 30700 22483 30740 22492
rect 30604 21776 30644 21785
rect 30796 21776 30836 23071
rect 31180 22289 31220 23155
rect 31276 23045 31316 23752
rect 31467 23792 31509 23801
rect 31467 23752 31468 23792
rect 31508 23752 31509 23792
rect 31467 23743 31509 23752
rect 33100 23792 33140 23801
rect 33484 23792 33524 23801
rect 33140 23752 33484 23792
rect 33100 23743 33140 23752
rect 31372 23624 31412 23633
rect 31412 23584 31604 23624
rect 31372 23575 31412 23584
rect 31564 23120 31604 23584
rect 31851 23204 31893 23213
rect 31851 23164 31852 23204
rect 31892 23164 31893 23204
rect 31851 23155 31893 23164
rect 31564 23071 31604 23080
rect 31755 23120 31797 23129
rect 31755 23080 31756 23120
rect 31796 23080 31797 23120
rect 31755 23071 31797 23080
rect 31852 23120 31892 23155
rect 31275 23036 31317 23045
rect 31275 22996 31276 23036
rect 31316 22996 31317 23036
rect 31275 22987 31317 22996
rect 31756 22986 31796 23071
rect 31852 23069 31892 23080
rect 32908 23120 32948 23129
rect 32044 22952 32084 22961
rect 31564 22868 31604 22877
rect 31179 22280 31221 22289
rect 31179 22240 31180 22280
rect 31220 22240 31221 22280
rect 31179 22231 31221 22240
rect 31564 22280 31604 22828
rect 31564 22231 31604 22240
rect 31948 22280 31988 22289
rect 32044 22280 32084 22912
rect 32908 22541 32948 23080
rect 33484 22868 33524 23752
rect 33580 23120 33620 23129
rect 33868 23120 33908 23129
rect 33620 23080 33868 23120
rect 33580 23071 33620 23080
rect 33868 23071 33908 23080
rect 34156 22952 34196 25003
rect 34252 22961 34292 25012
rect 34347 23876 34389 23885
rect 34347 23836 34348 23876
rect 34388 23836 34389 23876
rect 34347 23827 34389 23836
rect 34444 23876 34484 26608
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34539 25640 34581 25649
rect 35020 25640 35060 27607
rect 35212 27522 35252 27607
rect 35308 27581 35348 28456
rect 35692 28328 35732 28337
rect 35596 28244 35636 28253
rect 35500 28204 35596 28244
rect 35307 27572 35349 27581
rect 35307 27532 35308 27572
rect 35348 27532 35349 27572
rect 35307 27523 35349 27532
rect 35500 26984 35540 28204
rect 35596 28195 35636 28204
rect 35692 27833 35732 28288
rect 35980 28328 36020 28337
rect 36172 28328 36212 28792
rect 36460 28496 36500 28960
rect 36460 28447 36500 28456
rect 36020 28288 36116 28328
rect 36172 28288 36500 28328
rect 35980 28279 36020 28288
rect 35691 27824 35733 27833
rect 35691 27784 35692 27824
rect 35732 27784 35733 27824
rect 35691 27775 35733 27784
rect 36076 27656 36116 28288
rect 36363 27740 36405 27749
rect 36363 27700 36364 27740
rect 36404 27700 36405 27740
rect 36363 27691 36405 27700
rect 36268 27656 36308 27665
rect 36116 27616 36268 27656
rect 36076 27607 36116 27616
rect 35595 27404 35637 27413
rect 35595 27364 35596 27404
rect 35636 27364 35637 27404
rect 35595 27355 35637 27364
rect 35308 26944 35540 26984
rect 35212 26732 35252 26741
rect 35212 25985 35252 26692
rect 35211 25976 35253 25985
rect 35211 25936 35212 25976
rect 35252 25936 35253 25976
rect 35211 25927 35253 25936
rect 34539 25600 34540 25640
rect 34580 25600 34581 25640
rect 34539 25591 34581 25600
rect 34636 25600 35060 25640
rect 34540 25481 34580 25591
rect 34539 25472 34581 25481
rect 34539 25432 34540 25472
rect 34580 25432 34581 25472
rect 34539 25423 34581 25432
rect 34636 25145 34676 25600
rect 34923 25472 34965 25481
rect 34923 25432 34924 25472
rect 34964 25432 34965 25472
rect 34923 25423 34965 25432
rect 35115 25472 35157 25481
rect 35115 25432 35116 25472
rect 35156 25432 35157 25472
rect 35115 25423 35157 25432
rect 34827 25388 34869 25397
rect 34827 25348 34828 25388
rect 34868 25348 34869 25388
rect 34827 25339 34869 25348
rect 34732 25304 34772 25315
rect 34732 25229 34772 25264
rect 34828 25304 34868 25339
rect 34828 25253 34868 25264
rect 34924 25304 34964 25423
rect 34924 25255 34964 25264
rect 34731 25220 34773 25229
rect 34731 25180 34732 25220
rect 34772 25180 34773 25220
rect 34731 25171 34773 25180
rect 35019 25220 35061 25229
rect 35019 25180 35020 25220
rect 35060 25180 35061 25220
rect 35019 25171 35061 25180
rect 34635 25136 34677 25145
rect 34635 25096 34636 25136
rect 34676 25096 34677 25136
rect 34635 25087 34677 25096
rect 35020 25086 35060 25171
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 35116 23960 35156 25423
rect 35308 25397 35348 26944
rect 35500 26816 35540 26825
rect 35403 26648 35445 26657
rect 35403 26608 35404 26648
rect 35444 26608 35445 26648
rect 35403 26599 35445 26608
rect 35404 26514 35444 26599
rect 35500 25481 35540 26776
rect 35596 26816 35636 27355
rect 36172 26825 36212 26910
rect 36268 26909 36308 27616
rect 36364 27606 36404 27691
rect 36460 27656 36500 28288
rect 36940 27656 36980 32992
rect 37036 32780 37076 33664
rect 37228 32957 37268 34336
rect 37323 34040 37365 34049
rect 37323 34000 37324 34040
rect 37364 34000 37365 34040
rect 37323 33991 37365 34000
rect 37227 32948 37269 32957
rect 37227 32908 37228 32948
rect 37268 32908 37269 32948
rect 37227 32899 37269 32908
rect 37324 32864 37364 33991
rect 37515 33620 37557 33629
rect 37515 33580 37516 33620
rect 37556 33580 37557 33620
rect 37515 33571 37557 33580
rect 37324 32815 37364 32824
rect 37228 32780 37268 32789
rect 37036 32740 37228 32780
rect 37228 32731 37268 32740
rect 37516 32192 37556 33571
rect 37612 32864 37652 34411
rect 38380 34208 38420 34217
rect 38380 34049 38420 34168
rect 38379 34040 38421 34049
rect 38379 34000 38380 34040
rect 38420 34000 38421 34040
rect 38379 33991 38421 34000
rect 37996 33704 38036 33713
rect 37612 32369 37652 32824
rect 37708 33664 37996 33704
rect 37611 32360 37653 32369
rect 37611 32320 37612 32360
rect 37652 32320 37653 32360
rect 37611 32311 37653 32320
rect 37708 32360 37748 33664
rect 37996 33655 38036 33664
rect 38092 33704 38132 33715
rect 38092 33629 38132 33664
rect 38284 33704 38324 33713
rect 38476 33704 38516 34495
rect 38572 34217 38612 35176
rect 38668 35216 38708 35251
rect 38668 35165 38708 35176
rect 39052 35166 39092 35251
rect 39148 35216 39188 35419
rect 39724 35384 39764 36688
rect 40012 36679 40052 36688
rect 41068 36728 41108 36737
rect 40396 36476 40436 36485
rect 40300 35888 40340 35897
rect 40300 35393 40340 35848
rect 40396 35477 40436 36436
rect 40395 35468 40437 35477
rect 40395 35428 40396 35468
rect 40436 35428 40437 35468
rect 40395 35419 40437 35428
rect 39436 35344 39764 35384
rect 40299 35384 40341 35393
rect 40299 35344 40300 35384
rect 40340 35344 40341 35384
rect 39436 35300 39476 35344
rect 40299 35335 40341 35344
rect 39436 35251 39476 35260
rect 39340 35216 39380 35225
rect 39148 35167 39188 35176
rect 39244 35176 39340 35216
rect 38955 35132 38997 35141
rect 38955 35092 38956 35132
rect 38996 35092 38997 35132
rect 38955 35083 38997 35092
rect 38860 34376 38900 34385
rect 38860 34217 38900 34336
rect 38956 34376 38996 35083
rect 39051 34628 39093 34637
rect 39051 34588 39052 34628
rect 39092 34588 39093 34628
rect 39051 34579 39093 34588
rect 38956 34327 38996 34336
rect 39052 34376 39092 34579
rect 39052 34327 39092 34336
rect 39148 34376 39188 34385
rect 39244 34376 39284 35176
rect 39340 35167 39380 35176
rect 39532 35216 39572 35225
rect 39532 34880 39572 35176
rect 39188 34336 39284 34376
rect 39340 34840 39572 34880
rect 39628 35216 39668 35225
rect 39340 34376 39380 34840
rect 39435 34712 39477 34721
rect 39435 34672 39436 34712
rect 39476 34672 39477 34712
rect 39435 34663 39477 34672
rect 39148 34327 39188 34336
rect 39340 34217 39380 34336
rect 39436 34376 39476 34663
rect 39531 34628 39573 34637
rect 39531 34588 39532 34628
rect 39572 34588 39573 34628
rect 39531 34579 39573 34588
rect 39436 34301 39476 34336
rect 39532 34376 39572 34579
rect 39628 34553 39668 35176
rect 40108 35216 40148 35225
rect 40108 34712 40148 35176
rect 40300 35216 40340 35227
rect 40300 35141 40340 35176
rect 40876 35216 40916 35225
rect 40299 35132 40341 35141
rect 40299 35092 40300 35132
rect 40340 35092 40341 35132
rect 40299 35083 40341 35092
rect 40683 35048 40725 35057
rect 40683 35008 40684 35048
rect 40724 35008 40725 35048
rect 40683 34999 40725 35008
rect 40204 34964 40244 34973
rect 40244 34924 40436 34964
rect 40204 34915 40244 34924
rect 40108 34672 40244 34712
rect 39627 34544 39669 34553
rect 39627 34504 39628 34544
rect 39668 34504 39669 34544
rect 39627 34495 39669 34504
rect 40107 34460 40149 34469
rect 40107 34420 40108 34460
rect 40148 34420 40149 34460
rect 40107 34411 40149 34420
rect 39435 34292 39477 34301
rect 39435 34252 39436 34292
rect 39476 34252 39477 34292
rect 39435 34243 39477 34252
rect 38571 34208 38613 34217
rect 38571 34168 38572 34208
rect 38612 34168 38613 34208
rect 38571 34159 38613 34168
rect 38859 34208 38901 34217
rect 38859 34168 38860 34208
rect 38900 34168 38901 34208
rect 38859 34159 38901 34168
rect 39051 34208 39093 34217
rect 39051 34168 39052 34208
rect 39092 34168 39093 34208
rect 39051 34159 39093 34168
rect 39339 34208 39381 34217
rect 39436 34212 39476 34243
rect 39339 34168 39340 34208
rect 39380 34168 39381 34208
rect 39339 34159 39381 34168
rect 38859 33872 38901 33881
rect 38859 33832 38860 33872
rect 38900 33832 38901 33872
rect 38859 33823 38901 33832
rect 38324 33664 38420 33704
rect 38284 33655 38324 33664
rect 38091 33620 38133 33629
rect 38074 33580 38092 33620
rect 38132 33580 38133 33620
rect 38074 33571 38133 33580
rect 38074 33536 38114 33571
rect 37996 33496 38114 33536
rect 37899 33452 37941 33461
rect 37899 33412 37900 33452
rect 37940 33412 37941 33452
rect 37899 33403 37941 33412
rect 37900 32864 37940 33403
rect 37900 32815 37940 32824
rect 37708 32311 37748 32320
rect 37803 32360 37845 32369
rect 37803 32320 37804 32360
rect 37844 32320 37845 32360
rect 37803 32311 37845 32320
rect 37612 32192 37652 32201
rect 37804 32192 37844 32311
rect 37516 32152 37612 32192
rect 37612 32143 37652 32152
rect 37708 32152 37844 32192
rect 37996 32192 38036 33496
rect 38283 33452 38325 33461
rect 38283 33412 38284 33452
rect 38324 33412 38325 33452
rect 38380 33452 38420 33664
rect 38476 33655 38516 33664
rect 38571 33704 38613 33713
rect 38571 33664 38572 33704
rect 38612 33664 38613 33704
rect 38571 33655 38613 33664
rect 38764 33704 38804 33713
rect 38572 33570 38612 33655
rect 38764 33452 38804 33664
rect 38380 33412 38804 33452
rect 38860 33704 38900 33823
rect 38283 33403 38325 33412
rect 38284 33318 38324 33403
rect 38284 32864 38324 32873
rect 38324 32824 38420 32864
rect 38284 32815 38324 32824
rect 37420 31184 37460 31193
rect 37036 31144 37420 31184
rect 37036 30689 37076 31144
rect 37420 31135 37460 31144
rect 37708 30689 37748 32152
rect 37996 32143 38036 32152
rect 38188 32192 38228 32201
rect 38228 32152 38324 32192
rect 38188 32143 38228 32152
rect 38284 31352 38324 32152
rect 38380 32024 38420 32824
rect 38860 32780 38900 33664
rect 38955 33704 38997 33713
rect 38955 33664 38956 33704
rect 38996 33664 38997 33704
rect 38955 33655 38997 33664
rect 39052 33704 39092 34159
rect 39243 34040 39285 34049
rect 39243 34000 39244 34040
rect 39284 34000 39285 34040
rect 39243 33991 39285 34000
rect 39052 33655 39092 33664
rect 39244 33704 39284 33991
rect 39532 33881 39572 34336
rect 39628 34376 39668 34385
rect 39820 34376 39860 34385
rect 39668 34336 39820 34376
rect 39628 34327 39668 34336
rect 39820 34327 39860 34336
rect 40012 34376 40052 34385
rect 39915 34292 39957 34301
rect 39915 34252 39916 34292
rect 39956 34252 39957 34292
rect 39915 34243 39957 34252
rect 39916 34158 39956 34243
rect 40012 34217 40052 34336
rect 40108 34376 40148 34411
rect 40204 34385 40244 34672
rect 40108 34325 40148 34336
rect 40203 34376 40245 34385
rect 40203 34336 40204 34376
rect 40244 34336 40245 34376
rect 40203 34327 40245 34336
rect 40396 34376 40436 34924
rect 40684 34914 40724 34999
rect 40876 34637 40916 35176
rect 40971 35216 41013 35225
rect 40971 35176 40972 35216
rect 41012 35176 41013 35216
rect 40971 35167 41013 35176
rect 40875 34628 40917 34637
rect 40875 34588 40876 34628
rect 40916 34588 40917 34628
rect 40875 34579 40917 34588
rect 40587 34460 40629 34469
rect 40587 34420 40588 34460
rect 40628 34420 40629 34460
rect 40587 34411 40629 34420
rect 40396 34327 40436 34336
rect 40491 34376 40533 34385
rect 40491 34336 40492 34376
rect 40532 34336 40533 34376
rect 40491 34327 40533 34336
rect 40588 34376 40628 34411
rect 40492 34242 40532 34327
rect 40588 34325 40628 34336
rect 40780 34376 40820 34387
rect 40780 34301 40820 34336
rect 40779 34292 40821 34301
rect 40779 34252 40780 34292
rect 40820 34252 40821 34292
rect 40779 34243 40821 34252
rect 40011 34208 40053 34217
rect 40011 34168 40012 34208
rect 40052 34168 40053 34208
rect 40011 34159 40053 34168
rect 40300 34208 40340 34217
rect 40340 34168 40436 34208
rect 40300 34159 40340 34168
rect 39531 33872 39573 33881
rect 39531 33832 39532 33872
rect 39572 33832 39573 33872
rect 39531 33823 39573 33832
rect 40012 33797 40052 34159
rect 40011 33788 40053 33797
rect 40011 33748 40012 33788
rect 40052 33748 40053 33788
rect 40011 33739 40053 33748
rect 39244 33655 39284 33664
rect 40107 33704 40149 33713
rect 40107 33664 40108 33704
rect 40148 33664 40149 33704
rect 40107 33655 40149 33664
rect 38956 33570 38996 33655
rect 40108 33570 40148 33655
rect 39915 33536 39957 33545
rect 39915 33496 39916 33536
rect 39956 33496 40052 33536
rect 39915 33487 39957 33496
rect 39916 33402 39956 33487
rect 39147 32864 39189 32873
rect 39147 32824 39148 32864
rect 39188 32824 39189 32864
rect 39147 32815 39189 32824
rect 38860 32740 38996 32780
rect 38475 32192 38517 32201
rect 38475 32152 38476 32192
rect 38516 32152 38517 32192
rect 38475 32143 38517 32152
rect 38380 31975 38420 31984
rect 38188 30689 38228 30774
rect 37035 30680 37077 30689
rect 37035 30640 37036 30680
rect 37076 30640 37077 30680
rect 37035 30631 37077 30640
rect 37227 30680 37269 30689
rect 37227 30640 37228 30680
rect 37268 30640 37269 30680
rect 37227 30631 37269 30640
rect 37707 30680 37749 30689
rect 37707 30640 37708 30680
rect 37748 30640 37749 30680
rect 37707 30631 37749 30640
rect 38092 30680 38132 30689
rect 37036 30546 37076 30631
rect 37228 30546 37268 30631
rect 37132 30428 37172 30437
rect 37172 30388 37652 30428
rect 37132 30379 37172 30388
rect 37515 30260 37557 30269
rect 37515 30220 37516 30260
rect 37556 30220 37557 30260
rect 37515 30211 37557 30220
rect 37131 30092 37173 30101
rect 37131 30052 37132 30092
rect 37172 30052 37173 30092
rect 37131 30043 37173 30052
rect 37132 29840 37172 30043
rect 37419 29924 37461 29933
rect 37419 29884 37420 29924
rect 37460 29884 37461 29924
rect 37419 29875 37461 29884
rect 37132 29791 37172 29800
rect 37323 29840 37365 29849
rect 37323 29800 37324 29840
rect 37364 29800 37365 29840
rect 37323 29791 37365 29800
rect 37420 29840 37460 29875
rect 37227 29168 37269 29177
rect 37227 29128 37228 29168
rect 37268 29128 37269 29168
rect 37227 29119 37269 29128
rect 37131 29084 37173 29093
rect 37131 29044 37132 29084
rect 37172 29044 37173 29084
rect 37131 29035 37173 29044
rect 37132 28328 37172 29035
rect 37228 29034 37268 29119
rect 37227 28916 37269 28925
rect 37227 28876 37228 28916
rect 37268 28876 37269 28916
rect 37227 28867 37269 28876
rect 37228 28664 37268 28867
rect 37324 28748 37364 29791
rect 37420 29789 37460 29800
rect 37516 29840 37556 30211
rect 37516 29791 37556 29800
rect 37612 29840 37652 30388
rect 37708 30269 37748 30631
rect 37707 30260 37749 30269
rect 37707 30220 37708 30260
rect 37748 30220 37749 30260
rect 37707 30211 37749 30220
rect 37612 29791 37652 29800
rect 37707 29672 37749 29681
rect 37707 29632 37708 29672
rect 37748 29632 37749 29672
rect 37707 29623 37749 29632
rect 37708 29538 37748 29623
rect 37324 28708 37460 28748
rect 37228 28624 37364 28664
rect 37132 28279 37172 28288
rect 37227 28328 37269 28337
rect 37227 28288 37228 28328
rect 37268 28288 37269 28328
rect 37227 28279 37269 28288
rect 37324 28328 37364 28624
rect 37324 28279 37364 28288
rect 37420 28328 37460 28708
rect 38092 28673 38132 30640
rect 38187 30680 38229 30689
rect 38187 30640 38188 30680
rect 38228 30640 38229 30680
rect 38187 30631 38229 30640
rect 38284 30512 38324 31312
rect 38379 30680 38421 30689
rect 38379 30640 38380 30680
rect 38420 30640 38421 30680
rect 38379 30631 38421 30640
rect 38380 30546 38420 30631
rect 38188 30472 38324 30512
rect 38188 29261 38228 30472
rect 38380 30428 38420 30437
rect 38476 30428 38516 32143
rect 38956 31856 38996 32740
rect 39148 32730 39188 32815
rect 39244 32201 39284 32286
rect 39243 32192 39285 32201
rect 39243 32152 39244 32192
rect 39284 32152 39285 32192
rect 40012 32192 40052 33496
rect 40299 32948 40341 32957
rect 40299 32908 40300 32948
rect 40340 32908 40341 32948
rect 40299 32899 40341 32908
rect 40300 32814 40340 32899
rect 40203 32528 40245 32537
rect 40203 32488 40204 32528
rect 40244 32488 40245 32528
rect 40203 32479 40245 32488
rect 40204 32360 40244 32479
rect 40204 32311 40244 32320
rect 40108 32192 40148 32201
rect 40012 32152 40108 32192
rect 39243 32143 39285 32152
rect 40108 32143 40148 32152
rect 39052 32024 39092 32033
rect 39092 31984 39764 32024
rect 39052 31975 39092 31984
rect 38956 31816 39092 31856
rect 38668 31184 38708 31193
rect 38708 31144 38804 31184
rect 38668 31135 38708 31144
rect 38668 30857 38708 30942
rect 38667 30848 38709 30857
rect 38667 30808 38668 30848
rect 38708 30808 38709 30848
rect 38667 30799 38709 30808
rect 38572 30680 38612 30689
rect 38764 30680 38804 31144
rect 39052 30848 39092 31816
rect 39724 31352 39764 31984
rect 39724 31303 39764 31312
rect 39916 31940 39956 31949
rect 39340 31268 39380 31277
rect 39340 31184 39380 31228
rect 39916 31184 39956 31900
rect 39340 31144 39956 31184
rect 40299 31184 40341 31193
rect 40299 31144 40300 31184
rect 40340 31144 40341 31184
rect 40299 31135 40341 31144
rect 39243 31016 39285 31025
rect 39243 30976 39244 31016
rect 39284 30976 39285 31016
rect 39243 30967 39285 30976
rect 38956 30808 39188 30848
rect 38612 30640 38708 30680
rect 38572 30631 38612 30640
rect 38420 30388 38516 30428
rect 38380 30379 38420 30388
rect 38283 30344 38325 30353
rect 38283 30304 38284 30344
rect 38324 30304 38325 30344
rect 38283 30295 38325 30304
rect 38284 29840 38324 30295
rect 38379 30008 38421 30017
rect 38379 29968 38380 30008
rect 38420 29968 38421 30008
rect 38379 29959 38421 29968
rect 38284 29791 38324 29800
rect 38380 29840 38420 29959
rect 38380 29791 38420 29800
rect 38476 29840 38516 29849
rect 38187 29252 38229 29261
rect 38187 29212 38188 29252
rect 38228 29212 38229 29252
rect 38187 29203 38229 29212
rect 38476 29093 38516 29800
rect 38572 29840 38612 29849
rect 38668 29840 38708 30640
rect 38764 30605 38804 30640
rect 38860 30680 38900 30689
rect 38763 30596 38805 30605
rect 38763 30556 38764 30596
rect 38804 30556 38805 30596
rect 38763 30547 38805 30556
rect 38764 30353 38804 30547
rect 38763 30344 38805 30353
rect 38763 30304 38764 30344
rect 38804 30304 38805 30344
rect 38763 30295 38805 30304
rect 38612 29800 38708 29840
rect 38764 30008 38804 30017
rect 38572 29791 38612 29800
rect 38475 29084 38517 29093
rect 38475 29044 38476 29084
rect 38516 29044 38517 29084
rect 38475 29035 38517 29044
rect 38380 28916 38420 28925
rect 38091 28664 38133 28673
rect 38091 28624 38092 28664
rect 38132 28624 38133 28664
rect 38091 28615 38133 28624
rect 38380 28337 38420 28876
rect 37420 28279 37460 28288
rect 38379 28328 38421 28337
rect 38379 28288 38380 28328
rect 38420 28288 38421 28328
rect 38379 28279 38421 28288
rect 37228 28194 37268 28279
rect 38188 28160 38228 28169
rect 36460 27607 36500 27616
rect 36844 27616 36980 27656
rect 37804 28120 38188 28160
rect 37804 27656 37844 28120
rect 38188 28111 38228 28120
rect 38764 27992 38804 29968
rect 38860 28589 38900 30640
rect 38956 29093 38996 30808
rect 39051 30680 39093 30689
rect 39051 30640 39052 30680
rect 39092 30640 39093 30680
rect 39051 30631 39093 30640
rect 39148 30680 39188 30808
rect 39148 30631 39188 30640
rect 39244 30680 39284 30967
rect 39531 30848 39573 30857
rect 39531 30808 39532 30848
rect 39572 30808 39573 30848
rect 39531 30799 39573 30808
rect 39244 30631 39284 30640
rect 39340 30680 39380 30691
rect 39052 30546 39092 30631
rect 39340 30605 39380 30640
rect 39532 30680 39572 30799
rect 39532 30631 39572 30640
rect 39339 30596 39381 30605
rect 39339 30556 39340 30596
rect 39380 30556 39381 30596
rect 39339 30547 39381 30556
rect 40300 30521 40340 31135
rect 39147 30512 39189 30521
rect 39147 30472 39148 30512
rect 39188 30472 39189 30512
rect 39147 30463 39189 30472
rect 40299 30512 40341 30521
rect 40299 30472 40300 30512
rect 40340 30472 40341 30512
rect 40299 30463 40341 30472
rect 39051 29840 39093 29849
rect 39051 29800 39052 29840
rect 39092 29800 39093 29840
rect 39051 29791 39093 29800
rect 39148 29840 39188 30463
rect 40204 30428 40244 30437
rect 39724 30388 40204 30428
rect 39435 30260 39477 30269
rect 39435 30220 39436 30260
rect 39476 30220 39477 30260
rect 39435 30211 39477 30220
rect 39148 29791 39188 29800
rect 39436 29840 39476 30211
rect 39052 29706 39092 29791
rect 38955 29084 38997 29093
rect 38955 29044 38956 29084
rect 38996 29044 38997 29084
rect 38955 29035 38997 29044
rect 39051 28664 39093 28673
rect 39051 28624 39052 28664
rect 39092 28624 39093 28664
rect 39051 28615 39093 28624
rect 38859 28580 38901 28589
rect 38859 28540 38860 28580
rect 38900 28540 38901 28580
rect 38859 28531 38901 28540
rect 39052 28580 39092 28615
rect 39052 28529 39092 28540
rect 39339 28580 39381 28589
rect 39339 28540 39340 28580
rect 39380 28540 39381 28580
rect 39339 28531 39381 28540
rect 39340 28446 39380 28531
rect 39436 28505 39476 29800
rect 39724 29840 39764 30388
rect 40204 30379 40244 30388
rect 39724 29791 39764 29800
rect 40108 29840 40148 29849
rect 39819 29336 39861 29345
rect 39819 29296 39820 29336
rect 39860 29296 39861 29336
rect 39819 29287 39861 29296
rect 39820 29168 39860 29287
rect 39820 29119 39860 29128
rect 40108 29093 40148 29800
rect 40107 29084 40149 29093
rect 40107 29044 40108 29084
rect 40148 29044 40149 29084
rect 40107 29035 40149 29044
rect 39435 28496 39477 28505
rect 39435 28456 39436 28496
rect 39476 28456 39477 28496
rect 39435 28447 39477 28456
rect 38859 28328 38901 28337
rect 38859 28288 38860 28328
rect 38900 28288 38901 28328
rect 38859 28279 38901 28288
rect 39148 28328 39188 28337
rect 38860 28194 38900 28279
rect 38668 27952 38804 27992
rect 38379 27740 38421 27749
rect 38379 27700 38380 27740
rect 38420 27700 38421 27740
rect 38379 27691 38421 27700
rect 36844 27077 36884 27616
rect 37804 27607 37844 27616
rect 38188 27656 38228 27665
rect 36940 27488 36980 27497
rect 36843 27068 36885 27077
rect 36843 27028 36844 27068
rect 36884 27028 36885 27068
rect 36843 27019 36885 27028
rect 36267 26900 36309 26909
rect 36267 26860 36268 26900
rect 36308 26860 36309 26900
rect 36267 26851 36309 26860
rect 35596 26767 35636 26776
rect 35691 26816 35733 26825
rect 35691 26776 35692 26816
rect 35732 26776 35733 26816
rect 35691 26767 35733 26776
rect 35884 26816 35924 26825
rect 35692 26682 35732 26767
rect 35884 26657 35924 26776
rect 35979 26816 36021 26825
rect 36076 26816 36116 26825
rect 35979 26776 35980 26816
rect 36020 26776 36076 26816
rect 35979 26767 36021 26776
rect 36076 26767 36116 26776
rect 36171 26816 36213 26825
rect 36171 26776 36172 26816
rect 36212 26776 36213 26816
rect 36171 26767 36213 26776
rect 35883 26648 35925 26657
rect 35883 26608 35884 26648
rect 35924 26608 35925 26648
rect 35883 26599 35925 26608
rect 35980 26648 36020 26657
rect 36075 26648 36117 26657
rect 36020 26608 36076 26648
rect 36116 26608 36117 26648
rect 35980 26599 36020 26608
rect 36075 26599 36117 26608
rect 35980 26144 36020 26153
rect 35692 26104 35980 26144
rect 35499 25472 35541 25481
rect 35499 25432 35500 25472
rect 35540 25432 35541 25472
rect 35499 25423 35541 25432
rect 35307 25388 35349 25397
rect 35307 25348 35308 25388
rect 35348 25348 35349 25388
rect 35307 25339 35349 25348
rect 35211 25304 35253 25313
rect 35211 25264 35212 25304
rect 35252 25264 35253 25304
rect 35211 25255 35253 25264
rect 35212 24800 35252 25255
rect 35595 25220 35637 25229
rect 35595 25180 35596 25220
rect 35636 25180 35637 25220
rect 35595 25171 35637 25180
rect 35212 24751 35252 24760
rect 35596 24632 35636 25171
rect 35692 24800 35732 26104
rect 35980 26095 36020 26104
rect 36075 25304 36117 25313
rect 36075 25264 36076 25304
rect 36116 25264 36117 25304
rect 36075 25255 36117 25264
rect 36076 25170 36116 25255
rect 35884 25136 35924 25145
rect 35924 25096 36020 25136
rect 35884 25087 35924 25096
rect 35692 24751 35732 24760
rect 35596 24583 35636 24592
rect 35788 24632 35828 24641
rect 35116 23920 35252 23960
rect 34636 23876 34676 23885
rect 34444 23836 34636 23876
rect 34348 23742 34388 23827
rect 34444 23624 34484 23836
rect 34636 23827 34676 23836
rect 34828 23633 34868 23718
rect 34348 23584 34484 23624
rect 34827 23624 34869 23633
rect 34827 23584 34828 23624
rect 34868 23584 34869 23624
rect 34156 22903 34196 22912
rect 34251 22952 34293 22961
rect 34251 22912 34252 22952
rect 34292 22912 34293 22952
rect 34251 22903 34293 22912
rect 33484 22828 33812 22868
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 32907 22532 32949 22541
rect 32907 22492 32908 22532
rect 32948 22492 32949 22532
rect 32907 22483 32949 22492
rect 31988 22240 32084 22280
rect 32812 22280 32852 22289
rect 31948 22231 31988 22240
rect 30891 22112 30933 22121
rect 30891 22072 30892 22112
rect 30932 22072 30933 22112
rect 30891 22063 30933 22072
rect 30892 21978 30932 22063
rect 30644 21736 30836 21776
rect 30604 21727 30644 21736
rect 30987 21608 31029 21617
rect 30987 21568 30988 21608
rect 31028 21568 31029 21608
rect 30987 21559 31029 21568
rect 30508 20140 30644 20180
rect 29836 20096 29876 20105
rect 28972 20047 29012 20056
rect 29740 20056 29836 20096
rect 28683 19340 28725 19349
rect 28683 19300 28684 19340
rect 28724 19300 28725 19340
rect 28683 19291 28725 19300
rect 28684 19256 28724 19291
rect 28684 19205 28724 19216
rect 29164 19256 29204 19265
rect 28780 19088 28820 19099
rect 28780 19013 28820 19048
rect 29068 19088 29108 19097
rect 28779 19004 28821 19013
rect 28779 18964 28780 19004
rect 28820 18964 28821 19004
rect 28779 18955 28821 18964
rect 28203 18920 28245 18929
rect 28203 18880 28204 18920
rect 28244 18880 28245 18920
rect 28203 18871 28245 18880
rect 28587 18920 28629 18929
rect 28587 18880 28588 18920
rect 28628 18880 28629 18920
rect 28587 18871 28629 18880
rect 28971 18920 29013 18929
rect 28971 18880 28972 18920
rect 29012 18880 29013 18920
rect 28971 18871 29013 18880
rect 28395 18584 28437 18593
rect 28395 18544 28396 18584
rect 28436 18544 28437 18584
rect 28395 18535 28437 18544
rect 28396 18450 28436 18535
rect 28972 17996 29012 18871
rect 29068 18005 29108 19048
rect 28972 17947 29012 17956
rect 29067 17996 29109 18005
rect 29067 17956 29068 17996
rect 29108 17956 29109 17996
rect 29067 17947 29109 17956
rect 29164 17921 29204 19216
rect 29260 19256 29300 19265
rect 27916 17912 27956 17921
rect 29163 17912 29205 17921
rect 27956 17872 28052 17912
rect 27916 17863 27956 17872
rect 27916 17744 27956 17753
rect 27916 17249 27956 17704
rect 27915 17240 27957 17249
rect 27915 17200 27916 17240
rect 27956 17200 27957 17240
rect 27915 17191 27957 17200
rect 27724 17116 27860 17156
rect 27380 17032 27486 17072
rect 27532 17032 27668 17072
rect 27340 17023 27380 17032
rect 27243 16988 27285 16997
rect 27243 16948 27244 16988
rect 27284 16948 27285 16988
rect 27446 16988 27486 17032
rect 27446 16948 27572 16988
rect 27243 16939 27285 16948
rect 27147 16820 27189 16829
rect 27147 16780 27148 16820
rect 27188 16780 27189 16820
rect 27147 16771 27189 16780
rect 27244 16661 27284 16939
rect 27435 16820 27477 16829
rect 27340 16780 27436 16820
rect 27476 16780 27477 16820
rect 27243 16652 27285 16661
rect 27243 16612 27244 16652
rect 27284 16612 27285 16652
rect 27243 16603 27285 16612
rect 27243 16400 27285 16409
rect 27243 16360 27244 16400
rect 27284 16360 27285 16400
rect 27243 16351 27285 16360
rect 26956 16183 26996 16192
rect 27051 16232 27093 16241
rect 27051 16192 27052 16232
rect 27092 16192 27093 16232
rect 27051 16183 27093 16192
rect 26859 16064 26901 16073
rect 26859 16024 26860 16064
rect 26900 16024 26901 16064
rect 26859 16015 26901 16024
rect 27244 15821 27284 16351
rect 27243 15812 27285 15821
rect 27243 15772 27244 15812
rect 27284 15772 27285 15812
rect 27243 15763 27285 15772
rect 26667 15728 26709 15737
rect 26667 15688 26668 15728
rect 26708 15688 26709 15728
rect 26667 15679 26709 15688
rect 27244 15569 27284 15763
rect 27243 15560 27285 15569
rect 27243 15520 27244 15560
rect 27284 15520 27285 15560
rect 27243 15511 27285 15520
rect 27340 15392 27380 16780
rect 27435 16771 27477 16780
rect 27436 16686 27476 16771
rect 27435 16400 27477 16409
rect 27435 16360 27436 16400
rect 27476 16360 27477 16400
rect 27435 16351 27477 16360
rect 27436 16232 27476 16351
rect 27532 16325 27572 16948
rect 27628 16913 27668 17032
rect 27627 16904 27669 16913
rect 27627 16864 27628 16904
rect 27668 16864 27669 16904
rect 27627 16855 27669 16864
rect 27724 16484 27764 17116
rect 27916 17072 27956 17081
rect 28012 17072 28052 17872
rect 29163 17872 29164 17912
rect 29204 17872 29205 17912
rect 29163 17863 29205 17872
rect 28300 17744 28340 17753
rect 29164 17744 29204 17753
rect 28340 17704 28628 17744
rect 28300 17695 28340 17704
rect 27820 17030 27860 17039
rect 27820 16913 27860 16990
rect 27956 17032 28052 17072
rect 28108 17576 28148 17585
rect 27819 16904 27861 16913
rect 27819 16864 27820 16904
rect 27860 16864 27861 16904
rect 27819 16855 27861 16864
rect 27820 16493 27860 16855
rect 27628 16444 27764 16484
rect 27819 16484 27861 16493
rect 27819 16444 27820 16484
rect 27860 16444 27861 16484
rect 27531 16316 27573 16325
rect 27531 16276 27532 16316
rect 27572 16276 27573 16316
rect 27531 16267 27573 16276
rect 27436 16183 27476 16192
rect 27532 16232 27572 16267
rect 27532 16182 27572 16192
rect 27628 16148 27668 16444
rect 27819 16435 27861 16444
rect 27724 16316 27764 16325
rect 27916 16316 27956 17032
rect 28108 16409 28148 17536
rect 28204 16820 28244 16829
rect 28244 16780 28436 16820
rect 28204 16771 28244 16780
rect 28203 16484 28245 16493
rect 28203 16444 28204 16484
rect 28244 16444 28245 16484
rect 28203 16435 28245 16444
rect 28107 16400 28149 16409
rect 28107 16360 28108 16400
rect 28148 16360 28149 16400
rect 28107 16351 28149 16360
rect 27764 16276 27956 16316
rect 27724 16267 27764 16276
rect 27916 16232 27956 16276
rect 27916 16183 27956 16192
rect 28011 16232 28053 16241
rect 28011 16192 28012 16232
rect 28052 16192 28053 16232
rect 28011 16183 28053 16192
rect 28204 16232 28244 16435
rect 28204 16183 28244 16192
rect 28396 16232 28436 16780
rect 28396 16183 28436 16192
rect 28492 16232 28532 16241
rect 27628 16108 27764 16148
rect 27435 16064 27477 16073
rect 27435 16024 27436 16064
rect 27476 16024 27477 16064
rect 27435 16015 27477 16024
rect 27436 15728 27476 16015
rect 27627 15980 27669 15989
rect 27627 15940 27628 15980
rect 27668 15940 27669 15980
rect 27627 15931 27669 15940
rect 27436 15679 27476 15688
rect 27628 15560 27668 15931
rect 27724 15653 27764 16108
rect 28012 16098 28052 16183
rect 28204 16064 28244 16073
rect 28492 16064 28532 16192
rect 28244 16024 28532 16064
rect 28204 16015 28244 16024
rect 27916 15772 28436 15812
rect 27916 15728 27956 15772
rect 27916 15679 27956 15688
rect 27723 15644 27765 15653
rect 28107 15644 28149 15653
rect 27723 15604 27724 15644
rect 27764 15604 27860 15644
rect 27723 15595 27765 15604
rect 27628 15511 27668 15520
rect 27628 15392 27668 15401
rect 27340 15352 27628 15392
rect 27628 15343 27668 15352
rect 26571 15224 26613 15233
rect 26571 15184 26572 15224
rect 26612 15184 26613 15224
rect 26571 15175 26613 15184
rect 26283 15056 26325 15065
rect 26283 15016 26284 15056
rect 26324 15016 26325 15056
rect 26283 15007 26325 15016
rect 26379 14804 26421 14813
rect 26379 14764 26380 14804
rect 26420 14764 26421 14804
rect 26379 14755 26421 14764
rect 25996 14671 26036 14680
rect 26380 14720 26420 14755
rect 26380 14669 26420 14680
rect 26572 14720 26612 15175
rect 26859 14804 26901 14813
rect 26859 14764 26860 14804
rect 26900 14764 26901 14804
rect 26859 14755 26901 14764
rect 26572 14671 26612 14680
rect 26860 14720 26900 14755
rect 26860 14669 26900 14680
rect 25899 14636 25941 14645
rect 25899 14596 25900 14636
rect 25940 14596 25941 14636
rect 25899 14587 25941 14596
rect 25900 14502 25940 14587
rect 26091 14552 26133 14561
rect 26091 14512 26092 14552
rect 26132 14512 26133 14552
rect 26091 14503 26133 14512
rect 26667 14552 26709 14561
rect 26667 14512 26668 14552
rect 26708 14512 26709 14552
rect 26667 14503 26709 14512
rect 25900 14216 25940 14225
rect 25804 14176 25900 14216
rect 25420 14048 25460 14057
rect 25420 13217 25460 14008
rect 25515 14048 25557 14057
rect 25515 14008 25516 14048
rect 25556 14008 25557 14048
rect 25515 13999 25557 14008
rect 25708 14048 25748 14057
rect 25804 14048 25844 14176
rect 25900 14167 25940 14176
rect 25748 14008 25844 14048
rect 26092 14048 26132 14503
rect 26668 14418 26708 14503
rect 27052 14225 27092 14310
rect 27243 14300 27285 14309
rect 27243 14260 27244 14300
rect 27284 14260 27285 14300
rect 27243 14251 27285 14260
rect 27051 14216 27093 14225
rect 27051 14176 27052 14216
rect 27092 14176 27093 14216
rect 27051 14167 27093 14176
rect 27244 14216 27284 14251
rect 27244 14165 27284 14176
rect 26187 14132 26229 14141
rect 26187 14092 26188 14132
rect 26228 14092 26229 14132
rect 26187 14083 26229 14092
rect 25708 13999 25748 14008
rect 26092 13999 26132 14008
rect 26188 14048 26228 14083
rect 25516 13914 25556 13999
rect 26188 13973 26228 14008
rect 26283 14048 26325 14057
rect 26283 14008 26284 14048
rect 26324 14008 26325 14048
rect 26283 13999 26325 14008
rect 26764 14048 26804 14057
rect 26187 13964 26229 13973
rect 26187 13924 26188 13964
rect 26228 13924 26229 13964
rect 26187 13915 26229 13924
rect 25707 13880 25749 13889
rect 26188 13884 26228 13915
rect 25707 13840 25708 13880
rect 25748 13840 25749 13880
rect 25707 13831 25749 13840
rect 25708 13746 25748 13831
rect 25707 13292 25749 13301
rect 25707 13252 25708 13292
rect 25748 13252 25749 13292
rect 25707 13243 25749 13252
rect 26091 13292 26133 13301
rect 26091 13252 26092 13292
rect 26132 13252 26133 13292
rect 26091 13243 26133 13252
rect 25419 13208 25461 13217
rect 25419 13168 25420 13208
rect 25460 13168 25461 13208
rect 25419 13159 25461 13168
rect 25420 13040 25460 13049
rect 25460 13000 25652 13040
rect 25420 12991 25460 13000
rect 25612 12536 25652 13000
rect 25612 12487 25652 12496
rect 25708 11948 25748 13243
rect 26092 13208 26132 13243
rect 26092 13157 26132 13168
rect 26284 12713 26324 13999
rect 26475 13628 26517 13637
rect 26475 13588 26476 13628
rect 26516 13588 26517 13628
rect 26475 13579 26517 13588
rect 26476 13385 26516 13579
rect 26764 13553 26804 14008
rect 26860 14048 26900 14057
rect 27436 14048 27476 14057
rect 26900 14008 26996 14048
rect 26860 13999 26900 14008
rect 26763 13544 26805 13553
rect 26763 13504 26764 13544
rect 26804 13504 26805 13544
rect 26763 13495 26805 13504
rect 26475 13376 26517 13385
rect 26475 13336 26476 13376
rect 26516 13336 26517 13376
rect 26475 13327 26517 13336
rect 26668 13376 26708 13385
rect 26476 13166 26516 13327
rect 26476 13117 26516 13126
rect 26572 13292 26612 13301
rect 26572 12872 26612 13252
rect 26380 12832 26612 12872
rect 26283 12704 26325 12713
rect 26283 12664 26284 12704
rect 26324 12664 26325 12704
rect 26283 12655 26325 12664
rect 25899 12620 25941 12629
rect 25899 12580 25900 12620
rect 25940 12580 25941 12620
rect 25899 12571 25941 12580
rect 25612 11908 25748 11948
rect 25612 11537 25652 11908
rect 25900 11696 25940 12571
rect 25996 12536 26036 12545
rect 25996 12377 26036 12496
rect 26187 12536 26229 12545
rect 26187 12496 26188 12536
rect 26228 12496 26229 12536
rect 26187 12487 26229 12496
rect 26380 12536 26420 12832
rect 26668 12797 26708 13336
rect 26764 13301 26804 13386
rect 26763 13292 26805 13301
rect 26763 13252 26764 13292
rect 26804 13252 26805 13292
rect 26763 13243 26805 13252
rect 26860 13208 26900 13217
rect 26763 13124 26805 13133
rect 26763 13084 26764 13124
rect 26804 13084 26805 13124
rect 26763 13075 26805 13084
rect 26764 12965 26804 13075
rect 26763 12956 26805 12965
rect 26763 12916 26764 12956
rect 26804 12916 26805 12956
rect 26763 12907 26805 12916
rect 26667 12788 26709 12797
rect 26667 12748 26668 12788
rect 26708 12748 26709 12788
rect 26667 12739 26709 12748
rect 26571 12704 26613 12713
rect 26571 12664 26572 12704
rect 26612 12664 26613 12704
rect 26571 12655 26613 12664
rect 26572 12536 26612 12655
rect 26764 12620 26804 12907
rect 26860 12881 26900 13168
rect 26859 12872 26901 12881
rect 26859 12832 26860 12872
rect 26900 12832 26901 12872
rect 26859 12823 26901 12832
rect 26764 12580 26900 12620
rect 26668 12536 26708 12545
rect 26572 12496 26668 12536
rect 26860 12536 26900 12580
rect 26091 12452 26133 12461
rect 26091 12412 26092 12452
rect 26132 12412 26133 12452
rect 26091 12403 26133 12412
rect 25995 12368 26037 12377
rect 25995 12328 25996 12368
rect 26036 12328 26037 12368
rect 25995 12319 26037 12328
rect 26092 12318 26132 12403
rect 26188 12368 26228 12487
rect 26188 12319 26228 12328
rect 26284 12452 26324 12461
rect 26284 12209 26324 12412
rect 26283 12200 26325 12209
rect 26283 12160 26284 12200
rect 26324 12160 26325 12200
rect 26283 12151 26325 12160
rect 26380 11873 26420 12496
rect 26571 12368 26613 12377
rect 26571 12328 26572 12368
rect 26612 12328 26613 12368
rect 26571 12319 26613 12328
rect 26379 11864 26421 11873
rect 26379 11824 26380 11864
rect 26420 11824 26421 11864
rect 26379 11815 26421 11824
rect 25801 11685 25841 11694
rect 25900 11647 25940 11656
rect 26092 11696 26132 11705
rect 25801 11621 25841 11645
rect 25801 11612 25845 11621
rect 25801 11572 25804 11612
rect 25844 11572 25846 11612
rect 25803 11563 25846 11572
rect 25611 11528 25653 11537
rect 25611 11488 25612 11528
rect 25652 11488 25653 11528
rect 25611 11479 25653 11488
rect 25804 11528 25846 11563
rect 26092 11537 26132 11656
rect 26187 11696 26229 11705
rect 26187 11656 26188 11696
rect 26228 11656 26229 11696
rect 26187 11647 26229 11656
rect 26284 11696 26324 11705
rect 26188 11562 26228 11647
rect 26091 11528 26133 11537
rect 25804 11488 25940 11528
rect 25804 11478 25844 11488
rect 25803 11276 25845 11285
rect 25803 11236 25804 11276
rect 25844 11236 25845 11276
rect 25803 11227 25845 11236
rect 25707 11192 25749 11201
rect 25707 11152 25708 11192
rect 25748 11152 25749 11192
rect 25707 11143 25749 11152
rect 25708 11058 25748 11143
rect 25804 11024 25844 11227
rect 25804 10975 25844 10984
rect 25419 10184 25461 10193
rect 25419 10144 25420 10184
rect 25460 10144 25461 10184
rect 25419 10135 25461 10144
rect 25323 10016 25365 10025
rect 25323 9976 25324 10016
rect 25364 9976 25365 10016
rect 25323 9967 25365 9976
rect 25324 9882 25364 9967
rect 25228 9437 25268 9472
rect 25227 9428 25269 9437
rect 25227 9388 25228 9428
rect 25268 9388 25269 9428
rect 25227 9379 25269 9388
rect 25324 9260 25364 9269
rect 25132 9220 25324 9260
rect 24844 8833 24884 8842
rect 25035 8840 25077 8849
rect 24651 8791 24693 8800
rect 25035 8800 25036 8840
rect 25076 8800 25077 8840
rect 25035 8791 25077 8800
rect 24652 8672 24692 8791
rect 24652 8623 24692 8632
rect 24748 8756 24788 8765
rect 24940 8756 24980 8765
rect 24748 8597 24788 8716
rect 24844 8716 24940 8756
rect 24747 8588 24789 8597
rect 24747 8548 24748 8588
rect 24788 8548 24789 8588
rect 24747 8539 24789 8548
rect 24844 8429 24884 8716
rect 24940 8707 24980 8716
rect 25036 8672 25076 8681
rect 25036 8513 25076 8632
rect 25132 8597 25172 9220
rect 25324 9211 25364 9220
rect 25324 8672 25364 8681
rect 25420 8672 25460 10135
rect 25364 8632 25460 8672
rect 25516 8800 25748 8840
rect 25324 8623 25364 8632
rect 25131 8588 25173 8597
rect 25131 8548 25132 8588
rect 25172 8548 25173 8588
rect 25131 8539 25173 8548
rect 25035 8504 25077 8513
rect 25035 8464 25036 8504
rect 25076 8464 25077 8504
rect 25035 8455 25077 8464
rect 24843 8420 24885 8429
rect 24843 8380 24844 8420
rect 24884 8380 24885 8420
rect 24843 8371 24885 8380
rect 25036 8261 25076 8455
rect 25035 8252 25077 8261
rect 25035 8212 25036 8252
rect 25076 8212 25077 8252
rect 25132 8252 25172 8539
rect 25227 8504 25269 8513
rect 25227 8464 25228 8504
rect 25268 8464 25269 8504
rect 25227 8455 25269 8464
rect 25228 8370 25268 8455
rect 25132 8212 25364 8252
rect 25035 8203 25077 8212
rect 24748 8000 24788 8009
rect 25036 8000 25076 8011
rect 25228 8009 25268 8094
rect 24788 7960 24884 8000
rect 24748 7951 24788 7960
rect 24712 7328 24754 7337
rect 24712 7288 24713 7328
rect 24753 7288 24754 7328
rect 24712 7279 24754 7288
rect 24555 7244 24597 7253
rect 24555 7204 24556 7244
rect 24596 7204 24597 7244
rect 24555 7195 24597 7204
rect 24172 7160 24212 7169
rect 24076 7120 24172 7160
rect 23979 7111 24021 7120
rect 24172 7111 24212 7120
rect 24268 7160 24308 7169
rect 23883 7076 23925 7085
rect 23883 7036 23884 7076
rect 23924 7036 23925 7076
rect 23883 7027 23925 7036
rect 24268 7001 24308 7120
rect 24460 7160 24500 7169
rect 23787 6992 23829 7001
rect 23787 6952 23788 6992
rect 23828 6952 23829 6992
rect 23787 6943 23829 6952
rect 23980 6992 24020 7001
rect 23691 6572 23733 6581
rect 23691 6532 23692 6572
rect 23732 6532 23733 6572
rect 23691 6523 23733 6532
rect 23595 6488 23637 6497
rect 23595 6448 23596 6488
rect 23636 6448 23637 6488
rect 23595 6439 23637 6448
rect 23692 6488 23732 6523
rect 23692 6437 23732 6448
rect 23308 6355 23348 6364
rect 23308 5900 23348 5909
rect 23212 5860 23308 5900
rect 23308 5851 23348 5860
rect 23788 5732 23828 6943
rect 23980 6824 24020 6952
rect 24267 6992 24309 7001
rect 24267 6952 24268 6992
rect 24308 6952 24309 6992
rect 24267 6943 24309 6952
rect 24460 6824 24500 7120
rect 24556 7160 24596 7195
rect 24713 7175 24753 7279
rect 24713 7126 24753 7135
rect 24556 7109 24596 7120
rect 23980 6784 24500 6824
rect 23883 6656 23925 6665
rect 24460 6656 24500 6665
rect 23883 6616 23884 6656
rect 23924 6616 23925 6656
rect 23883 6607 23925 6616
rect 23980 6616 24212 6656
rect 23884 6522 23924 6607
rect 23980 6488 24020 6616
rect 23980 6439 24020 6448
rect 24075 6488 24117 6497
rect 24075 6448 24076 6488
rect 24116 6448 24117 6488
rect 24075 6439 24117 6448
rect 24172 6488 24212 6616
rect 24500 6616 24788 6656
rect 24460 6607 24500 6616
rect 23788 5683 23828 5692
rect 23307 5648 23349 5657
rect 23307 5608 23308 5648
rect 23348 5608 23349 5648
rect 23307 5599 23349 5608
rect 23404 5648 23444 5657
rect 23692 5648 23732 5657
rect 23444 5608 23692 5648
rect 23404 5599 23444 5608
rect 23692 5599 23732 5608
rect 23980 5648 24020 5657
rect 24076 5648 24116 6439
rect 24020 5608 24116 5648
rect 23980 5599 24020 5608
rect 23211 5060 23253 5069
rect 23211 5020 23212 5060
rect 23252 5020 23253 5060
rect 23211 5011 23253 5020
rect 23019 4976 23061 4985
rect 23019 4936 23020 4976
rect 23060 4936 23061 4976
rect 23019 4927 23061 4936
rect 23020 4842 23060 4927
rect 23212 4388 23252 5011
rect 23308 4976 23348 5599
rect 23308 4927 23348 4936
rect 23691 4976 23733 4985
rect 23691 4936 23692 4976
rect 23732 4936 23733 4976
rect 23691 4927 23733 4936
rect 23595 4892 23637 4901
rect 23595 4852 23596 4892
rect 23636 4852 23637 4892
rect 23595 4843 23637 4852
rect 23308 4388 23348 4397
rect 23212 4348 23308 4388
rect 23308 4339 23348 4348
rect 23596 4136 23636 4843
rect 23596 3893 23636 4096
rect 23692 4136 23732 4927
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23924 4220
rect 23787 4171 23829 4180
rect 23692 4087 23732 4096
rect 23884 4136 23924 4180
rect 23884 4087 23924 4096
rect 23883 3968 23925 3977
rect 23883 3928 23884 3968
rect 23924 3928 23925 3968
rect 23883 3919 23925 3928
rect 23595 3884 23637 3893
rect 23595 3844 23596 3884
rect 23636 3844 23637 3884
rect 23595 3835 23637 3844
rect 23884 3834 23924 3919
rect 23020 3464 23060 3473
rect 23308 3464 23348 3473
rect 22924 3424 23020 3464
rect 23060 3424 23308 3464
rect 23020 3415 23060 3424
rect 23308 3415 23348 3424
rect 23979 3212 24021 3221
rect 23979 3172 23980 3212
rect 24020 3172 24021 3212
rect 23979 3163 24021 3172
rect 23980 3078 24020 3163
rect 23979 2876 24021 2885
rect 23979 2836 23980 2876
rect 24020 2836 24021 2876
rect 23979 2827 24021 2836
rect 23116 2633 23156 2718
rect 23307 2708 23349 2717
rect 23307 2668 23308 2708
rect 23348 2668 23349 2708
rect 23307 2659 23349 2668
rect 23595 2708 23637 2717
rect 23595 2668 23596 2708
rect 23636 2668 23637 2708
rect 23595 2659 23637 2668
rect 23115 2624 23157 2633
rect 23115 2584 23116 2624
rect 23156 2584 23157 2624
rect 23115 2575 23157 2584
rect 21292 1903 21332 1912
rect 22251 1952 22293 1961
rect 22251 1912 22252 1952
rect 22292 1912 22293 1952
rect 22251 1903 22293 1912
rect 22539 1952 22581 1961
rect 22539 1912 22540 1952
rect 22580 1912 22581 1952
rect 22539 1903 22581 1912
rect 21004 1818 21044 1903
rect 22540 1818 22580 1903
rect 17451 1700 17493 1709
rect 17451 1660 17452 1700
rect 17492 1660 17493 1700
rect 17451 1651 17493 1660
rect 17452 1566 17492 1651
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 15532 1280 15572 1289
rect 15436 1240 15532 1280
rect 15532 1231 15572 1240
rect 11924 1072 12116 1112
rect 23308 1112 23348 2659
rect 23596 1952 23636 2659
rect 23980 2624 24020 2827
rect 24172 2801 24212 6448
rect 24267 6488 24309 6497
rect 24267 6448 24268 6488
rect 24308 6448 24309 6488
rect 24267 6439 24309 6448
rect 24652 6488 24692 6497
rect 24268 6354 24308 6439
rect 24652 5984 24692 6448
rect 24748 6488 24788 6616
rect 24748 6439 24788 6448
rect 24844 6161 24884 7960
rect 25036 7925 25076 7960
rect 25227 8000 25269 8009
rect 25227 7960 25228 8000
rect 25268 7960 25269 8000
rect 25227 7951 25269 7960
rect 25324 8000 25364 8212
rect 25516 8168 25556 8800
rect 25708 8714 25748 8800
rect 25612 8672 25652 8681
rect 25708 8665 25748 8674
rect 25804 8672 25844 8681
rect 25612 8597 25652 8632
rect 25900 8672 25940 11488
rect 26091 11488 26092 11528
rect 26132 11488 26133 11528
rect 26091 11479 26133 11488
rect 26284 11360 26324 11656
rect 26379 11696 26421 11705
rect 26379 11656 26380 11696
rect 26420 11656 26421 11696
rect 26379 11647 26421 11656
rect 26572 11696 26612 12319
rect 26668 12284 26708 12496
rect 26764 12494 26804 12503
rect 26763 12454 26764 12461
rect 26860 12487 26900 12496
rect 26804 12454 26805 12461
rect 26763 12452 26805 12454
rect 26763 12412 26764 12452
rect 26804 12412 26805 12452
rect 26763 12403 26805 12412
rect 26764 12359 26804 12403
rect 26668 12244 26900 12284
rect 26763 11864 26805 11873
rect 26763 11824 26764 11864
rect 26804 11824 26805 11864
rect 26763 11815 26805 11824
rect 26667 11780 26709 11789
rect 26667 11740 26668 11780
rect 26708 11740 26709 11780
rect 26667 11731 26709 11740
rect 26572 11647 26612 11656
rect 26668 11696 26708 11731
rect 26380 11562 26420 11647
rect 26668 11645 26708 11656
rect 26764 11696 26804 11815
rect 26764 11647 26804 11656
rect 26860 11696 26900 12244
rect 26956 12209 26996 14008
rect 27052 14008 27436 14048
rect 27052 13208 27092 14008
rect 27436 13999 27476 14008
rect 27532 14048 27572 14057
rect 27147 13880 27189 13889
rect 27147 13840 27148 13880
rect 27188 13840 27189 13880
rect 27147 13831 27189 13840
rect 27052 13159 27092 13168
rect 27148 13208 27188 13831
rect 27532 13469 27572 14008
rect 27628 14048 27668 14057
rect 27628 13880 27668 14008
rect 27724 14048 27764 14057
rect 27820 14048 27860 15604
rect 28107 15604 28108 15644
rect 28148 15604 28149 15644
rect 28107 15595 28149 15604
rect 28011 15560 28053 15569
rect 28011 15520 28012 15560
rect 28052 15520 28053 15560
rect 28011 15511 28053 15520
rect 28108 15560 28148 15595
rect 28012 15426 28052 15511
rect 28108 15509 28148 15520
rect 28203 15560 28245 15569
rect 28203 15520 28204 15560
rect 28244 15520 28245 15560
rect 28203 15511 28245 15520
rect 28396 15560 28436 15772
rect 28396 15511 28436 15520
rect 28204 15426 28244 15511
rect 28107 15224 28149 15233
rect 28107 15184 28108 15224
rect 28148 15184 28149 15224
rect 28107 15175 28149 15184
rect 28108 14720 28148 15175
rect 28588 14888 28628 17704
rect 29068 17704 29164 17744
rect 28774 17240 28816 17249
rect 28774 17200 28775 17240
rect 28815 17200 28816 17240
rect 28774 17191 28816 17200
rect 28775 17081 28815 17191
rect 28972 17081 29012 17166
rect 28774 17072 28816 17081
rect 28774 17032 28775 17072
rect 28815 17032 28816 17072
rect 28774 17023 28816 17032
rect 28876 17072 28916 17081
rect 28775 16938 28815 17023
rect 28876 16661 28916 17032
rect 28971 17072 29013 17081
rect 28971 17032 28972 17072
rect 29012 17032 29013 17072
rect 28971 17023 29013 17032
rect 28971 16820 29013 16829
rect 28971 16780 28972 16820
rect 29012 16780 29013 16820
rect 28971 16771 29013 16780
rect 28875 16652 28917 16661
rect 28875 16612 28876 16652
rect 28916 16612 28917 16652
rect 28875 16603 28917 16612
rect 28684 16232 28724 16241
rect 28972 16232 29012 16771
rect 29068 16400 29108 17704
rect 29164 17695 29204 17704
rect 29260 17501 29300 19216
rect 29356 19256 29396 19265
rect 29548 19256 29588 19265
rect 29396 19216 29492 19256
rect 29356 19207 29396 19216
rect 29355 17996 29397 18005
rect 29355 17956 29356 17996
rect 29396 17956 29397 17996
rect 29355 17947 29397 17956
rect 29259 17492 29301 17501
rect 29259 17452 29260 17492
rect 29300 17452 29301 17492
rect 29259 17443 29301 17452
rect 29259 17324 29301 17333
rect 29259 17284 29260 17324
rect 29300 17284 29301 17324
rect 29259 17275 29301 17284
rect 29163 17072 29205 17081
rect 29163 17032 29164 17072
rect 29204 17032 29205 17072
rect 29163 17023 29205 17032
rect 29260 17072 29300 17275
rect 29260 17023 29300 17032
rect 29164 16938 29204 17023
rect 29259 16820 29301 16829
rect 29259 16780 29260 16820
rect 29300 16780 29301 16820
rect 29259 16771 29301 16780
rect 29260 16686 29300 16771
rect 29068 16360 29204 16400
rect 28724 16192 28820 16232
rect 28684 16183 28724 16192
rect 28683 16064 28725 16073
rect 28683 16024 28684 16064
rect 28724 16024 28725 16064
rect 28683 16015 28725 16024
rect 28684 15930 28724 16015
rect 28780 15905 28820 16192
rect 28972 16183 29012 16192
rect 29068 16232 29108 16241
rect 29068 16073 29108 16192
rect 29164 16148 29204 16360
rect 29260 16232 29300 16241
rect 29356 16232 29396 17947
rect 29452 17912 29492 19216
rect 29588 19216 29684 19256
rect 29548 19207 29588 19216
rect 29547 18668 29589 18677
rect 29547 18628 29548 18668
rect 29588 18628 29589 18668
rect 29547 18619 29589 18628
rect 29548 18584 29588 18619
rect 29548 18533 29588 18544
rect 29644 17996 29684 19216
rect 29740 18593 29780 20056
rect 29836 20047 29876 20056
rect 30315 20096 30357 20105
rect 30315 20056 30316 20096
rect 30356 20056 30357 20096
rect 30315 20047 30357 20056
rect 29931 19928 29973 19937
rect 29931 19888 29932 19928
rect 29972 19888 29973 19928
rect 29931 19879 29973 19888
rect 29932 19256 29972 19879
rect 29932 19207 29972 19216
rect 29836 18677 29876 18762
rect 29835 18668 29877 18677
rect 29835 18628 29836 18668
rect 29876 18628 29972 18668
rect 29835 18619 29877 18628
rect 29739 18584 29781 18593
rect 29739 18544 29740 18584
rect 29780 18544 29781 18584
rect 29739 18535 29781 18544
rect 29836 18584 29876 18619
rect 29836 18535 29876 18544
rect 29836 17996 29876 18005
rect 29644 17956 29836 17996
rect 29836 17947 29876 17956
rect 29452 17872 29684 17912
rect 29451 17156 29493 17165
rect 29451 17116 29452 17156
rect 29492 17116 29493 17156
rect 29451 17107 29493 17116
rect 29452 16577 29492 17107
rect 29547 16988 29589 16997
rect 29547 16948 29548 16988
rect 29588 16948 29589 16988
rect 29547 16939 29589 16948
rect 29548 16854 29588 16939
rect 29451 16568 29493 16577
rect 29451 16528 29452 16568
rect 29492 16528 29493 16568
rect 29451 16519 29493 16528
rect 29451 16400 29493 16409
rect 29451 16360 29452 16400
rect 29492 16360 29493 16400
rect 29451 16351 29493 16360
rect 29300 16192 29396 16232
rect 29260 16183 29300 16192
rect 29452 16148 29492 16351
rect 29644 16157 29684 17872
rect 29932 17660 29972 18628
rect 30316 17996 30356 20047
rect 30604 19097 30644 20140
rect 30988 19844 31028 21559
rect 31468 20096 31508 20105
rect 31028 19804 31220 19844
rect 30988 19795 31028 19804
rect 30795 19256 30837 19265
rect 30795 19216 30796 19256
rect 30836 19216 30837 19256
rect 30795 19207 30837 19216
rect 30796 19122 30836 19207
rect 30603 19088 30645 19097
rect 30603 19048 30604 19088
rect 30644 19048 30645 19088
rect 30603 19039 30645 19048
rect 30316 17947 30356 17956
rect 30508 18332 30548 18341
rect 29932 17620 30068 17660
rect 29931 16316 29973 16325
rect 29931 16276 29932 16316
rect 29972 16276 29973 16316
rect 29931 16267 29973 16276
rect 29932 16232 29972 16267
rect 29164 16099 29204 16108
rect 29356 16108 29492 16148
rect 29643 16148 29685 16157
rect 29643 16108 29644 16148
rect 29684 16108 29685 16148
rect 29067 16064 29109 16073
rect 29067 16024 29068 16064
rect 29108 16024 29109 16064
rect 29067 16015 29109 16024
rect 29259 15980 29301 15989
rect 29259 15940 29260 15980
rect 29300 15940 29301 15980
rect 29259 15931 29301 15940
rect 28779 15896 28821 15905
rect 28779 15856 28780 15896
rect 28820 15856 28821 15896
rect 28779 15847 28821 15856
rect 28780 15485 28820 15847
rect 29260 15560 29300 15931
rect 29260 15511 29300 15520
rect 29356 15560 29396 16108
rect 29643 16099 29685 16108
rect 29836 16064 29876 16073
rect 29740 16024 29836 16064
rect 29740 15728 29780 16024
rect 29836 16015 29876 16024
rect 29932 15989 29972 16192
rect 30028 16232 30068 17620
rect 30219 17576 30261 17585
rect 30219 17536 30220 17576
rect 30260 17536 30261 17576
rect 30219 17527 30261 17536
rect 30220 17333 30260 17527
rect 30219 17324 30261 17333
rect 30219 17284 30220 17324
rect 30260 17284 30261 17324
rect 30219 17275 30261 17284
rect 30220 16493 30260 17275
rect 30411 17072 30453 17081
rect 30508 17072 30548 18292
rect 30604 17753 30644 19039
rect 31083 18584 31125 18593
rect 31083 18544 31084 18584
rect 31124 18544 31125 18584
rect 31180 18584 31220 19804
rect 31468 19172 31508 20056
rect 31852 20096 31892 20105
rect 31659 19340 31701 19349
rect 31659 19300 31660 19340
rect 31700 19300 31701 19340
rect 31659 19291 31701 19300
rect 31468 19132 31604 19172
rect 31467 19004 31509 19013
rect 31467 18964 31468 19004
rect 31508 18964 31509 19004
rect 31467 18955 31509 18964
rect 31372 18584 31412 18593
rect 31180 18544 31372 18584
rect 31083 18535 31125 18544
rect 31372 18535 31412 18544
rect 30700 18332 30740 18341
rect 30603 17744 30645 17753
rect 30603 17704 30604 17744
rect 30644 17704 30645 17744
rect 30603 17695 30645 17704
rect 30411 17032 30412 17072
rect 30452 17032 30548 17072
rect 30411 17023 30453 17032
rect 30412 16938 30452 17023
rect 30219 16484 30261 16493
rect 30219 16444 30220 16484
rect 30260 16444 30261 16484
rect 30219 16435 30261 16444
rect 30028 16183 30068 16192
rect 30123 16232 30165 16241
rect 30123 16192 30124 16232
rect 30164 16192 30165 16232
rect 30123 16183 30165 16192
rect 30507 16232 30549 16241
rect 30507 16192 30508 16232
rect 30548 16192 30549 16232
rect 30507 16183 30549 16192
rect 30124 16098 30164 16183
rect 30508 16098 30548 16183
rect 29931 15980 29973 15989
rect 29931 15940 29932 15980
rect 29972 15940 29973 15980
rect 29931 15931 29973 15940
rect 30603 15812 30645 15821
rect 30603 15772 30604 15812
rect 30644 15772 30645 15812
rect 30603 15763 30645 15772
rect 29356 15511 29396 15520
rect 29452 15688 29780 15728
rect 29931 15728 29973 15737
rect 29931 15688 29932 15728
rect 29972 15688 29973 15728
rect 29452 15560 29492 15688
rect 29931 15679 29973 15688
rect 30507 15728 30549 15737
rect 30507 15688 30508 15728
rect 30548 15688 30549 15728
rect 30507 15679 30549 15688
rect 29452 15511 29492 15520
rect 29548 15560 29588 15569
rect 28779 15476 28821 15485
rect 28779 15436 28780 15476
rect 28820 15436 28821 15476
rect 28779 15427 28821 15436
rect 29068 15308 29108 15317
rect 29068 15140 29108 15268
rect 29548 15149 29588 15520
rect 29740 15560 29780 15569
rect 28780 15100 29108 15140
rect 29547 15140 29589 15149
rect 29547 15100 29548 15140
rect 29588 15100 29589 15140
rect 28588 14848 28724 14888
rect 28299 14804 28341 14813
rect 28299 14764 28300 14804
rect 28340 14764 28341 14804
rect 28299 14755 28341 14764
rect 28108 14671 28148 14680
rect 28300 14720 28340 14755
rect 28300 14669 28340 14680
rect 28492 14720 28532 14729
rect 28204 14552 28244 14561
rect 28204 14393 28244 14512
rect 27915 14384 27957 14393
rect 27915 14344 27916 14384
rect 27956 14344 27957 14384
rect 27915 14335 27957 14344
rect 28203 14384 28245 14393
rect 28203 14344 28204 14384
rect 28244 14344 28245 14384
rect 28203 14335 28245 14344
rect 27764 14008 27860 14048
rect 27724 13999 27764 14008
rect 27628 13840 27764 13880
rect 27531 13460 27573 13469
rect 27531 13420 27532 13460
rect 27572 13420 27573 13460
rect 27531 13411 27573 13420
rect 27724 13460 27764 13840
rect 27724 13411 27764 13420
rect 27916 13250 27956 14335
rect 28492 14309 28532 14680
rect 28587 14720 28629 14729
rect 28587 14680 28588 14720
rect 28628 14680 28629 14720
rect 28587 14671 28629 14680
rect 28588 14586 28628 14671
rect 28684 14636 28724 14848
rect 28780 14720 28820 15100
rect 29547 15091 29589 15100
rect 29740 14813 29780 15520
rect 29932 15560 29972 15679
rect 30508 15594 30548 15679
rect 29932 15511 29972 15520
rect 30028 15560 30068 15569
rect 29836 15392 29876 15401
rect 29739 14804 29781 14813
rect 29739 14764 29740 14804
rect 29780 14764 29781 14804
rect 29739 14755 29781 14764
rect 28780 14671 28820 14680
rect 29068 14720 29108 14729
rect 28684 14587 28724 14596
rect 28972 14552 29012 14561
rect 28491 14300 28533 14309
rect 28491 14260 28492 14300
rect 28532 14260 28533 14300
rect 28491 14251 28533 14260
rect 28587 14216 28629 14225
rect 28587 14176 28588 14216
rect 28628 14176 28629 14216
rect 28587 14167 28629 14176
rect 28395 14132 28437 14141
rect 28395 14092 28396 14132
rect 28436 14092 28437 14132
rect 28395 14083 28437 14092
rect 28204 14048 28244 14057
rect 28108 14008 28204 14048
rect 27148 13159 27188 13168
rect 27244 13208 27284 13217
rect 27244 12872 27284 13168
rect 27340 13208 27380 13217
rect 27340 12881 27380 13168
rect 27724 13208 27764 13217
rect 28012 13217 28052 13302
rect 27916 13201 27956 13210
rect 28011 13208 28053 13217
rect 27052 12832 27284 12872
rect 27339 12872 27381 12881
rect 27339 12832 27340 12872
rect 27380 12832 27381 12872
rect 27052 12704 27092 12832
rect 27339 12823 27381 12832
rect 27724 12713 27764 13168
rect 28011 13168 28012 13208
rect 28052 13168 28053 13208
rect 28011 13159 28053 13168
rect 27819 12956 27861 12965
rect 27819 12916 27820 12956
rect 27860 12916 27861 12956
rect 27819 12907 27861 12916
rect 27052 12655 27092 12664
rect 27244 12704 27284 12713
rect 26955 12200 26997 12209
rect 27244 12200 27284 12664
rect 27339 12704 27381 12713
rect 27339 12664 27340 12704
rect 27380 12664 27381 12704
rect 27339 12655 27381 12664
rect 27723 12704 27765 12713
rect 27723 12664 27724 12704
rect 27764 12664 27765 12704
rect 27723 12655 27765 12664
rect 26955 12160 26956 12200
rect 26996 12160 26997 12200
rect 26955 12151 26997 12160
rect 27148 12160 27284 12200
rect 26955 11948 26997 11957
rect 26955 11908 26956 11948
rect 26996 11908 26997 11948
rect 26955 11899 26997 11908
rect 26860 11647 26900 11656
rect 26956 11360 26996 11899
rect 27148 11873 27188 12160
rect 27243 12032 27285 12041
rect 27243 11992 27244 12032
rect 27284 11992 27285 12032
rect 27243 11983 27285 11992
rect 27147 11864 27189 11873
rect 27147 11824 27148 11864
rect 27188 11824 27189 11864
rect 27147 11815 27189 11824
rect 25996 11320 26324 11360
rect 26860 11320 26996 11360
rect 27052 11696 27092 11705
rect 25996 11192 26036 11320
rect 25996 11143 26036 11152
rect 26475 11192 26517 11201
rect 26475 11152 26476 11192
rect 26516 11152 26517 11192
rect 26475 11143 26517 11152
rect 26667 11192 26709 11201
rect 26667 11152 26668 11192
rect 26708 11152 26709 11192
rect 26667 11143 26709 11152
rect 26284 11033 26324 11118
rect 26476 11033 26516 11143
rect 26092 11024 26132 11033
rect 26092 10781 26132 10984
rect 26188 11024 26228 11033
rect 26188 10856 26228 10984
rect 26283 11024 26325 11033
rect 26283 10984 26284 11024
rect 26324 10984 26325 11024
rect 26283 10975 26325 10984
rect 26475 11024 26517 11033
rect 26475 10984 26476 11024
rect 26516 10984 26517 11024
rect 26475 10975 26517 10984
rect 26668 11024 26708 11143
rect 26860 11045 26900 11320
rect 27052 11192 27092 11656
rect 27147 11696 27189 11705
rect 27147 11656 27148 11696
rect 27188 11656 27189 11696
rect 27147 11647 27189 11656
rect 27244 11696 27284 11983
rect 27244 11647 27284 11656
rect 27340 11696 27380 12655
rect 27627 12620 27669 12629
rect 27627 12580 27628 12620
rect 27668 12580 27669 12620
rect 27627 12578 27669 12580
rect 27820 12620 27860 12907
rect 27915 12872 27957 12881
rect 27915 12832 27916 12872
rect 27956 12832 27957 12872
rect 27915 12823 27957 12832
rect 27627 12571 27764 12578
rect 27820 12571 27860 12580
rect 27436 12536 27476 12547
rect 27436 12461 27476 12496
rect 27531 12536 27573 12545
rect 27628 12538 27764 12571
rect 27916 12545 27956 12823
rect 27531 12496 27532 12536
rect 27572 12496 27573 12536
rect 27531 12487 27573 12496
rect 27724 12536 27764 12538
rect 27724 12487 27764 12496
rect 27915 12536 27957 12545
rect 27915 12496 27916 12536
rect 27956 12496 27957 12536
rect 27915 12487 27957 12496
rect 27435 12452 27477 12461
rect 27435 12412 27436 12452
rect 27476 12412 27477 12452
rect 27435 12403 27477 12412
rect 27340 11647 27380 11656
rect 27148 11562 27188 11647
rect 27436 11621 27476 12403
rect 27532 12402 27572 12487
rect 27916 12402 27956 12487
rect 28108 12293 28148 14008
rect 28204 13999 28244 14008
rect 28300 14048 28340 14057
rect 28300 13721 28340 14008
rect 28299 13712 28341 13721
rect 28299 13672 28300 13712
rect 28340 13672 28341 13712
rect 28299 13663 28341 13672
rect 28204 13385 28244 13470
rect 28203 13376 28245 13385
rect 28203 13336 28204 13376
rect 28244 13336 28245 13376
rect 28203 13327 28245 13336
rect 28204 13166 28244 13219
rect 28203 13126 28204 13133
rect 28244 13126 28245 13133
rect 28203 13124 28245 13126
rect 28203 13084 28204 13124
rect 28244 13084 28245 13124
rect 28203 13075 28245 13084
rect 28300 12377 28340 13663
rect 28396 13208 28436 14083
rect 28588 14082 28628 14167
rect 28972 14141 29012 14512
rect 28971 14132 29013 14141
rect 28971 14092 28972 14132
rect 29012 14092 29013 14132
rect 28971 14083 29013 14092
rect 29068 14048 29108 14680
rect 29356 14720 29396 14729
rect 29259 14384 29301 14393
rect 29259 14344 29260 14384
rect 29300 14344 29301 14384
rect 29259 14335 29301 14344
rect 28875 13964 28917 13973
rect 28875 13924 28876 13964
rect 28916 13924 28917 13964
rect 28875 13915 28917 13924
rect 28779 13880 28821 13889
rect 28779 13840 28780 13880
rect 28820 13840 28821 13880
rect 28779 13831 28821 13840
rect 28587 13628 28629 13637
rect 28587 13588 28588 13628
rect 28628 13588 28629 13628
rect 28587 13579 28629 13588
rect 28396 12965 28436 13168
rect 28492 13208 28532 13217
rect 28395 12956 28437 12965
rect 28395 12916 28396 12956
rect 28436 12916 28437 12956
rect 28395 12907 28437 12916
rect 28492 12545 28532 13168
rect 28588 12956 28628 13579
rect 28683 13376 28725 13385
rect 28683 13336 28684 13376
rect 28724 13336 28725 13376
rect 28683 13327 28725 13336
rect 28684 13208 28724 13327
rect 28684 13159 28724 13168
rect 28780 13208 28820 13831
rect 28780 13159 28820 13168
rect 28876 13124 28916 13915
rect 28971 13880 29013 13889
rect 28971 13840 28972 13880
rect 29012 13840 29013 13880
rect 28971 13831 29013 13840
rect 28972 13746 29012 13831
rect 29068 13637 29108 14008
rect 29164 14048 29204 14057
rect 29164 13805 29204 14008
rect 29163 13796 29205 13805
rect 29163 13756 29164 13796
rect 29204 13756 29205 13796
rect 29163 13747 29205 13756
rect 29067 13628 29109 13637
rect 29067 13588 29068 13628
rect 29108 13588 29109 13628
rect 29260 13628 29300 14335
rect 29356 14141 29396 14680
rect 29548 14720 29588 14729
rect 29451 14636 29493 14645
rect 29451 14596 29452 14636
rect 29492 14596 29493 14636
rect 29451 14587 29493 14596
rect 29452 14502 29492 14587
rect 29355 14132 29397 14141
rect 29355 14092 29356 14132
rect 29396 14092 29397 14132
rect 29355 14083 29397 14092
rect 29548 13880 29588 14680
rect 29644 14720 29684 14731
rect 29836 14729 29876 15352
rect 30028 14888 30068 15520
rect 30604 15560 30644 15763
rect 30700 15653 30740 18292
rect 30987 17744 31029 17753
rect 30987 17704 30988 17744
rect 31028 17704 31029 17744
rect 30987 17695 31029 17704
rect 30988 17610 31028 17695
rect 30892 16157 30932 16188
rect 30891 16148 30933 16157
rect 30891 16108 30892 16148
rect 30932 16108 30933 16148
rect 30891 16099 30933 16108
rect 30892 16064 30932 16099
rect 30699 15644 30741 15653
rect 30699 15604 30700 15644
rect 30740 15604 30741 15644
rect 30699 15595 30741 15604
rect 30604 15233 30644 15520
rect 30603 15224 30645 15233
rect 30603 15184 30604 15224
rect 30644 15184 30645 15224
rect 30603 15175 30645 15184
rect 29932 14848 30068 14888
rect 29644 14645 29684 14680
rect 29835 14720 29877 14729
rect 29835 14680 29836 14720
rect 29876 14680 29877 14720
rect 29835 14671 29877 14680
rect 29643 14636 29685 14645
rect 29643 14596 29644 14636
rect 29684 14596 29685 14636
rect 29643 14587 29685 14596
rect 29932 14384 29972 14848
rect 30027 14720 30069 14729
rect 30027 14680 30028 14720
rect 30068 14680 30069 14720
rect 30027 14671 30069 14680
rect 30124 14720 30164 14729
rect 30164 14680 30260 14720
rect 30124 14671 30164 14680
rect 30028 14552 30068 14671
rect 30028 14503 30068 14512
rect 29932 14344 30068 14384
rect 29643 14216 29685 14225
rect 29643 14176 29644 14216
rect 29684 14176 29685 14216
rect 29643 14167 29685 14176
rect 29931 14216 29973 14225
rect 29931 14176 29932 14216
rect 29972 14176 29973 14216
rect 29931 14167 29973 14176
rect 29644 14048 29684 14167
rect 29740 14057 29780 14142
rect 29836 14132 29876 14141
rect 29644 13999 29684 14008
rect 29739 14048 29781 14057
rect 29739 14008 29740 14048
rect 29780 14008 29781 14048
rect 29739 13999 29781 14008
rect 29836 13889 29876 14092
rect 29932 14082 29972 14167
rect 29740 13880 29780 13889
rect 29548 13840 29740 13880
rect 29740 13831 29780 13840
rect 29835 13880 29877 13889
rect 29835 13840 29836 13880
rect 29876 13840 29877 13880
rect 29835 13831 29877 13840
rect 29260 13588 29396 13628
rect 29067 13579 29109 13588
rect 29259 13460 29301 13469
rect 29259 13420 29260 13460
rect 29300 13420 29301 13460
rect 29259 13411 29301 13420
rect 29260 13326 29300 13411
rect 28876 13075 28916 13084
rect 28972 13208 29012 13217
rect 28972 13049 29012 13168
rect 29259 13124 29301 13133
rect 29259 13084 29260 13124
rect 29300 13084 29301 13124
rect 29259 13075 29301 13084
rect 29356 13124 29396 13588
rect 30028 13217 30068 14344
rect 30220 13973 30260 14680
rect 30315 14636 30357 14645
rect 30315 14596 30316 14636
rect 30356 14596 30357 14636
rect 30315 14587 30357 14596
rect 30316 14502 30356 14587
rect 30219 13964 30261 13973
rect 30219 13924 30220 13964
rect 30260 13924 30261 13964
rect 30219 13915 30261 13924
rect 30795 13796 30837 13805
rect 30795 13756 30796 13796
rect 30836 13756 30837 13796
rect 30795 13747 30837 13756
rect 30411 13712 30453 13721
rect 30411 13672 30412 13712
rect 30452 13672 30453 13712
rect 30411 13663 30453 13672
rect 30220 13385 30260 13470
rect 30219 13376 30261 13385
rect 30219 13336 30220 13376
rect 30260 13336 30261 13376
rect 30219 13327 30261 13336
rect 29356 13075 29396 13084
rect 29452 13208 29492 13217
rect 28971 13040 29013 13049
rect 28971 13000 28972 13040
rect 29012 13000 29013 13040
rect 28971 12991 29013 13000
rect 29260 13040 29300 13075
rect 29260 12989 29300 13000
rect 28588 12916 28916 12956
rect 28684 12704 28724 12713
rect 28396 12536 28436 12545
rect 28299 12368 28341 12377
rect 28299 12328 28300 12368
rect 28340 12328 28341 12368
rect 28299 12319 28341 12328
rect 28396 12293 28436 12496
rect 28491 12536 28533 12545
rect 28491 12496 28492 12536
rect 28532 12496 28533 12536
rect 28491 12487 28533 12496
rect 28684 12461 28724 12664
rect 28876 12536 28916 12916
rect 29452 12713 29492 13168
rect 29548 13208 29588 13217
rect 29740 13208 29780 13217
rect 29588 13168 29684 13208
rect 29548 13159 29588 13168
rect 29547 12956 29589 12965
rect 29547 12916 29548 12956
rect 29588 12916 29589 12956
rect 29547 12907 29589 12916
rect 29067 12704 29109 12713
rect 29067 12664 29068 12704
rect 29108 12664 29109 12704
rect 29067 12655 29109 12664
rect 29451 12704 29493 12713
rect 29451 12664 29452 12704
rect 29492 12664 29493 12704
rect 29548 12704 29588 12907
rect 29548 12664 29593 12704
rect 29451 12655 29493 12664
rect 28971 12620 29013 12629
rect 28971 12580 28972 12620
rect 29012 12580 29013 12620
rect 28971 12571 29013 12580
rect 28876 12487 28916 12496
rect 28972 12536 29012 12571
rect 28972 12485 29012 12496
rect 28683 12452 28725 12461
rect 28683 12412 28684 12452
rect 28724 12412 28725 12452
rect 28683 12403 28725 12412
rect 28491 12368 28533 12377
rect 29068 12368 29108 12655
rect 29163 12620 29205 12629
rect 29163 12580 29164 12620
rect 29204 12580 29205 12620
rect 29163 12571 29205 12580
rect 29356 12578 29396 12587
rect 29553 12578 29593 12664
rect 29644 12620 29684 13168
rect 29740 12965 29780 13168
rect 29835 13208 29877 13217
rect 29835 13168 29836 13208
rect 29876 13168 29877 13208
rect 29835 13159 29877 13168
rect 30027 13208 30069 13217
rect 30027 13168 30028 13208
rect 30068 13168 30069 13208
rect 30027 13159 30069 13168
rect 30220 13208 30260 13217
rect 29836 13074 29876 13159
rect 30028 13040 30068 13049
rect 29932 13000 30028 13040
rect 29739 12956 29781 12965
rect 29739 12916 29740 12956
rect 29780 12916 29781 12956
rect 29739 12907 29781 12916
rect 29164 12536 29204 12571
rect 29164 12485 29204 12496
rect 29355 12538 29356 12545
rect 29396 12538 29397 12545
rect 29355 12536 29397 12538
rect 29355 12496 29356 12536
rect 29396 12496 29397 12536
rect 29355 12487 29397 12496
rect 29548 12538 29593 12578
rect 29643 12580 29684 12620
rect 29548 12536 29588 12538
rect 29548 12487 29588 12496
rect 29260 12452 29300 12463
rect 29356 12443 29396 12487
rect 29452 12452 29492 12461
rect 29260 12377 29300 12412
rect 29643 12452 29683 12580
rect 29835 12536 29877 12545
rect 29835 12496 29836 12536
rect 29876 12496 29877 12536
rect 29835 12487 29877 12496
rect 29932 12536 29972 13000
rect 30028 12991 30068 13000
rect 30220 12788 30260 13168
rect 30412 13208 30452 13663
rect 30796 13301 30836 13747
rect 30795 13292 30837 13301
rect 30795 13252 30796 13292
rect 30836 13252 30837 13292
rect 30795 13243 30837 13252
rect 30412 12965 30452 13168
rect 30604 13208 30644 13217
rect 30411 12956 30453 12965
rect 30411 12916 30412 12956
rect 30452 12916 30453 12956
rect 30411 12907 30453 12916
rect 30604 12881 30644 13168
rect 30796 13208 30836 13243
rect 30796 13158 30836 13168
rect 30699 13040 30741 13049
rect 30699 13000 30700 13040
rect 30740 13000 30741 13040
rect 30699 12991 30741 13000
rect 30700 12906 30740 12991
rect 30603 12872 30645 12881
rect 30603 12832 30604 12872
rect 30644 12832 30645 12872
rect 30603 12823 30645 12832
rect 30220 12748 30452 12788
rect 29932 12487 29972 12496
rect 30028 12536 30068 12545
rect 29643 12412 29684 12452
rect 28491 12328 28492 12368
rect 28532 12328 28533 12368
rect 28491 12319 28533 12328
rect 28972 12328 29108 12368
rect 29259 12368 29301 12377
rect 29452 12368 29492 12412
rect 29259 12328 29260 12368
rect 29300 12328 29301 12368
rect 28107 12284 28149 12293
rect 28107 12244 28108 12284
rect 28148 12244 28149 12284
rect 28107 12235 28149 12244
rect 28395 12284 28437 12293
rect 28395 12244 28396 12284
rect 28436 12244 28437 12284
rect 28395 12235 28437 12244
rect 28492 12234 28532 12319
rect 28972 11696 29012 12328
rect 29259 12319 29301 12328
rect 29356 12328 29492 12368
rect 29067 11948 29109 11957
rect 29067 11908 29068 11948
rect 29108 11908 29109 11948
rect 29067 11899 29109 11908
rect 28972 11647 29012 11656
rect 29068 11696 29108 11899
rect 29356 11789 29396 12328
rect 29644 12284 29684 12412
rect 29452 12244 29684 12284
rect 29740 12368 29780 12377
rect 29355 11780 29397 11789
rect 29355 11740 29356 11780
rect 29396 11740 29397 11780
rect 29355 11731 29397 11740
rect 29068 11647 29108 11656
rect 29164 11696 29204 11705
rect 27435 11612 27477 11621
rect 27435 11572 27436 11612
rect 27476 11572 27477 11612
rect 27435 11563 27477 11572
rect 29164 11537 29204 11656
rect 29260 11696 29300 11705
rect 29163 11528 29205 11537
rect 29163 11488 29164 11528
rect 29204 11488 29205 11528
rect 29163 11479 29205 11488
rect 26860 10996 26900 11005
rect 26956 11152 27092 11192
rect 28780 11192 28820 11201
rect 28820 11152 29108 11192
rect 26668 10949 26708 10984
rect 26667 10940 26709 10949
rect 26956 10940 26996 11152
rect 28780 11143 28820 11152
rect 27339 11108 27381 11117
rect 27339 11068 27340 11108
rect 27380 11068 27381 11108
rect 27339 11059 27381 11068
rect 27051 11024 27093 11033
rect 27051 10984 27052 11024
rect 27092 10984 27093 11024
rect 27051 10975 27093 10984
rect 27244 11024 27284 11033
rect 26667 10900 26668 10940
rect 26708 10900 26709 10940
rect 26667 10891 26709 10900
rect 26860 10900 26996 10940
rect 26476 10856 26516 10865
rect 26188 10816 26476 10856
rect 26476 10807 26516 10816
rect 26091 10772 26133 10781
rect 26091 10732 26092 10772
rect 26132 10732 26133 10772
rect 26091 10723 26133 10732
rect 26379 10688 26421 10697
rect 26379 10648 26380 10688
rect 26420 10648 26421 10688
rect 26379 10639 26421 10648
rect 26187 10520 26229 10529
rect 26187 10480 26188 10520
rect 26228 10480 26229 10520
rect 26187 10471 26229 10480
rect 26188 10193 26228 10471
rect 26283 10352 26325 10361
rect 26283 10312 26284 10352
rect 26324 10312 26325 10352
rect 26283 10303 26325 10312
rect 26187 10184 26229 10193
rect 26187 10144 26188 10184
rect 26228 10144 26229 10184
rect 26187 10135 26229 10144
rect 26284 10184 26324 10303
rect 26284 10135 26324 10144
rect 26380 10184 26420 10639
rect 26668 10436 26708 10445
rect 26860 10436 26900 10900
rect 27052 10890 27092 10975
rect 26955 10772 26997 10781
rect 26955 10732 26956 10772
rect 26996 10732 26997 10772
rect 26955 10723 26997 10732
rect 26956 10638 26996 10723
rect 26708 10396 26900 10436
rect 26668 10387 26708 10396
rect 27152 10352 27194 10361
rect 27244 10352 27284 10984
rect 27340 10974 27380 11059
rect 27436 11024 27476 11033
rect 27152 10312 27153 10352
rect 27193 10312 27284 10352
rect 27152 10303 27194 10312
rect 26380 10135 26420 10144
rect 26476 10184 26516 10193
rect 26668 10184 26708 10193
rect 26516 10144 26668 10184
rect 26476 10135 26516 10144
rect 26668 10135 26708 10144
rect 26764 10184 26804 10193
rect 26188 10050 26228 10135
rect 26283 10016 26325 10025
rect 26283 9976 26284 10016
rect 26324 9976 26325 10016
rect 26283 9967 26325 9976
rect 26092 8681 26132 8766
rect 26091 8672 26133 8681
rect 25900 8632 26036 8672
rect 25611 8588 25653 8597
rect 25611 8548 25612 8588
rect 25652 8548 25653 8588
rect 25611 8539 25653 8548
rect 25612 8429 25652 8539
rect 25611 8420 25653 8429
rect 25611 8380 25612 8420
rect 25652 8380 25653 8420
rect 25611 8371 25653 8380
rect 25611 8252 25653 8261
rect 25611 8212 25612 8252
rect 25652 8212 25653 8252
rect 25804 8252 25844 8632
rect 25899 8504 25941 8513
rect 25899 8464 25900 8504
rect 25940 8464 25941 8504
rect 25899 8455 25941 8464
rect 25900 8370 25940 8455
rect 25804 8212 25940 8252
rect 25611 8203 25653 8212
rect 25324 7925 25364 7960
rect 25420 8128 25556 8168
rect 24940 7916 24980 7925
rect 24940 6488 24980 7876
rect 25035 7916 25077 7925
rect 25035 7876 25036 7916
rect 25076 7876 25077 7916
rect 25035 7867 25077 7876
rect 25323 7916 25365 7925
rect 25323 7876 25324 7916
rect 25364 7876 25365 7916
rect 25323 7867 25365 7876
rect 25227 7748 25269 7757
rect 25227 7708 25228 7748
rect 25268 7708 25269 7748
rect 25227 7699 25269 7708
rect 25228 7614 25268 7699
rect 25420 7337 25460 8128
rect 25516 8000 25556 8009
rect 25516 7421 25556 7960
rect 25612 8000 25652 8203
rect 25767 8009 25807 8094
rect 25612 7951 25652 7960
rect 25766 8000 25808 8009
rect 25766 7960 25767 8000
rect 25807 7960 25808 8000
rect 25766 7951 25808 7960
rect 25900 7832 25940 8212
rect 25996 8168 26036 8632
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 26187 8504 26229 8513
rect 26187 8464 26188 8504
rect 26228 8464 26229 8504
rect 26187 8455 26229 8464
rect 25996 8128 26132 8168
rect 25995 8000 26037 8009
rect 25995 7960 25996 8000
rect 26036 7960 26037 8000
rect 25995 7951 26037 7960
rect 25708 7792 25940 7832
rect 25515 7412 25557 7421
rect 25515 7372 25516 7412
rect 25556 7372 25557 7412
rect 25515 7363 25557 7372
rect 25419 7328 25461 7337
rect 25419 7288 25420 7328
rect 25460 7288 25461 7328
rect 25419 7279 25461 7288
rect 25035 7160 25077 7169
rect 25035 7120 25036 7160
rect 25076 7120 25077 7160
rect 25035 7111 25077 7120
rect 25228 7160 25268 7171
rect 25036 6917 25076 7111
rect 25228 7085 25268 7120
rect 25419 7160 25461 7169
rect 25419 7120 25420 7160
rect 25460 7120 25461 7160
rect 25419 7111 25461 7120
rect 25516 7160 25556 7169
rect 25556 7120 25652 7160
rect 25516 7111 25556 7120
rect 25227 7076 25269 7085
rect 25227 7036 25228 7076
rect 25268 7036 25269 7076
rect 25227 7027 25269 7036
rect 25420 7026 25460 7111
rect 25035 6908 25077 6917
rect 25035 6868 25036 6908
rect 25076 6868 25077 6908
rect 25035 6859 25077 6868
rect 24940 6439 24980 6448
rect 25132 6488 25172 6497
rect 24939 6320 24981 6329
rect 24939 6280 24940 6320
rect 24980 6280 24981 6320
rect 24939 6271 24981 6280
rect 24940 6186 24980 6271
rect 25132 6236 25172 6448
rect 25227 6488 25269 6497
rect 25227 6448 25228 6488
rect 25268 6448 25269 6488
rect 25227 6439 25269 6448
rect 25516 6488 25556 6497
rect 25228 6404 25268 6439
rect 25228 6353 25268 6364
rect 25419 6404 25461 6413
rect 25419 6364 25420 6404
rect 25460 6364 25461 6404
rect 25419 6355 25461 6364
rect 25324 6320 25364 6329
rect 25132 6196 25268 6236
rect 24843 6152 24885 6161
rect 24843 6112 24844 6152
rect 24884 6112 24885 6152
rect 24843 6103 24885 6112
rect 25131 6068 25173 6077
rect 25131 6028 25132 6068
rect 25172 6028 25173 6068
rect 25131 6019 25173 6028
rect 24652 5944 25076 5984
rect 24939 5816 24981 5825
rect 24939 5776 24940 5816
rect 24980 5776 24981 5816
rect 24939 5767 24981 5776
rect 24267 5648 24309 5657
rect 24267 5608 24268 5648
rect 24308 5608 24309 5648
rect 24267 5599 24309 5608
rect 24268 5514 24308 5599
rect 24460 4976 24500 4985
rect 24171 2792 24213 2801
rect 24171 2752 24172 2792
rect 24212 2752 24213 2792
rect 24171 2743 24213 2752
rect 24460 2633 24500 4936
rect 24843 4136 24885 4145
rect 24843 4096 24844 4136
rect 24884 4096 24885 4136
rect 24940 4136 24980 5767
rect 25036 5480 25076 5944
rect 25132 5657 25172 6019
rect 25131 5648 25173 5657
rect 25131 5608 25132 5648
rect 25172 5608 25173 5648
rect 25131 5599 25173 5608
rect 25132 5480 25172 5489
rect 25036 5440 25132 5480
rect 25132 5431 25172 5440
rect 25228 4388 25268 6196
rect 25324 5909 25364 6280
rect 25420 6270 25460 6355
rect 25323 5900 25365 5909
rect 25323 5860 25324 5900
rect 25364 5860 25365 5900
rect 25323 5851 25365 5860
rect 25324 5648 25364 5657
rect 25324 5489 25364 5608
rect 25419 5648 25461 5657
rect 25419 5608 25420 5648
rect 25460 5608 25461 5648
rect 25419 5599 25461 5608
rect 25420 5514 25460 5599
rect 25323 5480 25365 5489
rect 25323 5440 25324 5480
rect 25364 5440 25365 5480
rect 25323 5431 25365 5440
rect 25324 4976 25364 4985
rect 25324 4649 25364 4936
rect 25323 4640 25365 4649
rect 25323 4600 25324 4640
rect 25364 4600 25365 4640
rect 25323 4591 25365 4600
rect 25228 4339 25268 4348
rect 25132 4136 25172 4145
rect 24940 4096 25132 4136
rect 24843 4087 24885 4096
rect 25132 4087 25172 4096
rect 24555 2708 24597 2717
rect 24555 2668 24556 2708
rect 24596 2668 24597 2708
rect 24555 2659 24597 2668
rect 23980 2575 24020 2584
rect 24364 2624 24404 2633
rect 23979 2036 24021 2045
rect 23979 1996 23980 2036
rect 24020 1996 24021 2036
rect 23979 1987 24021 1996
rect 23596 1903 23636 1912
rect 23980 1952 24020 1987
rect 23980 1901 24020 1912
rect 24364 1280 24404 2584
rect 24459 2624 24501 2633
rect 24459 2584 24460 2624
rect 24500 2584 24501 2624
rect 24459 2575 24501 2584
rect 24556 2574 24596 2659
rect 24844 1952 24884 4087
rect 25324 3968 25364 4591
rect 25516 4388 25556 6448
rect 25612 6161 25652 7120
rect 25708 6992 25748 7792
rect 25996 7664 26036 7951
rect 25900 7624 26036 7664
rect 25900 7160 25940 7624
rect 25995 7328 26037 7337
rect 25995 7288 25996 7328
rect 26036 7288 26037 7328
rect 25995 7279 26037 7288
rect 25900 7111 25940 7120
rect 25996 7160 26036 7279
rect 25996 7111 26036 7120
rect 25708 6943 25748 6952
rect 26092 6824 26132 8128
rect 26188 7832 26228 8455
rect 26284 8000 26324 9967
rect 26764 9773 26804 10144
rect 26956 10184 26996 10193
rect 26763 9764 26805 9773
rect 26763 9724 26764 9764
rect 26804 9724 26805 9764
rect 26763 9715 26805 9724
rect 26380 8840 26420 8849
rect 26420 8800 26612 8840
rect 26380 8791 26420 8800
rect 26572 8681 26612 8800
rect 26380 8672 26420 8681
rect 26380 8429 26420 8632
rect 26571 8672 26613 8681
rect 26571 8632 26572 8672
rect 26612 8632 26613 8672
rect 26571 8623 26613 8632
rect 26764 8672 26804 8681
rect 26668 8504 26708 8513
rect 26476 8464 26668 8504
rect 26379 8420 26421 8429
rect 26379 8380 26380 8420
rect 26420 8380 26421 8420
rect 26379 8371 26421 8380
rect 26380 8000 26420 8009
rect 26284 7960 26380 8000
rect 26188 7792 26324 7832
rect 26188 7160 26228 7169
rect 26188 6833 26228 7120
rect 26284 7160 26324 7792
rect 26380 7337 26420 7960
rect 26379 7328 26421 7337
rect 26379 7288 26380 7328
rect 26420 7288 26421 7328
rect 26379 7279 26421 7288
rect 26284 7111 26324 7120
rect 26380 7160 26420 7169
rect 26476 7160 26516 8464
rect 26668 8455 26708 8464
rect 26764 8252 26804 8632
rect 26572 8212 26804 8252
rect 26860 8672 26900 8681
rect 26572 8168 26612 8212
rect 26860 8168 26900 8632
rect 26956 8336 26996 10144
rect 27051 10184 27093 10193
rect 27051 10144 27052 10184
rect 27092 10144 27093 10184
rect 27051 10135 27093 10144
rect 27153 10184 27193 10303
rect 27436 10193 27476 10984
rect 28684 11024 28724 11033
rect 28684 10865 28724 10984
rect 28876 11024 28916 11033
rect 28876 10865 28916 10984
rect 29068 11024 29108 11152
rect 29260 11117 29300 11656
rect 29452 11528 29492 12244
rect 29740 11957 29780 12328
rect 29739 11948 29781 11957
rect 29739 11908 29740 11948
rect 29780 11908 29781 11948
rect 29739 11899 29781 11908
rect 29643 11864 29685 11873
rect 29643 11824 29644 11864
rect 29684 11824 29685 11864
rect 29643 11815 29685 11824
rect 29644 11696 29684 11815
rect 29644 11647 29684 11656
rect 29740 11696 29780 11705
rect 29836 11696 29876 12487
rect 29780 11656 29876 11696
rect 29740 11647 29780 11656
rect 29452 11479 29492 11488
rect 29643 11528 29685 11537
rect 29643 11488 29644 11528
rect 29684 11488 29685 11528
rect 29643 11479 29685 11488
rect 29932 11528 29972 11537
rect 30028 11528 30068 12496
rect 30124 12536 30164 12547
rect 30124 12461 30164 12496
rect 30219 12536 30261 12545
rect 30219 12496 30220 12536
rect 30260 12496 30261 12536
rect 30219 12487 30261 12496
rect 30123 12452 30165 12461
rect 30123 12412 30124 12452
rect 30164 12412 30165 12452
rect 30123 12403 30165 12412
rect 30124 11873 30164 12403
rect 30220 12402 30260 12487
rect 30412 12377 30452 12748
rect 30411 12368 30453 12377
rect 30411 12328 30412 12368
rect 30452 12328 30453 12368
rect 30411 12319 30453 12328
rect 30123 11864 30165 11873
rect 30123 11824 30124 11864
rect 30164 11824 30165 11864
rect 30123 11815 30165 11824
rect 29972 11488 30068 11528
rect 30124 11696 30164 11705
rect 29932 11479 29972 11488
rect 29355 11360 29397 11369
rect 29355 11320 29356 11360
rect 29396 11320 29397 11360
rect 29355 11311 29397 11320
rect 29356 11192 29396 11311
rect 29356 11143 29396 11152
rect 29259 11108 29301 11117
rect 29644 11108 29684 11479
rect 30124 11201 30164 11656
rect 30220 11696 30260 11707
rect 30220 11621 30260 11656
rect 30412 11696 30452 11705
rect 30219 11612 30261 11621
rect 30219 11572 30220 11612
rect 30260 11572 30261 11612
rect 30219 11563 30261 11572
rect 30028 11192 30068 11201
rect 29259 11068 29260 11108
rect 29300 11068 29301 11108
rect 29259 11059 29301 11068
rect 29548 11068 29684 11108
rect 29068 10975 29108 10984
rect 29164 11024 29204 11033
rect 29355 11024 29397 11033
rect 28683 10856 28725 10865
rect 28683 10816 28684 10856
rect 28724 10816 28725 10856
rect 28683 10807 28725 10816
rect 28875 10856 28917 10865
rect 28875 10816 28876 10856
rect 28916 10816 28917 10856
rect 28875 10807 28917 10816
rect 29164 10529 29204 10984
rect 29260 10982 29300 10991
rect 29259 10942 29260 10949
rect 29355 10984 29356 11024
rect 29396 10984 29397 11024
rect 29355 10975 29397 10984
rect 29548 11024 29588 11068
rect 29836 11033 29876 11118
rect 29740 11024 29780 11033
rect 29548 10975 29588 10984
rect 29644 10982 29684 10991
rect 29300 10942 29301 10949
rect 29259 10940 29301 10942
rect 29259 10900 29260 10940
rect 29300 10900 29301 10940
rect 29259 10891 29301 10900
rect 29260 10847 29300 10891
rect 29163 10520 29205 10529
rect 29163 10480 29164 10520
rect 29204 10480 29205 10520
rect 29163 10471 29205 10480
rect 29356 10436 29396 10975
rect 29644 10781 29684 10942
rect 29643 10772 29685 10781
rect 29643 10732 29644 10772
rect 29684 10732 29685 10772
rect 29643 10723 29685 10732
rect 29547 10520 29589 10529
rect 29547 10480 29548 10520
rect 29588 10480 29589 10520
rect 29740 10520 29780 10984
rect 29835 11024 29877 11033
rect 29835 10984 29836 11024
rect 29876 10984 29877 11024
rect 29835 10975 29877 10984
rect 30028 10781 30068 11152
rect 30123 11192 30165 11201
rect 30123 11152 30124 11192
rect 30164 11152 30165 11192
rect 30123 11143 30165 11152
rect 30123 11024 30165 11033
rect 30123 10984 30124 11024
rect 30164 10984 30165 11024
rect 30123 10975 30165 10984
rect 30220 11024 30260 11563
rect 30315 11192 30357 11201
rect 30315 11152 30316 11192
rect 30356 11152 30357 11192
rect 30315 11143 30357 11152
rect 30220 10975 30260 10984
rect 30316 11024 30356 11143
rect 30316 10975 30356 10984
rect 30027 10772 30069 10781
rect 30027 10732 30028 10772
rect 30068 10732 30069 10772
rect 30027 10723 30069 10732
rect 29740 10480 29881 10520
rect 29547 10471 29589 10480
rect 29356 10387 29396 10396
rect 29164 10352 29204 10361
rect 29204 10312 29300 10352
rect 29164 10303 29204 10312
rect 27052 10050 27092 10135
rect 27153 10025 27193 10144
rect 27435 10184 27477 10193
rect 27435 10144 27436 10184
rect 27476 10144 27477 10184
rect 27435 10135 27477 10144
rect 28203 10184 28245 10193
rect 28203 10144 28204 10184
rect 28244 10144 28245 10184
rect 28203 10135 28245 10144
rect 28876 10184 28916 10195
rect 27152 10016 27194 10025
rect 27152 9976 27153 10016
rect 27193 9976 27194 10016
rect 27152 9967 27194 9976
rect 27339 9764 27381 9773
rect 27339 9724 27340 9764
rect 27380 9724 27381 9764
rect 27339 9715 27381 9724
rect 27340 9680 27380 9715
rect 27340 9629 27380 9640
rect 27435 9680 27477 9689
rect 27435 9640 27436 9680
rect 27476 9640 27477 9680
rect 27435 9631 27477 9640
rect 27819 9680 27861 9689
rect 27819 9640 27820 9680
rect 27860 9640 27861 9680
rect 27819 9631 27861 9640
rect 28204 9680 28244 10135
rect 28876 10109 28916 10144
rect 29068 10184 29108 10193
rect 28875 10100 28917 10109
rect 28875 10060 28876 10100
rect 28916 10060 28917 10100
rect 28875 10051 28917 10060
rect 28587 9932 28629 9941
rect 28587 9892 28588 9932
rect 28628 9892 28629 9932
rect 28587 9883 28629 9892
rect 28204 9631 28244 9640
rect 27244 9512 27284 9521
rect 27148 9472 27244 9512
rect 27148 8840 27188 9472
rect 27244 9463 27284 9472
rect 27436 9512 27476 9631
rect 27820 9546 27860 9631
rect 27436 9463 27476 9472
rect 27532 9512 27572 9521
rect 27339 8924 27381 8933
rect 27339 8884 27340 8924
rect 27380 8884 27381 8924
rect 27339 8875 27381 8884
rect 27148 8791 27188 8800
rect 27340 8765 27380 8875
rect 27339 8756 27381 8765
rect 27339 8716 27340 8756
rect 27380 8716 27381 8756
rect 27339 8707 27381 8716
rect 27051 8672 27093 8681
rect 27051 8632 27052 8672
rect 27092 8632 27093 8672
rect 27051 8623 27093 8632
rect 27148 8672 27188 8681
rect 27052 8538 27092 8623
rect 27148 8513 27188 8632
rect 27340 8672 27380 8707
rect 27243 8588 27285 8597
rect 27243 8548 27244 8588
rect 27284 8548 27285 8588
rect 27243 8539 27285 8548
rect 27147 8504 27189 8513
rect 27147 8464 27148 8504
rect 27188 8464 27189 8504
rect 27147 8455 27189 8464
rect 26956 8296 27092 8336
rect 26956 8168 26996 8177
rect 26860 8128 26956 8168
rect 26572 8119 26612 8128
rect 26956 8119 26996 8128
rect 26668 8009 26708 8094
rect 26667 8000 26709 8009
rect 26667 7960 26668 8000
rect 26708 7960 26804 8000
rect 26667 7951 26709 7960
rect 26667 7832 26709 7841
rect 26667 7792 26668 7832
rect 26708 7792 26709 7832
rect 26667 7783 26709 7792
rect 26571 7496 26613 7505
rect 26571 7456 26572 7496
rect 26612 7456 26613 7496
rect 26571 7447 26613 7456
rect 26420 7120 26516 7160
rect 26380 7111 26420 7120
rect 26476 6992 26516 7001
rect 26572 6992 26612 7447
rect 26668 7412 26708 7783
rect 26764 7673 26804 7960
rect 26763 7664 26805 7673
rect 26763 7624 26764 7664
rect 26804 7624 26805 7664
rect 26763 7615 26805 7624
rect 27052 7505 27092 8296
rect 27148 8000 27188 8009
rect 27148 7505 27188 7960
rect 27244 7589 27284 8539
rect 27340 8000 27380 8632
rect 27532 8429 27572 9472
rect 27916 9512 27956 9521
rect 27723 8840 27765 8849
rect 27723 8800 27724 8840
rect 27764 8800 27765 8840
rect 27723 8791 27765 8800
rect 27531 8420 27573 8429
rect 27531 8380 27532 8420
rect 27572 8380 27573 8420
rect 27531 8371 27573 8380
rect 27436 8000 27476 8009
rect 27340 7960 27436 8000
rect 27436 7951 27476 7960
rect 27243 7580 27285 7589
rect 27243 7540 27244 7580
rect 27284 7540 27285 7580
rect 27243 7531 27285 7540
rect 27051 7496 27093 7505
rect 27051 7456 27052 7496
rect 27092 7456 27093 7496
rect 27148 7496 27194 7505
rect 27148 7456 27153 7496
rect 27193 7456 27194 7496
rect 27051 7447 27093 7456
rect 27152 7447 27194 7456
rect 26668 7363 26708 7372
rect 27244 7328 27284 7531
rect 27141 7288 27284 7328
rect 27141 7244 27181 7288
rect 27052 7204 27181 7244
rect 26667 7160 26709 7169
rect 26667 7120 26668 7160
rect 26708 7120 26709 7160
rect 26667 7111 26709 7120
rect 26764 7160 26804 7169
rect 26668 7026 26708 7111
rect 26516 6952 26612 6992
rect 26476 6943 26516 6952
rect 26667 6908 26709 6917
rect 26667 6868 26668 6908
rect 26708 6868 26709 6908
rect 26667 6859 26709 6868
rect 25900 6784 26132 6824
rect 25900 6572 25940 6784
rect 25900 6523 25940 6532
rect 25996 6656 26036 6665
rect 25708 6488 25748 6497
rect 25611 6152 25653 6161
rect 25611 6112 25612 6152
rect 25652 6112 25653 6152
rect 25611 6103 25653 6112
rect 25611 5900 25653 5909
rect 25611 5860 25612 5900
rect 25652 5860 25653 5900
rect 25611 5851 25653 5860
rect 25612 5648 25652 5851
rect 25708 5825 25748 6448
rect 25804 6488 25844 6497
rect 25707 5816 25749 5825
rect 25707 5776 25708 5816
rect 25748 5776 25749 5816
rect 25707 5767 25749 5776
rect 25612 5599 25652 5608
rect 25611 5144 25653 5153
rect 25611 5104 25612 5144
rect 25652 5104 25653 5144
rect 25611 5095 25653 5104
rect 25516 4339 25556 4348
rect 25612 4220 25652 5095
rect 25707 5060 25749 5069
rect 25707 5020 25708 5060
rect 25748 5020 25749 5060
rect 25707 5011 25749 5020
rect 25708 4976 25748 5011
rect 25708 4925 25748 4936
rect 25804 4304 25844 6448
rect 25996 6404 26036 6616
rect 25900 6364 26036 6404
rect 25900 5153 25940 6364
rect 25995 6236 26037 6245
rect 25995 6196 25996 6236
rect 26036 6196 26037 6236
rect 25995 6187 26037 6196
rect 25996 6102 26036 6187
rect 25899 5144 25941 5153
rect 25899 5104 25900 5144
rect 25940 5104 25941 5144
rect 26092 5144 26132 6784
rect 26187 6824 26229 6833
rect 26187 6784 26188 6824
rect 26228 6784 26229 6824
rect 26187 6775 26229 6784
rect 26475 6824 26517 6833
rect 26475 6784 26476 6824
rect 26516 6784 26517 6824
rect 26475 6775 26517 6784
rect 26476 6572 26516 6775
rect 26571 6740 26613 6749
rect 26571 6700 26572 6740
rect 26612 6700 26613 6740
rect 26571 6691 26613 6700
rect 26572 6656 26612 6691
rect 26572 6581 26612 6616
rect 26476 6523 26516 6532
rect 26571 6572 26613 6581
rect 26571 6532 26572 6572
rect 26612 6532 26613 6572
rect 26571 6523 26613 6532
rect 26284 6488 26324 6499
rect 26284 6413 26324 6448
rect 26380 6488 26420 6497
rect 26572 6492 26612 6523
rect 26668 6497 26708 6859
rect 26764 6665 26804 7120
rect 26956 7160 26996 7169
rect 26859 7076 26901 7085
rect 26859 7036 26860 7076
rect 26900 7036 26901 7076
rect 26859 7027 26901 7036
rect 26763 6656 26805 6665
rect 26763 6616 26764 6656
rect 26804 6616 26805 6656
rect 26763 6607 26805 6616
rect 26283 6404 26325 6413
rect 26283 6364 26284 6404
rect 26324 6364 26325 6404
rect 26283 6355 26325 6364
rect 26284 5480 26324 5489
rect 26092 5104 26228 5144
rect 25899 5095 25941 5104
rect 25996 4976 26036 4985
rect 25516 4180 25652 4220
rect 25708 4264 25844 4304
rect 25900 4936 25996 4976
rect 25516 3968 25556 4180
rect 25708 4145 25748 4264
rect 25707 4136 25749 4145
rect 25707 4096 25708 4136
rect 25748 4096 25749 4136
rect 25707 4087 25749 4096
rect 25804 4136 25844 4145
rect 25611 4052 25653 4061
rect 25611 4012 25612 4052
rect 25652 4012 25653 4052
rect 25611 4003 25653 4012
rect 25228 3928 25364 3968
rect 25420 3928 25516 3968
rect 25131 3716 25173 3725
rect 25131 3676 25132 3716
rect 25172 3676 25173 3716
rect 25131 3667 25173 3676
rect 24940 3548 24980 3557
rect 24940 2624 24980 3508
rect 25132 3464 25172 3667
rect 25132 3415 25172 3424
rect 25228 2885 25268 3928
rect 25420 3464 25460 3928
rect 25516 3919 25556 3928
rect 25612 3918 25652 4003
rect 25708 4002 25748 4087
rect 25515 3800 25557 3809
rect 25515 3760 25516 3800
rect 25556 3760 25557 3800
rect 25515 3751 25557 3760
rect 25420 3389 25460 3424
rect 25419 3380 25461 3389
rect 25419 3340 25420 3380
rect 25460 3340 25461 3380
rect 25419 3331 25461 3340
rect 25420 3300 25460 3331
rect 25516 3128 25556 3751
rect 25804 3725 25844 4096
rect 25803 3716 25845 3725
rect 25612 3690 25804 3716
rect 25652 3676 25804 3690
rect 25844 3676 25845 3716
rect 25803 3667 25845 3676
rect 25612 3641 25652 3650
rect 25804 3464 25844 3473
rect 25708 3422 25748 3431
rect 25707 3382 25708 3389
rect 25748 3382 25749 3389
rect 25707 3380 25749 3382
rect 25707 3340 25708 3380
rect 25748 3340 25749 3380
rect 25707 3331 25749 3340
rect 25708 3287 25748 3331
rect 25515 3088 25556 3128
rect 25227 2876 25269 2885
rect 25227 2836 25228 2876
rect 25268 2836 25269 2876
rect 25515 2876 25555 3088
rect 25804 2885 25844 3424
rect 25803 2876 25845 2885
rect 25515 2836 25556 2876
rect 25227 2827 25269 2836
rect 25516 2792 25556 2836
rect 25803 2836 25804 2876
rect 25844 2836 25845 2876
rect 25803 2827 25845 2836
rect 25516 2743 25556 2752
rect 25420 2633 25460 2718
rect 25228 2624 25268 2633
rect 24940 2584 25228 2624
rect 25228 2575 25268 2584
rect 25419 2624 25461 2633
rect 25419 2584 25420 2624
rect 25460 2584 25461 2624
rect 25419 2575 25461 2584
rect 25708 2624 25748 2633
rect 25900 2624 25940 4936
rect 25996 4927 26036 4936
rect 26091 4976 26133 4985
rect 26091 4936 26092 4976
rect 26132 4936 26133 4976
rect 26091 4927 26133 4936
rect 26092 4842 26132 4927
rect 26188 4313 26228 5104
rect 26284 5069 26324 5440
rect 26380 5153 26420 6448
rect 26667 6488 26709 6497
rect 26860 6488 26900 7027
rect 26956 6656 26996 7120
rect 27052 7160 27092 7204
rect 27052 7111 27092 7120
rect 27206 7160 27248 7169
rect 27206 7120 27207 7160
rect 27247 7120 27248 7160
rect 27206 7111 27248 7120
rect 27207 7026 27247 7111
rect 27339 6824 27381 6833
rect 27339 6784 27340 6824
rect 27380 6784 27381 6824
rect 27339 6775 27381 6784
rect 27148 6656 27188 6665
rect 26956 6616 27148 6656
rect 27148 6607 27188 6616
rect 26667 6448 26668 6488
rect 26708 6448 26804 6488
rect 26667 6439 26709 6448
rect 26475 6320 26517 6329
rect 26475 6280 26476 6320
rect 26516 6280 26517 6320
rect 26475 6271 26517 6280
rect 26572 6320 26612 6329
rect 26667 6320 26709 6329
rect 26612 6280 26668 6320
rect 26708 6280 26709 6320
rect 26572 6271 26612 6280
rect 26667 6271 26709 6280
rect 26379 5144 26421 5153
rect 26379 5104 26380 5144
rect 26420 5104 26421 5144
rect 26379 5095 26421 5104
rect 26283 5060 26325 5069
rect 26283 5020 26284 5060
rect 26324 5020 26325 5060
rect 26283 5011 26325 5020
rect 26476 4976 26516 6271
rect 26668 5144 26708 5153
rect 26764 5144 26804 6448
rect 26860 6439 26900 6448
rect 26956 6488 26996 6497
rect 26956 6161 26996 6448
rect 27051 6488 27093 6497
rect 27051 6448 27052 6488
rect 27092 6448 27093 6488
rect 27051 6439 27093 6448
rect 26955 6152 26997 6161
rect 26955 6112 26956 6152
rect 26996 6112 26997 6152
rect 26955 6103 26997 6112
rect 27052 5732 27092 6439
rect 26956 5692 27092 5732
rect 26708 5104 26804 5144
rect 26860 5480 26900 5489
rect 26668 5095 26708 5104
rect 26476 4927 26516 4936
rect 26667 4976 26709 4985
rect 26667 4936 26668 4976
rect 26708 4936 26709 4976
rect 26667 4927 26709 4936
rect 26764 4976 26804 4985
rect 26860 4976 26900 5440
rect 26956 5480 26996 5692
rect 27143 5643 27183 5652
rect 26956 5431 26996 5440
rect 27052 5564 27092 5573
rect 27143 5564 27183 5603
rect 27244 5648 27284 5657
rect 27143 5524 27188 5564
rect 27052 5405 27092 5524
rect 27051 5396 27093 5405
rect 27051 5356 27052 5396
rect 27092 5356 27093 5396
rect 27051 5347 27093 5356
rect 27051 5144 27093 5153
rect 27051 5104 27052 5144
rect 27092 5104 27093 5144
rect 27051 5095 27093 5104
rect 26804 4936 26900 4976
rect 26764 4927 26804 4936
rect 26187 4304 26229 4313
rect 26187 4264 26188 4304
rect 26228 4264 26324 4304
rect 26187 4255 26229 4264
rect 25996 4136 26036 4145
rect 25996 3977 26036 4096
rect 26187 4136 26229 4145
rect 26187 4096 26188 4136
rect 26228 4096 26229 4136
rect 26187 4087 26229 4096
rect 26091 4052 26133 4061
rect 26091 4012 26092 4052
rect 26132 4012 26133 4052
rect 26091 4003 26133 4012
rect 25995 3968 26037 3977
rect 25995 3928 25996 3968
rect 26036 3928 26037 3968
rect 25995 3919 26037 3928
rect 26092 3918 26132 4003
rect 26188 4002 26228 4087
rect 25748 2584 25940 2624
rect 25708 2575 25748 2584
rect 25900 1952 25940 2584
rect 26092 3212 26132 3221
rect 25996 1952 26036 1961
rect 25900 1912 25996 1952
rect 24844 1903 24884 1912
rect 25996 1903 26036 1912
rect 24364 1231 24404 1240
rect 25228 1196 25268 1205
rect 25036 1156 25228 1196
rect 11884 1063 11924 1072
rect 23308 1063 23348 1072
rect 23979 1112 24021 1121
rect 23979 1072 23980 1112
rect 24020 1072 24021 1112
rect 23979 1063 24021 1072
rect 25036 1112 25076 1156
rect 25228 1147 25268 1156
rect 25036 1063 25076 1072
rect 25515 1112 25557 1121
rect 25515 1072 25516 1112
rect 25556 1072 25557 1112
rect 25515 1063 25557 1072
rect 25612 1112 25652 1121
rect 23980 978 24020 1063
rect 25516 978 25556 1063
rect 25612 953 25652 1072
rect 26092 1112 26132 3172
rect 26284 2633 26324 4264
rect 26668 4145 26708 4927
rect 26476 4136 26516 4145
rect 26476 3809 26516 4096
rect 26667 4136 26709 4145
rect 26667 4096 26668 4136
rect 26708 4096 26709 4136
rect 26860 4136 26900 4936
rect 26955 4976 26997 4985
rect 26955 4936 26956 4976
rect 26996 4936 26997 4976
rect 26955 4927 26997 4936
rect 26956 4842 26996 4927
rect 26956 4136 26996 4145
rect 26860 4096 26956 4136
rect 26667 4087 26709 4096
rect 26956 4087 26996 4096
rect 26668 4002 26708 4087
rect 26764 3968 26804 3977
rect 26571 3884 26613 3893
rect 26571 3844 26572 3884
rect 26612 3844 26613 3884
rect 26571 3835 26613 3844
rect 26475 3800 26517 3809
rect 26475 3760 26476 3800
rect 26516 3760 26517 3800
rect 26475 3751 26517 3760
rect 26572 3632 26612 3835
rect 26764 3725 26804 3928
rect 26859 3800 26901 3809
rect 26859 3760 26860 3800
rect 26900 3760 26901 3800
rect 26859 3751 26901 3760
rect 26763 3716 26805 3725
rect 26763 3676 26764 3716
rect 26804 3676 26805 3716
rect 26763 3667 26805 3676
rect 26572 3583 26612 3592
rect 26476 3464 26516 3473
rect 26379 3380 26421 3389
rect 26379 3340 26380 3380
rect 26420 3340 26421 3380
rect 26379 3331 26421 3340
rect 26380 2876 26420 3331
rect 26476 3212 26516 3424
rect 26667 3464 26709 3473
rect 26667 3424 26668 3464
rect 26708 3424 26709 3464
rect 26667 3415 26709 3424
rect 26668 3330 26708 3415
rect 26764 3212 26804 3667
rect 26860 3464 26900 3751
rect 26860 3415 26900 3424
rect 27052 3221 27092 5095
rect 27148 4817 27188 5524
rect 27244 4901 27284 5608
rect 27340 5405 27380 6775
rect 27627 5984 27669 5993
rect 27627 5944 27628 5984
rect 27668 5944 27669 5984
rect 27627 5935 27669 5944
rect 27339 5396 27381 5405
rect 27339 5356 27340 5396
rect 27380 5356 27381 5396
rect 27339 5347 27381 5356
rect 27340 5153 27380 5238
rect 27339 5144 27381 5153
rect 27339 5104 27340 5144
rect 27380 5104 27381 5144
rect 27339 5095 27381 5104
rect 27435 5060 27477 5069
rect 27435 5020 27436 5060
rect 27476 5020 27477 5060
rect 27435 5011 27477 5020
rect 27339 4976 27381 4985
rect 27339 4936 27340 4976
rect 27380 4936 27381 4976
rect 27339 4927 27381 4936
rect 27243 4892 27285 4901
rect 27243 4852 27244 4892
rect 27284 4852 27285 4892
rect 27243 4843 27285 4852
rect 27147 4808 27189 4817
rect 27147 4768 27148 4808
rect 27188 4768 27189 4808
rect 27147 4759 27189 4768
rect 27340 4808 27380 4927
rect 27436 4926 27476 5011
rect 27531 4976 27573 4985
rect 27531 4936 27532 4976
rect 27572 4936 27573 4976
rect 27531 4927 27573 4936
rect 27628 4976 27668 5935
rect 27628 4927 27668 4936
rect 27532 4842 27572 4927
rect 27340 4759 27380 4768
rect 27627 4808 27669 4817
rect 27627 4768 27628 4808
rect 27668 4768 27669 4808
rect 27627 4759 27669 4768
rect 27339 4136 27381 4145
rect 27339 4096 27340 4136
rect 27380 4096 27381 4136
rect 27339 4087 27381 4096
rect 27243 3968 27285 3977
rect 27243 3928 27244 3968
rect 27284 3928 27285 3968
rect 27243 3919 27285 3928
rect 27244 3464 27284 3919
rect 27340 3632 27380 4087
rect 27340 3583 27380 3592
rect 27532 3968 27572 3977
rect 27244 3415 27284 3424
rect 26476 3172 26804 3212
rect 27051 3212 27093 3221
rect 27051 3172 27052 3212
rect 27092 3172 27093 3212
rect 26380 2827 26420 2836
rect 26571 2876 26613 2885
rect 26571 2836 26572 2876
rect 26612 2836 26613 2876
rect 26571 2827 26613 2836
rect 26572 2742 26612 2827
rect 26283 2624 26325 2633
rect 26283 2584 26284 2624
rect 26324 2584 26325 2624
rect 26283 2575 26325 2584
rect 26668 2540 26708 3172
rect 27051 3163 27093 3172
rect 27244 2633 27284 2718
rect 27243 2624 27285 2633
rect 27243 2584 27244 2624
rect 27284 2584 27285 2624
rect 27243 2575 27285 2584
rect 27436 2624 27476 2633
rect 27532 2624 27572 3928
rect 27628 3809 27668 4759
rect 27627 3800 27669 3809
rect 27627 3760 27628 3800
rect 27668 3760 27669 3800
rect 27627 3751 27669 3760
rect 27628 3632 27668 3751
rect 27628 3583 27668 3592
rect 27476 2584 27572 2624
rect 27724 2624 27764 8791
rect 27916 8681 27956 9472
rect 28300 9512 28340 9521
rect 28300 9269 28340 9472
rect 28396 9512 28436 9521
rect 28299 9260 28341 9269
rect 28299 9220 28300 9260
rect 28340 9220 28341 9260
rect 28299 9211 28341 9220
rect 28396 8765 28436 9472
rect 28492 9512 28532 9521
rect 28492 8849 28532 9472
rect 28491 8840 28533 8849
rect 28491 8800 28492 8840
rect 28532 8800 28533 8840
rect 28491 8791 28533 8800
rect 28395 8756 28437 8765
rect 28395 8716 28396 8756
rect 28436 8716 28437 8756
rect 28395 8707 28437 8716
rect 27915 8672 27957 8681
rect 27915 8632 27916 8672
rect 27956 8632 27957 8672
rect 27915 8623 27957 8632
rect 27916 8345 27956 8623
rect 28396 8345 28436 8707
rect 27915 8336 27957 8345
rect 27915 8296 27916 8336
rect 27956 8296 27957 8336
rect 27915 8287 27957 8296
rect 28395 8336 28437 8345
rect 28395 8296 28396 8336
rect 28436 8296 28437 8336
rect 28395 8287 28437 8296
rect 28396 8168 28436 8177
rect 28588 8168 28628 9883
rect 28875 9680 28917 9689
rect 28875 9640 28876 9680
rect 28916 9640 28917 9680
rect 28875 9631 28917 9640
rect 28683 9512 28725 9521
rect 28683 9472 28684 9512
rect 28724 9472 28725 9512
rect 28683 9463 28725 9472
rect 28780 9512 28820 9521
rect 28684 9378 28724 9463
rect 28780 9353 28820 9472
rect 28876 9512 28916 9631
rect 29068 9521 29108 10144
rect 29163 10184 29205 10193
rect 29163 10144 29164 10184
rect 29204 10144 29205 10184
rect 29163 10135 29205 10144
rect 29164 10050 29204 10135
rect 29260 9764 29300 10312
rect 29355 10184 29397 10193
rect 29355 10144 29356 10184
rect 29396 10144 29397 10184
rect 29355 10135 29397 10144
rect 29452 10184 29492 10193
rect 29356 10050 29396 10135
rect 29452 9941 29492 10144
rect 29451 9932 29493 9941
rect 29451 9892 29452 9932
rect 29492 9892 29493 9932
rect 29451 9883 29493 9892
rect 29260 9724 29492 9764
rect 28876 9463 28916 9472
rect 28972 9512 29012 9521
rect 28779 9344 28821 9353
rect 28779 9304 28780 9344
rect 28820 9304 28821 9344
rect 28779 9295 28821 9304
rect 28972 9185 29012 9472
rect 29067 9512 29109 9521
rect 29067 9472 29068 9512
rect 29108 9472 29109 9512
rect 29067 9463 29109 9472
rect 29255 9512 29295 9521
rect 29255 9353 29295 9472
rect 29355 9512 29397 9521
rect 29355 9472 29356 9512
rect 29396 9472 29397 9512
rect 29355 9463 29397 9472
rect 29452 9512 29492 9724
rect 29548 9680 29588 10471
rect 29643 10436 29685 10445
rect 29643 10396 29644 10436
rect 29684 10396 29780 10436
rect 29643 10387 29685 10396
rect 29644 10184 29684 10193
rect 29644 9773 29684 10144
rect 29740 10142 29780 10396
rect 29841 10193 29881 10480
rect 30124 10445 30164 10975
rect 30412 10520 30452 11656
rect 30507 11192 30549 11201
rect 30507 11152 30508 11192
rect 30548 11152 30549 11192
rect 30507 11143 30549 11152
rect 30508 11024 30548 11143
rect 30508 10975 30548 10984
rect 30699 11024 30741 11033
rect 30699 10984 30700 11024
rect 30740 10984 30741 11024
rect 30699 10975 30741 10984
rect 30603 10940 30645 10949
rect 30603 10900 30604 10940
rect 30644 10900 30645 10940
rect 30603 10891 30645 10900
rect 30604 10806 30644 10891
rect 30700 10890 30740 10975
rect 30412 10480 30548 10520
rect 30123 10436 30165 10445
rect 30123 10396 30124 10436
rect 30164 10396 30165 10436
rect 30123 10387 30165 10396
rect 29840 10184 29882 10193
rect 29840 10144 29841 10184
rect 29881 10144 29882 10184
rect 29840 10135 29882 10144
rect 30124 10184 30164 10387
rect 30411 10268 30453 10277
rect 30411 10228 30412 10268
rect 30452 10228 30453 10268
rect 30411 10219 30453 10228
rect 30124 10135 30164 10144
rect 30412 10184 30452 10219
rect 29740 10093 29780 10102
rect 29841 10050 29881 10135
rect 30412 10133 30452 10144
rect 30315 10100 30357 10109
rect 30315 10060 30316 10100
rect 30356 10060 30357 10100
rect 30315 10051 30357 10060
rect 29739 10016 29781 10025
rect 29739 9976 29740 10016
rect 29780 9976 29781 10016
rect 29739 9967 29781 9976
rect 29643 9764 29685 9773
rect 29643 9724 29644 9764
rect 29684 9724 29685 9764
rect 29643 9715 29685 9724
rect 29548 9631 29588 9640
rect 29452 9463 29492 9472
rect 29643 9512 29685 9521
rect 29643 9472 29644 9512
rect 29684 9472 29685 9512
rect 29643 9463 29685 9472
rect 29740 9512 29780 9967
rect 30316 9966 30356 10051
rect 29835 9932 29877 9941
rect 29835 9892 29836 9932
rect 29876 9892 29877 9932
rect 29835 9883 29877 9892
rect 29740 9463 29780 9472
rect 29356 9378 29396 9463
rect 29547 9428 29589 9437
rect 29547 9388 29548 9428
rect 29588 9388 29589 9428
rect 29547 9379 29589 9388
rect 29254 9344 29296 9353
rect 29254 9304 29255 9344
rect 29295 9304 29296 9344
rect 29254 9295 29296 9304
rect 28971 9176 29013 9185
rect 28971 9136 28972 9176
rect 29012 9136 29013 9176
rect 28971 9127 29013 9136
rect 29163 9176 29205 9185
rect 29163 9136 29164 9176
rect 29204 9136 29205 9176
rect 29255 9176 29295 9295
rect 29255 9136 29396 9176
rect 29163 9127 29205 9136
rect 28780 8672 28820 8681
rect 28780 8252 28820 8632
rect 29067 8672 29109 8681
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 29164 8672 29204 9127
rect 29164 8623 29204 8632
rect 29068 8538 29108 8623
rect 28876 8504 28916 8513
rect 28960 8504 29000 8532
rect 29356 8504 29396 9136
rect 28916 8464 29012 8504
rect 28876 8455 28916 8464
rect 28972 8420 29012 8464
rect 29356 8455 29396 8464
rect 29548 8504 29588 9379
rect 29644 9378 29684 9463
rect 29836 8840 29876 9883
rect 30123 9764 30165 9773
rect 30123 9724 30124 9764
rect 30164 9724 30165 9764
rect 30123 9715 30165 9724
rect 29931 9680 29973 9689
rect 29931 9640 29932 9680
rect 29972 9640 29973 9680
rect 29931 9631 29973 9640
rect 29932 9521 29972 9631
rect 29931 9512 29973 9521
rect 29931 9472 29932 9512
rect 29972 9472 29973 9512
rect 29931 9463 29973 9472
rect 29932 9378 29972 9463
rect 30028 9428 30068 9437
rect 30028 9008 30068 9388
rect 30124 9344 30164 9715
rect 30508 9680 30548 10480
rect 30603 10352 30645 10361
rect 30603 10312 30604 10352
rect 30644 10312 30645 10352
rect 30603 10303 30645 10312
rect 30412 9640 30548 9680
rect 30604 9680 30644 10303
rect 30795 10268 30837 10277
rect 30795 10228 30796 10268
rect 30836 10228 30837 10268
rect 30795 10219 30837 10228
rect 30796 10184 30836 10219
rect 30796 10133 30836 10144
rect 30315 9596 30357 9605
rect 30315 9556 30316 9596
rect 30356 9556 30357 9596
rect 30315 9547 30357 9556
rect 30316 9512 30356 9547
rect 30316 9461 30356 9472
rect 30124 9295 30164 9304
rect 30220 9428 30260 9437
rect 30220 9101 30260 9388
rect 30219 9092 30261 9101
rect 30219 9052 30220 9092
rect 30260 9052 30261 9092
rect 30219 9043 30261 9052
rect 30028 8968 30164 9008
rect 30124 8924 30164 8968
rect 30124 8884 30356 8924
rect 30027 8840 30069 8849
rect 29836 8800 29972 8840
rect 29548 8455 29588 8464
rect 29740 8672 29780 8681
rect 28972 8380 29204 8420
rect 29067 8252 29109 8261
rect 28780 8212 29012 8252
rect 28436 8128 28628 8168
rect 28396 8119 28436 8128
rect 28875 8084 28917 8093
rect 28875 8044 28876 8084
rect 28916 8044 28917 8084
rect 28875 8035 28917 8044
rect 28108 8000 28148 8009
rect 28108 7841 28148 7960
rect 28204 8000 28244 8009
rect 28107 7832 28149 7841
rect 28107 7792 28108 7832
rect 28148 7792 28149 7832
rect 28107 7783 28149 7792
rect 28011 7580 28053 7589
rect 28011 7540 28012 7580
rect 28052 7540 28053 7580
rect 28011 7531 28053 7540
rect 28012 7160 28052 7531
rect 28204 7496 28244 7960
rect 28299 8000 28341 8009
rect 28299 7960 28300 8000
rect 28340 7960 28341 8000
rect 28299 7951 28341 7960
rect 28588 8000 28628 8009
rect 28300 7866 28340 7951
rect 28491 7916 28533 7925
rect 28588 7916 28628 7960
rect 28491 7876 28492 7916
rect 28532 7876 28628 7916
rect 28684 8000 28724 8009
rect 28491 7867 28533 7876
rect 28684 7505 28724 7960
rect 28780 8000 28820 8009
rect 28780 7841 28820 7960
rect 28876 7950 28916 8035
rect 28779 7832 28821 7841
rect 28972 7832 29012 8212
rect 29067 8212 29068 8252
rect 29108 8212 29109 8252
rect 29067 8203 29109 8212
rect 29068 8000 29108 8203
rect 29068 7951 29108 7960
rect 29164 7916 29204 8380
rect 29740 8345 29780 8632
rect 29836 8672 29876 8683
rect 29836 8597 29876 8632
rect 29835 8588 29877 8597
rect 29835 8548 29836 8588
rect 29876 8548 29877 8588
rect 29835 8539 29877 8548
rect 29739 8336 29781 8345
rect 29739 8296 29740 8336
rect 29780 8296 29781 8336
rect 29739 8287 29781 8296
rect 29259 8000 29301 8009
rect 29259 7960 29260 8000
rect 29300 7960 29301 8000
rect 29259 7951 29301 7960
rect 29452 8000 29492 8009
rect 29740 8000 29780 8009
rect 29164 7867 29204 7876
rect 28779 7792 28780 7832
rect 28820 7792 28821 7832
rect 28779 7783 28821 7792
rect 28876 7792 29012 7832
rect 29260 7832 29300 7951
rect 28779 7580 28821 7589
rect 28779 7540 28780 7580
rect 28820 7540 28821 7580
rect 28779 7531 28821 7540
rect 28683 7496 28725 7505
rect 28204 7456 28340 7496
rect 28012 7111 28052 7120
rect 28107 7160 28149 7169
rect 28107 7120 28108 7160
rect 28148 7120 28149 7160
rect 28107 7111 28149 7120
rect 28204 7160 28244 7169
rect 28108 6656 28148 7111
rect 28204 7001 28244 7120
rect 28203 6992 28245 7001
rect 28203 6952 28204 6992
rect 28244 6952 28245 6992
rect 28203 6943 28245 6952
rect 28300 6992 28340 7456
rect 28683 7456 28684 7496
rect 28724 7456 28725 7496
rect 28683 7447 28725 7456
rect 28684 7328 28724 7447
rect 28588 7288 28724 7328
rect 28492 7001 28532 7086
rect 28300 6943 28340 6952
rect 28491 6992 28533 7001
rect 28491 6952 28492 6992
rect 28532 6952 28533 6992
rect 28491 6943 28533 6952
rect 28588 6824 28628 7288
rect 28780 7253 28820 7531
rect 28779 7244 28821 7253
rect 28779 7204 28780 7244
rect 28820 7204 28821 7244
rect 28779 7195 28821 7204
rect 28683 7160 28725 7169
rect 28683 7120 28684 7160
rect 28724 7120 28725 7160
rect 28683 7111 28725 7120
rect 28780 7160 28820 7195
rect 28876 7169 28916 7792
rect 29260 7783 29300 7792
rect 29356 7916 29396 7925
rect 29356 7589 29396 7876
rect 29452 7757 29492 7960
rect 29644 7960 29740 8000
rect 29451 7748 29493 7757
rect 29451 7708 29452 7748
rect 29492 7708 29493 7748
rect 29451 7699 29493 7708
rect 29355 7580 29397 7589
rect 29355 7540 29356 7580
rect 29396 7540 29397 7580
rect 29355 7531 29397 7540
rect 28971 7496 29013 7505
rect 28971 7456 28972 7496
rect 29012 7456 29013 7496
rect 28971 7447 29013 7456
rect 28684 7026 28724 7111
rect 28780 7109 28820 7120
rect 28875 7160 28917 7169
rect 28875 7120 28876 7160
rect 28916 7120 28917 7160
rect 28875 7111 28917 7120
rect 28972 7160 29012 7447
rect 29260 7337 29300 7422
rect 29259 7328 29301 7337
rect 29259 7288 29260 7328
rect 29300 7288 29301 7328
rect 29259 7279 29301 7288
rect 29644 7244 29684 7960
rect 29740 7951 29780 7960
rect 29836 8000 29876 8009
rect 29836 7337 29876 7960
rect 29835 7328 29877 7337
rect 29835 7288 29836 7328
rect 29876 7288 29877 7328
rect 29835 7279 29877 7288
rect 29644 7195 29684 7204
rect 28972 7111 29012 7120
rect 29259 7160 29301 7169
rect 29259 7120 29260 7160
rect 29300 7120 29301 7160
rect 29259 7111 29301 7120
rect 29452 7160 29492 7171
rect 29260 7026 29300 7111
rect 29452 7085 29492 7120
rect 29739 7160 29781 7169
rect 29932 7160 29972 8800
rect 30027 8800 30028 8840
rect 30068 8800 30069 8840
rect 30027 8791 30069 8800
rect 30028 8420 30068 8791
rect 30124 8672 30164 8683
rect 30124 8597 30164 8632
rect 30123 8588 30165 8597
rect 30123 8548 30124 8588
rect 30164 8548 30165 8588
rect 30123 8539 30165 8548
rect 30028 8380 30164 8420
rect 30028 8000 30068 8009
rect 30028 7841 30068 7960
rect 30124 8000 30164 8380
rect 30220 8177 30260 8262
rect 30219 8168 30261 8177
rect 30219 8128 30220 8168
rect 30260 8128 30261 8168
rect 30219 8119 30261 8128
rect 30316 8000 30356 8884
rect 30124 7951 30164 7960
rect 30281 7985 30356 8000
rect 30321 7960 30356 7985
rect 30281 7841 30321 7945
rect 30027 7832 30069 7841
rect 30027 7792 30028 7832
rect 30068 7792 30069 7832
rect 30027 7783 30069 7792
rect 30280 7832 30322 7841
rect 30280 7792 30281 7832
rect 30321 7792 30322 7832
rect 30280 7783 30322 7792
rect 29739 7120 29740 7160
rect 29780 7120 29781 7160
rect 29739 7111 29781 7120
rect 29836 7120 29972 7160
rect 29451 7076 29493 7085
rect 29451 7036 29452 7076
rect 29492 7036 29493 7076
rect 29451 7027 29493 7036
rect 29740 7026 29780 7111
rect 28396 6784 28628 6824
rect 28300 6656 28340 6665
rect 28108 6616 28300 6656
rect 28300 6607 28340 6616
rect 28396 6488 28436 6784
rect 29067 6572 29109 6581
rect 29067 6532 29068 6572
rect 29108 6532 29109 6572
rect 29067 6523 29109 6532
rect 29451 6572 29493 6581
rect 29451 6532 29452 6572
rect 29492 6532 29493 6572
rect 29451 6523 29493 6532
rect 28396 6439 28436 6448
rect 28588 6488 28628 6497
rect 28299 6404 28341 6413
rect 28299 6364 28300 6404
rect 28340 6364 28341 6404
rect 28299 6355 28341 6364
rect 28203 6320 28245 6329
rect 28203 6280 28204 6320
rect 28244 6280 28245 6320
rect 28203 6271 28245 6280
rect 27820 5648 27860 5657
rect 27820 5489 27860 5608
rect 27916 5648 27956 5657
rect 28108 5648 28148 5657
rect 27956 5608 28108 5648
rect 28204 5648 28244 6271
rect 28300 5900 28340 6355
rect 28300 5851 28340 5860
rect 28300 5648 28340 5657
rect 28204 5608 28300 5648
rect 27916 5599 27956 5608
rect 28108 5599 28148 5608
rect 27819 5480 27861 5489
rect 27819 5440 27820 5480
rect 27860 5440 27861 5480
rect 27819 5431 27861 5440
rect 27820 5069 27860 5431
rect 27915 5144 27957 5153
rect 27915 5104 27916 5144
rect 27956 5104 27957 5144
rect 27915 5095 27957 5104
rect 27819 5060 27861 5069
rect 27819 5020 27820 5060
rect 27860 5020 27861 5060
rect 27819 5011 27861 5020
rect 27916 4976 27956 5095
rect 27916 3977 27956 4936
rect 28012 4976 28052 4985
rect 28012 4817 28052 4936
rect 28204 4976 28244 4987
rect 28300 4976 28340 5608
rect 28492 5648 28532 5657
rect 28396 5144 28436 5153
rect 28492 5144 28532 5608
rect 28588 5153 28628 6448
rect 28779 6488 28821 6497
rect 28779 6448 28780 6488
rect 28820 6448 28821 6488
rect 28779 6439 28821 6448
rect 28972 6488 29012 6499
rect 28780 6354 28820 6439
rect 28972 6413 29012 6448
rect 29068 6488 29108 6523
rect 28971 6404 29013 6413
rect 28971 6364 28972 6404
rect 29012 6364 29013 6404
rect 28971 6355 29013 6364
rect 28780 6236 28820 6245
rect 28683 5480 28725 5489
rect 28683 5440 28684 5480
rect 28724 5440 28725 5480
rect 28683 5431 28725 5440
rect 28436 5104 28532 5144
rect 28587 5144 28629 5153
rect 28587 5104 28588 5144
rect 28628 5104 28629 5144
rect 28396 5095 28436 5104
rect 28587 5095 28629 5104
rect 28588 4976 28628 4985
rect 28300 4936 28588 4976
rect 28204 4901 28244 4936
rect 28588 4927 28628 4936
rect 28684 4976 28724 5431
rect 28684 4927 28724 4936
rect 28203 4892 28245 4901
rect 28203 4852 28204 4892
rect 28244 4852 28245 4892
rect 28203 4843 28245 4852
rect 28011 4808 28053 4817
rect 28011 4768 28012 4808
rect 28052 4768 28053 4808
rect 28011 4759 28053 4768
rect 28204 4724 28244 4733
rect 28244 4684 28340 4724
rect 28204 4675 28244 4684
rect 28203 4136 28245 4145
rect 28203 4096 28204 4136
rect 28244 4096 28245 4136
rect 28203 4087 28245 4096
rect 28204 4002 28244 4087
rect 27915 3968 27957 3977
rect 27915 3928 27916 3968
rect 27956 3928 27957 3968
rect 27915 3919 27957 3928
rect 28300 3809 28340 4684
rect 28780 4145 28820 6196
rect 29068 4985 29108 6448
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 29260 6488 29300 6497
rect 29452 6488 29492 6523
rect 29300 6448 29396 6488
rect 29260 6439 29300 6448
rect 29164 5900 29204 6439
rect 29259 6236 29301 6245
rect 29259 6196 29260 6236
rect 29300 6196 29301 6236
rect 29259 6187 29301 6196
rect 29260 6102 29300 6187
rect 29356 6077 29396 6448
rect 29452 6437 29492 6448
rect 29739 6488 29781 6497
rect 29739 6448 29740 6488
rect 29780 6448 29781 6488
rect 29739 6439 29781 6448
rect 29740 6354 29780 6439
rect 29355 6068 29397 6077
rect 29355 6028 29356 6068
rect 29396 6028 29397 6068
rect 29355 6019 29397 6028
rect 29356 5900 29396 5909
rect 29164 5860 29356 5900
rect 29356 5851 29396 5860
rect 29164 5480 29204 5489
rect 29067 4976 29109 4985
rect 29067 4936 29068 4976
rect 29108 4936 29109 4976
rect 29067 4927 29109 4936
rect 29164 4976 29204 5440
rect 29164 4927 29204 4936
rect 29548 4976 29588 4985
rect 29548 4649 29588 4936
rect 29547 4640 29589 4649
rect 29547 4600 29548 4640
rect 29588 4600 29589 4640
rect 29547 4591 29589 4600
rect 29739 4640 29781 4649
rect 29739 4600 29740 4640
rect 29780 4600 29781 4640
rect 29739 4591 29781 4600
rect 29068 4304 29108 4313
rect 29108 4264 29396 4304
rect 29068 4255 29108 4264
rect 28396 4136 28436 4145
rect 28396 3893 28436 4096
rect 28779 4136 28821 4145
rect 28779 4096 28780 4136
rect 28820 4096 28821 4136
rect 28779 4087 28821 4096
rect 29259 4136 29301 4145
rect 29259 4096 29260 4136
rect 29300 4096 29301 4136
rect 29259 4087 29301 4096
rect 29260 4002 29300 4087
rect 28395 3884 28437 3893
rect 28395 3844 28396 3884
rect 28436 3844 28437 3884
rect 28395 3835 28437 3844
rect 28299 3800 28341 3809
rect 28299 3760 28300 3800
rect 28340 3760 28341 3800
rect 28299 3751 28341 3760
rect 29163 3800 29205 3809
rect 29163 3760 29164 3800
rect 29204 3760 29205 3800
rect 29163 3751 29205 3760
rect 28300 3464 28340 3473
rect 28300 2885 28340 3424
rect 28491 3464 28533 3473
rect 28491 3424 28492 3464
rect 28532 3424 28533 3464
rect 28491 3415 28533 3424
rect 28683 3464 28725 3473
rect 28683 3424 28684 3464
rect 28724 3424 28725 3464
rect 28683 3415 28725 3424
rect 29164 3464 29204 3751
rect 29164 3415 29204 3424
rect 29356 3464 29396 4264
rect 29740 4145 29780 4591
rect 29739 4136 29781 4145
rect 29739 4096 29740 4136
rect 29780 4096 29781 4136
rect 29739 4087 29781 4096
rect 29356 3415 29396 3424
rect 29740 3464 29780 4087
rect 29740 3415 29780 3424
rect 28492 3330 28532 3415
rect 28299 2876 28341 2885
rect 28299 2836 28300 2876
rect 28340 2836 28341 2876
rect 28299 2827 28341 2836
rect 27820 2624 27860 2652
rect 27724 2584 27820 2624
rect 27436 2575 27476 2584
rect 26668 2500 26804 2540
rect 26380 2456 26420 2465
rect 26284 1952 26324 1961
rect 26284 1364 26324 1912
rect 26284 1315 26324 1324
rect 26380 1280 26420 2416
rect 26572 2456 26612 2465
rect 26380 1240 26516 1280
rect 26092 1063 26132 1072
rect 26476 1112 26516 1240
rect 26572 1112 26612 2416
rect 26667 2036 26709 2045
rect 26667 1996 26668 2036
rect 26708 1996 26709 2036
rect 26667 1987 26709 1996
rect 26668 1952 26708 1987
rect 26668 1901 26708 1912
rect 26668 1112 26708 1121
rect 26572 1072 26668 1112
rect 26476 1063 26516 1072
rect 26668 1063 26708 1072
rect 26764 1112 26804 2500
rect 27724 2045 27764 2584
rect 27820 2575 27860 2584
rect 28684 2624 28724 3415
rect 29836 3053 29876 7120
rect 29932 6992 29972 7001
rect 30028 6992 30068 7783
rect 30123 7160 30165 7169
rect 30123 7120 30124 7160
rect 30164 7120 30165 7160
rect 30123 7111 30165 7120
rect 30220 7160 30260 7171
rect 30124 7026 30164 7111
rect 30220 7085 30260 7120
rect 30219 7076 30261 7085
rect 30219 7036 30220 7076
rect 30260 7036 30261 7076
rect 30219 7027 30261 7036
rect 29972 6952 30068 6992
rect 29932 6943 29972 6952
rect 29932 6572 29972 6581
rect 29972 6532 30260 6572
rect 29932 6523 29972 6532
rect 30220 6488 30260 6532
rect 30220 6439 30260 6448
rect 30027 6236 30069 6245
rect 30027 6196 30028 6236
rect 30068 6196 30069 6236
rect 30027 6187 30069 6196
rect 30028 5648 30068 6187
rect 30028 5599 30068 5608
rect 30219 5480 30261 5489
rect 30219 5440 30220 5480
rect 30260 5440 30261 5480
rect 30219 5431 30261 5440
rect 30220 5346 30260 5431
rect 30412 4976 30452 9640
rect 30604 9631 30644 9640
rect 30699 9596 30741 9605
rect 30699 9556 30700 9596
rect 30740 9556 30741 9596
rect 30699 9547 30741 9556
rect 30507 9512 30549 9521
rect 30507 9472 30508 9512
rect 30548 9472 30549 9512
rect 30507 9463 30549 9472
rect 30700 9512 30740 9547
rect 30508 9378 30548 9463
rect 30700 9461 30740 9472
rect 30795 8756 30837 8765
rect 30795 8716 30796 8756
rect 30836 8716 30837 8756
rect 30795 8707 30837 8716
rect 30699 8168 30741 8177
rect 30699 8128 30700 8168
rect 30740 8128 30741 8168
rect 30699 8119 30741 8128
rect 30796 8168 30836 8707
rect 30796 8119 30836 8128
rect 30507 8000 30549 8009
rect 30507 7960 30508 8000
rect 30548 7960 30549 8000
rect 30507 7951 30549 7960
rect 30604 8000 30644 8009
rect 30508 7866 30548 7951
rect 30604 7589 30644 7960
rect 30700 8000 30740 8119
rect 30700 7951 30740 7960
rect 30892 7925 30932 16024
rect 31084 11948 31124 18535
rect 31372 17744 31412 17753
rect 31468 17744 31508 18955
rect 31564 18425 31604 19132
rect 31660 18584 31700 19291
rect 31852 19013 31892 20056
rect 32331 20096 32373 20105
rect 32331 20056 32332 20096
rect 32372 20056 32373 20096
rect 32331 20047 32373 20056
rect 32332 19962 32372 20047
rect 31947 19844 31989 19853
rect 31947 19804 31948 19844
rect 31988 19804 31989 19844
rect 31947 19795 31989 19804
rect 31948 19710 31988 19795
rect 32812 19265 32852 22240
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 33772 21020 33812 22828
rect 33963 22532 34005 22541
rect 33963 22492 33964 22532
rect 34004 22492 34005 22532
rect 33963 22483 34005 22492
rect 33964 22398 34004 22483
rect 34348 21617 34388 23584
rect 34827 23575 34869 23584
rect 35020 23624 35060 23633
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 35020 23288 35060 23584
rect 35115 23372 35157 23381
rect 35115 23332 35116 23372
rect 35156 23332 35157 23372
rect 35115 23323 35157 23332
rect 34444 23248 35060 23288
rect 34444 22280 34484 23248
rect 35020 23120 35060 23129
rect 35020 22961 35060 23080
rect 35116 23120 35156 23323
rect 35116 23071 35156 23080
rect 35212 23120 35252 23920
rect 35788 23801 35828 24592
rect 35884 24632 35924 24643
rect 35980 24632 36020 25096
rect 36076 24632 36116 24641
rect 35980 24592 36076 24632
rect 35884 24557 35924 24592
rect 36076 24583 36116 24592
rect 35883 24548 35925 24557
rect 35883 24508 35884 24548
rect 35924 24508 35925 24548
rect 35883 24499 35925 24508
rect 36171 24548 36213 24557
rect 36171 24508 36172 24548
rect 36212 24508 36213 24548
rect 36171 24499 36213 24508
rect 36172 24414 36212 24499
rect 36268 23960 36308 26851
rect 36651 26816 36693 26825
rect 36651 26776 36652 26816
rect 36692 26776 36693 26816
rect 36651 26767 36693 26776
rect 36748 26816 36788 26825
rect 36940 26816 36980 27448
rect 37708 27404 37748 27413
rect 37708 27245 37748 27364
rect 38188 27245 38228 27616
rect 38284 27656 38324 27665
rect 37707 27236 37749 27245
rect 37707 27196 37708 27236
rect 37748 27196 37749 27236
rect 37707 27187 37749 27196
rect 38187 27236 38229 27245
rect 38187 27196 38188 27236
rect 38228 27196 38229 27236
rect 38187 27187 38229 27196
rect 37612 26816 37652 26825
rect 36788 26776 36980 26816
rect 37324 26776 37612 26816
rect 36748 26767 36788 26776
rect 36364 26732 36404 26743
rect 36364 26657 36404 26692
rect 36363 26648 36405 26657
rect 36363 26608 36364 26648
rect 36404 26608 36405 26648
rect 36363 26599 36405 26608
rect 36652 26060 36692 26767
rect 36652 26020 36788 26060
rect 36459 25976 36501 25985
rect 36459 25936 36460 25976
rect 36500 25936 36501 25976
rect 36459 25927 36501 25936
rect 36460 25304 36500 25927
rect 36652 25892 36692 25901
rect 36555 25808 36597 25817
rect 36555 25768 36556 25808
rect 36596 25768 36597 25808
rect 36555 25759 36597 25768
rect 36460 25255 36500 25264
rect 36556 24632 36596 25759
rect 36652 25313 36692 25852
rect 36651 25304 36693 25313
rect 36651 25264 36652 25304
rect 36692 25264 36693 25304
rect 36651 25255 36693 25264
rect 36748 25136 36788 26020
rect 36843 25976 36885 25985
rect 36843 25936 36844 25976
rect 36884 25936 36885 25976
rect 36843 25927 36885 25936
rect 36844 25842 36884 25927
rect 37324 25304 37364 26776
rect 37612 26767 37652 26776
rect 38284 26489 38324 27616
rect 38380 27656 38420 27691
rect 38380 27605 38420 27616
rect 38476 27656 38516 27665
rect 38283 26480 38325 26489
rect 38283 26440 38284 26480
rect 38324 26440 38325 26480
rect 38283 26431 38325 26440
rect 37364 25264 37460 25304
rect 37324 25255 37364 25264
rect 36748 25096 36884 25136
rect 36748 24632 36788 24641
rect 36556 24592 36748 24632
rect 36748 24583 36788 24592
rect 36844 24632 36884 25096
rect 36844 24305 36884 24592
rect 37228 24548 37268 24557
rect 36843 24296 36885 24305
rect 36843 24256 36844 24296
rect 36884 24256 36885 24296
rect 36843 24247 36885 24256
rect 37132 24044 37172 24053
rect 37228 24044 37268 24508
rect 37323 24548 37365 24557
rect 37323 24508 37324 24548
rect 37364 24508 37365 24548
rect 37323 24499 37365 24508
rect 37324 24414 37364 24499
rect 37172 24004 37268 24044
rect 37132 23995 37172 24004
rect 37420 23960 37460 25264
rect 36172 23920 36308 23960
rect 37324 23920 37460 23960
rect 37804 24632 37844 24641
rect 35692 23792 35732 23801
rect 35692 23297 35732 23752
rect 35787 23792 35829 23801
rect 35787 23752 35788 23792
rect 35828 23752 35829 23792
rect 35787 23743 35829 23752
rect 35788 23633 35828 23743
rect 35980 23708 36020 23717
rect 35787 23624 35829 23633
rect 35787 23584 35788 23624
rect 35828 23584 35829 23624
rect 35787 23575 35829 23584
rect 35787 23456 35829 23465
rect 35787 23416 35788 23456
rect 35828 23416 35829 23456
rect 35787 23407 35829 23416
rect 35691 23288 35733 23297
rect 35691 23248 35692 23288
rect 35732 23248 35733 23288
rect 35691 23239 35733 23248
rect 35788 23204 35828 23407
rect 35788 23155 35828 23164
rect 35883 23204 35925 23213
rect 35883 23164 35884 23204
rect 35924 23164 35925 23204
rect 35883 23155 35925 23164
rect 35212 23071 35252 23080
rect 35307 23120 35349 23129
rect 35307 23080 35308 23120
rect 35348 23080 35349 23120
rect 35307 23071 35349 23080
rect 35884 23120 35924 23155
rect 35308 22986 35348 23071
rect 35884 23069 35924 23080
rect 35691 23036 35733 23045
rect 35691 22996 35692 23036
rect 35732 22996 35733 23036
rect 35691 22987 35733 22996
rect 35019 22952 35061 22961
rect 35019 22912 35020 22952
rect 35060 22912 35061 22952
rect 35019 22903 35061 22912
rect 35499 22868 35541 22877
rect 35499 22828 35500 22868
rect 35540 22828 35541 22868
rect 35499 22819 35541 22828
rect 35500 22734 35540 22819
rect 34444 22231 34484 22240
rect 34828 22280 34868 22289
rect 35692 22280 35732 22987
rect 35980 22961 36020 23668
rect 36172 23120 36212 23920
rect 36748 23801 36788 23886
rect 36747 23792 36789 23801
rect 36652 23752 36748 23792
rect 36788 23752 36789 23792
rect 36555 23288 36597 23297
rect 36555 23248 36556 23288
rect 36596 23248 36597 23288
rect 36555 23239 36597 23248
rect 36556 23154 36596 23239
rect 36172 23071 36212 23080
rect 36459 23120 36501 23129
rect 36459 23080 36460 23120
rect 36500 23080 36501 23120
rect 36459 23071 36501 23080
rect 36652 23120 36692 23752
rect 36747 23743 36789 23752
rect 37228 23792 37268 23801
rect 37132 23624 37172 23633
rect 36652 23071 36692 23080
rect 36748 23584 37132 23624
rect 36748 23120 36788 23584
rect 37132 23575 37172 23584
rect 37131 23372 37173 23381
rect 37131 23332 37132 23372
rect 37172 23332 37173 23372
rect 37131 23323 37173 23332
rect 37132 23288 37172 23323
rect 37228 23297 37268 23752
rect 37132 23237 37172 23248
rect 37227 23288 37269 23297
rect 37227 23248 37228 23288
rect 37268 23248 37269 23288
rect 37227 23239 37269 23248
rect 36748 23071 36788 23080
rect 36843 23120 36885 23129
rect 36843 23080 36844 23120
rect 36884 23080 36885 23120
rect 36843 23071 36885 23080
rect 36460 22986 36500 23071
rect 35979 22952 36021 22961
rect 35979 22912 35980 22952
rect 36020 22912 36021 22952
rect 35979 22903 36021 22912
rect 36844 22532 36884 23071
rect 37324 23045 37364 23920
rect 37420 23792 37460 23801
rect 37420 23381 37460 23752
rect 37515 23792 37557 23801
rect 37515 23752 37516 23792
rect 37556 23752 37557 23792
rect 37515 23743 37557 23752
rect 37707 23792 37749 23801
rect 37707 23752 37708 23792
rect 37748 23752 37749 23792
rect 37707 23743 37749 23752
rect 37516 23658 37556 23743
rect 37708 23658 37748 23743
rect 37611 23624 37653 23633
rect 37611 23584 37612 23624
rect 37652 23584 37653 23624
rect 37611 23575 37653 23584
rect 37612 23490 37652 23575
rect 37804 23381 37844 24592
rect 38284 24627 38324 26431
rect 38476 26321 38516 27616
rect 38668 26993 38708 27952
rect 38763 27824 38805 27833
rect 38763 27784 38764 27824
rect 38804 27784 38805 27824
rect 38763 27775 38805 27784
rect 38955 27824 38997 27833
rect 38955 27784 38956 27824
rect 38996 27784 38997 27824
rect 38955 27775 38997 27784
rect 38764 27068 38804 27775
rect 38956 27656 38996 27775
rect 38956 27607 38996 27616
rect 39148 27413 39188 28288
rect 39436 28328 39476 28337
rect 40012 28333 40052 28342
rect 39476 28288 39572 28328
rect 39436 28279 39476 28288
rect 39147 27404 39189 27413
rect 39147 27364 39148 27404
rect 39188 27364 39189 27404
rect 39147 27355 39189 27364
rect 39532 27068 39572 28288
rect 39820 28160 39860 28169
rect 39627 27404 39669 27413
rect 39627 27364 39628 27404
rect 39668 27364 39669 27404
rect 39627 27355 39669 27364
rect 39628 27270 39668 27355
rect 39820 27161 39860 28120
rect 40012 28085 40052 28293
rect 40011 28076 40053 28085
rect 40011 28036 40012 28076
rect 40052 28036 40053 28076
rect 40011 28027 40053 28036
rect 39915 27656 39957 27665
rect 39915 27616 39916 27656
rect 39956 27616 39957 27656
rect 39915 27607 39957 27616
rect 40108 27656 40148 27665
rect 39916 27522 39956 27607
rect 39819 27152 39861 27161
rect 39819 27112 39820 27152
rect 39860 27112 39861 27152
rect 39819 27103 39861 27112
rect 39628 27068 39668 27077
rect 39532 27028 39628 27068
rect 38764 27019 38804 27028
rect 39628 27019 39668 27028
rect 38667 26984 38709 26993
rect 38667 26944 38668 26984
rect 38708 26944 38709 26984
rect 38667 26935 38709 26944
rect 40108 26825 40148 27616
rect 38956 26816 38996 26825
rect 38475 26312 38517 26321
rect 38475 26272 38476 26312
rect 38516 26272 38517 26312
rect 38475 26263 38517 26272
rect 38859 25724 38901 25733
rect 38859 25684 38860 25724
rect 38900 25684 38901 25724
rect 38859 25675 38901 25684
rect 38475 25388 38517 25397
rect 38475 25348 38476 25388
rect 38516 25348 38517 25388
rect 38475 25339 38517 25348
rect 38476 25254 38516 25339
rect 38860 25229 38900 25675
rect 38956 25481 38996 26776
rect 40107 26816 40149 26825
rect 40107 26776 40108 26816
rect 40148 26776 40149 26816
rect 40107 26767 40149 26776
rect 40299 26816 40341 26825
rect 40299 26776 40300 26816
rect 40340 26776 40341 26816
rect 40299 26767 40341 26776
rect 40300 26682 40340 26767
rect 39147 26228 39189 26237
rect 39147 26188 39148 26228
rect 39188 26188 39189 26228
rect 39147 26179 39189 26188
rect 39148 26094 39188 26179
rect 39339 26144 39381 26153
rect 39339 26099 39340 26144
rect 39380 26099 39381 26144
rect 39339 26095 39381 26099
rect 39819 26144 39861 26153
rect 39819 26104 39820 26144
rect 39860 26104 39861 26144
rect 39819 26095 39861 26104
rect 40299 26144 40341 26153
rect 40299 26104 40300 26144
rect 40340 26104 40341 26144
rect 40299 26095 40341 26104
rect 40396 26144 40436 34168
rect 40780 33704 40820 33713
rect 40588 33664 40780 33704
rect 40491 32948 40533 32957
rect 40588 32948 40628 33664
rect 40780 33655 40820 33664
rect 40491 32908 40492 32948
rect 40532 32908 40628 32948
rect 40684 32992 40916 33032
rect 40491 32899 40533 32908
rect 40492 32864 40532 32899
rect 40492 32814 40532 32824
rect 40684 32864 40724 32992
rect 40684 32815 40724 32824
rect 40779 32864 40821 32873
rect 40779 32824 40780 32864
rect 40820 32824 40821 32864
rect 40779 32815 40821 32824
rect 40587 32780 40629 32789
rect 40587 32740 40588 32780
rect 40628 32740 40629 32780
rect 40587 32731 40629 32740
rect 40588 32646 40628 32731
rect 40491 32276 40533 32285
rect 40491 32236 40492 32276
rect 40532 32236 40533 32276
rect 40491 32227 40533 32236
rect 40492 32192 40532 32227
rect 40492 30680 40532 32152
rect 40492 30631 40532 30640
rect 40588 31352 40628 31361
rect 40780 31352 40820 32815
rect 40628 31312 40820 31352
rect 40588 29840 40628 31312
rect 40876 30269 40916 32992
rect 40972 32285 41012 35167
rect 41068 35141 41108 36688
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 41452 35720 41492 35729
rect 41260 35216 41300 35225
rect 41067 35132 41109 35141
rect 41067 35092 41068 35132
rect 41108 35092 41109 35132
rect 41067 35083 41109 35092
rect 41260 35057 41300 35176
rect 41452 35141 41492 35680
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 42124 35216 42164 35225
rect 42028 35176 42124 35216
rect 41451 35132 41493 35141
rect 41451 35092 41452 35132
rect 41492 35092 41493 35132
rect 41451 35083 41493 35092
rect 41259 35048 41301 35057
rect 41259 35008 41260 35048
rect 41300 35008 41301 35048
rect 41259 34999 41301 35008
rect 41451 34628 41493 34637
rect 41451 34588 41452 34628
rect 41492 34588 41493 34628
rect 41451 34579 41493 34588
rect 41452 34494 41492 34579
rect 41644 34376 41684 34385
rect 41548 34336 41644 34376
rect 41163 34208 41205 34217
rect 41163 34168 41164 34208
rect 41204 34168 41205 34208
rect 41163 34159 41205 34168
rect 41164 33704 41204 34159
rect 41259 33788 41301 33797
rect 41259 33748 41260 33788
rect 41300 33748 41301 33788
rect 41259 33739 41301 33748
rect 41164 33655 41204 33664
rect 41067 33032 41109 33041
rect 41067 32992 41068 33032
rect 41108 32992 41109 33032
rect 41067 32983 41109 32992
rect 41068 32898 41108 32983
rect 41260 32864 41300 33739
rect 41355 33200 41397 33209
rect 41355 33160 41356 33200
rect 41396 33160 41397 33200
rect 41355 33151 41397 33160
rect 41260 32815 41300 32824
rect 41356 32864 41396 33151
rect 41451 32948 41493 32957
rect 41451 32908 41452 32948
rect 41492 32908 41493 32948
rect 41451 32899 41493 32908
rect 41356 32815 41396 32824
rect 41452 32864 41492 32899
rect 41452 32813 41492 32824
rect 41548 32864 41588 34336
rect 41644 34327 41684 34336
rect 41836 34376 41876 34385
rect 41739 34208 41781 34217
rect 41739 34168 41740 34208
rect 41780 34168 41781 34208
rect 41739 34159 41781 34168
rect 41740 34074 41780 34159
rect 41836 33797 41876 34336
rect 41932 34376 41972 34385
rect 41835 33788 41877 33797
rect 41835 33748 41836 33788
rect 41876 33748 41877 33788
rect 41835 33739 41877 33748
rect 41836 33452 41876 33461
rect 41548 32815 41588 32824
rect 41740 32864 41780 32873
rect 41836 32864 41876 33412
rect 41780 32824 41876 32864
rect 41740 32815 41780 32824
rect 41643 32780 41685 32789
rect 41643 32740 41644 32780
rect 41684 32740 41685 32780
rect 41643 32731 41685 32740
rect 40971 32276 41013 32285
rect 40971 32236 40972 32276
rect 41012 32236 41013 32276
rect 40971 32227 41013 32236
rect 40972 30848 41012 32227
rect 41451 32192 41493 32201
rect 41451 32152 41452 32192
rect 41492 32152 41493 32192
rect 41451 32143 41493 32152
rect 41452 32058 41492 32143
rect 41644 31016 41684 32731
rect 41932 32537 41972 34336
rect 42028 32873 42068 35176
rect 42124 35167 42164 35176
rect 44427 35216 44469 35225
rect 44427 35176 44428 35216
rect 44468 35176 44469 35216
rect 44427 35167 44469 35176
rect 45963 35216 46005 35225
rect 45963 35176 45964 35216
rect 46004 35176 46005 35216
rect 45963 35167 46005 35176
rect 44428 35082 44468 35167
rect 42891 34964 42933 34973
rect 42891 34924 42892 34964
rect 42932 34924 42933 34964
rect 42891 34915 42933 34924
rect 43276 34964 43316 34973
rect 42604 34544 42644 34553
rect 42123 34460 42165 34469
rect 42123 34420 42124 34460
rect 42164 34420 42165 34460
rect 42123 34411 42165 34420
rect 42124 34326 42164 34411
rect 42219 34376 42261 34385
rect 42219 34336 42220 34376
rect 42260 34336 42261 34376
rect 42219 34327 42261 34336
rect 42220 34242 42260 34327
rect 42123 33788 42165 33797
rect 42123 33748 42124 33788
rect 42164 33748 42165 33788
rect 42123 33739 42165 33748
rect 42124 33654 42164 33739
rect 42219 33116 42261 33125
rect 42219 33076 42220 33116
rect 42260 33076 42261 33116
rect 42219 33067 42261 33076
rect 42123 33032 42165 33041
rect 42123 32992 42124 33032
rect 42164 32992 42165 33032
rect 42123 32983 42165 32992
rect 42027 32864 42069 32873
rect 42027 32824 42028 32864
rect 42068 32824 42069 32864
rect 42027 32815 42069 32824
rect 42124 32864 42164 32983
rect 42124 32815 42164 32824
rect 42123 32696 42165 32705
rect 42123 32656 42124 32696
rect 42164 32656 42165 32696
rect 42123 32647 42165 32656
rect 41931 32528 41973 32537
rect 41931 32488 41932 32528
rect 41972 32488 41973 32528
rect 41931 32479 41973 32488
rect 42027 32444 42069 32453
rect 42027 32404 42028 32444
rect 42068 32404 42069 32444
rect 42027 32395 42069 32404
rect 41931 32360 41973 32369
rect 41931 32320 41932 32360
rect 41972 32320 41973 32360
rect 41931 32311 41973 32320
rect 41932 32192 41972 32311
rect 41836 32152 41932 32192
rect 41740 31193 41780 31278
rect 41739 31184 41781 31193
rect 41739 31144 41740 31184
rect 41780 31144 41781 31184
rect 41836 31184 41876 32152
rect 41932 32143 41972 32152
rect 42028 32192 42068 32395
rect 42124 32360 42164 32647
rect 42124 32311 42164 32320
rect 42028 32143 42068 32152
rect 42220 32192 42260 33067
rect 42412 32192 42452 32201
rect 42220 32143 42260 32152
rect 42316 32152 42412 32192
rect 42028 31604 42068 31613
rect 42316 31604 42356 32152
rect 42412 32143 42452 32152
rect 42508 32192 42548 32201
rect 42508 32033 42548 32152
rect 42507 32024 42549 32033
rect 42507 31984 42508 32024
rect 42548 31984 42549 32024
rect 42507 31975 42549 31984
rect 42068 31564 42356 31604
rect 42028 31555 42068 31564
rect 41932 31352 41972 31361
rect 41972 31312 42068 31352
rect 41932 31303 41972 31312
rect 41836 31144 41972 31184
rect 41739 31135 41781 31144
rect 41644 30976 41780 31016
rect 40972 30799 41012 30808
rect 41644 30680 41684 30689
rect 40875 30260 40917 30269
rect 40875 30220 40876 30260
rect 40916 30220 40917 30260
rect 40875 30211 40917 30220
rect 41259 30260 41301 30269
rect 41259 30220 41260 30260
rect 41300 30220 41301 30260
rect 41259 30211 41301 30220
rect 40972 29840 41012 29849
rect 40588 29800 40972 29840
rect 40972 29791 41012 29800
rect 41067 29756 41109 29765
rect 41067 29716 41068 29756
rect 41108 29716 41109 29756
rect 41067 29707 41109 29716
rect 40876 29093 40916 29095
rect 40875 29084 40917 29093
rect 40875 29044 40876 29084
rect 40916 29044 40917 29084
rect 40875 29035 40917 29044
rect 40876 29000 40916 29035
rect 40876 28951 40916 28960
rect 41068 28412 41108 29707
rect 41260 29336 41300 30211
rect 41644 29765 41684 30640
rect 41740 30680 41780 30976
rect 41740 30631 41780 30640
rect 41836 30680 41876 30689
rect 41836 30269 41876 30640
rect 41932 30680 41972 31144
rect 41932 30631 41972 30640
rect 41835 30260 41877 30269
rect 41835 30220 41836 30260
rect 41876 30220 41877 30260
rect 41835 30211 41877 30220
rect 42028 30017 42068 31312
rect 42220 31184 42260 31193
rect 42220 30764 42260 31144
rect 42220 30715 42260 30724
rect 42604 30680 42644 34504
rect 42892 34385 42932 34915
rect 43276 34721 43316 34924
rect 43755 34964 43797 34973
rect 43755 34924 43756 34964
rect 43796 34924 43797 34964
rect 43755 34915 43797 34924
rect 43756 34830 43796 34915
rect 43275 34712 43317 34721
rect 43275 34672 43276 34712
rect 43316 34672 43317 34712
rect 43275 34663 43317 34672
rect 43660 34544 43700 34553
rect 42796 34376 42836 34385
rect 42796 33788 42836 34336
rect 42891 34376 42933 34385
rect 42891 34336 42892 34376
rect 42932 34336 42933 34376
rect 42891 34327 42933 34336
rect 42988 34376 43028 34385
rect 42892 34242 42932 34327
rect 42700 33748 42932 33788
rect 42700 33629 42740 33748
rect 42892 33704 42932 33748
rect 42892 33655 42932 33664
rect 42699 33620 42741 33629
rect 42699 33580 42700 33620
rect 42740 33580 42741 33620
rect 42699 33571 42741 33580
rect 42700 32453 42740 33571
rect 42988 33041 43028 34336
rect 43084 34208 43124 34217
rect 43084 33125 43124 34168
rect 43371 34208 43413 34217
rect 43371 34168 43372 34208
rect 43412 34168 43413 34208
rect 43371 34159 43413 34168
rect 43372 33704 43412 34159
rect 43372 33655 43412 33664
rect 43564 33704 43604 33713
rect 43660 33704 43700 34504
rect 44524 34376 44564 34385
rect 43851 34208 43893 34217
rect 43851 34168 43852 34208
rect 43892 34168 43893 34208
rect 43851 34159 43893 34168
rect 43852 34074 43892 34159
rect 43948 33704 43988 33713
rect 43660 33664 43948 33704
rect 43276 33452 43316 33461
rect 43083 33116 43125 33125
rect 43083 33076 43084 33116
rect 43124 33076 43125 33116
rect 43083 33067 43125 33076
rect 42987 33032 43029 33041
rect 42987 32992 42988 33032
rect 43028 32992 43029 33032
rect 42987 32983 43029 32992
rect 43083 32948 43125 32957
rect 43083 32908 43084 32948
rect 43124 32908 43125 32948
rect 43083 32899 43125 32908
rect 42987 32864 43029 32873
rect 42987 32824 42988 32864
rect 43028 32824 43029 32864
rect 42987 32815 43029 32824
rect 42988 32730 43028 32815
rect 43084 32612 43124 32899
rect 42988 32572 43124 32612
rect 42699 32444 42741 32453
rect 42699 32404 42700 32444
rect 42740 32404 42741 32444
rect 42699 32395 42741 32404
rect 42700 32192 42740 32201
rect 42892 32192 42932 32201
rect 42740 32152 42892 32192
rect 42700 32143 42740 32152
rect 42892 32143 42932 32152
rect 42988 32192 43028 32572
rect 43276 32369 43316 33412
rect 43564 32789 43604 33664
rect 43948 33655 43988 33664
rect 44524 33209 44564 34336
rect 45964 33872 46004 35167
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 45964 33823 46004 33832
rect 44812 33704 44852 33713
rect 44716 33664 44812 33704
rect 44139 33200 44181 33209
rect 44139 33160 44140 33200
rect 44180 33160 44181 33200
rect 44139 33151 44181 33160
rect 44523 33200 44565 33209
rect 44523 33160 44524 33200
rect 44564 33160 44565 33200
rect 44523 33151 44565 33160
rect 44140 33116 44180 33151
rect 44140 33065 44180 33076
rect 44716 32873 44756 33664
rect 44812 33655 44852 33664
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 44812 33032 44852 33041
rect 47884 33032 47924 33041
rect 44852 32992 45140 33032
rect 44812 32983 44852 32992
rect 43947 32864 43989 32873
rect 43947 32824 43948 32864
rect 43988 32824 43989 32864
rect 43947 32815 43989 32824
rect 44715 32864 44757 32873
rect 44715 32824 44716 32864
rect 44756 32824 44757 32864
rect 44715 32815 44757 32824
rect 43563 32780 43605 32789
rect 43563 32740 43564 32780
rect 43604 32740 43605 32780
rect 43563 32731 43605 32740
rect 43275 32360 43317 32369
rect 43275 32320 43276 32360
rect 43316 32320 43317 32360
rect 43275 32311 43317 32320
rect 43948 32360 43988 32815
rect 45004 32696 45044 32705
rect 43948 32311 43988 32320
rect 44716 32656 45004 32696
rect 43467 32276 43509 32285
rect 43467 32236 43468 32276
rect 43508 32236 43509 32276
rect 43467 32227 43509 32236
rect 44716 32276 44756 32656
rect 45004 32647 45044 32656
rect 44716 32227 44756 32236
rect 42700 31940 42740 31949
rect 42740 31900 42932 31940
rect 42700 31891 42740 31900
rect 42892 31352 42932 31900
rect 42988 31445 43028 32152
rect 43084 32192 43124 32201
rect 43084 31529 43124 32152
rect 43180 32192 43220 32201
rect 43180 32033 43220 32152
rect 43468 32192 43508 32227
rect 43468 32141 43508 32152
rect 44139 32192 44181 32201
rect 44139 32152 44140 32192
rect 44180 32152 44181 32192
rect 44139 32143 44181 32152
rect 45100 32192 45140 32992
rect 45100 32143 45140 32152
rect 45676 32864 45716 32873
rect 43179 32024 43221 32033
rect 43179 31984 43180 32024
rect 43220 31984 43221 32024
rect 43179 31975 43221 31984
rect 43083 31520 43125 31529
rect 43083 31480 43084 31520
rect 43124 31480 43125 31520
rect 43083 31471 43125 31480
rect 42987 31436 43029 31445
rect 42987 31396 42988 31436
rect 43028 31396 43029 31436
rect 42987 31387 43029 31396
rect 43180 31361 43220 31975
rect 43371 31436 43413 31445
rect 43371 31396 43372 31436
rect 43412 31396 43413 31436
rect 43371 31387 43413 31396
rect 42892 31303 42932 31312
rect 43084 31352 43124 31361
rect 43084 31193 43124 31312
rect 43179 31352 43221 31361
rect 43179 31312 43180 31352
rect 43220 31312 43221 31352
rect 43179 31303 43221 31312
rect 43372 31193 43412 31387
rect 43083 31184 43125 31193
rect 43083 31144 43084 31184
rect 43124 31144 43125 31184
rect 43083 31135 43125 31144
rect 43371 31184 43413 31193
rect 43371 31144 43372 31184
rect 43412 31144 43413 31184
rect 43371 31135 43413 31144
rect 43756 31184 43796 31193
rect 43948 31184 43988 31193
rect 42604 30631 42644 30640
rect 43179 30596 43221 30605
rect 43179 30556 43180 30596
rect 43220 30556 43221 30596
rect 43179 30547 43221 30556
rect 42027 30008 42069 30017
rect 42027 29968 42028 30008
rect 42068 29968 42069 30008
rect 42027 29959 42069 29968
rect 42315 30008 42357 30017
rect 42315 29968 42316 30008
rect 42356 29968 42357 30008
rect 42315 29959 42357 29968
rect 42124 29924 42164 29935
rect 42124 29849 42164 29884
rect 42316 29874 42356 29959
rect 42123 29840 42165 29849
rect 42123 29800 42124 29840
rect 42164 29800 42165 29840
rect 42123 29791 42165 29800
rect 42987 29840 43029 29849
rect 42987 29800 42988 29840
rect 43028 29800 43029 29840
rect 42987 29791 43029 29800
rect 43180 29840 43220 30547
rect 43180 29791 43220 29800
rect 43276 29840 43316 29851
rect 41643 29756 41685 29765
rect 41643 29716 41644 29756
rect 41684 29716 41685 29756
rect 41643 29707 41685 29716
rect 41835 29756 41877 29765
rect 41835 29716 41836 29756
rect 41876 29716 41877 29756
rect 41835 29707 41877 29716
rect 41355 29672 41397 29681
rect 41355 29632 41356 29672
rect 41396 29632 41397 29672
rect 41355 29623 41397 29632
rect 41260 29261 41300 29296
rect 41259 29252 41301 29261
rect 41259 29212 41260 29252
rect 41300 29212 41301 29252
rect 41259 29203 41301 29212
rect 41260 29172 41300 29203
rect 41068 28363 41108 28372
rect 40491 28328 40533 28337
rect 40491 28288 40492 28328
rect 40532 28288 40533 28328
rect 40491 28279 40533 28288
rect 40972 28328 41012 28337
rect 41356 28328 41396 29623
rect 41643 29252 41685 29261
rect 41643 29212 41644 29252
rect 41684 29212 41685 29252
rect 41643 29203 41685 29212
rect 41644 29168 41684 29203
rect 41644 29117 41684 29128
rect 41740 29093 41780 29178
rect 41836 29168 41876 29707
rect 42988 29706 43028 29791
rect 43276 29765 43316 29800
rect 43372 29840 43412 31135
rect 43756 31025 43796 31144
rect 43852 31144 43948 31184
rect 43755 31016 43797 31025
rect 43755 30976 43756 31016
rect 43796 30976 43797 31016
rect 43755 30967 43797 30976
rect 43468 30680 43508 30689
rect 43468 29849 43508 30640
rect 43563 30680 43605 30689
rect 43563 30640 43564 30680
rect 43604 30640 43605 30680
rect 43563 30631 43605 30640
rect 43275 29756 43317 29765
rect 43275 29716 43276 29756
rect 43316 29716 43317 29756
rect 43275 29707 43317 29716
rect 43372 29681 43412 29800
rect 43467 29840 43509 29849
rect 43467 29800 43468 29840
rect 43508 29800 43509 29840
rect 43467 29791 43509 29800
rect 42507 29672 42549 29681
rect 42507 29632 42508 29672
rect 42548 29632 42549 29672
rect 42507 29623 42549 29632
rect 43371 29672 43413 29681
rect 43371 29632 43372 29672
rect 43412 29632 43413 29672
rect 43371 29623 43413 29632
rect 43468 29672 43508 29681
rect 43564 29672 43604 30631
rect 43659 30428 43701 30437
rect 43659 30388 43660 30428
rect 43700 30388 43701 30428
rect 43659 30379 43701 30388
rect 43660 29840 43700 30379
rect 43660 29791 43700 29800
rect 43508 29632 43604 29672
rect 43468 29623 43508 29632
rect 42508 29336 42548 29623
rect 43852 29504 43892 31144
rect 43948 31135 43988 31144
rect 42988 29464 43892 29504
rect 42508 29287 42548 29296
rect 42891 29336 42933 29345
rect 42891 29296 42892 29336
rect 42932 29296 42933 29336
rect 42891 29287 42933 29296
rect 41836 29119 41876 29128
rect 42892 29168 42932 29287
rect 41452 29084 41492 29093
rect 41452 28496 41492 29044
rect 41739 29084 41781 29093
rect 41739 29044 41740 29084
rect 41780 29044 41781 29084
rect 41739 29035 41781 29044
rect 42220 28496 42260 28507
rect 41452 28456 41780 28496
rect 41452 28328 41492 28337
rect 41356 28288 41452 28328
rect 40492 28194 40532 28279
rect 40972 27749 41012 28288
rect 41452 28279 41492 28288
rect 41548 28328 41588 28337
rect 41740 28328 41780 28456
rect 42220 28421 42260 28456
rect 42219 28412 42261 28421
rect 42219 28372 42220 28412
rect 42260 28372 42261 28412
rect 42219 28363 42261 28372
rect 41932 28328 41972 28337
rect 41740 28288 41932 28328
rect 40971 27740 41013 27749
rect 40971 27700 40972 27740
rect 41012 27700 41013 27740
rect 40971 27691 41013 27700
rect 40684 26648 40724 26657
rect 40684 26489 40724 26608
rect 41548 26489 41588 28288
rect 41739 27404 41781 27413
rect 41739 27364 41740 27404
rect 41780 27364 41781 27404
rect 41739 27355 41781 27364
rect 41740 26816 41780 27355
rect 41932 26825 41972 28288
rect 42892 28001 42932 29128
rect 42891 27992 42933 28001
rect 42891 27952 42892 27992
rect 42932 27952 42933 27992
rect 42891 27943 42933 27952
rect 42891 27824 42933 27833
rect 42891 27784 42892 27824
rect 42932 27784 42933 27824
rect 42891 27775 42933 27784
rect 42892 27690 42932 27775
rect 42988 27656 43028 29464
rect 44043 29252 44085 29261
rect 44043 29212 44044 29252
rect 44084 29212 44085 29252
rect 44043 29203 44085 29212
rect 43275 29168 43317 29177
rect 43275 29128 43276 29168
rect 43316 29128 43317 29168
rect 43275 29119 43317 29128
rect 43179 28496 43221 28505
rect 43179 28456 43180 28496
rect 43220 28456 43221 28496
rect 43179 28447 43221 28456
rect 43180 28328 43220 28447
rect 43180 28279 43220 28288
rect 43084 28169 43124 28254
rect 43083 28160 43125 28169
rect 43083 28120 43084 28160
rect 43124 28120 43125 28160
rect 43083 28111 43125 28120
rect 43276 27992 43316 29119
rect 43467 29084 43509 29093
rect 43467 29044 43468 29084
rect 43508 29044 43509 29084
rect 43467 29035 43509 29044
rect 43371 28328 43413 28337
rect 43371 28288 43372 28328
rect 43412 28288 43413 28328
rect 43371 28279 43413 28288
rect 43468 28328 43508 29035
rect 43563 28412 43605 28421
rect 43563 28372 43564 28412
rect 43604 28372 43605 28412
rect 43563 28363 43605 28372
rect 43468 28279 43508 28288
rect 43564 28328 43604 28363
rect 43660 28337 43700 28422
rect 44044 28342 44084 29203
rect 44140 29168 44180 32143
rect 45100 31529 45140 31614
rect 45676 31529 45716 32824
rect 45963 32864 46005 32873
rect 45963 32824 45964 32864
rect 46004 32824 46005 32864
rect 45963 32815 46005 32824
rect 47692 32864 47732 32873
rect 45964 32192 46004 32815
rect 46539 32696 46581 32705
rect 46539 32656 46540 32696
rect 46580 32656 46581 32696
rect 46539 32647 46581 32656
rect 47019 32696 47061 32705
rect 47019 32656 47020 32696
rect 47060 32656 47061 32696
rect 47019 32647 47061 32656
rect 45964 32143 46004 32152
rect 45771 31940 45813 31949
rect 45771 31900 45772 31940
rect 45812 31900 45813 31940
rect 45771 31891 45813 31900
rect 44619 31520 44661 31529
rect 44619 31480 44620 31520
rect 44660 31480 44661 31520
rect 44619 31471 44661 31480
rect 45099 31520 45141 31529
rect 45099 31480 45100 31520
rect 45140 31480 45141 31520
rect 45099 31471 45141 31480
rect 45675 31520 45717 31529
rect 45675 31480 45676 31520
rect 45716 31480 45717 31520
rect 45675 31471 45717 31480
rect 44620 31352 44660 31471
rect 44620 30848 44660 31312
rect 44812 31352 44852 31363
rect 44812 31277 44852 31312
rect 44907 31352 44949 31361
rect 44907 31312 44908 31352
rect 44948 31312 44949 31352
rect 44907 31303 44949 31312
rect 45099 31352 45141 31361
rect 45099 31312 45100 31352
rect 45140 31312 45141 31352
rect 45099 31303 45141 31312
rect 45292 31352 45332 31361
rect 44811 31268 44853 31277
rect 44811 31228 44812 31268
rect 44852 31228 44853 31268
rect 44811 31219 44853 31228
rect 44908 31218 44948 31303
rect 45100 31218 45140 31303
rect 45292 31025 45332 31312
rect 45579 31352 45621 31361
rect 45579 31312 45580 31352
rect 45620 31312 45621 31352
rect 45579 31303 45621 31312
rect 45676 31352 45716 31361
rect 45387 31268 45429 31277
rect 45387 31228 45388 31268
rect 45428 31228 45429 31268
rect 45387 31219 45429 31228
rect 45388 31134 45428 31219
rect 45580 31218 45620 31303
rect 45676 31193 45716 31312
rect 45772 31352 45812 31891
rect 46444 31520 46484 31531
rect 46444 31445 46484 31480
rect 45867 31436 45909 31445
rect 45867 31396 45868 31436
rect 45908 31396 45909 31436
rect 45867 31387 45909 31396
rect 46443 31436 46485 31445
rect 46443 31396 46444 31436
rect 46484 31396 46485 31436
rect 46443 31387 46485 31396
rect 45772 31303 45812 31312
rect 45868 31352 45908 31387
rect 45868 31301 45908 31312
rect 46252 31352 46292 31361
rect 45675 31184 45717 31193
rect 45675 31144 45676 31184
rect 45716 31144 45717 31184
rect 45675 31135 45717 31144
rect 45291 31016 45333 31025
rect 45291 30976 45292 31016
rect 45332 30976 45333 31016
rect 45291 30967 45333 30976
rect 44620 30799 44660 30808
rect 45004 30689 45044 30774
rect 46252 30689 46292 31312
rect 44811 30680 44853 30689
rect 44811 30640 44812 30680
rect 44852 30640 44853 30680
rect 44811 30631 44853 30640
rect 45003 30680 45045 30689
rect 45003 30640 45004 30680
rect 45044 30640 45045 30680
rect 45003 30631 45045 30640
rect 45100 30680 45140 30689
rect 46251 30680 46293 30689
rect 45140 30640 45236 30680
rect 45100 30631 45140 30640
rect 44812 30546 44852 30631
rect 44907 30512 44949 30521
rect 44907 30472 44908 30512
rect 44948 30472 44949 30512
rect 44907 30463 44949 30472
rect 44811 30428 44853 30437
rect 44811 30388 44812 30428
rect 44852 30388 44853 30428
rect 44811 30379 44853 30388
rect 44812 30294 44852 30379
rect 44908 29840 44948 30463
rect 44908 29791 44948 29800
rect 45099 29840 45141 29849
rect 45099 29800 45100 29840
rect 45140 29800 45141 29840
rect 45099 29791 45141 29800
rect 44332 29756 44372 29765
rect 44524 29756 44564 29765
rect 44372 29716 44524 29756
rect 44332 29707 44372 29716
rect 44524 29707 44564 29716
rect 45100 29336 45140 29791
rect 45100 29287 45140 29296
rect 44620 29168 44660 29177
rect 44180 29128 44620 29168
rect 44140 29119 44180 29128
rect 44620 29119 44660 29128
rect 45196 29000 45236 30640
rect 46251 30640 46252 30680
rect 46292 30640 46293 30680
rect 46251 30631 46293 30640
rect 46540 30680 46580 32647
rect 47020 32562 47060 32647
rect 47692 32369 47732 32824
rect 47115 32360 47157 32369
rect 47115 32320 47116 32360
rect 47156 32320 47157 32360
rect 47115 32311 47157 32320
rect 47691 32360 47733 32369
rect 47691 32320 47692 32360
rect 47732 32320 47733 32360
rect 47691 32311 47733 32320
rect 47116 32226 47156 32311
rect 47211 32192 47253 32201
rect 47884 32192 47924 32992
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 47211 32152 47212 32192
rect 47252 32152 47253 32192
rect 47211 32143 47253 32152
rect 47788 32152 47924 32192
rect 48075 32192 48117 32201
rect 48075 32152 48076 32192
rect 48116 32152 48117 32192
rect 47115 31940 47157 31949
rect 47115 31900 47116 31940
rect 47156 31900 47157 31940
rect 47115 31891 47157 31900
rect 47116 31806 47156 31891
rect 46923 31436 46965 31445
rect 46923 31396 46924 31436
rect 46964 31396 46965 31436
rect 46923 31387 46965 31396
rect 46827 30764 46869 30773
rect 46827 30724 46828 30764
rect 46868 30724 46869 30764
rect 46827 30715 46869 30724
rect 46540 30631 46580 30640
rect 46828 30680 46868 30715
rect 46828 30629 46868 30640
rect 45291 30512 45333 30521
rect 45291 30472 45292 30512
rect 45332 30472 45333 30512
rect 45291 30463 45333 30472
rect 45292 30378 45332 30463
rect 45483 30428 45525 30437
rect 45483 30388 45484 30428
rect 45524 30388 45525 30428
rect 45483 30379 45525 30388
rect 46443 30428 46485 30437
rect 46443 30388 46444 30428
rect 46484 30388 46485 30428
rect 46443 30379 46485 30388
rect 46732 30428 46772 30437
rect 43372 28194 43412 28279
rect 43467 28160 43509 28169
rect 43467 28120 43468 28160
rect 43508 28120 43509 28160
rect 43564 28160 43604 28288
rect 43659 28328 43701 28337
rect 43659 28288 43660 28328
rect 43700 28288 43701 28328
rect 45004 28960 45236 29000
rect 44044 28293 44084 28302
rect 44524 28328 44564 28337
rect 43659 28279 43701 28288
rect 44524 28169 44564 28288
rect 45004 28328 45044 28960
rect 45099 28412 45141 28421
rect 45099 28372 45100 28412
rect 45140 28372 45141 28412
rect 45099 28363 45141 28372
rect 43852 28160 43892 28169
rect 44523 28160 44565 28169
rect 43564 28120 43796 28160
rect 43467 28111 43509 28120
rect 42988 27607 43028 27616
rect 43084 27952 43316 27992
rect 43371 27992 43413 28001
rect 43371 27952 43372 27992
rect 43412 27952 43413 27992
rect 42220 27488 42260 27497
rect 41740 26767 41780 26776
rect 41931 26816 41973 26825
rect 41931 26776 41932 26816
rect 41972 26776 41973 26816
rect 41931 26767 41973 26776
rect 42124 26816 42164 26825
rect 42220 26816 42260 27448
rect 43084 26825 43124 27952
rect 43371 27943 43413 27952
rect 43276 27656 43316 27665
rect 43180 27637 43220 27646
rect 43180 27581 43220 27597
rect 43179 27572 43221 27581
rect 43179 27532 43180 27572
rect 43220 27532 43221 27572
rect 43179 27523 43221 27532
rect 43180 27502 43220 27523
rect 42164 26776 42260 26816
rect 42411 26816 42453 26825
rect 42411 26776 42412 26816
rect 42452 26776 42453 26816
rect 42124 26767 42164 26776
rect 42411 26767 42453 26776
rect 42988 26816 43028 26825
rect 43083 26816 43125 26825
rect 43028 26776 43084 26816
rect 43124 26776 43125 26816
rect 42988 26767 43028 26776
rect 43083 26767 43125 26776
rect 40683 26480 40725 26489
rect 40683 26440 40684 26480
rect 40724 26440 40725 26480
rect 40683 26431 40725 26440
rect 40875 26480 40917 26489
rect 40875 26440 40876 26480
rect 40916 26440 40917 26480
rect 40875 26431 40917 26440
rect 41547 26480 41589 26489
rect 41547 26440 41548 26480
rect 41588 26440 41589 26480
rect 41547 26431 41589 26440
rect 40396 26095 40436 26104
rect 39340 26009 39380 26095
rect 39820 26010 39860 26095
rect 40300 26010 40340 26095
rect 40587 26060 40629 26069
rect 40587 26020 40588 26060
rect 40628 26020 40629 26060
rect 40587 26011 40629 26020
rect 39627 25808 39669 25817
rect 39627 25768 39628 25808
rect 39668 25768 39669 25808
rect 39627 25759 39669 25768
rect 39628 25556 39668 25759
rect 39628 25507 39668 25516
rect 38955 25472 38997 25481
rect 38955 25432 38956 25472
rect 38996 25432 38997 25472
rect 38955 25423 38997 25432
rect 40299 25472 40341 25481
rect 40299 25432 40300 25472
rect 40340 25432 40341 25472
rect 40299 25423 40341 25432
rect 39052 25304 39092 25313
rect 39340 25304 39380 25313
rect 38943 25293 38983 25302
rect 39092 25264 39340 25304
rect 39052 25255 39092 25264
rect 39340 25255 39380 25264
rect 39915 25304 39957 25313
rect 39915 25264 39916 25304
rect 39956 25264 39957 25304
rect 39915 25255 39957 25264
rect 40300 25304 40340 25423
rect 40300 25255 40340 25264
rect 40491 25304 40533 25313
rect 40491 25264 40492 25304
rect 40532 25264 40533 25304
rect 40491 25255 40533 25264
rect 40588 25304 40628 26011
rect 40684 25313 40724 26431
rect 40779 26312 40821 26321
rect 40779 26272 40780 26312
rect 40820 26272 40821 26312
rect 40779 26263 40821 26272
rect 40780 26144 40820 26263
rect 40780 26095 40820 26104
rect 40876 26144 40916 26431
rect 40779 25892 40821 25901
rect 40779 25852 40780 25892
rect 40820 25852 40821 25892
rect 40779 25843 40821 25852
rect 40588 25255 40628 25264
rect 40683 25304 40725 25313
rect 40683 25264 40684 25304
rect 40724 25264 40725 25304
rect 40683 25255 40725 25264
rect 38859 25220 38901 25229
rect 38943 25220 38983 25253
rect 38859 25180 38860 25220
rect 38900 25180 38983 25220
rect 38859 25171 38901 25180
rect 38860 25086 38900 25171
rect 39820 24800 39860 24809
rect 39916 24800 39956 25255
rect 40011 25220 40053 25229
rect 40011 25180 40012 25220
rect 40052 25180 40053 25220
rect 40011 25171 40053 25180
rect 39860 24760 39956 24800
rect 39820 24751 39860 24760
rect 38475 24716 38517 24725
rect 38475 24676 38476 24716
rect 38516 24676 38517 24716
rect 38475 24667 38517 24676
rect 38284 24578 38324 24587
rect 38476 24582 38516 24667
rect 40012 24627 40052 25171
rect 40492 25170 40532 25255
rect 40780 25136 40820 25843
rect 40876 25229 40916 26104
rect 42219 26144 42261 26153
rect 42219 26104 42220 26144
rect 42260 26104 42261 26144
rect 42219 26095 42261 26104
rect 42316 26144 42356 26153
rect 42220 26010 42260 26095
rect 41259 25556 41301 25565
rect 41259 25516 41260 25556
rect 41300 25516 41301 25556
rect 42316 25556 42356 26104
rect 42412 26144 42452 26767
rect 43084 26682 43124 26767
rect 42891 26648 42933 26657
rect 42891 26608 42892 26648
rect 42932 26608 42933 26648
rect 42891 26599 42933 26608
rect 42412 26095 42452 26104
rect 42508 26144 42548 26153
rect 42795 26144 42837 26153
rect 42548 26104 42796 26144
rect 42836 26104 42837 26144
rect 42508 26095 42548 26104
rect 42795 26095 42837 26104
rect 42892 26144 42932 26599
rect 43276 26489 43316 27616
rect 43275 26480 43317 26489
rect 43275 26440 43276 26480
rect 43316 26440 43317 26480
rect 43275 26431 43317 26440
rect 43372 26321 43412 27943
rect 43468 27824 43508 28111
rect 43468 27784 43700 27824
rect 43468 27656 43508 27665
rect 43660 27656 43700 27784
rect 43508 27616 43604 27656
rect 43468 27607 43508 27616
rect 43467 27404 43509 27413
rect 43467 27364 43468 27404
rect 43508 27364 43509 27404
rect 43467 27355 43509 27364
rect 43468 27270 43508 27355
rect 43371 26312 43413 26321
rect 43276 26272 43372 26312
rect 43412 26272 43413 26312
rect 42892 26095 42932 26104
rect 43083 26144 43125 26153
rect 43083 26104 43084 26144
rect 43124 26104 43125 26144
rect 43083 26095 43125 26104
rect 43180 26144 43220 26153
rect 42796 26010 42836 26095
rect 43084 26010 43124 26095
rect 42507 25976 42549 25985
rect 42507 25936 42508 25976
rect 42548 25936 42549 25976
rect 42507 25927 42549 25936
rect 42412 25556 42452 25565
rect 42316 25516 42412 25556
rect 41259 25507 41301 25516
rect 42412 25507 42452 25516
rect 41260 25422 41300 25507
rect 41931 25388 41973 25397
rect 41931 25348 41932 25388
rect 41972 25348 41973 25388
rect 41931 25339 41973 25348
rect 42315 25388 42357 25397
rect 42315 25348 42316 25388
rect 42356 25348 42357 25388
rect 42315 25339 42357 25348
rect 41355 25304 41397 25313
rect 41355 25264 41356 25304
rect 41396 25264 41397 25304
rect 41355 25255 41397 25264
rect 41644 25304 41684 25313
rect 41739 25304 41781 25313
rect 41684 25264 41740 25304
rect 41780 25264 41781 25304
rect 41644 25255 41684 25264
rect 41739 25255 41781 25264
rect 41932 25304 41972 25339
rect 40875 25220 40917 25229
rect 40875 25180 40876 25220
rect 40916 25180 40917 25220
rect 40875 25171 40917 25180
rect 40780 25087 40820 25096
rect 40012 24578 40052 24587
rect 40492 24632 40532 24641
rect 40492 24473 40532 24592
rect 40971 24548 41013 24557
rect 40971 24508 40972 24548
rect 41012 24508 41013 24548
rect 40971 24499 41013 24508
rect 41068 24548 41108 24557
rect 38860 24464 38900 24473
rect 38283 24296 38325 24305
rect 38283 24256 38284 24296
rect 38324 24256 38325 24296
rect 38283 24247 38325 24256
rect 37900 23792 37940 23803
rect 37900 23717 37940 23752
rect 37996 23792 38036 23801
rect 37899 23708 37941 23717
rect 37899 23668 37900 23708
rect 37940 23668 37941 23708
rect 37899 23659 37941 23668
rect 37996 23549 38036 23752
rect 38092 23792 38132 23801
rect 37995 23540 38037 23549
rect 37995 23500 37996 23540
rect 38036 23500 38037 23540
rect 37995 23491 38037 23500
rect 37419 23372 37461 23381
rect 37419 23332 37420 23372
rect 37460 23332 37461 23372
rect 37419 23323 37461 23332
rect 37803 23372 37845 23381
rect 37803 23332 37804 23372
rect 37844 23332 37845 23372
rect 37803 23323 37845 23332
rect 37803 23120 37845 23129
rect 37803 23080 37804 23120
rect 37844 23080 37845 23120
rect 37803 23071 37845 23080
rect 37323 23036 37365 23045
rect 37323 22996 37324 23036
rect 37364 22996 37365 23036
rect 37323 22987 37365 22996
rect 37804 22986 37844 23071
rect 37995 23036 38037 23045
rect 37995 22996 37996 23036
rect 38036 22996 38037 23036
rect 37995 22987 38037 22996
rect 37996 22902 38036 22987
rect 36844 22483 36884 22492
rect 37132 22868 37172 22877
rect 34868 22240 35060 22280
rect 34828 22231 34868 22240
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 34347 21608 34389 21617
rect 34347 21568 34348 21608
rect 34388 21568 34389 21608
rect 34347 21559 34389 21568
rect 34924 21440 34964 21449
rect 35020 21440 35060 22240
rect 35692 22231 35732 22240
rect 36267 22196 36309 22205
rect 36267 22156 36268 22196
rect 36308 22156 36309 22196
rect 36267 22147 36309 22156
rect 35691 22112 35733 22121
rect 35691 22072 35692 22112
rect 35732 22072 35733 22112
rect 35691 22063 35733 22072
rect 34964 21400 35060 21440
rect 34924 21391 34964 21400
rect 33772 20971 33812 20980
rect 33291 20936 33333 20945
rect 33291 20896 33292 20936
rect 33332 20896 33333 20936
rect 33291 20887 33333 20896
rect 34828 20936 34868 20945
rect 34868 20896 35060 20936
rect 34828 20887 34868 20896
rect 33292 20768 33332 20887
rect 33292 20719 33332 20728
rect 33291 20600 33333 20609
rect 33291 20560 33292 20600
rect 33332 20560 33333 20600
rect 33291 20551 33333 20560
rect 33771 20600 33813 20609
rect 33771 20560 33772 20600
rect 33812 20560 33813 20600
rect 33771 20551 33813 20560
rect 33292 20096 33332 20551
rect 33772 20466 33812 20551
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 34251 20264 34293 20273
rect 34251 20224 34252 20264
rect 34292 20224 34293 20264
rect 34251 20215 34293 20224
rect 33292 20047 33332 20056
rect 33099 20012 33141 20021
rect 33099 19972 33100 20012
rect 33140 19972 33141 20012
rect 33099 19963 33141 19972
rect 33579 20012 33621 20021
rect 33579 19972 33580 20012
rect 33620 19972 33621 20012
rect 33579 19963 33621 19972
rect 31948 19256 31988 19265
rect 31851 19004 31893 19013
rect 31851 18964 31852 19004
rect 31892 18964 31893 19004
rect 31851 18955 31893 18964
rect 31852 18845 31892 18889
rect 31851 18836 31893 18845
rect 31851 18796 31852 18836
rect 31892 18796 31893 18836
rect 31851 18794 31893 18796
rect 31851 18787 31852 18794
rect 31892 18787 31893 18794
rect 31852 18745 31892 18754
rect 31852 18584 31892 18593
rect 31660 18535 31700 18544
rect 31756 18544 31852 18584
rect 31756 18425 31796 18544
rect 31563 18416 31605 18425
rect 31563 18376 31564 18416
rect 31604 18376 31605 18416
rect 31563 18367 31605 18376
rect 31755 18416 31797 18425
rect 31755 18376 31756 18416
rect 31796 18376 31797 18416
rect 31755 18367 31797 18376
rect 31755 17828 31797 17837
rect 31755 17788 31756 17828
rect 31796 17788 31797 17828
rect 31755 17779 31797 17788
rect 31180 17704 31372 17744
rect 31412 17704 31508 17744
rect 31564 17744 31604 17753
rect 31180 17072 31220 17704
rect 31372 17695 31412 17704
rect 31564 17240 31604 17704
rect 31756 17694 31796 17779
rect 31852 17744 31892 18544
rect 31852 17576 31892 17704
rect 31468 17200 31604 17240
rect 31660 17536 31892 17576
rect 31180 17023 31220 17032
rect 31372 17072 31412 17081
rect 31372 15737 31412 17032
rect 31468 16820 31508 17200
rect 31660 17072 31700 17536
rect 31755 17408 31797 17417
rect 31755 17368 31756 17408
rect 31796 17368 31797 17408
rect 31755 17359 31797 17368
rect 31660 17023 31700 17032
rect 31564 16988 31604 16997
rect 31564 16904 31604 16948
rect 31659 16904 31701 16913
rect 31564 16864 31660 16904
rect 31700 16864 31701 16904
rect 31659 16855 31701 16864
rect 31468 16780 31604 16820
rect 31467 16400 31509 16409
rect 31467 16360 31468 16400
rect 31508 16360 31509 16400
rect 31467 16351 31509 16360
rect 31371 15728 31413 15737
rect 31371 15688 31372 15728
rect 31412 15688 31413 15728
rect 31371 15679 31413 15688
rect 31468 15056 31508 16351
rect 31564 15821 31604 16780
rect 31756 16409 31796 17359
rect 31948 17240 31988 19216
rect 32811 19256 32853 19265
rect 32811 19216 32812 19256
rect 32852 19216 32853 19256
rect 32811 19207 32853 19216
rect 33003 19256 33045 19265
rect 33003 19216 33004 19256
rect 33044 19216 33045 19256
rect 33003 19207 33045 19216
rect 32427 19172 32469 19181
rect 32427 19132 32428 19172
rect 32468 19132 32469 19172
rect 32427 19123 32469 19132
rect 32428 19038 32468 19123
rect 32043 18836 32085 18845
rect 32043 18796 32044 18836
rect 32084 18796 32085 18836
rect 32043 18787 32085 18796
rect 32044 18005 32084 18787
rect 32236 18584 32276 18593
rect 32139 18080 32181 18089
rect 32139 18040 32140 18080
rect 32180 18040 32181 18080
rect 32139 18031 32181 18040
rect 32043 17996 32085 18005
rect 32043 17956 32044 17996
rect 32084 17956 32085 17996
rect 32043 17947 32085 17956
rect 32140 17921 32180 18031
rect 32139 17912 32181 17921
rect 32139 17872 32140 17912
rect 32180 17872 32181 17912
rect 32139 17863 32181 17872
rect 32043 17492 32085 17501
rect 32043 17452 32044 17492
rect 32084 17452 32085 17492
rect 32043 17443 32085 17452
rect 31852 17200 31988 17240
rect 31755 16400 31797 16409
rect 31755 16360 31756 16400
rect 31796 16360 31797 16400
rect 31755 16351 31797 16360
rect 31852 16241 31892 17200
rect 31948 17072 31988 17081
rect 31948 16745 31988 17032
rect 32044 17072 32084 17443
rect 32044 17023 32084 17032
rect 32140 17072 32180 17863
rect 32236 17501 32276 18544
rect 32331 17744 32373 17753
rect 32331 17704 32332 17744
rect 32372 17704 32373 17744
rect 32331 17695 32373 17704
rect 32235 17492 32277 17501
rect 32235 17452 32236 17492
rect 32276 17452 32277 17492
rect 32235 17443 32277 17452
rect 32043 16904 32085 16913
rect 32043 16864 32044 16904
rect 32084 16864 32085 16904
rect 32140 16904 32180 17032
rect 32236 17072 32276 17081
rect 32332 17072 32372 17695
rect 32428 17660 32468 17669
rect 32428 17249 32468 17620
rect 32427 17240 32469 17249
rect 32427 17200 32428 17240
rect 32468 17200 32469 17240
rect 32427 17191 32469 17200
rect 32427 17072 32469 17081
rect 32332 17032 32428 17072
rect 32468 17032 32469 17072
rect 32236 16988 32276 17032
rect 32427 17023 32469 17032
rect 32236 16948 32372 16988
rect 32140 16864 32276 16904
rect 32043 16855 32085 16864
rect 31947 16736 31989 16745
rect 31947 16696 31948 16736
rect 31988 16696 31989 16736
rect 31947 16687 31989 16696
rect 31947 16484 31989 16493
rect 31947 16444 31948 16484
rect 31988 16444 31989 16484
rect 31947 16435 31989 16444
rect 31851 16232 31893 16241
rect 31851 16192 31852 16232
rect 31892 16192 31893 16232
rect 31851 16183 31893 16192
rect 31660 16148 31700 16157
rect 31700 16108 31796 16148
rect 31660 16099 31700 16108
rect 31659 15896 31701 15905
rect 31659 15856 31660 15896
rect 31700 15856 31701 15896
rect 31659 15847 31701 15856
rect 31563 15812 31605 15821
rect 31563 15772 31564 15812
rect 31604 15772 31605 15812
rect 31563 15763 31605 15772
rect 31563 15644 31605 15653
rect 31563 15604 31564 15644
rect 31604 15604 31605 15644
rect 31563 15595 31605 15604
rect 31564 15560 31604 15595
rect 31564 15509 31604 15520
rect 31660 15560 31700 15847
rect 31660 15511 31700 15520
rect 31563 15308 31605 15317
rect 31563 15268 31564 15308
rect 31604 15268 31605 15308
rect 31563 15259 31605 15268
rect 31564 15174 31604 15259
rect 31468 15016 31604 15056
rect 31467 14888 31509 14897
rect 31467 14848 31468 14888
rect 31508 14848 31509 14888
rect 31467 14839 31509 14848
rect 31371 14720 31413 14729
rect 31371 14680 31372 14720
rect 31412 14680 31413 14720
rect 31371 14671 31413 14680
rect 31468 14720 31508 14839
rect 31372 14586 31412 14671
rect 31468 13889 31508 14680
rect 31564 14720 31604 15016
rect 31659 14804 31701 14813
rect 31659 14764 31660 14804
rect 31700 14764 31701 14804
rect 31659 14755 31701 14764
rect 31564 14671 31604 14680
rect 31660 14720 31700 14755
rect 31660 14669 31700 14680
rect 31563 14552 31605 14561
rect 31563 14512 31564 14552
rect 31604 14512 31605 14552
rect 31563 14503 31605 14512
rect 31467 13880 31509 13889
rect 31467 13840 31468 13880
rect 31508 13840 31509 13880
rect 31467 13831 31509 13840
rect 31564 13628 31604 14503
rect 31468 13588 31604 13628
rect 31372 13208 31412 13219
rect 31468 13208 31508 13588
rect 31564 13385 31604 13470
rect 31563 13376 31605 13385
rect 31563 13336 31564 13376
rect 31604 13336 31605 13376
rect 31563 13327 31605 13336
rect 31564 13208 31604 13217
rect 31468 13168 31564 13208
rect 31372 13133 31412 13168
rect 31564 13159 31604 13168
rect 31660 13208 31700 13219
rect 31660 13133 31700 13168
rect 31371 13124 31413 13133
rect 31371 13084 31372 13124
rect 31412 13084 31413 13124
rect 31371 13075 31413 13084
rect 31659 13124 31701 13133
rect 31659 13084 31660 13124
rect 31700 13084 31701 13124
rect 31659 13075 31701 13084
rect 31467 12788 31509 12797
rect 31467 12748 31468 12788
rect 31508 12748 31509 12788
rect 31467 12739 31509 12748
rect 31084 11899 31124 11908
rect 31371 11696 31413 11705
rect 31371 11656 31372 11696
rect 31412 11656 31413 11696
rect 31371 11647 31413 11656
rect 31372 11562 31412 11647
rect 31468 11192 31508 12739
rect 31756 12545 31796 16108
rect 31852 15905 31892 16183
rect 31851 15896 31893 15905
rect 31851 15856 31852 15896
rect 31892 15856 31893 15896
rect 31851 15847 31893 15856
rect 31948 15644 31988 16435
rect 31852 15604 31988 15644
rect 31852 15560 31892 15604
rect 32044 15569 32084 16855
rect 32044 15560 32090 15569
rect 31852 15511 31892 15520
rect 31948 15531 31988 15540
rect 32044 15520 32049 15560
rect 32089 15520 32090 15560
rect 32048 15511 32090 15520
rect 31948 15401 31988 15491
rect 32049 15426 32089 15511
rect 31947 15392 31989 15401
rect 31947 15352 31948 15392
rect 31988 15352 31989 15392
rect 31947 15343 31989 15352
rect 31851 15308 31893 15317
rect 31851 15268 31852 15308
rect 31892 15268 31893 15308
rect 31851 15259 31893 15268
rect 31852 14720 31892 15259
rect 32236 15065 32276 16864
rect 32332 16241 32372 16948
rect 32331 16232 32373 16241
rect 32331 16192 32332 16232
rect 32372 16192 32373 16232
rect 32331 16183 32373 16192
rect 32428 16232 32468 17023
rect 32619 16820 32661 16829
rect 32619 16780 32620 16820
rect 32660 16780 32661 16820
rect 32619 16771 32661 16780
rect 32908 16820 32948 16829
rect 32428 16183 32468 16192
rect 32422 15560 32464 15569
rect 32422 15520 32423 15560
rect 32463 15520 32464 15560
rect 32422 15511 32464 15520
rect 32524 15560 32564 15569
rect 32423 15426 32463 15511
rect 32524 15317 32564 15520
rect 32620 15560 32660 16771
rect 32908 16400 32948 16780
rect 32716 16360 32948 16400
rect 33004 16400 33044 19207
rect 33100 18584 33140 19963
rect 33580 19878 33620 19963
rect 33195 19844 33237 19853
rect 33195 19804 33196 19844
rect 33236 19804 33237 19844
rect 33195 19795 33237 19804
rect 33772 19844 33812 19853
rect 33196 19256 33236 19795
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 33772 19256 33812 19804
rect 33963 19592 34005 19601
rect 33963 19552 33964 19592
rect 34004 19552 34005 19592
rect 33963 19543 34005 19552
rect 33964 19265 34004 19543
rect 34252 19424 34292 20215
rect 35020 20180 35060 20896
rect 35404 20768 35444 20777
rect 35308 20600 35348 20609
rect 35308 20180 35348 20560
rect 34732 20140 35060 20180
rect 35212 20140 35348 20180
rect 34348 20096 34388 20105
rect 34348 19508 34388 20056
rect 34732 20096 34772 20140
rect 34732 20047 34772 20056
rect 35115 19592 35157 19601
rect 35115 19552 35116 19592
rect 35156 19552 35157 19592
rect 35115 19543 35157 19552
rect 34924 19508 34964 19517
rect 34348 19468 34924 19508
rect 34924 19459 34964 19468
rect 34060 19384 34388 19424
rect 33196 19097 33236 19216
rect 33676 19216 33812 19256
rect 33868 19256 33908 19265
rect 33195 19088 33237 19097
rect 33195 19048 33196 19088
rect 33236 19048 33237 19088
rect 33195 19039 33237 19048
rect 33676 18761 33716 19216
rect 33772 19088 33812 19097
rect 33675 18752 33717 18761
rect 33675 18712 33676 18752
rect 33716 18712 33717 18752
rect 33675 18703 33717 18712
rect 33100 17669 33140 18544
rect 33580 18584 33620 18593
rect 33580 18341 33620 18544
rect 33676 18584 33716 18593
rect 33772 18584 33812 19048
rect 33868 18929 33908 19216
rect 33963 19256 34005 19265
rect 33963 19216 33964 19256
rect 34004 19216 34005 19256
rect 33963 19207 34005 19216
rect 34060 19256 34100 19384
rect 34252 19256 34292 19265
rect 34060 19207 34100 19216
rect 34156 19216 34252 19256
rect 33964 19122 34004 19207
rect 34059 19088 34101 19097
rect 34059 19048 34060 19088
rect 34100 19048 34101 19088
rect 34059 19039 34101 19048
rect 33963 19004 34005 19013
rect 33963 18964 33964 19004
rect 34004 18964 34005 19004
rect 33963 18955 34005 18964
rect 33867 18920 33909 18929
rect 33867 18880 33868 18920
rect 33908 18880 33909 18920
rect 33867 18871 33909 18880
rect 33868 18593 33908 18678
rect 33716 18544 33812 18584
rect 33867 18584 33909 18593
rect 33867 18544 33868 18584
rect 33908 18544 33909 18584
rect 33676 18535 33716 18544
rect 33867 18535 33909 18544
rect 33868 18416 33908 18425
rect 33964 18416 34004 18955
rect 33908 18376 34004 18416
rect 33868 18367 33908 18376
rect 33579 18332 33621 18341
rect 33579 18292 33580 18332
rect 33620 18292 33621 18332
rect 33579 18283 33621 18292
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 33387 17996 33429 18005
rect 33387 17956 33388 17996
rect 33428 17956 33429 17996
rect 33387 17947 33429 17956
rect 33195 17828 33237 17837
rect 33195 17788 33196 17828
rect 33236 17788 33237 17828
rect 33195 17779 33237 17788
rect 33196 17744 33236 17779
rect 33196 17693 33236 17704
rect 33099 17660 33141 17669
rect 33099 17620 33100 17660
rect 33140 17620 33141 17660
rect 33099 17611 33141 17620
rect 33388 17072 33428 17947
rect 34060 17744 34100 19039
rect 34156 19013 34196 19216
rect 34252 19207 34292 19216
rect 34155 19004 34197 19013
rect 34155 18964 34156 19004
rect 34196 18964 34197 19004
rect 34155 18955 34197 18964
rect 34251 18920 34293 18929
rect 34251 18880 34252 18920
rect 34292 18880 34293 18920
rect 34251 18871 34293 18880
rect 34252 18752 34292 18871
rect 34348 18761 34388 19384
rect 35116 19340 35156 19543
rect 35116 19291 35156 19300
rect 34443 19256 34485 19265
rect 34443 19216 34444 19256
rect 34484 19216 34485 19256
rect 34443 19207 34485 19216
rect 34156 18712 34292 18752
rect 34347 18752 34389 18761
rect 34347 18712 34348 18752
rect 34388 18712 34389 18752
rect 34156 17996 34196 18712
rect 34347 18703 34389 18712
rect 34252 18584 34292 18593
rect 34252 18509 34292 18544
rect 34348 18584 34388 18593
rect 34251 18500 34293 18509
rect 34251 18460 34252 18500
rect 34292 18460 34293 18500
rect 34251 18451 34293 18460
rect 34156 17947 34196 17956
rect 34156 17744 34196 17753
rect 34060 17704 34156 17744
rect 34156 17695 34196 17704
rect 34155 17240 34197 17249
rect 34155 17200 34156 17240
rect 34196 17200 34197 17240
rect 34155 17191 34197 17200
rect 33196 17032 33388 17072
rect 33196 16484 33236 17032
rect 33388 17023 33428 17032
rect 33772 17072 33812 17081
rect 33772 16829 33812 17032
rect 33771 16820 33813 16829
rect 33771 16780 33772 16820
rect 33812 16780 33813 16820
rect 33771 16771 33813 16780
rect 34060 16820 34100 16829
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 34060 16493 34100 16780
rect 34059 16484 34101 16493
rect 33196 16444 33332 16484
rect 33004 16360 33236 16400
rect 32716 15905 32756 16360
rect 32812 16232 32852 16241
rect 32715 15896 32757 15905
rect 32715 15856 32716 15896
rect 32756 15856 32757 15896
rect 32715 15847 32757 15856
rect 32716 15728 32756 15737
rect 32812 15728 32852 16192
rect 32908 16232 32948 16241
rect 32908 16073 32948 16192
rect 33099 16232 33141 16241
rect 33099 16192 33100 16232
rect 33140 16192 33141 16232
rect 33099 16183 33141 16192
rect 33003 16148 33045 16157
rect 33003 16108 33004 16148
rect 33044 16108 33045 16148
rect 33003 16099 33045 16108
rect 32907 16064 32949 16073
rect 32907 16024 32908 16064
rect 32948 16024 32949 16064
rect 32907 16015 32949 16024
rect 33004 16014 33044 16099
rect 33100 16098 33140 16183
rect 33003 15896 33045 15905
rect 33003 15856 33004 15896
rect 33044 15856 33045 15896
rect 33003 15847 33045 15856
rect 32756 15688 32852 15728
rect 32716 15679 32756 15688
rect 32907 15644 32949 15653
rect 32907 15604 32908 15644
rect 32948 15604 32949 15644
rect 32907 15595 32949 15604
rect 32620 15511 32660 15520
rect 32812 15560 32852 15569
rect 32523 15308 32565 15317
rect 32523 15268 32524 15308
rect 32564 15268 32565 15308
rect 32523 15259 32565 15268
rect 32427 15224 32469 15233
rect 32427 15184 32428 15224
rect 32468 15184 32469 15224
rect 32427 15175 32469 15184
rect 32235 15056 32277 15065
rect 32235 15016 32236 15056
rect 32276 15016 32277 15056
rect 32235 15007 32277 15016
rect 32332 14888 32372 14897
rect 32044 14848 32332 14888
rect 32044 14720 32084 14848
rect 32332 14839 32372 14848
rect 31852 14671 31892 14680
rect 31948 14706 32084 14720
rect 31988 14680 32084 14706
rect 32139 14720 32181 14729
rect 32139 14680 32140 14720
rect 32180 14680 32181 14720
rect 32139 14671 32181 14680
rect 32332 14720 32372 14729
rect 32428 14720 32468 15175
rect 32812 14813 32852 15520
rect 32908 15560 32948 15595
rect 32908 15509 32948 15520
rect 33004 15233 33044 15847
rect 33003 15224 33045 15233
rect 33003 15184 33004 15224
rect 33044 15184 33045 15224
rect 33003 15175 33045 15184
rect 33099 15140 33141 15149
rect 33099 15100 33100 15140
rect 33140 15100 33141 15140
rect 33099 15091 33141 15100
rect 32811 14804 32853 14813
rect 33003 14804 33045 14813
rect 32811 14764 32812 14804
rect 32852 14764 32948 14804
rect 32811 14755 32853 14764
rect 32372 14680 32468 14720
rect 32523 14720 32565 14729
rect 32523 14680 32524 14720
rect 32564 14680 32565 14720
rect 32332 14671 32372 14680
rect 32523 14671 32565 14680
rect 32620 14720 32660 14729
rect 31948 14657 31988 14666
rect 32140 14586 32180 14671
rect 32524 14586 32564 14671
rect 32044 14552 32084 14561
rect 32044 14393 32084 14512
rect 32620 14477 32660 14680
rect 32812 14552 32852 14563
rect 32812 14477 32852 14512
rect 32619 14468 32661 14477
rect 32619 14428 32620 14468
rect 32660 14428 32661 14468
rect 32619 14419 32661 14428
rect 32811 14468 32853 14477
rect 32811 14428 32812 14468
rect 32852 14428 32853 14468
rect 32811 14419 32853 14428
rect 32043 14384 32085 14393
rect 32043 14344 32044 14384
rect 32084 14344 32085 14384
rect 32043 14335 32085 14344
rect 32908 14225 32948 14764
rect 33003 14764 33004 14804
rect 33044 14764 33045 14804
rect 33003 14755 33045 14764
rect 33004 14720 33044 14755
rect 33004 14669 33044 14680
rect 33100 14720 33140 15091
rect 33100 14671 33140 14680
rect 32907 14216 32949 14225
rect 32907 14176 32908 14216
rect 32948 14176 32949 14216
rect 32907 14167 32949 14176
rect 32331 14132 32373 14141
rect 32331 14092 32332 14132
rect 32372 14092 32373 14132
rect 32331 14083 32373 14092
rect 31947 14048 31989 14057
rect 31947 14008 31948 14048
rect 31988 14008 31989 14048
rect 31947 13999 31989 14008
rect 31755 12536 31797 12545
rect 31755 12496 31756 12536
rect 31796 12496 31797 12536
rect 31948 12536 31988 13999
rect 32139 13880 32181 13889
rect 32139 13840 32140 13880
rect 32180 13840 32181 13880
rect 32139 13831 32181 13840
rect 32140 13746 32180 13831
rect 32235 13376 32277 13385
rect 32235 13336 32236 13376
rect 32276 13336 32277 13376
rect 32235 13327 32277 13336
rect 32236 13208 32276 13327
rect 32236 13159 32276 13168
rect 32332 13124 32372 14083
rect 32811 13376 32853 13385
rect 32811 13336 32812 13376
rect 32852 13336 32853 13376
rect 32811 13327 32853 13336
rect 32332 13075 32372 13084
rect 32428 13208 32468 13217
rect 32044 12536 32084 12545
rect 31948 12496 32044 12536
rect 31755 12487 31797 12496
rect 32044 12487 32084 12496
rect 31756 11705 31796 12487
rect 31851 12284 31893 12293
rect 31851 12244 31852 12284
rect 31892 12244 31893 12284
rect 31851 12235 31893 12244
rect 32331 12284 32373 12293
rect 32331 12244 32332 12284
rect 32372 12244 32373 12284
rect 32331 12235 32373 12244
rect 31755 11696 31797 11705
rect 31755 11656 31756 11696
rect 31796 11656 31797 11696
rect 31755 11647 31797 11656
rect 31852 11453 31892 12235
rect 32235 12200 32277 12209
rect 32235 12160 32236 12200
rect 32276 12160 32277 12200
rect 32235 12151 32277 12160
rect 32236 11696 32276 12151
rect 32332 12150 32372 12235
rect 32332 11696 32372 11705
rect 32236 11656 32332 11696
rect 32332 11647 32372 11656
rect 32236 11528 32276 11537
rect 31851 11444 31893 11453
rect 31851 11404 31852 11444
rect 31892 11404 31893 11444
rect 31851 11395 31893 11404
rect 31664 11276 31706 11285
rect 31664 11236 31665 11276
rect 31705 11236 31706 11276
rect 31664 11227 31706 11236
rect 31468 11143 31508 11152
rect 31563 11108 31605 11117
rect 31563 11068 31564 11108
rect 31604 11068 31605 11108
rect 31563 11059 31605 11068
rect 31180 11024 31220 11033
rect 30988 10436 31028 10445
rect 31180 10436 31220 10984
rect 31028 10396 31220 10436
rect 31276 11024 31316 11033
rect 31276 10436 31316 10984
rect 31467 11024 31509 11033
rect 31467 10984 31468 11024
rect 31508 10984 31509 11024
rect 31467 10975 31509 10984
rect 31564 11024 31604 11059
rect 31665 11024 31705 11227
rect 31468 10890 31508 10975
rect 31564 10973 31604 10984
rect 31660 10984 31665 11024
rect 31660 10975 31705 10984
rect 30988 10387 31028 10396
rect 31276 10387 31316 10396
rect 31371 10268 31413 10277
rect 31371 10228 31372 10268
rect 31412 10228 31413 10268
rect 31371 10219 31413 10228
rect 30995 10199 31035 10206
rect 30995 10197 31124 10199
rect 31035 10184 31124 10197
rect 31180 10184 31220 10193
rect 31035 10159 31180 10184
rect 30995 10148 31035 10157
rect 31084 10144 31180 10159
rect 31180 9941 31220 10144
rect 31372 10184 31412 10219
rect 31372 10133 31412 10144
rect 31179 9932 31221 9941
rect 31179 9892 31180 9932
rect 31220 9892 31221 9932
rect 31179 9883 31221 9892
rect 31660 9848 31700 10975
rect 31564 9808 31700 9848
rect 31467 9008 31509 9017
rect 31467 8968 31468 9008
rect 31508 8968 31509 9008
rect 31467 8959 31509 8968
rect 31468 8924 31508 8959
rect 31468 8873 31508 8884
rect 31564 8849 31604 9808
rect 31852 9764 31892 11395
rect 32236 11117 32276 11488
rect 32428 11360 32468 13168
rect 32524 13208 32564 13217
rect 32524 12713 32564 13168
rect 32812 13208 32852 13327
rect 33099 13292 33141 13301
rect 33099 13252 33100 13292
rect 33140 13252 33141 13292
rect 33099 13243 33141 13252
rect 32523 12704 32565 12713
rect 32523 12664 32524 12704
rect 32564 12664 32565 12704
rect 32523 12655 32565 12664
rect 32812 12629 32852 13168
rect 33003 13208 33045 13217
rect 33003 13168 33004 13208
rect 33044 13168 33045 13208
rect 33003 13159 33045 13168
rect 33100 13208 33140 13243
rect 33004 13074 33044 13159
rect 33100 13157 33140 13168
rect 32907 12788 32949 12797
rect 32907 12748 32908 12788
rect 32948 12748 32949 12788
rect 32907 12739 32949 12748
rect 32811 12620 32853 12629
rect 32811 12580 32812 12620
rect 32852 12580 32853 12620
rect 32811 12571 32853 12580
rect 32716 11873 32756 11958
rect 32715 11864 32757 11873
rect 32715 11824 32716 11864
rect 32756 11824 32757 11864
rect 32715 11815 32757 11824
rect 32332 11320 32468 11360
rect 32524 11696 32564 11705
rect 32235 11108 32277 11117
rect 32235 11068 32236 11108
rect 32276 11068 32277 11108
rect 32235 11059 32277 11068
rect 32043 11024 32085 11033
rect 32043 10984 32044 11024
rect 32084 10984 32085 11024
rect 32043 10975 32085 10984
rect 31660 9724 31892 9764
rect 31660 9260 31700 9724
rect 32044 9680 32084 10975
rect 32332 10688 32372 11320
rect 32524 11117 32564 11656
rect 32716 11696 32756 11707
rect 32716 11621 32756 11656
rect 32908 11696 32948 12739
rect 33099 12704 33141 12713
rect 33099 12664 33100 12704
rect 33140 12664 33141 12704
rect 33099 12655 33141 12664
rect 32908 11647 32948 11656
rect 32715 11612 32757 11621
rect 32715 11572 32716 11612
rect 32756 11572 32757 11612
rect 32715 11563 32757 11572
rect 33100 11528 33140 12655
rect 33196 12629 33236 16360
rect 33292 16232 33332 16444
rect 34059 16444 34060 16484
rect 34100 16444 34101 16484
rect 34059 16435 34101 16444
rect 33484 16232 33524 16241
rect 33292 16183 33332 16192
rect 33388 16192 33484 16232
rect 33291 16064 33333 16073
rect 33291 16024 33292 16064
rect 33332 16024 33333 16064
rect 33291 16015 33333 16024
rect 33292 15930 33332 16015
rect 33388 15392 33428 16192
rect 33484 16183 33524 16192
rect 33580 16232 33620 16241
rect 33580 16064 33620 16192
rect 33772 16232 33812 16241
rect 33964 16232 34004 16241
rect 33812 16192 33908 16232
rect 33772 16183 33812 16192
rect 33772 16064 33812 16073
rect 33580 16024 33772 16064
rect 33772 16015 33812 16024
rect 33868 15896 33908 16192
rect 33772 15856 33908 15896
rect 33675 15644 33717 15653
rect 33675 15604 33676 15644
rect 33716 15604 33717 15644
rect 33675 15595 33717 15604
rect 33676 15560 33716 15595
rect 33772 15569 33812 15856
rect 33964 15812 34004 16192
rect 33868 15772 34004 15812
rect 34060 16232 34100 16241
rect 33868 15732 33908 15772
rect 33676 15509 33716 15520
rect 33771 15560 33813 15569
rect 33771 15520 33772 15560
rect 33812 15520 33813 15560
rect 33771 15511 33813 15520
rect 33772 15426 33812 15511
rect 33388 15343 33428 15352
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 33868 14729 33908 15692
rect 34060 15653 34100 16192
rect 34059 15644 34101 15653
rect 34059 15604 34060 15644
rect 34100 15604 34101 15644
rect 34059 15595 34101 15604
rect 34156 14888 34196 17191
rect 34252 15989 34292 18451
rect 34348 18257 34388 18544
rect 34347 18248 34389 18257
rect 34347 18208 34348 18248
rect 34388 18208 34389 18248
rect 34347 18199 34389 18208
rect 34347 17912 34389 17921
rect 34347 17872 34348 17912
rect 34388 17872 34389 17912
rect 34347 17863 34389 17872
rect 34348 17744 34388 17863
rect 34348 17695 34388 17704
rect 34444 17744 34484 19207
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 34539 18752 34581 18761
rect 34539 18712 34540 18752
rect 34580 18712 34581 18752
rect 34539 18703 34581 18712
rect 34540 17921 34580 18703
rect 35020 18584 35060 18593
rect 34636 18544 35020 18584
rect 34636 18500 34676 18544
rect 35020 18535 35060 18544
rect 35116 18584 35156 18593
rect 35212 18584 35252 20140
rect 35404 19424 35444 20728
rect 35500 20768 35540 20777
rect 35500 19601 35540 20728
rect 35596 20768 35636 20777
rect 35596 20273 35636 20728
rect 35595 20264 35637 20273
rect 35595 20224 35596 20264
rect 35636 20224 35637 20264
rect 35595 20215 35637 20224
rect 35596 20096 35636 20105
rect 35692 20096 35732 22063
rect 36268 21776 36308 22147
rect 36268 21727 36308 21736
rect 36939 21776 36981 21785
rect 36939 21736 36940 21776
rect 36980 21736 36981 21776
rect 36939 21727 36981 21736
rect 36940 21642 36980 21727
rect 35787 21608 35829 21617
rect 35787 21568 35788 21608
rect 35828 21568 35829 21608
rect 35787 21559 35829 21568
rect 35788 21474 35828 21559
rect 37132 20768 37172 22828
rect 38092 22709 38132 23752
rect 38187 23792 38229 23801
rect 38187 23752 38188 23792
rect 38228 23752 38229 23792
rect 38187 23743 38229 23752
rect 38188 23658 38228 23743
rect 38091 22700 38133 22709
rect 38091 22660 38092 22700
rect 38132 22660 38133 22700
rect 38091 22651 38133 22660
rect 37324 22448 37364 22457
rect 37324 21617 37364 22408
rect 37515 22280 37557 22289
rect 38284 22280 38324 24247
rect 38860 23960 38900 24424
rect 40491 24464 40533 24473
rect 40491 24424 40492 24464
rect 40532 24424 40533 24464
rect 40491 24415 40533 24424
rect 40972 24414 41012 24499
rect 41068 24305 41108 24508
rect 41356 24464 41396 25255
rect 41932 25253 41972 25264
rect 42316 25304 42356 25339
rect 42316 25253 42356 25264
rect 42508 25304 42548 25927
rect 42508 25255 42548 25264
rect 41547 25220 41589 25229
rect 41547 25180 41548 25220
rect 41588 25180 41589 25220
rect 41547 25171 41589 25180
rect 41548 25086 41588 25171
rect 43180 25145 43220 26104
rect 42700 25136 42740 25145
rect 41932 25096 42700 25136
rect 41451 24968 41493 24977
rect 41451 24928 41452 24968
rect 41492 24928 41493 24968
rect 41451 24919 41493 24928
rect 41452 24632 41492 24919
rect 41452 24583 41492 24592
rect 41548 24632 41588 24641
rect 41548 24464 41588 24592
rect 41356 24424 41588 24464
rect 41067 24296 41109 24305
rect 41067 24256 41068 24296
rect 41108 24256 41109 24296
rect 41067 24247 41109 24256
rect 38764 23920 38900 23960
rect 38764 23792 38804 23920
rect 38764 23743 38804 23752
rect 39628 23792 39668 23801
rect 38380 23708 38420 23717
rect 38380 23288 38420 23668
rect 38955 23624 38997 23633
rect 38955 23584 38956 23624
rect 38996 23584 38997 23624
rect 38955 23575 38997 23584
rect 38859 23372 38901 23381
rect 38859 23332 38860 23372
rect 38900 23332 38901 23372
rect 38859 23323 38901 23332
rect 38380 23239 38420 23248
rect 38571 22700 38613 22709
rect 38571 22660 38572 22700
rect 38612 22660 38613 22700
rect 38571 22651 38613 22660
rect 37515 22240 37516 22280
rect 37556 22240 37557 22280
rect 37515 22231 37557 22240
rect 37804 22240 38324 22280
rect 38572 22280 38612 22651
rect 38763 22532 38805 22541
rect 38763 22492 38764 22532
rect 38804 22492 38805 22532
rect 38763 22483 38805 22492
rect 37516 21785 37556 22231
rect 37515 21776 37557 21785
rect 37515 21736 37516 21776
rect 37556 21736 37557 21776
rect 37515 21727 37557 21736
rect 37323 21608 37365 21617
rect 37323 21568 37324 21608
rect 37364 21568 37365 21608
rect 37323 21559 37365 21568
rect 37227 21020 37269 21029
rect 37227 20980 37228 21020
rect 37268 20980 37269 21020
rect 37227 20971 37269 20980
rect 37804 21020 37844 22240
rect 38572 22231 38612 22240
rect 38667 22280 38709 22289
rect 38667 22240 38668 22280
rect 38708 22240 38709 22280
rect 38667 22231 38709 22240
rect 38764 22280 38804 22483
rect 38764 22231 38804 22240
rect 38668 22146 38708 22231
rect 38188 22112 38228 22121
rect 37804 20971 37844 20980
rect 37900 22072 38188 22112
rect 37228 20886 37268 20971
rect 37132 20719 37172 20728
rect 37900 20768 37940 22072
rect 38188 22063 38228 22072
rect 38476 22112 38516 22121
rect 38476 21692 38516 22072
rect 38476 21652 38708 21692
rect 38092 21608 38132 21617
rect 38132 21568 38612 21608
rect 38092 21559 38132 21568
rect 37900 20719 37940 20728
rect 35636 20056 35732 20096
rect 36844 20096 36884 20105
rect 35596 20047 35636 20056
rect 35499 19592 35541 19601
rect 35499 19552 35500 19592
rect 35540 19552 35541 19592
rect 35499 19543 35541 19552
rect 36364 19424 36404 19433
rect 35404 19384 35540 19424
rect 35308 19256 35348 19265
rect 35308 19097 35348 19216
rect 35403 19256 35445 19265
rect 35403 19216 35404 19256
rect 35444 19216 35445 19256
rect 35403 19207 35445 19216
rect 35404 19122 35444 19207
rect 35307 19088 35349 19097
rect 35307 19048 35308 19088
rect 35348 19048 35349 19088
rect 35307 19039 35349 19048
rect 35500 18920 35540 19384
rect 36404 19384 36500 19424
rect 36364 19375 36404 19384
rect 36363 19256 36405 19265
rect 36363 19216 36364 19256
rect 36404 19216 36405 19256
rect 36363 19207 36405 19216
rect 35156 18544 35252 18584
rect 35308 18880 35540 18920
rect 35116 18535 35156 18544
rect 34636 18451 34676 18460
rect 34635 18332 34677 18341
rect 34635 18292 34636 18332
rect 34676 18292 34677 18332
rect 34635 18283 34677 18292
rect 34923 18332 34965 18341
rect 34923 18292 34924 18332
rect 34964 18292 34965 18332
rect 34923 18283 34965 18292
rect 34636 17996 34676 18283
rect 34636 17947 34676 17956
rect 34539 17912 34581 17921
rect 34539 17872 34540 17912
rect 34580 17872 34581 17912
rect 34539 17863 34581 17872
rect 34444 17695 34484 17704
rect 34636 17744 34676 17755
rect 34636 17669 34676 17704
rect 34731 17744 34773 17753
rect 34731 17704 34732 17744
rect 34772 17704 34773 17744
rect 34731 17695 34773 17704
rect 34924 17744 34964 18283
rect 35019 18248 35061 18257
rect 35019 18208 35020 18248
rect 35060 18208 35061 18248
rect 35019 18199 35061 18208
rect 34635 17660 34677 17669
rect 34635 17620 34636 17660
rect 34676 17620 34677 17660
rect 34635 17611 34677 17620
rect 34732 17610 34772 17695
rect 34924 17585 34964 17704
rect 35020 17996 35060 18199
rect 35020 17956 35252 17996
rect 35020 17744 35060 17956
rect 35120 17828 35162 17837
rect 35120 17788 35121 17828
rect 35161 17788 35162 17828
rect 35120 17779 35162 17788
rect 35020 17695 35060 17704
rect 35121 17744 35161 17779
rect 34443 17576 34485 17585
rect 34443 17536 34444 17576
rect 34484 17536 34485 17576
rect 34443 17527 34485 17536
rect 34923 17576 34965 17585
rect 34923 17536 34924 17576
rect 34964 17536 34965 17576
rect 34923 17527 34965 17536
rect 34444 16904 34484 17527
rect 35121 17501 35161 17704
rect 35120 17492 35162 17501
rect 35120 17452 35121 17492
rect 35161 17452 35162 17492
rect 35120 17443 35162 17452
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 35115 17240 35157 17249
rect 35115 17200 35116 17240
rect 35156 17200 35157 17240
rect 35115 17191 35157 17200
rect 35019 17156 35061 17165
rect 35019 17116 35020 17156
rect 35060 17116 35061 17156
rect 35019 17107 35061 17116
rect 34444 16855 34484 16864
rect 34924 17072 34964 17081
rect 34347 16568 34389 16577
rect 34347 16528 34348 16568
rect 34388 16528 34389 16568
rect 34347 16519 34389 16528
rect 34251 15980 34293 15989
rect 34251 15940 34252 15980
rect 34292 15940 34293 15980
rect 34251 15931 34293 15940
rect 34348 15737 34388 16519
rect 34636 16232 34676 16241
rect 34636 16073 34676 16192
rect 34924 16073 34964 17032
rect 35020 17022 35060 17107
rect 35116 17072 35156 17191
rect 35116 17023 35156 17032
rect 34635 16064 34677 16073
rect 34635 16024 34636 16064
rect 34676 16024 34677 16064
rect 34635 16015 34677 16024
rect 34923 16064 34965 16073
rect 34923 16024 34924 16064
rect 34964 16024 34965 16064
rect 34923 16015 34965 16024
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 34443 15812 34485 15821
rect 34443 15772 34444 15812
rect 34484 15772 34485 15812
rect 34443 15763 34485 15772
rect 35019 15812 35061 15821
rect 35019 15772 35020 15812
rect 35060 15772 35061 15812
rect 35019 15763 35061 15772
rect 34347 15728 34389 15737
rect 34347 15688 34348 15728
rect 34388 15688 34389 15728
rect 34347 15679 34389 15688
rect 34348 15560 34388 15679
rect 34060 14848 34196 14888
rect 34252 15520 34348 15560
rect 33292 14720 33332 14729
rect 33292 14393 33332 14680
rect 33867 14720 33909 14729
rect 33867 14680 33868 14720
rect 33908 14680 33909 14720
rect 33867 14671 33909 14680
rect 33964 14552 34004 14561
rect 33772 14512 33964 14552
rect 33291 14384 33333 14393
rect 33291 14344 33292 14384
rect 33332 14344 33333 14384
rect 33291 14335 33333 14344
rect 33675 14216 33717 14225
rect 33675 14176 33676 14216
rect 33716 14176 33717 14216
rect 33675 14167 33717 14176
rect 33676 14082 33716 14167
rect 33484 13889 33524 13974
rect 33483 13880 33525 13889
rect 33483 13840 33484 13880
rect 33524 13840 33525 13880
rect 33483 13831 33525 13840
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 33291 13208 33333 13217
rect 33291 13168 33292 13208
rect 33332 13168 33333 13208
rect 33291 13159 33333 13168
rect 33484 13208 33524 13217
rect 33292 13074 33332 13159
rect 33387 13124 33429 13133
rect 33387 13084 33388 13124
rect 33428 13084 33429 13124
rect 33387 13075 33429 13084
rect 33388 12990 33428 13075
rect 33484 12713 33524 13168
rect 33580 13208 33620 13217
rect 33772 13208 33812 14512
rect 33964 14503 34004 14512
rect 33620 13168 33716 13208
rect 33580 13159 33620 13168
rect 33483 12704 33525 12713
rect 33483 12664 33484 12704
rect 33524 12664 33525 12704
rect 33483 12655 33525 12664
rect 33195 12620 33237 12629
rect 33195 12580 33196 12620
rect 33236 12580 33237 12620
rect 33195 12571 33237 12580
rect 33579 12620 33621 12629
rect 33579 12580 33580 12620
rect 33620 12580 33621 12620
rect 33579 12571 33621 12580
rect 33291 12536 33333 12545
rect 33291 12496 33292 12536
rect 33332 12496 33333 12536
rect 33291 12487 33333 12496
rect 33292 12402 33332 12487
rect 33580 12368 33620 12571
rect 33676 12452 33716 13168
rect 33772 13159 33812 13168
rect 34060 12797 34100 14848
rect 34155 14720 34197 14729
rect 34155 14680 34156 14720
rect 34196 14680 34197 14720
rect 34155 14671 34197 14680
rect 34156 14552 34196 14671
rect 34156 14503 34196 14512
rect 34155 13880 34197 13889
rect 34155 13840 34156 13880
rect 34196 13840 34197 13880
rect 34155 13831 34197 13840
rect 34156 13208 34196 13831
rect 34156 13159 34196 13168
rect 34252 13040 34292 15520
rect 34348 15511 34388 15520
rect 34444 15560 34484 15763
rect 34827 15728 34869 15737
rect 34827 15688 34828 15728
rect 34868 15688 34869 15728
rect 34827 15679 34869 15688
rect 34444 15511 34484 15520
rect 34828 15560 34868 15679
rect 34635 15476 34677 15485
rect 34635 15436 34636 15476
rect 34676 15436 34677 15476
rect 34635 15427 34677 15436
rect 34636 15342 34676 15427
rect 34540 15308 34580 15317
rect 34444 15268 34540 15308
rect 34347 15224 34389 15233
rect 34347 15184 34348 15224
rect 34388 15184 34389 15224
rect 34347 15175 34389 15184
rect 34348 14720 34388 15175
rect 34444 14813 34484 15268
rect 34540 15259 34580 15268
rect 34443 14804 34485 14813
rect 34443 14764 34444 14804
rect 34484 14764 34485 14804
rect 34443 14755 34485 14764
rect 34348 14671 34388 14680
rect 34444 14720 34484 14755
rect 34444 14671 34484 14680
rect 34828 14636 34868 15520
rect 34923 15560 34965 15569
rect 34923 15520 34924 15560
rect 34964 15520 34965 15560
rect 34923 15511 34965 15520
rect 35020 15560 35060 15763
rect 35020 15511 35060 15520
rect 34924 15426 34964 15511
rect 34828 14596 35156 14636
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 34635 14216 34677 14225
rect 34635 14176 34636 14216
rect 34676 14176 34677 14216
rect 34635 14167 34677 14176
rect 35116 14216 35156 14596
rect 35116 14167 35156 14176
rect 34347 14048 34389 14057
rect 34347 14008 34348 14048
rect 34388 14008 34389 14048
rect 34347 13999 34389 14008
rect 34636 14048 34676 14167
rect 34636 13999 34676 14008
rect 34348 13914 34388 13999
rect 35212 13301 35252 17956
rect 35308 17165 35348 18880
rect 35404 18752 35444 18761
rect 36364 18752 36404 19207
rect 35444 18712 35924 18752
rect 35404 18703 35444 18712
rect 35403 18584 35445 18593
rect 35403 18544 35404 18584
rect 35444 18544 35445 18584
rect 35403 18535 35445 18544
rect 35595 18584 35637 18593
rect 35595 18544 35596 18584
rect 35636 18544 35637 18584
rect 35595 18535 35637 18544
rect 35687 18584 35727 18593
rect 35404 17744 35444 18535
rect 35499 18080 35541 18089
rect 35499 18040 35500 18080
rect 35540 18040 35541 18080
rect 35499 18031 35541 18040
rect 35404 17695 35444 17704
rect 35500 17744 35540 18031
rect 35500 17695 35540 17704
rect 35596 17744 35636 18535
rect 35687 18341 35727 18544
rect 35788 18584 35828 18593
rect 35788 18416 35828 18544
rect 35884 18584 35924 18712
rect 35884 18535 35924 18544
rect 35980 18712 36364 18752
rect 35980 18416 36020 18712
rect 36364 18703 36404 18712
rect 36075 18584 36117 18593
rect 36075 18544 36076 18584
rect 36116 18544 36117 18584
rect 36075 18535 36117 18544
rect 36172 18584 36212 18593
rect 36212 18544 36308 18584
rect 36172 18535 36212 18544
rect 35788 18376 36020 18416
rect 35686 18332 35728 18341
rect 35686 18292 35687 18332
rect 35727 18292 35728 18332
rect 35686 18283 35728 18292
rect 35596 17695 35636 17704
rect 35692 17744 35732 17753
rect 35788 17744 35828 18376
rect 36076 18005 36116 18535
rect 36172 18332 36212 18341
rect 36075 17996 36117 18005
rect 36075 17956 36076 17996
rect 36116 17956 36117 17996
rect 36075 17947 36117 17956
rect 35883 17912 35925 17921
rect 35883 17872 35884 17912
rect 35924 17872 35925 17912
rect 35883 17863 35925 17872
rect 35732 17704 35828 17744
rect 35692 17695 35732 17704
rect 35884 17660 35924 17863
rect 36172 17753 36212 18292
rect 36171 17744 36213 17753
rect 36171 17704 36172 17744
rect 36212 17704 36213 17744
rect 36171 17695 36213 17704
rect 36268 17669 36308 18544
rect 35788 17620 35924 17660
rect 36267 17660 36309 17669
rect 36267 17620 36268 17660
rect 36308 17620 36309 17660
rect 35691 17324 35733 17333
rect 35691 17284 35692 17324
rect 35732 17284 35733 17324
rect 35691 17275 35733 17284
rect 35307 17156 35349 17165
rect 35307 17116 35308 17156
rect 35348 17116 35349 17156
rect 35307 17107 35349 17116
rect 35596 16232 35636 16241
rect 35596 15821 35636 16192
rect 35595 15812 35637 15821
rect 35595 15772 35596 15812
rect 35636 15772 35637 15812
rect 35595 15763 35637 15772
rect 35692 15728 35732 17275
rect 35788 17156 35828 17620
rect 36267 17611 36309 17620
rect 35883 17324 35925 17333
rect 35883 17284 35884 17324
rect 35924 17284 35925 17324
rect 35883 17275 35925 17284
rect 36307 17324 36349 17333
rect 36307 17284 36308 17324
rect 36348 17284 36349 17324
rect 36307 17275 36349 17284
rect 35788 17116 35830 17156
rect 35790 16988 35830 17116
rect 35884 17072 35924 17275
rect 36308 17165 36348 17275
rect 36460 17249 36500 19384
rect 36844 18584 36884 20056
rect 37900 19928 37940 19937
rect 37708 19888 37900 19928
rect 36939 19256 36981 19265
rect 37324 19256 37364 19265
rect 36939 19216 36940 19256
rect 36980 19216 36981 19256
rect 36939 19207 36981 19216
rect 37132 19216 37324 19256
rect 36940 19122 36980 19207
rect 37036 18584 37076 18593
rect 36844 18544 37036 18584
rect 37036 18535 37076 18544
rect 37132 18416 37172 19216
rect 37324 19207 37364 19216
rect 37708 19256 37748 19888
rect 37900 19879 37940 19888
rect 37708 19207 37748 19216
rect 38572 19256 38612 21568
rect 38668 19937 38708 21652
rect 38860 21020 38900 23323
rect 38956 23120 38996 23575
rect 39052 23120 39092 23129
rect 38956 23080 39052 23120
rect 39052 23071 39092 23080
rect 39340 23120 39380 23131
rect 39340 23045 39380 23080
rect 39339 23036 39381 23045
rect 39339 22996 39340 23036
rect 39380 22996 39381 23036
rect 39339 22987 39381 22996
rect 39628 22952 39668 23752
rect 41740 23792 41780 23801
rect 40780 23624 40820 23633
rect 40587 23540 40629 23549
rect 40587 23500 40588 23540
rect 40628 23500 40629 23540
rect 40587 23491 40629 23500
rect 39628 22903 39668 22912
rect 40300 23120 40340 23129
rect 40011 22868 40053 22877
rect 40011 22828 40012 22868
rect 40052 22828 40053 22868
rect 40011 22819 40053 22828
rect 40012 22734 40052 22819
rect 39819 22700 39861 22709
rect 39819 22660 39820 22700
rect 39860 22660 39861 22700
rect 39819 22651 39861 22660
rect 39051 22532 39093 22541
rect 39051 22492 39052 22532
rect 39092 22492 39093 22532
rect 39051 22483 39093 22492
rect 38955 22280 38997 22289
rect 38955 22240 38956 22280
rect 38996 22240 38997 22280
rect 38955 22231 38997 22240
rect 39052 22280 39092 22483
rect 39052 22231 39092 22240
rect 39244 22280 39284 22289
rect 39284 22240 39764 22280
rect 39244 22231 39284 22240
rect 38956 22146 38996 22231
rect 39148 22112 39188 22121
rect 39148 21617 39188 22072
rect 39436 22112 39476 22121
rect 39340 21692 39380 21701
rect 39436 21692 39476 22072
rect 39380 21652 39476 21692
rect 39340 21643 39380 21652
rect 38955 21608 38997 21617
rect 38955 21568 38956 21608
rect 38996 21568 38997 21608
rect 38955 21559 38997 21568
rect 39147 21608 39189 21617
rect 39147 21568 39148 21608
rect 39188 21568 39189 21608
rect 39147 21559 39189 21568
rect 38956 21474 38996 21559
rect 39628 21356 39668 21365
rect 39244 21316 39628 21356
rect 38956 21020 38996 21029
rect 38860 20980 38956 21020
rect 38956 20971 38996 20980
rect 39051 20768 39093 20777
rect 39051 20728 39052 20768
rect 39092 20728 39093 20768
rect 39051 20719 39093 20728
rect 39244 20768 39284 21316
rect 39628 21307 39668 21316
rect 39628 20768 39668 20777
rect 39244 20719 39284 20728
rect 39532 20728 39628 20768
rect 39052 20634 39092 20719
rect 38667 19928 38709 19937
rect 38667 19888 38668 19928
rect 38708 19888 38709 19928
rect 38667 19879 38709 19888
rect 39532 19928 39572 20728
rect 39628 20719 39668 20728
rect 39724 20180 39764 22240
rect 39724 20131 39764 20140
rect 39820 20096 39860 22651
rect 40203 22532 40245 22541
rect 40203 22492 40204 22532
rect 40244 22492 40245 22532
rect 40203 22483 40245 22492
rect 40108 22280 40148 22289
rect 39915 21356 39957 21365
rect 39915 21316 39916 21356
rect 39956 21316 39957 21356
rect 39915 21307 39957 21316
rect 39916 20777 39956 21307
rect 39915 20768 39957 20777
rect 39915 20728 39916 20768
rect 39956 20728 39957 20768
rect 39915 20719 39957 20728
rect 39820 20047 39860 20056
rect 39916 20096 39956 20719
rect 39916 20047 39956 20056
rect 40011 20096 40053 20105
rect 40011 20056 40012 20096
rect 40052 20056 40053 20096
rect 40011 20047 40053 20056
rect 40012 19962 40052 20047
rect 40108 19928 40148 22240
rect 40204 21356 40244 22483
rect 40300 21776 40340 23080
rect 40588 23120 40628 23491
rect 40780 23465 40820 23584
rect 41068 23624 41108 23635
rect 41068 23549 41108 23584
rect 41067 23540 41109 23549
rect 41067 23500 41068 23540
rect 41108 23500 41109 23540
rect 41067 23491 41109 23500
rect 41740 23465 41780 23752
rect 41835 23792 41877 23801
rect 41835 23752 41836 23792
rect 41876 23752 41877 23792
rect 41835 23743 41877 23752
rect 41932 23792 41972 25096
rect 42700 25087 42740 25096
rect 43179 25136 43221 25145
rect 43179 25096 43180 25136
rect 43220 25096 43221 25136
rect 43179 25087 43221 25096
rect 43276 24632 43316 26272
rect 43371 26263 43413 26272
rect 43564 26312 43604 27616
rect 43660 27581 43700 27616
rect 43756 27656 43796 28120
rect 43892 28120 44084 28160
rect 43852 28111 43892 28120
rect 43851 27740 43893 27749
rect 43851 27700 43852 27740
rect 43892 27700 43893 27740
rect 43851 27691 43893 27700
rect 43756 27607 43796 27616
rect 43852 27656 43892 27691
rect 43852 27605 43892 27616
rect 43947 27656 43989 27665
rect 43947 27616 43948 27656
rect 43988 27616 43989 27656
rect 43947 27607 43989 27616
rect 43659 27572 43701 27581
rect 43659 27532 43660 27572
rect 43700 27532 43701 27572
rect 43659 27523 43701 27532
rect 43660 27492 43700 27523
rect 43948 27522 43988 27607
rect 44044 27329 44084 28120
rect 44523 28120 44524 28160
rect 44564 28120 44565 28160
rect 44523 28111 44565 28120
rect 45004 27833 45044 28288
rect 45100 28278 45140 28363
rect 45484 28328 45524 30379
rect 46444 30294 46484 30379
rect 45771 29840 45813 29849
rect 45771 29800 45772 29840
rect 45812 29800 45813 29840
rect 45771 29791 45813 29800
rect 45963 29840 46005 29849
rect 45963 29800 45964 29840
rect 46004 29800 46005 29840
rect 45963 29791 46005 29800
rect 45772 29706 45812 29791
rect 45867 29672 45909 29681
rect 45867 29632 45868 29672
rect 45908 29632 45909 29672
rect 45867 29623 45909 29632
rect 45868 29168 45908 29623
rect 45868 29119 45908 29128
rect 45964 29000 46004 29791
rect 46732 29000 46772 30388
rect 46924 30176 46964 31387
rect 47212 30848 47252 32143
rect 47404 31940 47444 31949
rect 47308 31352 47348 31361
rect 47404 31352 47444 31900
rect 47499 31940 47541 31949
rect 47499 31900 47500 31940
rect 47540 31900 47541 31940
rect 47499 31891 47541 31900
rect 47348 31312 47444 31352
rect 47308 31303 47348 31312
rect 47212 30799 47252 30808
rect 47020 30680 47060 30689
rect 47020 30437 47060 30640
rect 47115 30680 47157 30689
rect 47115 30640 47116 30680
rect 47156 30640 47157 30680
rect 47115 30631 47157 30640
rect 47308 30680 47348 30689
rect 47500 30680 47540 31891
rect 47692 31352 47732 31361
rect 47788 31352 47828 32152
rect 48075 32143 48117 32152
rect 48268 32192 48308 32201
rect 48076 32058 48116 32143
rect 47883 31520 47925 31529
rect 47883 31480 47884 31520
rect 47924 31480 47925 31520
rect 47883 31471 47925 31480
rect 47732 31312 47828 31352
rect 47692 31303 47732 31312
rect 47884 31277 47924 31471
rect 48268 31445 48308 32152
rect 48363 32192 48405 32201
rect 48363 32152 48364 32192
rect 48404 32152 48405 32192
rect 48363 32143 48405 32152
rect 48460 32192 48500 32201
rect 48364 32058 48404 32143
rect 48460 31940 48500 32152
rect 48556 32192 48596 32201
rect 48556 31949 48596 32152
rect 49803 32192 49845 32201
rect 49803 32152 49804 32192
rect 49844 32152 49845 32192
rect 49803 32143 49845 32152
rect 48364 31900 48500 31940
rect 48555 31940 48597 31949
rect 48555 31900 48556 31940
rect 48596 31900 48597 31940
rect 48364 31529 48404 31900
rect 48555 31891 48597 31900
rect 49132 31940 49172 31949
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 48363 31520 48405 31529
rect 48363 31480 48364 31520
rect 48404 31480 48405 31520
rect 48363 31471 48405 31480
rect 48267 31436 48309 31445
rect 48267 31396 48268 31436
rect 48308 31396 48309 31436
rect 48267 31387 48309 31396
rect 48556 31352 48596 31361
rect 48364 31312 48556 31352
rect 47883 31268 47925 31277
rect 47883 31228 47884 31268
rect 47924 31228 47925 31268
rect 47883 31219 47925 31228
rect 47691 30680 47733 30689
rect 47348 30640 47540 30680
rect 47596 30640 47692 30680
rect 47732 30640 47733 30680
rect 47308 30631 47348 30640
rect 47116 30546 47156 30631
rect 47019 30428 47061 30437
rect 47019 30388 47020 30428
rect 47060 30388 47061 30428
rect 47019 30379 47061 30388
rect 46924 30136 47060 30176
rect 46923 30008 46965 30017
rect 46923 29968 46924 30008
rect 46964 29968 46965 30008
rect 46923 29959 46965 29968
rect 46924 29765 46964 29959
rect 46923 29756 46965 29765
rect 46923 29716 46924 29756
rect 46964 29716 46965 29756
rect 46923 29707 46965 29716
rect 47020 29168 47060 30136
rect 47307 29756 47349 29765
rect 47307 29716 47308 29756
rect 47348 29716 47349 29756
rect 47307 29707 47349 29716
rect 47115 29672 47157 29681
rect 47115 29632 47116 29672
rect 47156 29632 47157 29672
rect 47115 29623 47157 29632
rect 47116 29538 47156 29623
rect 47116 29168 47156 29177
rect 47020 29128 47116 29168
rect 47156 29128 47252 29168
rect 47116 29119 47156 29128
rect 45868 28960 46004 29000
rect 46636 28960 46772 29000
rect 45772 28916 45812 28925
rect 45484 28279 45524 28288
rect 45580 28328 45620 28337
rect 45003 27824 45045 27833
rect 45003 27784 45004 27824
rect 45044 27784 45045 27824
rect 45003 27775 45045 27784
rect 45483 27824 45525 27833
rect 45483 27784 45484 27824
rect 45524 27784 45525 27824
rect 45483 27775 45525 27784
rect 44427 27740 44469 27749
rect 44427 27700 44428 27740
rect 44468 27700 44469 27740
rect 44427 27691 44469 27700
rect 44332 27656 44372 27665
rect 44043 27320 44085 27329
rect 44043 27280 44044 27320
rect 44084 27280 44085 27320
rect 44043 27271 44085 27280
rect 44139 26900 44181 26909
rect 44139 26860 44140 26900
rect 44180 26860 44181 26900
rect 44139 26851 44181 26860
rect 44140 26766 44180 26851
rect 44332 26816 44372 27616
rect 44428 27606 44468 27691
rect 44524 27656 44564 27665
rect 44524 27077 44564 27616
rect 45100 27656 45140 27665
rect 45100 27329 45140 27616
rect 45195 27656 45237 27665
rect 45195 27616 45196 27656
rect 45236 27616 45237 27656
rect 45195 27607 45237 27616
rect 45292 27656 45332 27665
rect 45196 27522 45236 27607
rect 45099 27320 45141 27329
rect 45099 27280 45100 27320
rect 45140 27280 45141 27320
rect 45099 27271 45141 27280
rect 44523 27068 44565 27077
rect 44523 27028 44524 27068
rect 44564 27028 44565 27068
rect 44523 27019 44565 27028
rect 45003 26900 45045 26909
rect 45003 26860 45004 26900
rect 45044 26860 45045 26900
rect 45003 26851 45045 26860
rect 45004 26816 45044 26851
rect 44332 26776 44468 26816
rect 43755 26648 43797 26657
rect 43755 26608 43756 26648
rect 43796 26608 43797 26648
rect 43755 26599 43797 26608
rect 44331 26648 44373 26657
rect 44331 26608 44332 26648
rect 44372 26608 44373 26648
rect 44331 26599 44373 26608
rect 43564 26263 43604 26272
rect 43659 26312 43701 26321
rect 43659 26272 43660 26312
rect 43700 26272 43701 26312
rect 43659 26263 43701 26272
rect 43372 26144 43412 26153
rect 43660 26144 43700 26263
rect 43412 26104 43604 26144
rect 43372 26095 43412 26104
rect 43372 25892 43412 25901
rect 43372 25304 43412 25852
rect 43467 25640 43509 25649
rect 43467 25600 43468 25640
rect 43508 25600 43509 25640
rect 43467 25591 43509 25600
rect 43372 25255 43412 25264
rect 43372 24632 43412 24641
rect 43276 24592 43372 24632
rect 43468 24632 43508 25591
rect 43564 25304 43604 26104
rect 43660 26095 43700 26104
rect 43756 26144 43796 26599
rect 44332 26514 44372 26599
rect 43851 26312 43893 26321
rect 43851 26272 43852 26312
rect 43892 26272 43893 26312
rect 43851 26263 43893 26272
rect 43756 26095 43796 26104
rect 43852 26144 43892 26263
rect 44235 26228 44277 26237
rect 44235 26188 44236 26228
rect 44276 26188 44277 26228
rect 44235 26179 44277 26188
rect 43852 25649 43892 26104
rect 44139 26144 44181 26153
rect 44139 26104 44140 26144
rect 44180 26104 44181 26144
rect 44139 26095 44181 26104
rect 43851 25640 43893 25649
rect 43851 25600 43852 25640
rect 43892 25600 43893 25640
rect 43851 25591 43893 25600
rect 44140 25481 44180 26095
rect 44236 26094 44276 26179
rect 44428 26153 44468 26776
rect 45004 26765 45044 26776
rect 45292 26405 45332 27616
rect 45387 27656 45429 27665
rect 45387 27616 45388 27656
rect 45428 27616 45429 27656
rect 45387 27607 45429 27616
rect 45388 27522 45428 27607
rect 45387 27404 45429 27413
rect 45387 27364 45388 27404
rect 45428 27364 45429 27404
rect 45387 27355 45429 27364
rect 45099 26396 45141 26405
rect 45099 26356 45100 26396
rect 45140 26356 45141 26396
rect 45099 26347 45141 26356
rect 45291 26396 45333 26405
rect 45291 26356 45292 26396
rect 45332 26356 45333 26396
rect 45291 26347 45333 26356
rect 44523 26312 44565 26321
rect 44523 26272 44524 26312
rect 44564 26272 44565 26312
rect 44523 26263 44565 26272
rect 44332 26144 44372 26153
rect 44332 25976 44372 26104
rect 44427 26144 44469 26153
rect 44427 26104 44428 26144
rect 44468 26104 44469 26144
rect 44427 26095 44469 26104
rect 44524 26144 44564 26263
rect 44716 26153 44756 26238
rect 44524 26095 44564 26104
rect 44715 26144 44757 26153
rect 44715 26104 44716 26144
rect 44756 26104 44757 26144
rect 44715 26095 44757 26104
rect 44907 26144 44949 26153
rect 44907 26104 44908 26144
rect 44948 26104 44949 26144
rect 44907 26095 44949 26104
rect 44908 26010 44948 26095
rect 44812 25976 44852 25985
rect 44332 25936 44812 25976
rect 44812 25927 44852 25936
rect 44523 25640 44565 25649
rect 44523 25600 44524 25640
rect 44564 25600 44565 25640
rect 44523 25591 44565 25600
rect 44332 25481 44372 25566
rect 44139 25472 44181 25481
rect 44139 25432 44140 25472
rect 44180 25432 44181 25472
rect 44139 25423 44181 25432
rect 44331 25472 44373 25481
rect 44331 25432 44332 25472
rect 44372 25432 44373 25472
rect 44331 25423 44373 25432
rect 43851 25388 43893 25397
rect 43851 25348 43852 25388
rect 43892 25348 43893 25388
rect 43851 25339 43893 25348
rect 43756 25304 43796 25313
rect 43564 25264 43756 25304
rect 43756 25255 43796 25264
rect 43852 25304 43892 25339
rect 43852 25253 43892 25264
rect 43948 25304 43988 25313
rect 43948 24977 43988 25264
rect 44044 25304 44084 25313
rect 44332 25304 44372 25313
rect 44044 25145 44084 25264
rect 44140 25264 44332 25304
rect 44043 25136 44085 25145
rect 44043 25096 44044 25136
rect 44084 25096 44085 25136
rect 44043 25087 44085 25096
rect 43947 24968 43989 24977
rect 43947 24928 43948 24968
rect 43988 24928 43989 24968
rect 43947 24919 43989 24928
rect 44140 24800 44180 25264
rect 44332 25255 44372 25264
rect 44524 25304 44564 25591
rect 44811 25472 44853 25481
rect 44811 25432 44812 25472
rect 44852 25432 44853 25472
rect 44811 25423 44853 25432
rect 44524 25255 44564 25264
rect 44619 25304 44661 25313
rect 44619 25264 44620 25304
rect 44660 25264 44661 25304
rect 44619 25255 44661 25264
rect 44812 25304 44852 25423
rect 45100 25397 45140 26347
rect 45292 25976 45332 25985
rect 45099 25388 45141 25397
rect 45099 25348 45100 25388
rect 45140 25348 45141 25388
rect 45099 25339 45141 25348
rect 44812 25255 44852 25264
rect 44620 25170 44660 25255
rect 44715 25220 44757 25229
rect 44715 25180 44716 25220
rect 44756 25180 44757 25220
rect 44715 25171 44757 25180
rect 44331 25136 44373 25145
rect 44331 25096 44332 25136
rect 44372 25096 44373 25136
rect 44331 25087 44373 25096
rect 44235 24968 44277 24977
rect 44235 24928 44236 24968
rect 44276 24928 44277 24968
rect 44235 24919 44277 24928
rect 44140 24751 44180 24760
rect 43947 24716 43989 24725
rect 43947 24676 43948 24716
rect 43988 24676 43989 24716
rect 43947 24667 43989 24676
rect 43852 24632 43892 24641
rect 43468 24592 43852 24632
rect 41932 23743 41972 23752
rect 42316 24464 42356 24473
rect 42316 23792 42356 24424
rect 42988 24380 43028 24389
rect 42988 23801 43028 24340
rect 43372 23885 43412 24592
rect 43852 24583 43892 24592
rect 43948 24632 43988 24667
rect 43948 24581 43988 24592
rect 44044 24632 44084 24641
rect 43371 23876 43413 23885
rect 43371 23836 43372 23876
rect 43412 23836 43413 23876
rect 43371 23827 43413 23836
rect 44044 23801 44084 24592
rect 44236 23960 44276 24919
rect 44332 24893 44372 25087
rect 44331 24884 44373 24893
rect 44331 24844 44332 24884
rect 44372 24844 44373 24884
rect 44331 24835 44373 24844
rect 44332 24632 44372 24835
rect 44523 24800 44565 24809
rect 44523 24760 44524 24800
rect 44564 24760 44565 24800
rect 44523 24751 44565 24760
rect 44620 24800 44660 24809
rect 44716 24800 44756 25171
rect 44811 25052 44853 25061
rect 44811 25012 44812 25052
rect 44852 25012 44853 25052
rect 44811 25003 44853 25012
rect 44660 24760 44756 24800
rect 44620 24751 44660 24760
rect 44332 24583 44372 24592
rect 44428 24632 44468 24641
rect 44332 23960 44372 23969
rect 44236 23920 44332 23960
rect 44332 23911 44372 23920
rect 42316 23743 42356 23752
rect 42987 23792 43029 23801
rect 42987 23752 42988 23792
rect 43028 23752 43029 23792
rect 42987 23743 43029 23752
rect 43180 23792 43220 23801
rect 40779 23456 40821 23465
rect 40779 23416 40780 23456
rect 40820 23416 40821 23456
rect 40779 23407 40821 23416
rect 41739 23456 41781 23465
rect 41739 23416 41740 23456
rect 41780 23416 41781 23456
rect 41739 23407 41781 23416
rect 40588 23071 40628 23080
rect 40684 23120 40724 23129
rect 41260 23120 41300 23129
rect 40724 23080 41260 23120
rect 40684 23071 40724 23080
rect 41260 23071 41300 23080
rect 41356 23120 41396 23129
rect 41068 22952 41108 22961
rect 40587 22868 40629 22877
rect 40587 22828 40588 22868
rect 40628 22828 40629 22868
rect 40587 22819 40629 22828
rect 40395 22448 40437 22457
rect 40395 22408 40396 22448
rect 40436 22408 40437 22448
rect 40395 22399 40437 22408
rect 40396 22280 40436 22399
rect 40396 22205 40436 22240
rect 40395 22196 40437 22205
rect 40395 22156 40396 22196
rect 40436 22156 40437 22196
rect 40395 22147 40437 22156
rect 40300 21736 40436 21776
rect 40299 21608 40341 21617
rect 40299 21568 40300 21608
rect 40340 21568 40341 21608
rect 40299 21559 40341 21568
rect 40300 21474 40340 21559
rect 40396 21449 40436 21736
rect 40395 21440 40437 21449
rect 40395 21400 40396 21440
rect 40436 21400 40437 21440
rect 40395 21391 40437 21400
rect 40491 21356 40533 21365
rect 40204 21316 40340 21356
rect 40300 21272 40340 21316
rect 40491 21316 40492 21356
rect 40532 21316 40533 21356
rect 40491 21307 40533 21316
rect 40300 21232 40436 21272
rect 40396 20105 40436 21232
rect 40492 21222 40532 21307
rect 40492 20768 40532 20777
rect 40588 20768 40628 22819
rect 41068 22793 41108 22912
rect 41067 22784 41109 22793
rect 41067 22744 41068 22784
rect 41108 22744 41109 22784
rect 41067 22735 41109 22744
rect 41356 22709 41396 23080
rect 41548 23120 41588 23129
rect 41740 23120 41780 23129
rect 41588 23080 41740 23120
rect 41548 23071 41588 23080
rect 41740 23071 41780 23080
rect 41836 23120 41876 23743
rect 41931 23540 41973 23549
rect 41931 23500 41932 23540
rect 41972 23500 41973 23540
rect 41931 23491 41973 23500
rect 41451 23036 41493 23045
rect 41451 22996 41452 23036
rect 41492 22996 41493 23036
rect 41451 22987 41493 22996
rect 41355 22700 41397 22709
rect 41355 22660 41356 22700
rect 41396 22660 41397 22700
rect 41355 22651 41397 22660
rect 40683 22532 40725 22541
rect 40683 22492 40684 22532
rect 40724 22492 40725 22532
rect 40683 22483 40725 22492
rect 40684 22398 40724 22483
rect 41356 22280 41396 22651
rect 41356 22231 41396 22240
rect 41163 21608 41205 21617
rect 41163 21568 41164 21608
rect 41204 21568 41205 21608
rect 41163 21559 41205 21568
rect 41452 21608 41492 22987
rect 41547 22952 41589 22961
rect 41836 22952 41876 23080
rect 41932 23120 41972 23491
rect 43083 23288 43125 23297
rect 43083 23248 43084 23288
rect 43124 23248 43125 23288
rect 43083 23239 43125 23248
rect 43084 23154 43124 23239
rect 41932 23071 41972 23080
rect 42028 23120 42068 23129
rect 41547 22912 41548 22952
rect 41588 22912 41589 22952
rect 41547 22903 41589 22912
rect 41644 22912 41876 22952
rect 41548 22818 41588 22903
rect 41644 22541 41684 22912
rect 42028 22709 42068 23080
rect 42220 23120 42260 23129
rect 42220 22961 42260 23080
rect 42219 22952 42261 22961
rect 42219 22912 42220 22952
rect 42260 22912 42261 22952
rect 42219 22903 42261 22912
rect 43180 22877 43220 23752
rect 44043 23792 44085 23801
rect 44043 23752 44044 23792
rect 44084 23752 44085 23792
rect 44043 23743 44085 23752
rect 43563 23120 43605 23129
rect 43563 23080 43564 23120
rect 43604 23080 43605 23120
rect 43563 23071 43605 23080
rect 43756 23120 43796 23129
rect 42892 22868 42932 22877
rect 42699 22784 42741 22793
rect 42699 22744 42700 22784
rect 42740 22744 42741 22784
rect 42699 22735 42741 22744
rect 42027 22700 42069 22709
rect 42027 22660 42028 22700
rect 42068 22660 42069 22700
rect 42027 22651 42069 22660
rect 42315 22700 42357 22709
rect 42315 22660 42316 22700
rect 42356 22660 42357 22700
rect 42315 22651 42357 22660
rect 41739 22616 41781 22625
rect 41739 22576 41740 22616
rect 41780 22576 41781 22616
rect 41739 22567 41781 22576
rect 41643 22532 41685 22541
rect 41643 22492 41644 22532
rect 41684 22492 41685 22532
rect 41643 22483 41685 22492
rect 41644 22280 41684 22483
rect 41644 22231 41684 22240
rect 41740 22280 41780 22567
rect 42028 22448 42068 22651
rect 42123 22532 42165 22541
rect 42123 22492 42124 22532
rect 42164 22492 42165 22532
rect 42123 22483 42165 22492
rect 41740 22231 41780 22240
rect 41836 22408 42068 22448
rect 41836 22280 41876 22408
rect 41547 22112 41589 22121
rect 41547 22072 41548 22112
rect 41588 22072 41589 22112
rect 41547 22063 41589 22072
rect 41548 21978 41588 22063
rect 41452 21559 41492 21568
rect 41547 21608 41589 21617
rect 41547 21568 41548 21608
rect 41588 21568 41589 21608
rect 41547 21559 41589 21568
rect 41644 21608 41684 21617
rect 41164 21474 41204 21559
rect 41451 21440 41493 21449
rect 41451 21400 41452 21440
rect 41492 21400 41493 21440
rect 41548 21440 41588 21559
rect 41548 21400 41600 21440
rect 41451 21391 41493 21400
rect 41356 21356 41396 21365
rect 40532 20728 40628 20768
rect 40684 21316 41356 21356
rect 40492 20719 40532 20728
rect 40684 20180 40724 21316
rect 41356 21307 41396 21316
rect 40492 20140 40724 20180
rect 40204 20096 40244 20105
rect 40395 20096 40437 20105
rect 40244 20056 40340 20096
rect 40204 20047 40244 20056
rect 40300 19937 40340 20056
rect 40395 20056 40396 20096
rect 40436 20056 40437 20096
rect 40395 20047 40437 20056
rect 40492 20096 40532 20140
rect 40492 20047 40532 20056
rect 40396 19962 40436 20047
rect 40204 19928 40244 19937
rect 40108 19888 40204 19928
rect 39532 19879 39572 19888
rect 40204 19879 40244 19888
rect 40299 19928 40341 19937
rect 40299 19888 40300 19928
rect 40340 19888 40341 19928
rect 40299 19879 40341 19888
rect 37419 18668 37461 18677
rect 37419 18628 37420 18668
rect 37460 18628 37461 18668
rect 37419 18619 37461 18628
rect 36652 18376 37172 18416
rect 37228 18584 37268 18593
rect 36652 17828 36692 18376
rect 37228 18248 37268 18544
rect 36652 17779 36692 17788
rect 36748 18208 37268 18248
rect 37324 18584 37364 18593
rect 36555 17744 36597 17753
rect 36555 17704 36556 17744
rect 36596 17704 36597 17744
rect 36555 17695 36597 17704
rect 36748 17744 36788 18208
rect 37324 18089 37364 18544
rect 37420 18584 37460 18619
rect 37035 18080 37077 18089
rect 37035 18040 37036 18080
rect 37076 18040 37077 18080
rect 37035 18031 37077 18040
rect 37323 18080 37365 18089
rect 37323 18040 37324 18080
rect 37364 18040 37365 18080
rect 37323 18031 37365 18040
rect 36748 17695 36788 17704
rect 37036 17744 37076 18031
rect 37131 17996 37173 18005
rect 37131 17956 37132 17996
rect 37172 17956 37173 17996
rect 37131 17947 37173 17956
rect 37036 17695 37076 17704
rect 37132 17723 37172 17947
rect 36556 17610 36596 17695
rect 37227 17744 37269 17753
rect 37227 17704 37228 17744
rect 37268 17704 37269 17744
rect 37227 17695 37269 17704
rect 36939 17660 36981 17669
rect 36939 17620 36940 17660
rect 36980 17620 36981 17660
rect 36939 17611 36981 17620
rect 36843 17576 36885 17585
rect 36843 17536 36844 17576
rect 36884 17536 36885 17576
rect 36843 17527 36885 17536
rect 36651 17492 36693 17501
rect 36651 17452 36652 17492
rect 36692 17452 36693 17492
rect 36651 17443 36693 17452
rect 36459 17240 36501 17249
rect 36459 17200 36460 17240
rect 36500 17200 36501 17240
rect 36459 17191 36501 17200
rect 36652 17240 36692 17443
rect 36652 17191 36692 17200
rect 36307 17156 36349 17165
rect 36307 17116 36308 17156
rect 36348 17116 36349 17156
rect 36307 17107 36349 17116
rect 35884 17023 35924 17032
rect 36076 17072 36116 17081
rect 36308 17072 36348 17107
rect 36116 17032 36212 17072
rect 36076 17023 36116 17032
rect 35788 16948 35830 16988
rect 35788 16652 35828 16948
rect 35980 16820 36020 16829
rect 35788 16612 35924 16652
rect 35787 16484 35829 16493
rect 35787 16444 35788 16484
rect 35828 16444 35829 16484
rect 35787 16435 35829 16444
rect 35788 16232 35828 16435
rect 35788 16183 35828 16192
rect 35884 16148 35924 16612
rect 35980 16493 36020 16780
rect 35979 16484 36021 16493
rect 35979 16444 35980 16484
rect 36020 16444 36021 16484
rect 35979 16435 36021 16444
rect 35884 16099 35924 16108
rect 35980 16232 36020 16241
rect 35980 16073 36020 16192
rect 36076 16232 36116 16241
rect 36172 16232 36212 17032
rect 36308 17022 36348 17032
rect 36460 17072 36500 17191
rect 36460 17023 36500 17032
rect 36556 17072 36596 17081
rect 36556 16997 36596 17032
rect 36748 17072 36788 17081
rect 36555 16988 36597 16997
rect 36555 16948 36556 16988
rect 36596 16948 36597 16988
rect 36555 16939 36597 16948
rect 36556 16829 36596 16939
rect 36555 16820 36597 16829
rect 36555 16780 36556 16820
rect 36596 16780 36597 16820
rect 36555 16771 36597 16780
rect 36748 16493 36788 17032
rect 36844 17072 36884 17527
rect 36940 17526 36980 17611
rect 37132 17324 37172 17683
rect 37228 17610 37268 17695
rect 36844 17023 36884 17032
rect 36940 17284 37172 17324
rect 37227 17324 37269 17333
rect 37227 17284 37228 17324
rect 37268 17284 37269 17324
rect 36940 16661 36980 17284
rect 37227 17275 37269 17284
rect 37072 17156 37114 17165
rect 37072 17116 37073 17156
rect 37113 17116 37114 17156
rect 37072 17107 37114 17116
rect 37073 17072 37113 17107
rect 37073 17021 37113 17032
rect 37228 17072 37268 17275
rect 37324 17249 37364 18031
rect 37420 18005 37460 18544
rect 37516 18584 37556 18593
rect 37516 18257 37556 18544
rect 37803 18584 37845 18593
rect 37803 18544 37804 18584
rect 37844 18544 37845 18584
rect 37803 18535 37845 18544
rect 37900 18584 37940 18593
rect 37515 18248 37557 18257
rect 37515 18208 37516 18248
rect 37556 18208 37557 18248
rect 37515 18199 37557 18208
rect 37419 17996 37461 18005
rect 37419 17956 37420 17996
rect 37460 17956 37461 17996
rect 37419 17947 37461 17956
rect 37708 17921 37748 18006
rect 37707 17912 37749 17921
rect 37707 17872 37708 17912
rect 37748 17872 37749 17912
rect 37707 17863 37749 17872
rect 37420 17744 37460 17753
rect 37420 17501 37460 17704
rect 37516 17744 37556 17753
rect 37708 17744 37748 17753
rect 37556 17704 37652 17744
rect 37516 17695 37556 17704
rect 37515 17576 37557 17585
rect 37515 17536 37516 17576
rect 37556 17536 37557 17576
rect 37515 17527 37557 17536
rect 37419 17492 37461 17501
rect 37419 17452 37420 17492
rect 37460 17452 37461 17492
rect 37419 17443 37461 17452
rect 37323 17240 37365 17249
rect 37323 17200 37324 17240
rect 37364 17200 37365 17240
rect 37323 17191 37365 17200
rect 37516 17156 37556 17527
rect 37612 17240 37652 17704
rect 37708 17585 37748 17704
rect 37707 17576 37749 17585
rect 37707 17536 37708 17576
rect 37748 17536 37749 17576
rect 37804 17576 37844 18535
rect 37900 18257 37940 18544
rect 37899 18248 37941 18257
rect 37899 18208 37900 18248
rect 37940 18208 37941 18248
rect 37899 18199 37941 18208
rect 37900 17872 38324 17912
rect 37900 17744 37940 17872
rect 37900 17695 37940 17704
rect 37995 17744 38037 17753
rect 37995 17704 37996 17744
rect 38036 17704 38037 17744
rect 37995 17695 38037 17704
rect 37804 17536 37940 17576
rect 37707 17527 37749 17536
rect 37612 17200 37748 17240
rect 37516 17116 37652 17156
rect 37612 17072 37652 17116
rect 37228 17023 37268 17032
rect 37324 17057 37364 17066
rect 37324 16997 37364 17017
rect 37516 17057 37556 17066
rect 37708 17072 37748 17200
rect 37708 17032 37844 17072
rect 37612 17023 37652 17032
rect 37323 16988 37365 16997
rect 37323 16948 37324 16988
rect 37364 16948 37365 16988
rect 37323 16939 37365 16948
rect 37324 16922 37364 16939
rect 36939 16652 36981 16661
rect 36939 16612 36940 16652
rect 36980 16612 36981 16652
rect 36939 16603 36981 16612
rect 37419 16652 37461 16661
rect 37419 16612 37420 16652
rect 37460 16612 37461 16652
rect 37419 16603 37461 16612
rect 36555 16484 36597 16493
rect 36555 16444 36556 16484
rect 36596 16444 36597 16484
rect 36555 16435 36597 16444
rect 36747 16484 36789 16493
rect 36747 16444 36748 16484
rect 36788 16444 36789 16484
rect 36747 16435 36789 16444
rect 37323 16484 37365 16493
rect 37323 16444 37324 16484
rect 37364 16444 37365 16484
rect 37323 16435 37365 16444
rect 36268 16232 36308 16241
rect 36172 16192 36268 16232
rect 35979 16064 36021 16073
rect 35979 16024 35980 16064
rect 36020 16024 36021 16064
rect 35979 16015 36021 16024
rect 35883 15812 35925 15821
rect 35883 15772 35884 15812
rect 35924 15772 35925 15812
rect 35883 15763 35925 15772
rect 35788 15728 35828 15737
rect 35692 15688 35788 15728
rect 35595 15644 35637 15653
rect 35595 15604 35596 15644
rect 35636 15604 35637 15644
rect 35595 15595 35637 15604
rect 35404 15560 35444 15571
rect 35404 15485 35444 15520
rect 35596 15560 35636 15595
rect 35596 15509 35636 15520
rect 35691 15560 35733 15569
rect 35691 15520 35692 15560
rect 35732 15520 35733 15560
rect 35691 15511 35733 15520
rect 35403 15476 35445 15485
rect 35403 15436 35404 15476
rect 35444 15436 35445 15476
rect 35403 15427 35445 15436
rect 35595 15392 35637 15401
rect 35595 15352 35596 15392
rect 35636 15352 35637 15392
rect 35595 15343 35637 15352
rect 35596 15258 35636 15343
rect 35692 14972 35732 15511
rect 35692 14923 35732 14932
rect 35788 14720 35828 15688
rect 35884 15560 35924 15763
rect 36076 15737 36116 16192
rect 36268 16183 36308 16192
rect 36364 16232 36404 16241
rect 36267 16064 36309 16073
rect 36267 16024 36268 16064
rect 36308 16024 36309 16064
rect 36267 16015 36309 16024
rect 36075 15728 36117 15737
rect 36075 15688 36076 15728
rect 36116 15688 36117 15728
rect 36075 15679 36117 15688
rect 36171 15644 36213 15653
rect 36171 15604 36172 15644
rect 36212 15604 36213 15644
rect 36268 15644 36308 16015
rect 36364 15821 36404 16192
rect 36459 16232 36501 16241
rect 36459 16192 36460 16232
rect 36500 16192 36501 16232
rect 36459 16183 36501 16192
rect 36556 16232 36596 16435
rect 36651 16400 36693 16409
rect 36651 16360 36652 16400
rect 36692 16360 36693 16400
rect 36651 16351 36693 16360
rect 37035 16400 37077 16409
rect 37035 16360 37036 16400
rect 37076 16360 37077 16400
rect 37035 16351 37077 16360
rect 36460 16098 36500 16183
rect 36556 15905 36596 16192
rect 36555 15896 36597 15905
rect 36555 15856 36556 15896
rect 36596 15856 36597 15896
rect 36555 15847 36597 15856
rect 36363 15812 36405 15821
rect 36363 15772 36364 15812
rect 36404 15772 36500 15812
rect 36363 15763 36405 15772
rect 36268 15604 36404 15644
rect 36171 15595 36213 15604
rect 35884 15511 35924 15520
rect 35980 15560 36020 15569
rect 35980 14720 36020 15520
rect 36076 15560 36116 15569
rect 36076 15149 36116 15520
rect 36075 15140 36117 15149
rect 36075 15100 36076 15140
rect 36116 15100 36117 15140
rect 36075 15091 36117 15100
rect 36076 14972 36116 14981
rect 36172 14972 36212 15595
rect 36364 15560 36404 15604
rect 36268 15541 36308 15550
rect 36268 15401 36308 15501
rect 36267 15392 36309 15401
rect 36267 15352 36268 15392
rect 36308 15352 36309 15392
rect 36267 15343 36309 15352
rect 36364 15233 36404 15520
rect 36363 15224 36405 15233
rect 36363 15184 36364 15224
rect 36404 15184 36405 15224
rect 36363 15175 36405 15184
rect 36267 15140 36309 15149
rect 36267 15100 36268 15140
rect 36308 15100 36309 15140
rect 36267 15091 36309 15100
rect 36116 14932 36212 14972
rect 36076 14923 36116 14932
rect 36268 14720 36308 15091
rect 35980 14680 36116 14720
rect 35788 14671 35828 14680
rect 36076 14057 36116 14680
rect 36268 14561 36308 14680
rect 36364 14720 36404 14729
rect 36460 14720 36500 15772
rect 36555 15560 36597 15569
rect 36555 15520 36556 15560
rect 36596 15520 36597 15560
rect 36555 15511 36597 15520
rect 36556 15426 36596 15511
rect 36555 15308 36597 15317
rect 36555 15268 36556 15308
rect 36596 15268 36597 15308
rect 36555 15259 36597 15268
rect 36556 15174 36596 15259
rect 36404 14680 36500 14720
rect 36652 14720 36692 16351
rect 37036 16266 37076 16351
rect 36940 16232 36980 16241
rect 36844 15737 36884 15822
rect 36843 15728 36885 15737
rect 36843 15688 36844 15728
rect 36884 15688 36885 15728
rect 36843 15679 36885 15688
rect 36940 15653 36980 16192
rect 37132 16232 37172 16241
rect 37132 16073 37172 16192
rect 37324 16232 37364 16435
rect 37324 16183 37364 16192
rect 37420 16232 37460 16603
rect 37516 16577 37556 17017
rect 37707 16904 37749 16913
rect 37707 16864 37708 16904
rect 37748 16864 37749 16904
rect 37707 16855 37749 16864
rect 37611 16820 37653 16829
rect 37611 16780 37612 16820
rect 37652 16780 37653 16820
rect 37611 16771 37653 16780
rect 37612 16686 37652 16771
rect 37515 16568 37557 16577
rect 37515 16528 37516 16568
rect 37556 16528 37557 16568
rect 37515 16519 37557 16528
rect 37420 16183 37460 16192
rect 37516 16232 37556 16241
rect 37516 16157 37556 16192
rect 37612 16232 37652 16241
rect 37708 16232 37748 16855
rect 37652 16192 37748 16232
rect 37612 16183 37652 16192
rect 37515 16148 37557 16157
rect 37515 16108 37516 16148
rect 37556 16108 37557 16148
rect 37515 16099 37557 16108
rect 37131 16064 37173 16073
rect 37131 16024 37132 16064
rect 37172 16024 37173 16064
rect 37131 16015 37173 16024
rect 37323 15896 37365 15905
rect 37323 15856 37324 15896
rect 37364 15856 37365 15896
rect 37323 15847 37365 15856
rect 37324 15653 37364 15847
rect 37516 15728 37556 16099
rect 37804 15905 37844 17032
rect 37803 15896 37845 15905
rect 37803 15856 37804 15896
rect 37844 15856 37845 15896
rect 37803 15847 37845 15856
rect 37420 15688 37556 15728
rect 36939 15644 36981 15653
rect 36939 15604 36940 15644
rect 36980 15604 36981 15644
rect 36939 15595 36981 15604
rect 37323 15644 37365 15653
rect 37323 15604 37324 15644
rect 37364 15604 37365 15644
rect 37323 15595 37365 15604
rect 36747 15560 36789 15569
rect 36747 15520 36748 15560
rect 36788 15520 36789 15560
rect 36747 15511 36789 15520
rect 36844 15560 36884 15569
rect 37420 15560 37460 15688
rect 37900 15569 37940 17536
rect 37996 16988 38036 17695
rect 38284 17240 38324 17872
rect 38572 17753 38612 19216
rect 39723 19256 39765 19265
rect 39723 19216 39724 19256
rect 39764 19216 39765 19256
rect 39723 19207 39765 19216
rect 40683 19256 40725 19265
rect 40683 19216 40684 19256
rect 40724 19216 40725 19256
rect 40683 19207 40725 19216
rect 38859 19088 38901 19097
rect 38859 19048 38860 19088
rect 38900 19048 38901 19088
rect 38859 19039 38901 19048
rect 38860 18584 38900 19039
rect 38860 18535 38900 18544
rect 39244 18584 39284 18593
rect 38763 17912 38805 17921
rect 38763 17872 38764 17912
rect 38804 17872 38805 17912
rect 38763 17863 38805 17872
rect 38571 17744 38613 17753
rect 38571 17704 38572 17744
rect 38612 17704 38613 17744
rect 38571 17695 38613 17704
rect 38764 17744 38804 17863
rect 39148 17744 39188 17753
rect 38764 17695 38804 17704
rect 39052 17704 39148 17744
rect 38571 17576 38613 17585
rect 38571 17536 38572 17576
rect 38612 17536 38613 17576
rect 38571 17527 38613 17536
rect 38572 17442 38612 17527
rect 38284 17191 38324 17200
rect 37996 16652 38036 16948
rect 38188 17072 38228 17081
rect 38188 16913 38228 17032
rect 38380 17072 38420 17081
rect 38187 16904 38229 16913
rect 38187 16864 38188 16904
rect 38228 16864 38229 16904
rect 38187 16855 38229 16864
rect 37996 16612 38324 16652
rect 38091 16232 38133 16241
rect 38091 16192 38092 16232
rect 38132 16192 38133 16232
rect 38091 16183 38133 16192
rect 38188 16232 38228 16241
rect 38092 16098 38132 16183
rect 37995 16064 38037 16073
rect 37995 16020 37996 16064
rect 38036 16020 38037 16064
rect 37995 16015 38037 16020
rect 37996 15929 38036 16015
rect 38188 15989 38228 16192
rect 38187 15980 38229 15989
rect 38187 15940 38188 15980
rect 38228 15940 38229 15980
rect 38187 15931 38229 15940
rect 38091 15728 38133 15737
rect 38091 15688 38092 15728
rect 38132 15688 38133 15728
rect 38091 15679 38133 15688
rect 37419 15541 37460 15560
rect 36748 15426 36788 15511
rect 36844 15401 36884 15520
rect 37324 15520 37460 15541
rect 37516 15560 37556 15569
rect 37899 15560 37941 15569
rect 37556 15520 37652 15560
rect 37324 15501 37459 15520
rect 37516 15511 37556 15520
rect 36939 15476 36981 15485
rect 36939 15436 36940 15476
rect 36980 15436 36981 15476
rect 36939 15427 36981 15436
rect 36843 15392 36885 15401
rect 36843 15352 36844 15392
rect 36884 15352 36885 15392
rect 36843 15343 36885 15352
rect 36940 15342 36980 15427
rect 37035 15392 37077 15401
rect 37035 15352 37036 15392
rect 37076 15352 37077 15392
rect 37035 15343 37077 15352
rect 37036 15258 37076 15343
rect 37132 14981 37172 15066
rect 37131 14972 37173 14981
rect 37131 14932 37132 14972
rect 37172 14932 37173 14972
rect 37131 14923 37173 14932
rect 37324 14888 37364 15501
rect 37612 15401 37652 15520
rect 37899 15520 37900 15560
rect 37940 15520 37941 15560
rect 37899 15511 37941 15520
rect 38092 15560 38132 15679
rect 38187 15644 38229 15653
rect 38187 15604 38188 15644
rect 38228 15604 38229 15644
rect 38187 15595 38229 15604
rect 37708 15485 37748 15487
rect 37707 15476 37749 15485
rect 37707 15436 37708 15476
rect 37748 15436 37749 15476
rect 37707 15427 37749 15436
rect 37516 15392 37556 15401
rect 37516 15233 37556 15352
rect 37611 15392 37653 15401
rect 37611 15352 37612 15392
rect 37652 15352 37653 15392
rect 37611 15343 37653 15352
rect 37708 15392 37748 15427
rect 37708 15343 37748 15352
rect 37515 15224 37557 15233
rect 37515 15184 37516 15224
rect 37556 15184 37557 15224
rect 37515 15175 37557 15184
rect 37228 14848 37364 14888
rect 36652 14706 37172 14720
rect 36652 14680 37132 14706
rect 36364 14671 36404 14680
rect 37132 14657 37172 14666
rect 36267 14552 36309 14561
rect 36267 14512 36268 14552
rect 36308 14512 36309 14552
rect 36267 14503 36309 14512
rect 36843 14552 36885 14561
rect 36843 14512 36844 14552
rect 36884 14512 36885 14552
rect 36843 14503 36885 14512
rect 36075 14048 36117 14057
rect 36075 14008 36076 14048
rect 36116 14008 36117 14048
rect 36075 13999 36117 14008
rect 36844 14048 36884 14503
rect 36844 13999 36884 14008
rect 36076 13460 36116 13999
rect 36747 13796 36789 13805
rect 36747 13756 36748 13796
rect 36788 13756 36789 13796
rect 36747 13747 36789 13756
rect 36172 13460 36212 13469
rect 36076 13420 36172 13460
rect 36172 13411 36212 13420
rect 35211 13292 35253 13301
rect 35211 13252 35212 13292
rect 35252 13252 35253 13292
rect 35211 13243 35253 13252
rect 34443 13208 34485 13217
rect 34443 13168 34444 13208
rect 34484 13168 34485 13208
rect 34443 13159 34485 13168
rect 35020 13208 35060 13217
rect 34156 13000 34292 13040
rect 34059 12788 34101 12797
rect 34059 12748 34060 12788
rect 34100 12748 34101 12788
rect 34059 12739 34101 12748
rect 33676 12412 34004 12452
rect 33580 12319 33620 12328
rect 33772 12284 33812 12293
rect 33812 12244 33908 12284
rect 33772 12235 33812 12244
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 33196 11948 33236 11957
rect 33483 11948 33525 11957
rect 33236 11908 33428 11948
rect 33196 11899 33236 11908
rect 33196 11705 33236 11790
rect 33195 11696 33237 11705
rect 33195 11656 33196 11696
rect 33236 11656 33237 11696
rect 33388 11696 33428 11908
rect 33483 11908 33484 11948
rect 33524 11908 33525 11948
rect 33483 11899 33525 11908
rect 33484 11864 33524 11899
rect 33580 11873 33620 11917
rect 33484 11813 33524 11824
rect 33579 11864 33621 11873
rect 33579 11824 33580 11864
rect 33620 11824 33621 11864
rect 33579 11822 33621 11824
rect 33579 11815 33580 11822
rect 33620 11815 33621 11822
rect 33771 11864 33813 11873
rect 33771 11824 33772 11864
rect 33812 11824 33813 11864
rect 33771 11815 33813 11824
rect 33580 11773 33620 11782
rect 33676 11696 33716 11705
rect 33388 11656 33676 11696
rect 33195 11647 33237 11656
rect 33676 11647 33716 11656
rect 33772 11696 33812 11815
rect 33772 11647 33812 11656
rect 33676 11528 33716 11537
rect 33100 11488 33676 11528
rect 33676 11479 33716 11488
rect 33099 11276 33141 11285
rect 33099 11236 33100 11276
rect 33140 11236 33141 11276
rect 33099 11227 33141 11236
rect 32523 11108 32565 11117
rect 32523 11068 32524 11108
rect 32564 11068 32565 11108
rect 32523 11059 32565 11068
rect 32715 11108 32757 11117
rect 32715 11068 32716 11108
rect 32756 11068 32757 11108
rect 32715 11059 32757 11068
rect 32427 11024 32469 11033
rect 32427 10984 32428 11024
rect 32468 10984 32469 11024
rect 32427 10975 32469 10984
rect 32716 11024 32756 11059
rect 32428 10890 32468 10975
rect 32716 10973 32756 10984
rect 33100 11024 33140 11227
rect 33100 10975 33140 10984
rect 32812 10940 32852 10949
rect 32523 10856 32565 10865
rect 32523 10816 32524 10856
rect 32564 10816 32565 10856
rect 32523 10807 32565 10816
rect 32524 10722 32564 10807
rect 32140 10648 32372 10688
rect 32140 10184 32180 10648
rect 32715 10604 32757 10613
rect 32715 10564 32716 10604
rect 32756 10564 32757 10604
rect 32715 10555 32757 10564
rect 32716 10436 32756 10555
rect 32812 10445 32852 10900
rect 33004 10940 33044 10951
rect 33004 10865 33044 10900
rect 32908 10856 32948 10865
rect 32716 10387 32756 10396
rect 32811 10436 32853 10445
rect 32811 10396 32812 10436
rect 32852 10396 32853 10436
rect 32811 10387 32853 10396
rect 32331 10352 32373 10361
rect 32331 10312 32332 10352
rect 32372 10312 32373 10352
rect 32331 10303 32373 10312
rect 32140 10135 32180 10144
rect 32235 10184 32277 10193
rect 32235 10144 32236 10184
rect 32276 10144 32277 10184
rect 32235 10135 32277 10144
rect 32332 10184 32372 10303
rect 32811 10268 32853 10277
rect 32811 10228 32812 10268
rect 32852 10228 32853 10268
rect 32811 10219 32853 10228
rect 32332 10135 32372 10144
rect 32428 10184 32468 10193
rect 32620 10184 32660 10195
rect 32468 10144 32564 10184
rect 32428 10135 32468 10144
rect 32236 10050 32276 10135
rect 32140 9680 32180 9689
rect 32044 9640 32140 9680
rect 32140 9631 32180 9640
rect 32331 9596 32373 9605
rect 32331 9556 32332 9596
rect 32372 9556 32373 9596
rect 32331 9547 32373 9556
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 31948 9512 31988 9521
rect 31852 9378 31892 9463
rect 31660 9220 31713 9260
rect 31673 9176 31713 9220
rect 31673 9136 31796 9176
rect 31563 8840 31605 8849
rect 31563 8800 31564 8840
rect 31604 8800 31605 8840
rect 31756 8840 31796 9136
rect 31948 9017 31988 9472
rect 32044 9512 32084 9521
rect 31947 9008 31989 9017
rect 31947 8968 31948 9008
rect 31988 8968 31989 9008
rect 31947 8959 31989 8968
rect 32044 8924 32084 9472
rect 32140 8924 32180 8933
rect 32044 8884 32140 8924
rect 32140 8875 32180 8884
rect 31756 8800 32084 8840
rect 31563 8791 31605 8800
rect 31660 8681 31700 8766
rect 31084 8672 31124 8681
rect 30988 8632 31084 8672
rect 30891 7916 30933 7925
rect 30891 7876 30892 7916
rect 30932 7876 30933 7916
rect 30891 7867 30933 7876
rect 30795 7664 30837 7673
rect 30795 7624 30796 7664
rect 30836 7624 30837 7664
rect 30795 7615 30837 7624
rect 30603 7580 30645 7589
rect 30603 7540 30604 7580
rect 30644 7540 30645 7580
rect 30603 7531 30645 7540
rect 30796 5648 30836 7615
rect 30892 7169 30932 7867
rect 30988 7673 31028 8632
rect 31084 8623 31124 8632
rect 31372 8672 31412 8681
rect 31083 8504 31125 8513
rect 31083 8464 31084 8504
rect 31124 8464 31125 8504
rect 31083 8455 31125 8464
rect 31180 8504 31220 8513
rect 31084 8000 31124 8455
rect 31180 8093 31220 8464
rect 31179 8084 31221 8093
rect 31372 8084 31412 8632
rect 31468 8672 31508 8681
rect 31659 8672 31701 8681
rect 31508 8632 31604 8672
rect 31468 8623 31508 8632
rect 31467 8504 31509 8513
rect 31467 8464 31468 8504
rect 31508 8464 31509 8504
rect 31564 8504 31604 8632
rect 31659 8632 31660 8672
rect 31700 8632 31701 8672
rect 31659 8623 31701 8632
rect 31852 8672 31892 8681
rect 31659 8504 31701 8513
rect 31564 8464 31660 8504
rect 31700 8464 31701 8504
rect 31467 8455 31509 8464
rect 31659 8455 31701 8464
rect 31179 8044 31180 8084
rect 31220 8044 31221 8084
rect 31179 8035 31221 8044
rect 31276 8044 31412 8084
rect 30987 7664 31029 7673
rect 30987 7624 30988 7664
rect 31028 7624 31029 7664
rect 30987 7615 31029 7624
rect 31084 7412 31124 7960
rect 31179 7916 31221 7925
rect 31179 7876 31180 7916
rect 31220 7876 31221 7916
rect 31179 7867 31221 7876
rect 31180 7782 31220 7867
rect 31276 7832 31316 8044
rect 31468 8009 31508 8455
rect 31852 8429 31892 8632
rect 31947 8672 31989 8681
rect 31947 8632 31948 8672
rect 31988 8632 31989 8672
rect 31947 8623 31989 8632
rect 31948 8538 31988 8623
rect 31851 8420 31893 8429
rect 31851 8380 31852 8420
rect 31892 8380 31893 8420
rect 31851 8371 31893 8380
rect 31851 8252 31893 8261
rect 31851 8212 31852 8252
rect 31892 8212 31893 8252
rect 31851 8203 31893 8212
rect 31852 8084 31892 8203
rect 31852 8035 31892 8044
rect 31467 8000 31509 8009
rect 31467 7960 31468 8000
rect 31508 7960 31509 8000
rect 31467 7951 31509 7960
rect 31756 8000 31796 8009
rect 31371 7916 31413 7925
rect 31371 7876 31372 7916
rect 31412 7876 31413 7916
rect 31371 7867 31413 7876
rect 31276 7783 31316 7792
rect 31372 7782 31412 7867
rect 31468 7866 31508 7951
rect 31659 7832 31701 7841
rect 31659 7792 31660 7832
rect 31700 7792 31701 7832
rect 31659 7783 31701 7792
rect 31563 7748 31605 7757
rect 31563 7708 31564 7748
rect 31604 7708 31605 7748
rect 31563 7699 31605 7708
rect 31180 7412 31220 7421
rect 31084 7372 31180 7412
rect 31180 7363 31220 7372
rect 31275 7412 31317 7421
rect 31275 7372 31276 7412
rect 31316 7372 31317 7412
rect 31275 7363 31317 7372
rect 31564 7412 31604 7699
rect 31564 7363 31604 7372
rect 30891 7160 30933 7169
rect 30891 7120 30892 7160
rect 30932 7120 30933 7160
rect 30891 7111 30933 7120
rect 31276 7160 31316 7363
rect 31660 7253 31700 7783
rect 31756 7757 31796 7960
rect 31947 8000 31989 8009
rect 31947 7960 31948 8000
rect 31988 7960 31989 8000
rect 31947 7951 31989 7960
rect 31948 7866 31988 7951
rect 31755 7748 31797 7757
rect 31755 7708 31756 7748
rect 31796 7708 31797 7748
rect 31755 7699 31797 7708
rect 31947 7748 31989 7757
rect 31947 7708 31948 7748
rect 31988 7708 31989 7748
rect 31947 7699 31989 7708
rect 31755 7580 31797 7589
rect 31755 7540 31756 7580
rect 31796 7540 31797 7580
rect 31755 7531 31797 7540
rect 31659 7244 31701 7253
rect 31659 7204 31660 7244
rect 31700 7204 31701 7244
rect 31659 7195 31701 7204
rect 31276 7111 31316 7120
rect 31660 7160 31700 7195
rect 31660 7109 31700 7120
rect 30892 6488 30932 6497
rect 31084 6488 31124 6497
rect 30932 6448 31084 6488
rect 30892 6439 30932 6448
rect 31084 6439 31124 6448
rect 31468 6488 31508 6497
rect 31563 6488 31605 6497
rect 31508 6448 31564 6488
rect 31604 6448 31605 6488
rect 31468 6439 31508 6448
rect 31563 6439 31605 6448
rect 31083 5900 31125 5909
rect 31083 5860 31084 5900
rect 31124 5860 31125 5900
rect 31083 5851 31125 5860
rect 31084 5766 31124 5851
rect 30891 5648 30933 5657
rect 30796 5608 30892 5648
rect 30932 5608 30933 5648
rect 30891 5599 30933 5608
rect 31563 5648 31605 5657
rect 31563 5608 31564 5648
rect 31604 5608 31605 5648
rect 31563 5599 31605 5608
rect 31756 5648 31796 7531
rect 31852 6992 31892 7001
rect 31852 6581 31892 6952
rect 31851 6572 31893 6581
rect 31851 6532 31852 6572
rect 31892 6532 31893 6572
rect 31851 6523 31893 6532
rect 31756 5599 31796 5608
rect 30892 5514 30932 5599
rect 30219 4892 30261 4901
rect 30219 4852 30220 4892
rect 30260 4852 30261 4892
rect 30219 4843 30261 4852
rect 29932 4136 29972 4145
rect 30124 4136 30164 4145
rect 29972 4096 30124 4136
rect 29932 4087 29972 4096
rect 30124 4087 30164 4096
rect 29355 3044 29397 3053
rect 29355 3004 29356 3044
rect 29396 3004 29397 3044
rect 29355 2995 29397 3004
rect 29835 3044 29877 3053
rect 29835 3004 29836 3044
rect 29876 3004 29877 3044
rect 29835 2995 29877 3004
rect 27723 2036 27765 2045
rect 27723 1996 27724 2036
rect 27764 1996 27765 2036
rect 27723 1987 27765 1996
rect 28684 1961 28724 2584
rect 28779 2624 28821 2633
rect 28779 2584 28780 2624
rect 28820 2584 28821 2624
rect 28779 2575 28821 2584
rect 27531 1952 27573 1961
rect 27531 1912 27532 1952
rect 27572 1912 27573 1952
rect 27531 1903 27573 1912
rect 28683 1952 28725 1961
rect 28683 1912 28684 1952
rect 28724 1912 28725 1952
rect 28683 1903 28725 1912
rect 28780 1952 28820 2575
rect 29356 2120 29396 2995
rect 29451 2876 29493 2885
rect 29451 2836 29452 2876
rect 29492 2836 29493 2876
rect 29451 2827 29493 2836
rect 29835 2876 29877 2885
rect 29835 2836 29836 2876
rect 29876 2836 29877 2876
rect 29835 2827 29877 2836
rect 30220 2876 30260 4843
rect 30412 3473 30452 4936
rect 31564 4976 31604 5599
rect 31564 4927 31604 4936
rect 30507 4136 30549 4145
rect 30507 4096 30508 4136
rect 30548 4096 30549 4136
rect 30507 4087 30549 4096
rect 31371 4136 31413 4145
rect 31371 4096 31372 4136
rect 31412 4096 31413 4136
rect 31371 4087 31413 4096
rect 30508 4002 30548 4087
rect 31372 4002 31412 4087
rect 30411 3464 30453 3473
rect 30604 3464 30644 3473
rect 30411 3424 30412 3464
rect 30452 3424 30604 3464
rect 30411 3415 30453 3424
rect 30604 3415 30644 3424
rect 31852 3464 31892 3473
rect 31948 3464 31988 7699
rect 32044 7337 32084 8800
rect 32140 8672 32180 8681
rect 32332 8672 32372 9547
rect 32524 8840 32564 10144
rect 32620 10109 32660 10144
rect 32812 10184 32852 10219
rect 32908 10193 32948 10816
rect 33003 10856 33045 10865
rect 33003 10816 33004 10856
rect 33044 10816 33045 10856
rect 33003 10807 33045 10816
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 33195 10352 33237 10361
rect 33195 10312 33196 10352
rect 33236 10312 33237 10352
rect 33195 10303 33237 10312
rect 32812 10133 32852 10144
rect 32907 10184 32949 10193
rect 32907 10144 32908 10184
rect 32948 10144 32949 10184
rect 32907 10135 32949 10144
rect 33099 10184 33141 10193
rect 33099 10144 33100 10184
rect 33140 10144 33141 10184
rect 33099 10135 33141 10144
rect 32619 10100 32661 10109
rect 32619 10060 32620 10100
rect 32660 10060 32661 10100
rect 32619 10051 32661 10060
rect 33003 10100 33045 10109
rect 33003 10060 33004 10100
rect 33044 10060 33045 10100
rect 33003 10051 33045 10060
rect 33004 9966 33044 10051
rect 33100 10050 33140 10135
rect 33196 9680 33236 10303
rect 33196 9631 33236 9640
rect 33003 9596 33045 9605
rect 33003 9556 33004 9596
rect 33044 9556 33045 9596
rect 33003 9547 33045 9556
rect 32619 9512 32661 9521
rect 32619 9472 32620 9512
rect 32660 9472 32661 9512
rect 32619 9463 32661 9472
rect 32908 9512 32948 9521
rect 32620 9185 32660 9463
rect 32716 9260 32756 9269
rect 32908 9260 32948 9472
rect 33004 9512 33044 9547
rect 33004 9461 33044 9472
rect 33099 9512 33141 9521
rect 33099 9472 33100 9512
rect 33140 9472 33141 9512
rect 33099 9463 33141 9472
rect 33100 9378 33140 9463
rect 32756 9220 32948 9260
rect 32619 9176 32661 9185
rect 32619 9136 32620 9176
rect 32660 9136 32661 9176
rect 32619 9127 32661 9136
rect 32524 8791 32564 8800
rect 32427 8756 32469 8765
rect 32427 8716 32428 8756
rect 32468 8716 32469 8756
rect 32427 8707 32469 8716
rect 32620 8756 32660 8765
rect 32180 8632 32276 8672
rect 32140 8623 32180 8632
rect 32139 8504 32181 8513
rect 32139 8464 32140 8504
rect 32180 8464 32181 8504
rect 32139 8455 32181 8464
rect 32140 8168 32180 8455
rect 32236 8252 32276 8632
rect 32332 8623 32372 8632
rect 32428 8622 32468 8707
rect 32620 8345 32660 8716
rect 32716 8681 32756 9220
rect 33003 9176 33045 9185
rect 33003 9136 33004 9176
rect 33044 9136 33045 9176
rect 33003 9127 33045 9136
rect 32715 8672 32757 8681
rect 32908 8672 32948 8681
rect 32715 8632 32716 8672
rect 32756 8632 32757 8672
rect 32715 8623 32757 8632
rect 32812 8632 32908 8672
rect 32716 8538 32756 8623
rect 32812 8429 32852 8632
rect 32908 8623 32948 8632
rect 33004 8672 33044 9127
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 33483 8840 33525 8849
rect 33483 8800 33484 8840
rect 33524 8800 33525 8840
rect 33483 8791 33525 8800
rect 33004 8623 33044 8632
rect 33484 8672 33524 8791
rect 33195 8588 33237 8597
rect 33195 8548 33196 8588
rect 33236 8548 33237 8588
rect 33195 8539 33237 8548
rect 32907 8504 32949 8513
rect 32907 8464 32908 8504
rect 32948 8464 32949 8504
rect 32907 8455 32949 8464
rect 33099 8504 33141 8513
rect 33099 8464 33100 8504
rect 33140 8464 33141 8504
rect 33099 8455 33141 8464
rect 33196 8504 33236 8539
rect 33484 8513 33524 8632
rect 33675 8672 33717 8681
rect 33675 8629 33676 8672
rect 33716 8629 33717 8672
rect 33675 8623 33717 8629
rect 32811 8420 32853 8429
rect 32811 8380 32812 8420
rect 32852 8380 32853 8420
rect 32811 8371 32853 8380
rect 32619 8336 32661 8345
rect 32619 8296 32620 8336
rect 32660 8296 32661 8336
rect 32619 8287 32661 8296
rect 32236 8212 32564 8252
rect 32524 8168 32564 8212
rect 32716 8168 32756 8177
rect 32524 8128 32716 8168
rect 32140 7925 32180 8128
rect 32716 8119 32756 8128
rect 32428 8009 32468 8094
rect 32332 8000 32372 8009
rect 32139 7916 32181 7925
rect 32139 7876 32140 7916
rect 32180 7876 32181 7916
rect 32139 7867 32181 7876
rect 32332 7832 32372 7960
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 32620 8000 32660 8011
rect 32620 7925 32660 7960
rect 32619 7916 32661 7925
rect 32619 7876 32620 7916
rect 32660 7876 32661 7916
rect 32619 7867 32661 7876
rect 32332 7792 32375 7832
rect 32335 7748 32375 7792
rect 32332 7708 32375 7748
rect 32332 7421 32372 7708
rect 32812 7589 32852 8371
rect 32908 8000 32948 8455
rect 32908 7951 32948 7960
rect 32619 7580 32661 7589
rect 32619 7540 32620 7580
rect 32660 7540 32661 7580
rect 32619 7531 32661 7540
rect 32811 7580 32853 7589
rect 32811 7540 32812 7580
rect 32852 7540 32853 7580
rect 32811 7531 32853 7540
rect 32331 7412 32373 7421
rect 32331 7372 32332 7412
rect 32372 7372 32373 7412
rect 32331 7363 32373 7372
rect 32523 7412 32565 7421
rect 32523 7372 32524 7412
rect 32564 7372 32565 7412
rect 32523 7363 32565 7372
rect 32043 7328 32085 7337
rect 32043 7288 32044 7328
rect 32084 7288 32085 7328
rect 32043 7279 32085 7288
rect 32044 6497 32084 7279
rect 32331 7160 32373 7169
rect 32331 7120 32332 7160
rect 32372 7120 32373 7160
rect 32331 7111 32373 7120
rect 32524 7160 32564 7363
rect 32524 7111 32564 7120
rect 32043 6488 32085 6497
rect 32043 6448 32044 6488
rect 32084 6448 32085 6488
rect 32043 6439 32085 6448
rect 32332 6488 32372 7111
rect 32332 4145 32372 6448
rect 32331 4136 32373 4145
rect 32331 4096 32332 4136
rect 32372 4096 32373 4136
rect 32331 4087 32373 4096
rect 32620 4136 32660 7531
rect 33100 6917 33140 8455
rect 33196 8453 33236 8464
rect 33483 8504 33525 8513
rect 33483 8464 33484 8504
rect 33524 8464 33525 8504
rect 33483 8455 33525 8464
rect 33291 8252 33333 8261
rect 33291 8212 33292 8252
rect 33332 8212 33333 8252
rect 33291 8203 33333 8212
rect 33292 8000 33332 8203
rect 33676 8084 33716 8623
rect 33580 8044 33716 8084
rect 33292 7951 33332 7960
rect 33483 8000 33525 8009
rect 33483 7960 33484 8000
rect 33524 7960 33525 8000
rect 33483 7951 33525 7960
rect 33580 8000 33620 8044
rect 33580 7951 33620 7960
rect 33484 7866 33524 7951
rect 33676 7757 33716 8044
rect 33771 8084 33813 8093
rect 33771 8044 33772 8084
rect 33812 8044 33813 8084
rect 33771 8035 33813 8044
rect 33772 8000 33812 8035
rect 33772 7949 33812 7960
rect 33771 7832 33813 7841
rect 33771 7792 33772 7832
rect 33812 7792 33813 7832
rect 33771 7783 33813 7792
rect 33196 7748 33236 7757
rect 33099 6908 33141 6917
rect 33099 6868 33100 6908
rect 33140 6868 33141 6908
rect 33099 6859 33141 6868
rect 33196 5657 33236 7708
rect 33675 7748 33717 7757
rect 33675 7708 33676 7748
rect 33716 7708 33717 7748
rect 33675 7699 33717 7708
rect 33772 7698 33812 7783
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 33483 7412 33525 7421
rect 33483 7372 33484 7412
rect 33524 7372 33525 7412
rect 33483 7363 33525 7372
rect 33771 7412 33813 7421
rect 33771 7372 33772 7412
rect 33812 7372 33813 7412
rect 33771 7363 33813 7372
rect 33484 6488 33524 7363
rect 33772 7278 33812 7363
rect 33868 7169 33908 12244
rect 33964 11957 34004 12412
rect 33963 11948 34005 11957
rect 33963 11908 33964 11948
rect 34004 11908 34005 11948
rect 33963 11899 34005 11908
rect 33964 11814 34004 11899
rect 33964 11696 34004 11705
rect 34060 11696 34100 12739
rect 34004 11656 34100 11696
rect 33964 11647 34004 11656
rect 34156 11360 34196 13000
rect 34444 12536 34484 13159
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 34539 12704 34581 12713
rect 34539 12664 34540 12704
rect 34580 12664 34581 12704
rect 34539 12655 34581 12664
rect 34732 12704 34772 12713
rect 34444 12487 34484 12496
rect 34540 12536 34580 12655
rect 34540 12487 34580 12496
rect 34732 11873 34772 12664
rect 35020 12629 35060 13168
rect 35596 12664 35828 12704
rect 35019 12620 35061 12629
rect 35019 12580 35020 12620
rect 35060 12580 35061 12620
rect 35019 12571 35061 12580
rect 35500 12620 35540 12629
rect 35596 12620 35636 12664
rect 35540 12580 35636 12620
rect 35500 12571 35540 12580
rect 35404 12536 35444 12545
rect 35404 11948 35444 12496
rect 35692 12536 35732 12545
rect 35404 11908 35540 11948
rect 34731 11864 34773 11873
rect 34731 11824 34732 11864
rect 34772 11824 34773 11864
rect 34731 11815 34773 11824
rect 35019 11864 35061 11873
rect 35019 11824 35020 11864
rect 35060 11824 35061 11864
rect 35019 11815 35061 11824
rect 34924 11780 34964 11789
rect 34251 11696 34293 11705
rect 34828 11696 34868 11705
rect 34251 11656 34252 11696
rect 34292 11656 34293 11696
rect 34251 11647 34293 11656
rect 34444 11656 34828 11696
rect 34252 11562 34292 11647
rect 34060 11320 34196 11360
rect 33963 9428 34005 9437
rect 33963 9388 33964 9428
rect 34004 9388 34005 9428
rect 33963 9379 34005 9388
rect 33964 8840 34004 9379
rect 34060 9101 34100 11320
rect 34347 11276 34389 11285
rect 34347 11236 34348 11276
rect 34388 11236 34389 11276
rect 34347 11227 34389 11236
rect 34348 11024 34388 11227
rect 34444 11192 34484 11656
rect 34828 11647 34868 11656
rect 34924 11528 34964 11740
rect 35020 11730 35060 11815
rect 35116 11782 35300 11822
rect 35116 11780 35156 11782
rect 35260 11780 35300 11782
rect 35260 11740 35348 11780
rect 35116 11731 35156 11740
rect 35212 11654 35252 11663
rect 34924 11488 35060 11528
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 35020 11192 35060 11488
rect 34444 11143 34484 11152
rect 34636 11152 35060 11192
rect 34388 10984 34484 11024
rect 34348 10975 34388 10984
rect 34347 10436 34389 10445
rect 34347 10396 34348 10436
rect 34388 10396 34389 10436
rect 34347 10387 34389 10396
rect 34348 10277 34388 10387
rect 34347 10268 34389 10277
rect 34347 10228 34348 10268
rect 34388 10228 34389 10268
rect 34347 10219 34389 10228
rect 34348 10016 34388 10219
rect 34444 10184 34484 10984
rect 34636 10436 34676 11152
rect 34731 11024 34773 11033
rect 34731 10984 34732 11024
rect 34772 10984 34773 11024
rect 34731 10975 34773 10984
rect 34828 11024 34868 11033
rect 34732 10890 34772 10975
rect 34828 10865 34868 10984
rect 34924 11024 34964 11033
rect 34827 10856 34869 10865
rect 34827 10816 34828 10856
rect 34868 10816 34869 10856
rect 34827 10807 34869 10816
rect 34636 10387 34676 10396
rect 34828 10184 34868 10193
rect 34444 10135 34484 10144
rect 34636 10144 34828 10184
rect 34924 10184 34964 10984
rect 35020 11024 35060 11152
rect 35060 10984 35156 11024
rect 35020 10975 35060 10984
rect 35020 10445 35060 10530
rect 35019 10436 35061 10445
rect 35019 10396 35020 10436
rect 35060 10396 35061 10436
rect 35019 10387 35061 10396
rect 35020 10184 35060 10193
rect 34924 10144 35020 10184
rect 34636 10016 34676 10144
rect 34828 10135 34868 10144
rect 35020 10025 35060 10144
rect 35116 10184 35156 10984
rect 35212 10940 35252 11614
rect 35308 11117 35348 11740
rect 35404 11528 35444 11537
rect 35404 11369 35444 11488
rect 35403 11360 35445 11369
rect 35403 11320 35404 11360
rect 35444 11320 35445 11360
rect 35403 11311 35445 11320
rect 35403 11192 35445 11201
rect 35403 11152 35404 11192
rect 35444 11152 35445 11192
rect 35403 11143 35445 11152
rect 35307 11108 35349 11117
rect 35307 11068 35308 11108
rect 35348 11068 35349 11108
rect 35307 11059 35349 11068
rect 35404 11024 35444 11143
rect 35500 11033 35540 11908
rect 35404 10975 35444 10984
rect 35499 11024 35541 11033
rect 35499 10984 35500 11024
rect 35540 10984 35541 11024
rect 35499 10975 35541 10984
rect 35212 10900 35348 10940
rect 35211 10772 35253 10781
rect 35211 10732 35212 10772
rect 35252 10732 35253 10772
rect 35211 10723 35253 10732
rect 35212 10638 35252 10723
rect 35308 10436 35348 10900
rect 35499 10856 35541 10865
rect 35499 10816 35500 10856
rect 35540 10816 35541 10856
rect 35499 10807 35541 10816
rect 35308 10387 35348 10396
rect 35307 10268 35349 10277
rect 35307 10228 35308 10268
rect 35348 10228 35349 10268
rect 35307 10219 35349 10228
rect 35116 10135 35156 10144
rect 35308 10184 35348 10219
rect 35308 10133 35348 10144
rect 35500 10184 35540 10807
rect 35692 10445 35732 12496
rect 35788 12536 35828 12664
rect 36267 12620 36309 12629
rect 36267 12580 36268 12620
rect 36308 12580 36309 12620
rect 36267 12571 36309 12580
rect 35980 12536 36020 12545
rect 35788 12487 35828 12496
rect 35884 12496 35980 12536
rect 36020 12496 36212 12536
rect 35787 11360 35829 11369
rect 35787 11320 35788 11360
rect 35828 11320 35829 11360
rect 35787 11311 35829 11320
rect 35788 11024 35828 11311
rect 35788 10975 35828 10984
rect 35884 10781 35924 12496
rect 35980 12487 36020 12496
rect 36172 12368 36212 12496
rect 36268 12486 36308 12571
rect 36364 12536 36404 12545
rect 36364 12368 36404 12496
rect 36748 12536 36788 13747
rect 36940 13208 36980 13217
rect 37228 13208 37268 14848
rect 37323 14720 37365 14729
rect 37323 14680 37324 14720
rect 37364 14680 37365 14720
rect 37323 14671 37365 14680
rect 37420 14720 37460 14729
rect 37516 14720 37556 15175
rect 37612 14804 37652 15343
rect 37899 15224 37941 15233
rect 37899 15184 37900 15224
rect 37940 15184 37941 15224
rect 37899 15175 37941 15184
rect 37612 14729 37652 14764
rect 37460 14680 37556 14720
rect 37611 14720 37653 14729
rect 37611 14680 37612 14720
rect 37652 14680 37653 14720
rect 37420 14671 37460 14680
rect 37611 14671 37653 14680
rect 37900 14720 37940 15175
rect 38092 15149 38132 15520
rect 38188 15560 38228 15595
rect 38188 15509 38228 15520
rect 38091 15140 38133 15149
rect 38091 15100 38092 15140
rect 38132 15100 38133 15140
rect 38091 15091 38133 15100
rect 37900 14671 37940 14680
rect 37996 14720 38036 14729
rect 38092 14720 38132 15091
rect 38036 14680 38132 14720
rect 38187 14720 38229 14729
rect 38284 14720 38324 16612
rect 38380 16409 38420 17032
rect 38476 17072 38516 17081
rect 38476 16829 38516 17032
rect 39052 16988 39092 17704
rect 39148 17695 39188 17704
rect 39148 17240 39188 17249
rect 39244 17240 39284 18544
rect 39435 17828 39477 17837
rect 39435 17788 39436 17828
rect 39476 17788 39477 17828
rect 39435 17779 39477 17788
rect 39188 17200 39284 17240
rect 39148 17191 39188 17200
rect 39052 16948 39380 16988
rect 38475 16820 38517 16829
rect 39148 16820 39188 16829
rect 38475 16780 38476 16820
rect 38516 16780 38517 16820
rect 38475 16771 38517 16780
rect 39052 16780 39148 16820
rect 38379 16400 38421 16409
rect 38379 16360 38380 16400
rect 38420 16360 38421 16400
rect 38379 16351 38421 16360
rect 38476 16400 38516 16409
rect 38516 16360 38804 16400
rect 38476 16351 38516 16360
rect 38571 16232 38613 16241
rect 38571 16192 38572 16232
rect 38612 16192 38613 16232
rect 38571 16183 38613 16192
rect 38379 15980 38421 15989
rect 38379 15940 38380 15980
rect 38420 15940 38421 15980
rect 38379 15931 38421 15940
rect 38380 15317 38420 15931
rect 38379 15308 38421 15317
rect 38379 15268 38380 15308
rect 38420 15268 38421 15308
rect 38379 15259 38421 15268
rect 38380 15174 38420 15259
rect 38187 14680 38188 14720
rect 38228 14680 38324 14720
rect 37996 14671 38036 14680
rect 38187 14671 38229 14680
rect 37324 14586 37364 14671
rect 37612 14640 37652 14671
rect 37803 14048 37845 14057
rect 37803 14008 37804 14048
rect 37844 14008 37845 14048
rect 37803 13999 37845 14008
rect 37804 13914 37844 13999
rect 38091 13796 38133 13805
rect 38091 13756 38092 13796
rect 38132 13756 38133 13796
rect 38091 13747 38133 13756
rect 38092 13662 38132 13747
rect 37324 13208 37364 13217
rect 37228 13168 37324 13208
rect 36940 12704 36980 13168
rect 37324 13159 37364 13168
rect 38188 13208 38228 14671
rect 38572 14552 38612 16183
rect 38667 15896 38709 15905
rect 38667 15856 38668 15896
rect 38708 15856 38709 15896
rect 38667 15847 38709 15856
rect 38668 15728 38708 15847
rect 38668 15679 38708 15688
rect 38667 15560 38709 15569
rect 38667 15520 38668 15560
rect 38708 15520 38709 15560
rect 38667 15511 38709 15520
rect 38668 15426 38708 15511
rect 38764 15392 38804 16360
rect 38956 16241 38996 16326
rect 38955 16232 38997 16241
rect 38955 16192 38956 16232
rect 38996 16192 38997 16232
rect 38955 16183 38997 16192
rect 38956 16064 38996 16073
rect 38860 16024 38956 16064
rect 38860 15560 38900 16024
rect 38956 16015 38996 16024
rect 38860 15511 38900 15520
rect 38956 15560 38996 15569
rect 38956 15392 38996 15520
rect 38764 15352 38996 15392
rect 38667 15140 38709 15149
rect 38667 15100 38668 15140
rect 38708 15100 38709 15140
rect 38667 15091 38709 15100
rect 38859 15140 38901 15149
rect 38859 15100 38860 15140
rect 38900 15100 38901 15140
rect 38859 15091 38901 15100
rect 38668 14720 38708 15091
rect 38668 14671 38708 14680
rect 38860 14720 38900 15091
rect 38860 14671 38900 14680
rect 38764 14636 38804 14645
rect 38764 14552 38804 14596
rect 38572 14512 38804 14552
rect 38956 14216 38996 14225
rect 38764 14048 38804 14059
rect 38764 13973 38804 14008
rect 38763 13964 38805 13973
rect 38763 13924 38764 13964
rect 38804 13924 38805 13964
rect 38763 13915 38805 13924
rect 38188 13159 38228 13168
rect 38956 12713 38996 14176
rect 36940 12655 36980 12664
rect 38955 12704 38997 12713
rect 38955 12664 38956 12704
rect 38996 12664 38997 12704
rect 38955 12655 38997 12664
rect 37611 12620 37653 12629
rect 37611 12580 37612 12620
rect 37652 12580 37653 12620
rect 37611 12571 37653 12580
rect 36748 12487 36788 12496
rect 37612 12536 37652 12571
rect 37612 12485 37652 12496
rect 39052 12536 39092 16780
rect 39148 16771 39188 16780
rect 39148 16232 39188 16241
rect 39148 16073 39188 16192
rect 39244 16232 39284 16241
rect 39147 16064 39189 16073
rect 39147 16024 39148 16064
rect 39188 16024 39189 16064
rect 39147 16015 39189 16024
rect 39244 15989 39284 16192
rect 39243 15980 39285 15989
rect 39243 15940 39244 15980
rect 39284 15940 39285 15980
rect 39243 15931 39285 15940
rect 39148 15392 39188 15401
rect 39340 15392 39380 16948
rect 39436 16400 39476 17779
rect 39627 17072 39669 17081
rect 39627 17032 39628 17072
rect 39668 17032 39669 17072
rect 39627 17023 39669 17032
rect 39628 16938 39668 17023
rect 39436 16351 39476 16360
rect 39724 15896 39764 19207
rect 40684 19122 40724 19207
rect 40011 19088 40053 19097
rect 40011 19048 40012 19088
rect 40052 19048 40053 19088
rect 40011 19039 40053 19048
rect 40012 18954 40052 19039
rect 40492 18584 40532 18593
rect 39916 18332 39956 18341
rect 39956 18292 40052 18332
rect 39916 18283 39956 18292
rect 40012 17753 40052 18292
rect 40011 17744 40053 17753
rect 40011 17704 40012 17744
rect 40052 17704 40053 17744
rect 40011 17695 40053 17704
rect 39915 17660 39957 17669
rect 39915 17620 39916 17660
rect 39956 17620 39957 17660
rect 39915 17611 39957 17620
rect 39916 17072 39956 17611
rect 40012 17610 40052 17695
rect 40492 17081 40532 18544
rect 41452 18584 41492 21391
rect 41560 20852 41600 21400
rect 41644 21029 41684 21568
rect 41740 21608 41780 21617
rect 41836 21608 41876 22240
rect 42027 22280 42069 22289
rect 42027 22240 42028 22280
rect 42068 22240 42069 22280
rect 42027 22231 42069 22240
rect 42124 22280 42164 22483
rect 42124 22231 42164 22240
rect 42316 22280 42356 22651
rect 42316 22231 42356 22240
rect 42700 22280 42740 22735
rect 42892 22709 42932 22828
rect 43179 22868 43221 22877
rect 43179 22828 43180 22868
rect 43220 22828 43221 22868
rect 43179 22819 43221 22828
rect 42891 22700 42933 22709
rect 42891 22660 42892 22700
rect 42932 22660 42933 22700
rect 42891 22651 42933 22660
rect 42700 22231 42740 22240
rect 43564 22280 43604 23071
rect 43756 22961 43796 23080
rect 44428 23045 44468 24592
rect 44524 24632 44564 24751
rect 44812 24632 44852 25003
rect 44907 24968 44949 24977
rect 44907 24928 44908 24968
rect 44948 24928 44949 24968
rect 44907 24919 44949 24928
rect 44908 24641 44948 24919
rect 45100 24809 45140 25339
rect 45196 25304 45236 25313
rect 45292 25304 45332 25936
rect 45388 25565 45428 27355
rect 45387 25556 45429 25565
rect 45387 25516 45388 25556
rect 45428 25516 45429 25556
rect 45387 25507 45429 25516
rect 45236 25264 45332 25304
rect 45196 25255 45236 25264
rect 45099 24800 45141 24809
rect 45099 24760 45100 24800
rect 45140 24760 45141 24800
rect 45099 24751 45141 24760
rect 45484 24800 45524 27775
rect 45580 27581 45620 28288
rect 45579 27572 45621 27581
rect 45579 27532 45580 27572
rect 45620 27532 45621 27572
rect 45579 27523 45621 27532
rect 45579 27404 45621 27413
rect 45579 27364 45580 27404
rect 45620 27364 45621 27404
rect 45579 27355 45621 27364
rect 45580 26816 45620 27355
rect 45580 26767 45620 26776
rect 45676 26312 45716 26323
rect 45676 26237 45716 26272
rect 45675 26228 45717 26237
rect 45675 26188 45676 26228
rect 45716 26188 45717 26228
rect 45675 26179 45717 26188
rect 45675 25724 45717 25733
rect 45675 25684 45676 25724
rect 45716 25684 45717 25724
rect 45675 25675 45717 25684
rect 45676 24893 45716 25675
rect 45772 25313 45812 28876
rect 45868 26648 45908 28960
rect 46444 28328 46484 28337
rect 46251 28160 46293 28169
rect 46251 28120 46252 28160
rect 46292 28120 46293 28160
rect 46251 28111 46293 28120
rect 46155 27908 46197 27917
rect 46155 27868 46156 27908
rect 46196 27868 46197 27908
rect 46155 27859 46197 27868
rect 45963 27656 46005 27665
rect 45963 27616 45964 27656
rect 46004 27616 46005 27656
rect 45963 27607 46005 27616
rect 46156 27656 46196 27859
rect 46156 27607 46196 27616
rect 46252 27656 46292 28111
rect 46444 27833 46484 28288
rect 46539 28328 46581 28337
rect 46539 28288 46540 28328
rect 46580 28288 46581 28328
rect 46539 28279 46581 28288
rect 46540 28194 46580 28279
rect 46636 28253 46676 28960
rect 47115 28916 47157 28925
rect 47115 28876 47116 28916
rect 47156 28876 47157 28916
rect 47115 28867 47157 28876
rect 46828 28328 46868 28339
rect 46828 28253 46868 28288
rect 47019 28328 47061 28337
rect 47019 28288 47020 28328
rect 47060 28288 47061 28328
rect 47019 28279 47061 28288
rect 47116 28328 47156 28867
rect 46635 28244 46677 28253
rect 46635 28204 46636 28244
rect 46676 28204 46677 28244
rect 46635 28195 46677 28204
rect 46827 28244 46869 28253
rect 46827 28204 46828 28244
rect 46868 28204 46869 28244
rect 46827 28195 46869 28204
rect 46636 27833 46676 28195
rect 47020 28194 47060 28279
rect 46731 28160 46773 28169
rect 46731 28120 46732 28160
rect 46772 28120 46773 28160
rect 46731 28111 46773 28120
rect 46732 28026 46772 28111
rect 47116 28076 47156 28288
rect 47020 28036 47156 28076
rect 47020 27917 47060 28036
rect 47212 27992 47252 29128
rect 47308 28580 47348 29707
rect 47596 29336 47636 30640
rect 47691 30631 47733 30640
rect 47788 30680 47828 30689
rect 47692 30546 47732 30631
rect 47788 30269 47828 30640
rect 47884 30680 47924 31219
rect 47787 30260 47829 30269
rect 47787 30220 47788 30260
rect 47828 30220 47829 30260
rect 47787 30211 47829 30220
rect 47787 30008 47829 30017
rect 47787 29968 47788 30008
rect 47828 29968 47829 30008
rect 47787 29959 47829 29968
rect 47788 29840 47828 29959
rect 47788 29791 47828 29800
rect 47596 29287 47636 29296
rect 47787 28916 47829 28925
rect 47787 28876 47788 28916
rect 47828 28876 47829 28916
rect 47787 28867 47829 28876
rect 47788 28782 47828 28867
rect 47308 28531 47348 28540
rect 47499 28496 47541 28505
rect 47499 28456 47500 28496
rect 47540 28456 47541 28496
rect 47499 28447 47541 28456
rect 47500 28362 47540 28447
rect 47884 28337 47924 30640
rect 47980 30680 48020 30689
rect 48268 30680 48308 30689
rect 48020 30640 48268 30680
rect 47980 30631 48020 30640
rect 48268 30631 48308 30640
rect 48267 30512 48309 30521
rect 48267 30472 48268 30512
rect 48308 30472 48309 30512
rect 48267 30463 48309 30472
rect 48268 30378 48308 30463
rect 48075 30260 48117 30269
rect 48075 30220 48076 30260
rect 48116 30220 48117 30260
rect 48075 30211 48117 30220
rect 48267 30260 48309 30269
rect 48267 30220 48268 30260
rect 48308 30220 48309 30260
rect 48267 30211 48309 30220
rect 48076 29345 48116 30211
rect 48171 29756 48213 29765
rect 48171 29716 48172 29756
rect 48212 29716 48213 29756
rect 48171 29707 48213 29716
rect 48172 29622 48212 29707
rect 48075 29336 48117 29345
rect 48075 29296 48076 29336
rect 48116 29296 48117 29336
rect 48075 29287 48117 29296
rect 48076 29000 48116 29287
rect 48076 28960 48212 29000
rect 47308 28328 47348 28337
rect 47308 28169 47348 28288
rect 47883 28328 47925 28337
rect 47883 28288 47884 28328
rect 47924 28288 47925 28328
rect 47883 28279 47925 28288
rect 48172 28328 48212 28960
rect 48268 28421 48308 30211
rect 48364 29849 48404 31312
rect 48556 31303 48596 31312
rect 49132 30773 49172 31900
rect 49708 31604 49748 31613
rect 49804 31604 49844 32143
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 49748 31564 49844 31604
rect 49708 31555 49748 31564
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 49131 30764 49173 30773
rect 49131 30724 49132 30764
rect 49172 30724 49173 30764
rect 49131 30715 49173 30724
rect 48459 30680 48501 30689
rect 48459 30640 48460 30680
rect 48500 30640 48501 30680
rect 48459 30631 48501 30640
rect 48556 30680 48596 30689
rect 48460 30546 48500 30631
rect 48556 30437 48596 30640
rect 48940 30680 48980 30689
rect 48940 30521 48980 30640
rect 48939 30512 48981 30521
rect 48939 30472 48940 30512
rect 48980 30472 48981 30512
rect 48939 30463 48981 30472
rect 49995 30512 50037 30521
rect 49995 30472 49996 30512
rect 50036 30472 50037 30512
rect 49995 30463 50037 30472
rect 50188 30512 50228 30521
rect 48555 30428 48597 30437
rect 48555 30388 48556 30428
rect 48596 30388 48597 30428
rect 48555 30379 48597 30388
rect 49611 30428 49653 30437
rect 49611 30388 49612 30428
rect 49652 30388 49653 30428
rect 49611 30379 49653 30388
rect 48939 30344 48981 30353
rect 48939 30304 48940 30344
rect 48980 30304 48981 30344
rect 48939 30295 48981 30304
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 48363 29840 48405 29849
rect 48363 29800 48364 29840
rect 48404 29800 48405 29840
rect 48363 29791 48405 29800
rect 48556 29840 48596 29849
rect 48940 29840 48980 30295
rect 49612 30294 49652 30379
rect 49996 30378 50036 30463
rect 50188 30353 50228 30472
rect 51243 30512 51285 30521
rect 51243 30472 51244 30512
rect 51284 30472 51285 30512
rect 51243 30463 51285 30472
rect 50187 30344 50229 30353
rect 50187 30304 50188 30344
rect 50228 30304 50229 30344
rect 50187 30295 50229 30304
rect 48596 29800 48980 29840
rect 49419 29840 49461 29849
rect 49419 29800 49420 29840
rect 49460 29800 49461 29840
rect 48556 29791 48596 29800
rect 49419 29791 49461 29800
rect 50379 29840 50421 29849
rect 50379 29800 50380 29840
rect 50420 29800 50421 29840
rect 50379 29791 50421 29800
rect 49420 29706 49460 29791
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 49227 29336 49269 29345
rect 49227 29296 49228 29336
rect 49268 29296 49269 29336
rect 49227 29287 49269 29296
rect 49228 29202 49268 29287
rect 49035 29168 49077 29177
rect 49035 29128 49036 29168
rect 49076 29128 49077 29168
rect 49035 29119 49077 29128
rect 50380 29168 50420 29791
rect 50572 29672 50612 29681
rect 50572 29177 50612 29632
rect 50380 29119 50420 29128
rect 50571 29168 50613 29177
rect 50571 29128 50572 29168
rect 50612 29128 50613 29168
rect 50571 29119 50613 29128
rect 51244 29168 51284 30463
rect 51627 30428 51669 30437
rect 51627 30388 51628 30428
rect 51668 30388 51669 30428
rect 51627 30379 51669 30388
rect 51628 29252 51668 30379
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 51628 29203 51668 29212
rect 51244 29119 51284 29128
rect 49036 29034 49076 29119
rect 48364 28916 48404 28925
rect 48364 28496 48404 28876
rect 48939 28916 48981 28925
rect 48939 28876 48940 28916
rect 48980 28876 48981 28916
rect 48939 28867 48981 28876
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 48364 28456 48884 28496
rect 48267 28412 48309 28421
rect 48267 28372 48268 28412
rect 48308 28372 48404 28412
rect 48267 28363 48309 28372
rect 48172 28279 48212 28288
rect 48364 28328 48404 28372
rect 48364 28279 48404 28288
rect 48460 28328 48500 28456
rect 48460 28279 48500 28288
rect 48747 28328 48789 28337
rect 48747 28288 48748 28328
rect 48788 28288 48789 28328
rect 48747 28279 48789 28288
rect 48844 28328 48884 28456
rect 48844 28279 48884 28288
rect 48940 28328 48980 28867
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 50860 28496 50900 28505
rect 48748 28194 48788 28279
rect 47307 28160 47349 28169
rect 47307 28120 47308 28160
rect 47348 28120 47349 28160
rect 47307 28111 47349 28120
rect 48651 28160 48693 28169
rect 48651 28120 48652 28160
rect 48692 28120 48693 28160
rect 48651 28111 48693 28120
rect 48652 28026 48692 28111
rect 47116 27952 47252 27992
rect 47019 27908 47061 27917
rect 47019 27868 47020 27908
rect 47060 27868 47061 27908
rect 47019 27859 47061 27868
rect 46443 27824 46485 27833
rect 46443 27784 46444 27824
rect 46484 27784 46485 27824
rect 46443 27775 46485 27784
rect 46635 27824 46677 27833
rect 46635 27784 46636 27824
rect 46676 27784 46677 27824
rect 46635 27775 46677 27784
rect 46252 27607 46292 27616
rect 46924 27656 46964 27665
rect 45964 27522 46004 27607
rect 46444 27488 46484 27497
rect 45963 27404 46005 27413
rect 45963 27364 45964 27404
rect 46004 27364 46005 27404
rect 45963 27355 46005 27364
rect 45964 27270 46004 27355
rect 45964 26816 46004 26825
rect 46444 26816 46484 27448
rect 46004 26776 46484 26816
rect 46827 26816 46869 26825
rect 46827 26776 46828 26816
rect 46868 26776 46869 26816
rect 45964 26767 46004 26776
rect 46827 26767 46869 26776
rect 46828 26682 46868 26767
rect 45868 26608 46004 26648
rect 45868 26060 45908 26069
rect 45868 25481 45908 26020
rect 45867 25472 45909 25481
rect 45867 25432 45868 25472
rect 45908 25432 45909 25472
rect 45867 25423 45909 25432
rect 45771 25304 45813 25313
rect 45771 25264 45772 25304
rect 45812 25264 45813 25304
rect 45964 25304 46004 26608
rect 46060 26144 46100 26153
rect 46060 25472 46100 26104
rect 46156 26144 46196 26153
rect 46348 26144 46388 26153
rect 46156 25733 46196 26104
rect 46252 26104 46348 26144
rect 46155 25724 46197 25733
rect 46155 25684 46156 25724
rect 46196 25684 46197 25724
rect 46155 25675 46197 25684
rect 46060 25432 46196 25472
rect 46060 25304 46100 25313
rect 45964 25264 46060 25304
rect 45771 25255 45813 25264
rect 46060 25255 46100 25264
rect 45771 24968 45813 24977
rect 45771 24928 45772 24968
rect 45812 24928 45813 24968
rect 45771 24919 45813 24928
rect 45675 24884 45717 24893
rect 45675 24844 45676 24884
rect 45716 24844 45717 24884
rect 45675 24835 45717 24844
rect 45484 24751 45524 24760
rect 44524 24583 44564 24592
rect 44620 24592 44812 24632
rect 44620 23960 44660 24592
rect 44812 24583 44852 24592
rect 44907 24632 44949 24641
rect 44907 24592 44908 24632
rect 44948 24592 44949 24632
rect 44907 24583 44949 24592
rect 44908 23960 44948 24583
rect 45003 24464 45045 24473
rect 45003 24424 45004 24464
rect 45044 24424 45045 24464
rect 45003 24415 45045 24424
rect 44524 23920 44660 23960
rect 44716 23920 44948 23960
rect 44139 23036 44181 23045
rect 44139 22996 44140 23036
rect 44180 22996 44181 23036
rect 44139 22987 44181 22996
rect 44427 23036 44469 23045
rect 44427 22996 44428 23036
rect 44468 22996 44469 23036
rect 44427 22987 44469 22996
rect 43755 22952 43797 22961
rect 43755 22912 43756 22952
rect 43796 22912 43797 22952
rect 43755 22903 43797 22912
rect 44140 22902 44180 22987
rect 44524 22364 44564 23920
rect 44619 23792 44661 23801
rect 44619 23752 44620 23792
rect 44660 23752 44661 23792
rect 44619 23743 44661 23752
rect 44620 23658 44660 23743
rect 44716 22532 44756 23920
rect 44907 23792 44949 23801
rect 44907 23752 44908 23792
rect 44948 23752 44949 23792
rect 44907 23743 44949 23752
rect 44811 23288 44853 23297
rect 44811 23248 44812 23288
rect 44852 23248 44853 23288
rect 44811 23239 44853 23248
rect 44812 23120 44852 23239
rect 44812 23071 44852 23080
rect 44811 22952 44853 22961
rect 44811 22912 44812 22952
rect 44852 22912 44853 22952
rect 44811 22903 44853 22912
rect 44716 22483 44756 22492
rect 44715 22364 44757 22373
rect 44524 22324 44660 22364
rect 42028 22146 42068 22231
rect 41931 22112 41973 22121
rect 41931 22072 41932 22112
rect 41972 22072 41973 22112
rect 41931 22063 41973 22072
rect 41780 21568 41876 21608
rect 41932 21608 41972 22063
rect 41740 21559 41780 21568
rect 41932 21559 41972 21568
rect 42124 21608 42164 21617
rect 41932 21440 41972 21449
rect 42124 21440 42164 21568
rect 43276 21608 43316 21617
rect 43276 21449 43316 21568
rect 41972 21400 42164 21440
rect 43275 21440 43317 21449
rect 43275 21400 43276 21440
rect 43316 21400 43317 21440
rect 41932 21391 41972 21400
rect 43275 21391 43317 21400
rect 43564 21440 43604 22240
rect 44523 21692 44565 21701
rect 44523 21652 44524 21692
rect 44564 21652 44565 21692
rect 44523 21643 44565 21652
rect 44427 21608 44469 21617
rect 44427 21568 44428 21608
rect 44468 21568 44469 21608
rect 44427 21559 44469 21568
rect 44524 21608 44564 21643
rect 44428 21474 44468 21559
rect 44524 21557 44564 21568
rect 42796 21356 42836 21365
rect 42220 21316 42796 21356
rect 41643 21020 41685 21029
rect 41643 20980 41644 21020
rect 41684 20980 41685 21020
rect 41643 20971 41685 20980
rect 41644 20852 41684 20861
rect 41560 20812 41644 20852
rect 41644 20803 41684 20812
rect 42220 20768 42260 21316
rect 42796 21307 42836 21316
rect 42220 20719 42260 20728
rect 42604 20768 42644 20777
rect 42604 20180 42644 20728
rect 43468 20768 43508 20777
rect 43564 20768 43604 21400
rect 44620 21020 44660 22324
rect 44715 22324 44716 22364
rect 44756 22324 44757 22364
rect 44715 22315 44757 22324
rect 44716 21785 44756 22315
rect 44715 21776 44757 21785
rect 44715 21736 44716 21776
rect 44756 21736 44757 21776
rect 44715 21727 44757 21736
rect 44716 21608 44756 21727
rect 44716 21559 44756 21568
rect 44812 21608 44852 22903
rect 44812 21559 44852 21568
rect 44908 21608 44948 23743
rect 45004 23297 45044 24415
rect 45100 24044 45140 24751
rect 45772 24725 45812 24919
rect 45771 24716 45813 24725
rect 45771 24676 45772 24716
rect 45812 24676 45813 24716
rect 45771 24667 45813 24676
rect 45675 24632 45717 24641
rect 45675 24592 45676 24632
rect 45716 24592 45717 24632
rect 45675 24583 45717 24592
rect 45676 24498 45716 24583
rect 45100 23995 45140 24004
rect 45484 24380 45524 24389
rect 45003 23288 45045 23297
rect 45003 23248 45004 23288
rect 45044 23248 45045 23288
rect 45003 23239 45045 23248
rect 45003 22952 45045 22961
rect 45003 22912 45004 22952
rect 45044 22912 45045 22952
rect 45003 22903 45045 22912
rect 45004 22818 45044 22903
rect 45484 22625 45524 24340
rect 45772 23792 45812 24667
rect 45868 23960 45908 23969
rect 46156 23960 46196 25432
rect 46252 25229 46292 26104
rect 46348 26095 46388 26104
rect 46347 25892 46389 25901
rect 46347 25852 46348 25892
rect 46388 25852 46389 25892
rect 46347 25843 46389 25852
rect 46540 25892 46580 25901
rect 46348 25758 46388 25843
rect 46251 25220 46293 25229
rect 46251 25180 46252 25220
rect 46292 25180 46293 25220
rect 46251 25171 46293 25180
rect 46251 25052 46293 25061
rect 46251 25012 46252 25052
rect 46292 25012 46293 25052
rect 46251 25003 46293 25012
rect 46252 24809 46292 25003
rect 46540 24977 46580 25852
rect 46731 25892 46773 25901
rect 46731 25852 46732 25892
rect 46772 25852 46773 25892
rect 46731 25843 46773 25852
rect 46539 24968 46581 24977
rect 46539 24928 46540 24968
rect 46580 24928 46581 24968
rect 46539 24919 46581 24928
rect 46347 24884 46389 24893
rect 46347 24844 46348 24884
rect 46388 24844 46389 24884
rect 46347 24835 46389 24844
rect 46251 24800 46293 24809
rect 46251 24760 46252 24800
rect 46292 24760 46293 24800
rect 46251 24751 46293 24760
rect 46348 24800 46388 24835
rect 45908 23920 46196 23960
rect 45868 23911 45908 23920
rect 45772 23743 45812 23752
rect 46156 23792 46196 23801
rect 46252 23792 46292 24751
rect 46348 24749 46388 24760
rect 46539 24800 46581 24809
rect 46539 24760 46540 24800
rect 46580 24760 46581 24800
rect 46539 24751 46581 24760
rect 46540 24666 46580 24751
rect 46196 23752 46292 23792
rect 46348 24380 46388 24389
rect 46156 23743 46196 23752
rect 46348 23549 46388 24340
rect 46540 24380 46580 24389
rect 46347 23540 46389 23549
rect 46347 23500 46348 23540
rect 46388 23500 46389 23540
rect 46347 23491 46389 23500
rect 45771 23204 45813 23213
rect 45771 23164 45772 23204
rect 45812 23164 45813 23204
rect 45771 23155 45813 23164
rect 45483 22616 45525 22625
rect 45483 22576 45484 22616
rect 45524 22576 45525 22616
rect 45483 22567 45525 22576
rect 45772 22532 45812 23155
rect 46155 23120 46197 23129
rect 46155 23080 46156 23120
rect 46196 23080 46197 23120
rect 46155 23071 46197 23080
rect 46156 22986 46196 23071
rect 46155 22700 46197 22709
rect 46155 22660 46156 22700
rect 46196 22660 46197 22700
rect 46155 22651 46197 22660
rect 45772 22483 45812 22492
rect 46156 22448 46196 22651
rect 46540 22541 46580 24340
rect 46539 22532 46581 22541
rect 46539 22492 46540 22532
rect 46580 22492 46581 22532
rect 46539 22483 46581 22492
rect 46156 22399 46196 22408
rect 45100 22280 45140 22289
rect 45100 21776 45140 22240
rect 46732 22280 46772 25843
rect 46827 25472 46869 25481
rect 46827 25432 46828 25472
rect 46868 25432 46869 25472
rect 46827 25423 46869 25432
rect 46828 23792 46868 25423
rect 46924 24893 46964 27616
rect 47116 27497 47156 27952
rect 48940 27908 48980 28288
rect 49132 28328 49172 28337
rect 49172 28288 49364 28328
rect 49132 28279 49172 28288
rect 48844 27868 48980 27908
rect 48651 27824 48693 27833
rect 48651 27784 48652 27824
rect 48692 27784 48693 27824
rect 47212 27749 47252 27780
rect 48651 27775 48693 27784
rect 47211 27740 47253 27749
rect 47211 27700 47212 27740
rect 47252 27700 47253 27740
rect 47211 27691 47253 27700
rect 47212 27656 47252 27691
rect 47115 27488 47157 27497
rect 47115 27448 47116 27488
rect 47156 27448 47157 27488
rect 47115 27439 47157 27448
rect 47019 27404 47061 27413
rect 47019 27364 47020 27404
rect 47060 27364 47061 27404
rect 47019 27355 47061 27364
rect 47020 27270 47060 27355
rect 47212 27329 47252 27616
rect 47500 27656 47540 27665
rect 47500 27497 47540 27616
rect 47596 27656 47636 27667
rect 47596 27581 47636 27616
rect 47692 27656 47732 27665
rect 47595 27572 47637 27581
rect 47595 27532 47596 27572
rect 47636 27532 47637 27572
rect 47595 27523 47637 27532
rect 47692 27497 47732 27616
rect 47788 27656 47828 27665
rect 47499 27488 47541 27497
rect 47499 27448 47500 27488
rect 47540 27448 47541 27488
rect 47499 27439 47541 27448
rect 47691 27488 47733 27497
rect 47691 27448 47692 27488
rect 47732 27448 47733 27488
rect 47691 27439 47733 27448
rect 47308 27404 47348 27413
rect 47211 27320 47253 27329
rect 47211 27280 47212 27320
rect 47252 27280 47253 27320
rect 47211 27271 47253 27280
rect 47308 26489 47348 27364
rect 47307 26480 47349 26489
rect 47307 26440 47308 26480
rect 47348 26440 47349 26480
rect 47307 26431 47349 26440
rect 47692 26405 47732 27439
rect 47788 26741 47828 27616
rect 48171 27656 48213 27665
rect 48171 27616 48172 27656
rect 48212 27616 48213 27656
rect 48171 27607 48213 27616
rect 48268 27656 48308 27665
rect 48172 27522 48212 27607
rect 48268 27497 48308 27616
rect 48364 27656 48404 27665
rect 48267 27488 48309 27497
rect 48267 27448 48268 27488
rect 48308 27448 48309 27488
rect 48267 27439 48309 27448
rect 48171 27320 48213 27329
rect 48171 27280 48172 27320
rect 48212 27280 48213 27320
rect 48171 27271 48213 27280
rect 47979 27068 48021 27077
rect 47979 27028 47980 27068
rect 48020 27028 48021 27068
rect 47979 27019 48021 27028
rect 48172 27068 48212 27271
rect 48172 27019 48212 27028
rect 47980 26934 48020 27019
rect 47787 26732 47829 26741
rect 47787 26692 47788 26732
rect 47828 26692 47829 26732
rect 47787 26683 47829 26692
rect 48171 26480 48213 26489
rect 48171 26440 48172 26480
rect 48212 26440 48213 26480
rect 48171 26431 48213 26440
rect 47691 26396 47733 26405
rect 47691 26356 47692 26396
rect 47732 26356 47733 26396
rect 47691 26347 47733 26356
rect 47211 26144 47253 26153
rect 47211 26104 47212 26144
rect 47252 26104 47253 26144
rect 47211 26095 47253 26104
rect 47404 26144 47444 26153
rect 47212 25556 47252 26095
rect 47212 25507 47252 25516
rect 47404 25304 47444 26104
rect 47500 26144 47540 26153
rect 47500 25985 47540 26104
rect 47595 26144 47637 26153
rect 47595 26104 47596 26144
rect 47636 26104 47637 26144
rect 47595 26095 47637 26104
rect 47692 26144 47732 26153
rect 47884 26144 47924 26153
rect 47732 26104 47884 26144
rect 47692 26095 47732 26104
rect 47884 26095 47924 26104
rect 48075 26144 48117 26153
rect 48075 26104 48076 26144
rect 48116 26104 48117 26144
rect 48075 26095 48117 26104
rect 48172 26144 48212 26431
rect 48364 26153 48404 27616
rect 48460 27656 48500 27665
rect 48460 27497 48500 27616
rect 48652 27656 48692 27775
rect 48652 27607 48692 27616
rect 48748 27656 48788 27665
rect 48844 27656 48884 27868
rect 48940 27665 48980 27750
rect 48788 27616 48884 27656
rect 48939 27656 48981 27665
rect 48939 27616 48940 27656
rect 48980 27616 48981 27656
rect 48748 27497 48788 27616
rect 48939 27607 48981 27616
rect 49227 27572 49269 27581
rect 49227 27532 49228 27572
rect 49268 27532 49269 27572
rect 49227 27523 49269 27532
rect 48459 27488 48501 27497
rect 48459 27448 48460 27488
rect 48500 27448 48501 27488
rect 48459 27439 48501 27448
rect 48747 27488 48789 27497
rect 48747 27448 48748 27488
rect 48788 27448 48789 27488
rect 48747 27439 48789 27448
rect 49131 27488 49173 27497
rect 49131 27448 49132 27488
rect 49172 27448 49173 27488
rect 49131 27439 49173 27448
rect 48940 27404 48980 27413
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 48843 27068 48885 27077
rect 48843 27028 48844 27068
rect 48884 27028 48885 27068
rect 48843 27019 48885 27028
rect 48844 26816 48884 27019
rect 48940 26909 48980 27364
rect 49035 27404 49077 27413
rect 49035 27364 49036 27404
rect 49076 27364 49077 27404
rect 49035 27355 49077 27364
rect 48939 26900 48981 26909
rect 48939 26860 48940 26900
rect 48980 26860 48981 26900
rect 48939 26851 48981 26860
rect 48844 26767 48884 26776
rect 49036 26816 49076 27355
rect 49036 26767 49076 26776
rect 49132 26816 49172 27439
rect 49228 27438 49268 27523
rect 49324 27068 49364 28288
rect 49804 28169 49844 28254
rect 49996 28253 50036 28338
rect 50668 28328 50708 28337
rect 49995 28244 50037 28253
rect 49995 28204 49996 28244
rect 50036 28204 50037 28244
rect 49995 28195 50037 28204
rect 49803 28160 49845 28169
rect 49803 28120 49804 28160
rect 49844 28120 49845 28160
rect 49803 28111 49845 28120
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 49995 27824 50037 27833
rect 49995 27784 49996 27824
rect 50036 27784 50037 27824
rect 49995 27775 50037 27784
rect 49324 27019 49364 27028
rect 49611 26900 49653 26909
rect 49611 26860 49612 26900
rect 49652 26860 49653 26900
rect 49611 26851 49653 26860
rect 49132 26767 49172 26776
rect 49324 26816 49364 26827
rect 49324 26741 49364 26776
rect 49612 26816 49652 26851
rect 49612 26765 49652 26776
rect 49996 26816 50036 27775
rect 50380 27656 50420 27665
rect 50380 26825 50420 27616
rect 50668 27581 50708 28288
rect 50860 27833 50900 28456
rect 51244 28496 51284 28505
rect 50859 27824 50901 27833
rect 50859 27784 50860 27824
rect 50900 27784 50901 27824
rect 50859 27775 50901 27784
rect 51244 27656 51284 28456
rect 51627 28160 51669 28169
rect 51627 28120 51628 28160
rect 51668 28120 51669 28160
rect 51627 28111 51669 28120
rect 51628 27740 51668 28111
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 51628 27691 51668 27700
rect 51244 27607 51284 27616
rect 50667 27572 50709 27581
rect 50667 27532 50668 27572
rect 50708 27532 50709 27572
rect 50667 27523 50709 27532
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 49996 26767 50036 26776
rect 50187 26816 50229 26825
rect 50187 26776 50188 26816
rect 50228 26776 50229 26816
rect 50187 26767 50229 26776
rect 50379 26816 50421 26825
rect 50379 26776 50380 26816
rect 50420 26776 50421 26816
rect 50379 26767 50421 26776
rect 50859 26816 50901 26825
rect 50859 26776 50860 26816
rect 50900 26776 50901 26816
rect 50859 26767 50901 26776
rect 49323 26732 49365 26741
rect 49323 26692 49324 26732
rect 49364 26692 49365 26732
rect 49323 26683 49365 26692
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 49227 26312 49269 26321
rect 49227 26272 49228 26312
rect 49268 26272 49269 26312
rect 49227 26263 49269 26272
rect 49803 26312 49845 26321
rect 49803 26272 49804 26312
rect 49844 26272 49845 26312
rect 49803 26263 49845 26272
rect 48172 26095 48212 26104
rect 48363 26144 48405 26153
rect 48363 26104 48364 26144
rect 48404 26104 48405 26144
rect 48363 26095 48405 26104
rect 48940 26144 48980 26153
rect 47499 25976 47541 25985
rect 47499 25936 47500 25976
rect 47540 25936 47541 25976
rect 47499 25927 47541 25936
rect 47404 25061 47444 25264
rect 47500 25304 47540 25313
rect 47403 25052 47445 25061
rect 47403 25012 47404 25052
rect 47444 25012 47445 25052
rect 47403 25003 47445 25012
rect 46923 24884 46965 24893
rect 46923 24844 46924 24884
rect 46964 24844 46965 24884
rect 46923 24835 46965 24844
rect 47500 24809 47540 25264
rect 47596 25304 47636 26095
rect 48076 26010 48116 26095
rect 48748 25985 48788 26070
rect 48747 25976 48789 25985
rect 48747 25936 48748 25976
rect 48788 25936 48789 25976
rect 48747 25927 48789 25936
rect 47499 24800 47541 24809
rect 47499 24760 47500 24800
rect 47540 24760 47541 24800
rect 47499 24751 47541 24760
rect 47211 24632 47253 24641
rect 47211 24592 47212 24632
rect 47252 24592 47253 24632
rect 47211 24583 47253 24592
rect 47404 24632 47444 24641
rect 47212 24498 47252 24583
rect 46924 23792 46964 23801
rect 47404 23792 47444 24592
rect 47500 24632 47540 24641
rect 47500 24044 47540 24592
rect 47596 24632 47636 25264
rect 47884 25892 47924 25901
rect 47884 25304 47924 25852
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 47884 25255 47924 25264
rect 47691 25220 47733 25229
rect 47691 25180 47692 25220
rect 47732 25180 47733 25220
rect 47691 25171 47733 25180
rect 48459 25220 48501 25229
rect 48459 25180 48460 25220
rect 48500 25180 48501 25220
rect 48459 25171 48501 25180
rect 48556 25220 48596 25229
rect 48748 25220 48788 25229
rect 48596 25180 48748 25220
rect 48556 25171 48596 25180
rect 48748 25171 48788 25180
rect 47692 25086 47732 25171
rect 48171 25052 48213 25061
rect 48171 25012 48172 25052
rect 48212 25012 48213 25052
rect 48171 25003 48213 25012
rect 47596 24583 47636 24592
rect 47692 24632 47732 24641
rect 47980 24632 48020 24641
rect 47732 24592 47980 24632
rect 47692 24583 47732 24592
rect 47980 24583 48020 24592
rect 48172 24632 48212 25003
rect 48267 24716 48309 24725
rect 48267 24676 48268 24716
rect 48308 24676 48309 24716
rect 48267 24667 48309 24676
rect 48172 24557 48212 24592
rect 48268 24632 48308 24667
rect 48268 24581 48308 24592
rect 48460 24632 48500 25171
rect 48940 25052 48980 26104
rect 49131 25976 49173 25985
rect 49131 25936 49132 25976
rect 49172 25936 49173 25976
rect 49131 25927 49173 25936
rect 49035 25892 49077 25901
rect 49035 25852 49036 25892
rect 49076 25852 49077 25892
rect 49035 25843 49077 25852
rect 48460 24583 48500 24592
rect 48556 25012 48980 25052
rect 48171 24548 48213 24557
rect 48171 24508 48172 24548
rect 48212 24508 48213 24548
rect 48171 24499 48213 24508
rect 48172 24468 48212 24499
rect 48460 24464 48500 24473
rect 48556 24464 48596 25012
rect 48939 24716 48981 24725
rect 48939 24676 48940 24716
rect 48980 24676 48981 24716
rect 48939 24667 48981 24676
rect 48652 24632 48692 24643
rect 48652 24557 48692 24592
rect 48748 24632 48788 24641
rect 48651 24548 48693 24557
rect 48651 24508 48652 24548
rect 48692 24508 48693 24548
rect 48651 24499 48693 24508
rect 48500 24424 48596 24464
rect 48748 24464 48788 24592
rect 48940 24582 48980 24667
rect 49036 24632 49076 25843
rect 49132 25304 49172 25927
rect 49132 25255 49172 25264
rect 49036 24583 49076 24592
rect 49228 24464 49268 26263
rect 49804 26178 49844 26263
rect 49899 26144 49941 26153
rect 49899 26104 49900 26144
rect 49940 26104 49941 26144
rect 49899 26095 49941 26104
rect 49900 26010 49940 26095
rect 49612 25892 49652 25901
rect 49420 25852 49612 25892
rect 49420 24632 49460 25852
rect 49612 25843 49652 25852
rect 50091 25892 50133 25901
rect 50091 25852 50092 25892
rect 50132 25852 50133 25892
rect 50091 25843 50133 25852
rect 50092 25758 50132 25843
rect 49996 25304 50036 25313
rect 50188 25304 50228 26767
rect 50860 26682 50900 26767
rect 51627 26648 51669 26657
rect 51627 26608 51628 26648
rect 51668 26608 51669 26648
rect 51627 26599 51669 26608
rect 52011 26648 52053 26657
rect 52011 26608 52012 26648
rect 52052 26608 52053 26648
rect 52011 26599 52053 26608
rect 50764 26144 50804 26155
rect 50764 26069 50804 26104
rect 50955 26144 50997 26153
rect 50955 26104 50956 26144
rect 50996 26104 50997 26144
rect 50955 26095 50997 26104
rect 51628 26144 51668 26599
rect 52012 26514 52052 26599
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 51628 26095 51668 26104
rect 50763 26060 50805 26069
rect 50763 26020 50764 26060
rect 50804 26020 50805 26060
rect 50763 26011 50805 26020
rect 50956 26010 50996 26095
rect 51147 26060 51189 26069
rect 51147 26020 51148 26060
rect 51188 26020 51189 26060
rect 51147 26011 51189 26020
rect 51148 25556 51188 26011
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 51148 25507 51188 25516
rect 50036 25264 50228 25304
rect 49996 25255 50036 25264
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 49420 24583 49460 24592
rect 49804 24632 49844 24641
rect 50668 24632 50708 24641
rect 49844 24592 49940 24632
rect 49804 24583 49844 24592
rect 48748 24424 49268 24464
rect 48460 24415 48500 24424
rect 47980 24380 48020 24389
rect 48020 24340 48404 24380
rect 47980 24331 48020 24340
rect 48267 24212 48309 24221
rect 48267 24172 48268 24212
rect 48308 24172 48309 24212
rect 48267 24163 48309 24172
rect 47596 24044 47636 24053
rect 47500 24004 47596 24044
rect 47596 23995 47636 24004
rect 46828 23752 46924 23792
rect 46964 23752 47444 23792
rect 48268 23792 48308 24163
rect 48364 23792 48404 24340
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 49515 23960 49557 23969
rect 49515 23920 49516 23960
rect 49556 23920 49557 23960
rect 49515 23911 49557 23920
rect 49900 23960 49940 24592
rect 49900 23911 49940 23920
rect 49516 23826 49556 23911
rect 48460 23792 48500 23801
rect 48364 23752 48460 23792
rect 46924 22457 46964 23752
rect 47596 23624 47636 23633
rect 47636 23584 47732 23624
rect 47596 23575 47636 23584
rect 47403 23204 47445 23213
rect 47403 23164 47404 23204
rect 47444 23164 47445 23204
rect 47403 23155 47445 23164
rect 47020 23120 47060 23129
rect 47020 22709 47060 23080
rect 47404 23070 47444 23155
rect 47596 22952 47636 22961
rect 47116 22912 47596 22952
rect 47019 22700 47061 22709
rect 47019 22660 47020 22700
rect 47060 22660 47061 22700
rect 47019 22651 47061 22660
rect 46923 22448 46965 22457
rect 46923 22408 46924 22448
rect 46964 22408 46965 22448
rect 46923 22399 46965 22408
rect 46732 22231 46772 22240
rect 47116 22280 47156 22912
rect 47596 22903 47636 22912
rect 47116 22231 47156 22240
rect 45292 21776 45332 21785
rect 45100 21736 45292 21776
rect 45292 21727 45332 21736
rect 45387 21776 45429 21785
rect 45387 21736 45388 21776
rect 45428 21736 45429 21776
rect 45387 21727 45429 21736
rect 44908 21559 44948 21568
rect 45004 21608 45044 21617
rect 45196 21608 45236 21617
rect 45044 21568 45196 21608
rect 45004 21559 45044 21568
rect 45196 21559 45236 21568
rect 45388 21608 45428 21727
rect 47692 21701 47732 23584
rect 47979 23120 48021 23129
rect 47979 23080 47980 23120
rect 48020 23080 48021 23120
rect 48268 23120 48308 23752
rect 48460 23743 48500 23752
rect 49131 23624 49173 23633
rect 49131 23584 49132 23624
rect 49172 23584 49173 23624
rect 49131 23575 49173 23584
rect 49132 23490 49172 23575
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 49131 23288 49173 23297
rect 49131 23248 49132 23288
rect 49172 23248 49173 23288
rect 49131 23239 49173 23248
rect 48652 23120 48692 23129
rect 48268 23080 48652 23120
rect 47979 23071 48021 23080
rect 48652 23071 48692 23080
rect 47980 22280 48020 23071
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 49132 22532 49172 23239
rect 50668 23129 50708 24592
rect 51819 24632 51861 24641
rect 51819 24592 51820 24632
rect 51860 24592 51861 24632
rect 51819 24583 51861 24592
rect 51820 24498 51860 24583
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 50763 23960 50805 23969
rect 50763 23920 50764 23960
rect 50804 23920 50805 23960
rect 50763 23911 50805 23920
rect 49899 23120 49941 23129
rect 49899 23080 49900 23120
rect 49940 23080 49941 23120
rect 49899 23071 49941 23080
rect 50667 23120 50709 23129
rect 50667 23080 50668 23120
rect 50708 23080 50709 23120
rect 50667 23071 50709 23080
rect 50764 23120 50804 23911
rect 51147 23624 51189 23633
rect 51147 23584 51148 23624
rect 51188 23584 51189 23624
rect 51147 23575 51189 23584
rect 50764 23071 50804 23080
rect 51148 23120 51188 23575
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 51148 23071 51188 23080
rect 49900 22986 49940 23071
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 49132 22483 49172 22492
rect 47980 22231 48020 22240
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 47691 21692 47733 21701
rect 47691 21652 47692 21692
rect 47732 21652 47733 21692
rect 47691 21643 47733 21652
rect 45388 21559 45428 21568
rect 45483 21608 45525 21617
rect 45483 21568 45484 21608
rect 45524 21568 45525 21608
rect 45483 21559 45525 21568
rect 45484 21474 45524 21559
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 44620 20971 44660 20980
rect 43508 20728 43604 20768
rect 43468 20719 43508 20728
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 42604 20140 42836 20180
rect 42796 19928 42836 20140
rect 42796 19879 42836 19888
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 41452 18535 41492 18544
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 41067 17744 41109 17753
rect 41067 17704 41068 17744
rect 41108 17704 41109 17744
rect 41067 17695 41109 17704
rect 41260 17744 41300 17753
rect 39916 17023 39956 17032
rect 40300 17072 40340 17081
rect 40300 16400 40340 17032
rect 40491 17072 40533 17081
rect 40491 17032 40492 17072
rect 40532 17032 40533 17072
rect 41068 17072 41108 17695
rect 41164 17072 41204 17081
rect 41068 17032 41164 17072
rect 40491 17023 40533 17032
rect 41164 17023 41204 17032
rect 41164 16400 41204 16409
rect 40300 16360 41164 16400
rect 41164 16351 41204 16360
rect 39819 16316 39861 16325
rect 39819 16276 39820 16316
rect 39860 16276 39861 16316
rect 39819 16267 39861 16276
rect 39188 15352 39380 15392
rect 39436 15856 39764 15896
rect 39148 15343 39188 15352
rect 39147 15224 39189 15233
rect 39147 15184 39148 15224
rect 39188 15184 39189 15224
rect 39147 15175 39189 15184
rect 39148 14720 39188 15175
rect 39148 14671 39188 14680
rect 39436 14552 39476 15856
rect 39532 15560 39572 15569
rect 39532 15149 39572 15520
rect 39820 15233 39860 16267
rect 40108 16232 40148 16241
rect 40108 16073 40148 16192
rect 40299 16232 40341 16241
rect 40299 16192 40300 16232
rect 40340 16192 40341 16232
rect 40299 16183 40341 16192
rect 40491 16232 40533 16241
rect 40491 16192 40492 16232
rect 40532 16192 40533 16232
rect 40491 16183 40533 16192
rect 40972 16232 41012 16243
rect 40107 16064 40149 16073
rect 40107 16024 40108 16064
rect 40148 16024 40149 16064
rect 40107 16015 40149 16024
rect 40108 15653 40148 16015
rect 40107 15644 40149 15653
rect 40107 15604 40108 15644
rect 40148 15604 40149 15644
rect 40107 15595 40149 15604
rect 40300 15560 40340 16183
rect 40396 15560 40436 15569
rect 40300 15520 40396 15560
rect 40396 15511 40436 15520
rect 39819 15224 39861 15233
rect 39819 15184 39820 15224
rect 39860 15184 39861 15224
rect 39819 15175 39861 15184
rect 39531 15140 39573 15149
rect 39531 15100 39532 15140
rect 39572 15100 39573 15140
rect 39531 15091 39573 15100
rect 40492 14981 40532 16183
rect 40972 16157 41012 16192
rect 40971 16148 41013 16157
rect 40971 16108 40972 16148
rect 41012 16108 41013 16148
rect 40971 16099 41013 16108
rect 41260 16073 41300 17704
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 42316 16820 42356 16829
rect 42316 16157 42356 16780
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 42315 16148 42357 16157
rect 42315 16108 42316 16148
rect 42356 16108 42357 16148
rect 42315 16099 42357 16108
rect 41259 16064 41301 16073
rect 41259 16024 41260 16064
rect 41300 16024 41301 16064
rect 41259 16015 41301 16024
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 40491 14972 40533 14981
rect 40491 14932 40492 14972
rect 40532 14932 40533 14972
rect 40491 14923 40533 14932
rect 41547 14972 41589 14981
rect 41547 14932 41548 14972
rect 41588 14932 41589 14972
rect 41547 14923 41589 14932
rect 39148 14512 39476 14552
rect 39532 14720 39572 14729
rect 39148 14048 39188 14512
rect 39148 13999 39188 14008
rect 39244 14048 39284 14057
rect 39244 13973 39284 14008
rect 39243 13964 39285 13973
rect 39243 13924 39244 13964
rect 39284 13924 39285 13964
rect 39243 13915 39285 13924
rect 39244 13376 39284 13915
rect 39532 13880 39572 14680
rect 40395 14720 40437 14729
rect 40395 14680 40396 14720
rect 40436 14680 40437 14720
rect 40395 14671 40437 14680
rect 40396 14586 40436 14671
rect 39819 14048 39861 14057
rect 39819 14008 39820 14048
rect 39860 14008 39861 14048
rect 39819 13999 39861 14008
rect 40492 14048 40532 14923
rect 41548 14838 41588 14923
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 40492 13999 40532 14008
rect 39820 13914 39860 13999
rect 39628 13880 39668 13889
rect 39532 13840 39628 13880
rect 39628 13831 39668 13840
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 39339 13376 39381 13385
rect 39244 13336 39340 13376
rect 39380 13336 39381 13376
rect 39339 13327 39381 13336
rect 39340 13242 39380 13327
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 39052 12487 39092 12496
rect 36172 12328 36404 12368
rect 35980 12284 36020 12293
rect 38380 12284 38420 12293
rect 36020 12244 36308 12284
rect 35980 12235 36020 12244
rect 36076 11696 36116 11707
rect 36076 11621 36116 11656
rect 36268 11696 36308 12244
rect 36268 11647 36308 11656
rect 36940 11696 36980 11705
rect 37132 11696 37172 11705
rect 36980 11656 37132 11696
rect 36940 11647 36980 11656
rect 37132 11647 37172 11656
rect 37516 11696 37556 11705
rect 36075 11612 36117 11621
rect 36075 11572 36076 11612
rect 36116 11572 36117 11612
rect 36075 11563 36117 11572
rect 37516 11453 37556 11656
rect 38380 11696 38420 12244
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 37803 11612 37845 11621
rect 37803 11572 37804 11612
rect 37844 11572 37845 11612
rect 37803 11563 37845 11572
rect 37515 11444 37557 11453
rect 37515 11404 37516 11444
rect 37556 11404 37557 11444
rect 37515 11395 37557 11404
rect 37707 11444 37749 11453
rect 37707 11404 37708 11444
rect 37748 11404 37749 11444
rect 37707 11395 37749 11404
rect 36075 11108 36117 11117
rect 36075 11068 36076 11108
rect 36116 11068 36117 11108
rect 36075 11059 36117 11068
rect 35883 10772 35925 10781
rect 35883 10732 35884 10772
rect 35924 10732 35925 10772
rect 35883 10723 35925 10732
rect 35691 10436 35733 10445
rect 35691 10396 35692 10436
rect 35732 10396 35733 10436
rect 35691 10387 35733 10396
rect 35787 10268 35829 10277
rect 35787 10228 35788 10268
rect 35828 10228 35829 10268
rect 35787 10219 35829 10228
rect 34348 9967 34388 9976
rect 34444 9976 34676 10016
rect 35019 10016 35061 10025
rect 35019 9976 35020 10016
rect 35060 9976 35061 10016
rect 34444 9848 34484 9976
rect 35019 9967 35061 9976
rect 34348 9808 34484 9848
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34251 9512 34293 9521
rect 34251 9472 34252 9512
rect 34292 9472 34293 9512
rect 34251 9463 34293 9472
rect 34252 9378 34292 9463
rect 34155 9260 34197 9269
rect 34155 9220 34156 9260
rect 34196 9220 34197 9260
rect 34155 9211 34197 9220
rect 34156 9126 34196 9211
rect 34348 9101 34388 9808
rect 34592 9799 34960 9808
rect 34443 9680 34485 9689
rect 34443 9640 34444 9680
rect 34484 9640 34485 9680
rect 34443 9631 34485 9640
rect 34444 9512 34484 9631
rect 34444 9437 34484 9472
rect 34540 9512 34676 9526
rect 34540 9486 34636 9512
rect 34540 9437 34580 9486
rect 34636 9463 34676 9472
rect 34732 9512 34772 9521
rect 34817 9512 34868 9526
rect 34772 9472 34868 9512
rect 34732 9463 34772 9472
rect 34443 9428 34485 9437
rect 34443 9388 34444 9428
rect 34484 9388 34485 9428
rect 34540 9428 34586 9437
rect 34540 9388 34545 9428
rect 34585 9388 34586 9428
rect 34443 9379 34485 9388
rect 34544 9379 34586 9388
rect 34444 9260 34484 9269
rect 34484 9220 34676 9260
rect 34444 9211 34484 9220
rect 34059 9092 34101 9101
rect 34059 9052 34060 9092
rect 34100 9052 34101 9092
rect 34059 9043 34101 9052
rect 34347 9092 34389 9101
rect 34347 9052 34348 9092
rect 34388 9052 34389 9092
rect 34347 9043 34389 9052
rect 34539 9092 34581 9101
rect 34539 9052 34540 9092
rect 34580 9052 34581 9092
rect 34539 9043 34581 9052
rect 33964 8800 34100 8840
rect 33963 8672 34005 8681
rect 33963 8632 33964 8672
rect 34004 8632 34005 8672
rect 33963 8623 34005 8632
rect 33964 8538 34004 8623
rect 34060 8093 34100 8800
rect 34155 8756 34197 8765
rect 34155 8716 34156 8756
rect 34196 8716 34197 8756
rect 34155 8707 34197 8716
rect 34156 8622 34196 8707
rect 34252 8672 34292 8681
rect 34444 8672 34484 8681
rect 34540 8672 34580 9043
rect 34636 8933 34676 9220
rect 34828 9101 34868 9472
rect 34924 9512 34964 9521
rect 35020 9512 35060 9967
rect 35212 9689 35252 9774
rect 35211 9680 35253 9689
rect 35211 9640 35212 9680
rect 35252 9640 35253 9680
rect 35500 9680 35540 10144
rect 35596 10184 35636 10193
rect 35596 10025 35636 10144
rect 35788 10184 35828 10219
rect 36076 10184 36116 11059
rect 36652 11024 36692 11033
rect 36652 10193 36692 10984
rect 36556 10184 36596 10193
rect 35788 10133 35828 10144
rect 35884 10144 36076 10184
rect 35595 10016 35637 10025
rect 35595 9976 35596 10016
rect 35636 9976 35732 10016
rect 35595 9967 35637 9976
rect 35596 9680 35636 9689
rect 35500 9640 35596 9680
rect 35211 9631 35253 9640
rect 34964 9472 35060 9512
rect 35116 9512 35156 9521
rect 34924 9463 34964 9472
rect 35116 9101 35156 9472
rect 35211 9512 35253 9521
rect 35211 9472 35212 9512
rect 35252 9472 35253 9512
rect 35211 9463 35253 9472
rect 35212 9378 35252 9463
rect 35596 9353 35636 9640
rect 35692 9512 35732 9976
rect 35884 9680 35924 10144
rect 36076 10135 36116 10144
rect 36268 10144 36556 10184
rect 36268 10100 36308 10144
rect 36556 10135 36596 10144
rect 36651 10184 36693 10193
rect 36651 10144 36652 10184
rect 36692 10144 36693 10184
rect 36651 10135 36693 10144
rect 37228 10184 37268 10193
rect 37420 10184 37460 10193
rect 37268 10144 37420 10184
rect 37708 10184 37748 11395
rect 37804 11024 37844 11563
rect 37804 10975 37844 10984
rect 38091 11024 38133 11033
rect 38091 10984 38092 11024
rect 38132 10984 38133 11024
rect 38091 10975 38133 10984
rect 38092 10890 38132 10975
rect 38187 10352 38229 10361
rect 38187 10312 38188 10352
rect 38228 10312 38229 10352
rect 38187 10303 38229 10312
rect 37804 10184 37844 10193
rect 37708 10144 37804 10184
rect 37228 10135 37268 10144
rect 37420 10135 37460 10144
rect 37804 10135 37844 10144
rect 37899 10184 37941 10193
rect 37899 10144 37900 10184
rect 37940 10144 37941 10184
rect 37899 10135 37941 10144
rect 36268 10051 36308 10060
rect 35884 9631 35924 9640
rect 35692 9463 35732 9472
rect 36268 9512 36308 9521
rect 35595 9344 35637 9353
rect 35595 9304 35596 9344
rect 35636 9304 35637 9344
rect 35595 9295 35637 9304
rect 35403 9260 35445 9269
rect 35403 9220 35404 9260
rect 35444 9220 35445 9260
rect 35403 9211 35445 9220
rect 35884 9260 35924 9269
rect 34827 9092 34869 9101
rect 34827 9052 34828 9092
rect 34868 9052 34869 9092
rect 34827 9043 34869 9052
rect 35115 9092 35157 9101
rect 35115 9052 35116 9092
rect 35156 9052 35157 9092
rect 35115 9043 35157 9052
rect 34635 8924 34677 8933
rect 34635 8884 34636 8924
rect 34676 8884 34677 8924
rect 34635 8875 34677 8884
rect 34732 8716 35060 8756
rect 34732 8697 34772 8716
rect 34252 8177 34292 8632
rect 34348 8632 34444 8672
rect 34484 8632 34580 8672
rect 34636 8672 34676 8681
rect 34732 8648 34772 8657
rect 34251 8168 34293 8177
rect 34251 8128 34252 8168
rect 34292 8128 34293 8168
rect 34251 8119 34293 8128
rect 34059 8084 34101 8093
rect 34059 8044 34060 8084
rect 34100 8044 34101 8084
rect 34059 8035 34101 8044
rect 34348 8009 34388 8632
rect 34444 8623 34484 8632
rect 34636 8588 34676 8632
rect 34827 8588 34869 8597
rect 34636 8548 34828 8588
rect 34868 8548 34869 8588
rect 34827 8539 34869 8548
rect 34444 8464 34772 8504
rect 34444 8168 34484 8464
rect 34732 8462 34772 8464
rect 34732 8413 34772 8422
rect 35020 8345 35060 8716
rect 35307 8672 35349 8681
rect 35307 8632 35308 8672
rect 35348 8632 35349 8672
rect 35307 8623 35349 8632
rect 35404 8672 35444 9211
rect 35596 8840 35636 8849
rect 35636 8800 35828 8840
rect 35596 8791 35636 8800
rect 35404 8623 35444 8632
rect 35596 8672 35636 8681
rect 35308 8538 35348 8623
rect 35596 8504 35636 8632
rect 35788 8672 35828 8800
rect 35788 8623 35828 8632
rect 35884 8504 35924 9220
rect 36268 8765 36308 9472
rect 37323 9512 37365 9521
rect 37323 9472 37324 9512
rect 37364 9472 37365 9512
rect 37323 9463 37365 9472
rect 37324 9378 37364 9463
rect 36940 9260 36980 9269
rect 36748 9220 36940 9260
rect 36267 8756 36309 8765
rect 36267 8716 36268 8756
rect 36308 8716 36309 8756
rect 36267 8707 36309 8716
rect 36460 8672 36500 8681
rect 36652 8672 36692 8681
rect 36500 8632 36652 8672
rect 36460 8623 36500 8632
rect 36652 8623 36692 8632
rect 36748 8504 36788 9220
rect 36940 9211 36980 9220
rect 37036 8672 37076 8681
rect 37900 8672 37940 10135
rect 38188 9680 38228 10303
rect 38380 10193 38420 11656
rect 38763 11696 38805 11705
rect 38763 11656 38764 11696
rect 38804 11656 38805 11696
rect 38763 11647 38805 11656
rect 39531 11696 39573 11705
rect 39531 11656 39532 11696
rect 39572 11656 39573 11696
rect 39531 11647 39573 11656
rect 38764 11024 38804 11647
rect 39532 11562 39572 11647
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 38764 10975 38804 10984
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 38379 10184 38421 10193
rect 38379 10144 38380 10184
rect 38420 10144 38421 10184
rect 38379 10135 38421 10144
rect 38667 10184 38709 10193
rect 38667 10144 38668 10184
rect 38708 10144 38709 10184
rect 38667 10135 38709 10144
rect 39820 10184 39860 10195
rect 38668 10050 38708 10135
rect 39820 10109 39860 10144
rect 38859 10100 38901 10109
rect 38859 10060 38860 10100
rect 38900 10060 38901 10100
rect 38859 10051 38901 10060
rect 39819 10100 39861 10109
rect 39819 10060 39820 10100
rect 39860 10060 39861 10100
rect 39819 10051 39861 10060
rect 38188 9631 38228 9640
rect 37996 9512 38036 9521
rect 37996 9437 38036 9472
rect 38860 9512 38900 10051
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 38860 9463 38900 9472
rect 37995 9428 38037 9437
rect 37995 9388 37996 9428
rect 38036 9388 38037 9428
rect 37995 9379 38037 9388
rect 37996 8933 38036 9379
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 37995 8924 38037 8933
rect 37995 8884 37996 8924
rect 38036 8884 38037 8924
rect 37995 8875 38037 8884
rect 39051 8924 39093 8933
rect 39051 8884 39052 8924
rect 39092 8884 39093 8924
rect 39051 8875 39093 8884
rect 39052 8790 39092 8875
rect 35596 8464 35924 8504
rect 36556 8464 36788 8504
rect 36940 8632 37036 8672
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 35019 8336 35061 8345
rect 35019 8296 35020 8336
rect 35060 8296 35061 8336
rect 35019 8287 35061 8296
rect 34636 8168 34676 8177
rect 34444 8128 34636 8168
rect 33964 8000 34004 8009
rect 33964 7421 34004 7960
rect 34347 8000 34389 8009
rect 34347 7960 34348 8000
rect 34388 7960 34389 8000
rect 34347 7951 34389 7960
rect 34059 7748 34101 7757
rect 34059 7708 34060 7748
rect 34100 7708 34101 7748
rect 34059 7699 34101 7708
rect 33963 7412 34005 7421
rect 33963 7372 33964 7412
rect 34004 7372 34005 7412
rect 33963 7363 34005 7372
rect 33867 7160 33909 7169
rect 33867 7120 33868 7160
rect 33908 7120 33909 7160
rect 33867 7111 33909 7120
rect 34060 7076 34100 7699
rect 34348 7589 34388 7951
rect 34347 7580 34389 7589
rect 34347 7540 34348 7580
rect 34388 7540 34389 7580
rect 34347 7531 34389 7540
rect 33964 7036 34100 7076
rect 33484 6439 33524 6448
rect 33867 6488 33909 6497
rect 33867 6448 33868 6488
rect 33908 6448 33909 6488
rect 33867 6439 33909 6448
rect 33772 6236 33812 6245
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 33195 5648 33237 5657
rect 33195 5608 33196 5648
rect 33236 5608 33237 5648
rect 33195 5599 33237 5608
rect 33484 5648 33524 5657
rect 33484 5489 33524 5608
rect 33772 5648 33812 6196
rect 33772 5599 33812 5608
rect 33483 5480 33525 5489
rect 33483 5440 33484 5480
rect 33524 5440 33525 5480
rect 33483 5431 33525 5440
rect 33676 5480 33716 5489
rect 33868 5480 33908 6439
rect 33964 5741 34004 7036
rect 34444 6656 34484 8128
rect 34636 8119 34676 8128
rect 35691 8168 35733 8177
rect 35691 8128 35692 8168
rect 35732 8128 35733 8168
rect 35691 8119 35733 8128
rect 35692 8034 35732 8119
rect 34828 8000 34868 8009
rect 36364 8000 36404 8009
rect 34868 7960 35156 8000
rect 34828 7951 34868 7960
rect 34923 7160 34965 7169
rect 34923 7120 34924 7160
rect 34964 7120 34965 7160
rect 34923 7111 34965 7120
rect 34924 7026 34964 7111
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 34444 6616 34580 6656
rect 34444 6488 34484 6497
rect 34252 5900 34292 5909
rect 34444 5900 34484 6448
rect 34292 5860 34484 5900
rect 34252 5851 34292 5860
rect 33963 5732 34005 5741
rect 33963 5692 33964 5732
rect 34004 5692 34005 5732
rect 33963 5683 34005 5692
rect 33964 5648 34004 5683
rect 33964 5598 34004 5608
rect 34060 5648 34100 5659
rect 34060 5573 34100 5608
rect 34252 5648 34292 5657
rect 34444 5648 34484 5657
rect 34540 5648 34580 6616
rect 34635 6488 34677 6497
rect 34635 6448 34636 6488
rect 34676 6448 34677 6488
rect 34635 6439 34677 6448
rect 34636 6354 34676 6439
rect 35116 5816 35156 7960
rect 36364 7841 36404 7960
rect 36556 8000 36596 8464
rect 36651 8336 36693 8345
rect 36651 8296 36652 8336
rect 36692 8296 36693 8336
rect 36651 8287 36693 8296
rect 36556 7951 36596 7960
rect 36363 7832 36405 7841
rect 36363 7792 36364 7832
rect 36404 7792 36405 7832
rect 36363 7783 36405 7792
rect 35500 7748 35540 7757
rect 35211 7580 35253 7589
rect 35211 7540 35212 7580
rect 35252 7540 35253 7580
rect 35211 7531 35253 7540
rect 35116 5767 35156 5776
rect 34731 5732 34773 5741
rect 34731 5692 34732 5732
rect 34772 5692 34773 5732
rect 34731 5683 34773 5692
rect 35019 5732 35061 5741
rect 35019 5692 35020 5732
rect 35060 5692 35061 5732
rect 35019 5683 35061 5692
rect 35212 5732 35252 7531
rect 35307 6656 35349 6665
rect 35307 6616 35308 6656
rect 35348 6616 35349 6656
rect 35307 6607 35349 6616
rect 35308 6522 35348 6607
rect 35500 6488 35540 7708
rect 36556 7412 36596 7421
rect 36652 7412 36692 8287
rect 36747 8000 36789 8009
rect 36747 7960 36748 8000
rect 36788 7960 36789 8000
rect 36747 7951 36789 7960
rect 36940 8000 36980 8632
rect 37036 8623 37076 8632
rect 37804 8632 37900 8672
rect 37419 8084 37461 8093
rect 37419 8044 37420 8084
rect 37460 8044 37461 8084
rect 37419 8035 37461 8044
rect 36596 7372 36692 7412
rect 36556 7363 36596 7372
rect 35787 7328 35829 7337
rect 35787 7288 35788 7328
rect 35828 7288 35829 7328
rect 35787 7279 35829 7288
rect 35788 7160 35828 7279
rect 35788 6488 35828 7120
rect 36172 7160 36212 7169
rect 36172 6665 36212 7120
rect 36171 6656 36213 6665
rect 36171 6616 36172 6656
rect 36212 6616 36213 6656
rect 36171 6607 36213 6616
rect 35884 6488 35924 6497
rect 35788 6448 35884 6488
rect 35500 6439 35540 6448
rect 35884 6439 35924 6448
rect 36748 6488 36788 7951
rect 36940 7337 36980 7960
rect 37420 7412 37460 8035
rect 37804 8009 37844 8632
rect 37900 8623 37940 8632
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 37803 8000 37845 8009
rect 37803 7960 37804 8000
rect 37844 7960 37845 8000
rect 37803 7951 37845 7960
rect 37804 7866 37844 7951
rect 37420 7363 37460 7372
rect 38956 7748 38996 7757
rect 36939 7328 36981 7337
rect 36939 7288 36940 7328
rect 36980 7288 36981 7328
rect 36939 7279 36981 7288
rect 38956 7253 38996 7708
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 38091 7244 38133 7253
rect 38091 7204 38092 7244
rect 38132 7204 38133 7244
rect 38091 7195 38133 7204
rect 38955 7244 38997 7253
rect 38955 7204 38956 7244
rect 38996 7204 38997 7244
rect 38955 7195 38997 7204
rect 37228 7160 37268 7171
rect 37228 7085 37268 7120
rect 38092 7160 38132 7195
rect 38092 7109 38132 7120
rect 37227 7076 37269 7085
rect 37227 7036 37228 7076
rect 37268 7036 37269 7076
rect 37227 7027 37269 7036
rect 37899 7076 37941 7085
rect 37899 7036 37900 7076
rect 37940 7036 37941 7076
rect 37899 7027 37941 7036
rect 36748 6439 36788 6448
rect 37900 6488 37940 7027
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 37900 6439 37940 6448
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 35212 5683 35252 5692
rect 34292 5608 34444 5648
rect 34484 5608 34580 5648
rect 34636 5648 34676 5659
rect 34252 5599 34292 5608
rect 34444 5599 34484 5608
rect 34636 5573 34676 5608
rect 34732 5648 34772 5683
rect 34732 5597 34772 5608
rect 34924 5648 34964 5657
rect 34059 5564 34101 5573
rect 34059 5524 34060 5564
rect 34100 5524 34101 5564
rect 34059 5515 34101 5524
rect 34635 5564 34677 5573
rect 34635 5524 34636 5564
rect 34676 5524 34677 5564
rect 34635 5515 34677 5524
rect 34924 5489 34964 5608
rect 35020 5598 35060 5683
rect 35307 5648 35349 5657
rect 35307 5608 35308 5648
rect 35348 5608 35349 5648
rect 35307 5599 35349 5608
rect 35308 5514 35348 5599
rect 33716 5440 33908 5480
rect 34443 5480 34485 5489
rect 34443 5440 34444 5480
rect 34484 5440 34485 5480
rect 33676 5431 33716 5440
rect 34443 5431 34485 5440
rect 34923 5480 34965 5489
rect 34923 5440 34924 5480
rect 34964 5440 34965 5480
rect 34923 5431 34965 5440
rect 34444 5346 34484 5431
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 32620 4087 32660 4096
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 31892 3424 31988 3464
rect 30412 3330 30452 3415
rect 30220 2827 30260 2836
rect 29356 2071 29396 2080
rect 28780 1903 28820 1912
rect 29452 1952 29492 2827
rect 29836 2742 29876 2827
rect 30892 2633 30932 2718
rect 31852 2633 31892 3424
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 30891 2624 30933 2633
rect 30891 2584 30892 2624
rect 30932 2584 30933 2624
rect 30891 2575 30933 2584
rect 31851 2624 31893 2633
rect 31851 2584 31852 2624
rect 31892 2584 31893 2624
rect 31851 2575 31893 2584
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 29452 1903 29492 1912
rect 27532 1818 27572 1903
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 26764 1063 26804 1072
rect 25611 944 25653 953
rect 25611 904 25612 944
rect 25652 904 25653 944
rect 25611 895 25653 904
rect 25995 944 26037 953
rect 25995 904 25996 944
rect 26036 904 26037 944
rect 25995 895 26037 904
rect 26475 944 26517 953
rect 26475 904 26476 944
rect 26516 904 26517 944
rect 26475 895 26517 904
rect 25996 810 26036 895
rect 26476 810 26516 895
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 268 37528 308 37568
rect 27436 37528 27476 37568
rect 27820 37528 27860 37568
rect 26572 37192 26612 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 12652 36436 12692 36476
rect 13132 36520 13172 36560
rect 13900 36520 13940 36560
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 5932 35260 5972 35300
rect 6988 35260 7028 35300
rect 4780 35176 4820 35216
rect 5356 35176 5396 35216
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 1324 33076 1364 33116
rect 3628 34336 3668 34376
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3244 33916 3284 33956
rect 5452 35092 5492 35132
rect 5644 34336 5684 34376
rect 4972 34084 5012 34124
rect 4876 34000 4916 34040
rect 6028 35092 6068 35132
rect 5836 34084 5876 34124
rect 5740 34000 5780 34040
rect 5068 33832 5108 33872
rect 4684 33664 4724 33704
rect 2764 33580 2804 33620
rect 4396 33580 4436 33620
rect 2380 32992 2420 33032
rect 1996 32908 2036 32948
rect 2188 32824 2228 32864
rect 4204 33496 4244 33536
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 3724 32992 3764 33032
rect 3052 32908 3092 32948
rect 2860 32824 2900 32864
rect 2668 32740 2708 32780
rect 4012 32824 4052 32864
rect 5164 33748 5204 33788
rect 6028 34588 6068 34628
rect 5356 33664 5396 33704
rect 5932 33664 5972 33704
rect 6028 33580 6068 33620
rect 4972 33496 5012 33536
rect 4492 33076 4532 33116
rect 4780 33076 4820 33116
rect 4684 32824 4724 32864
rect 4204 32740 4244 32780
rect 1228 31144 1268 31184
rect 1036 29968 1076 30008
rect 2092 31480 2132 31520
rect 3724 32152 3764 32192
rect 3532 31900 3572 31940
rect 4108 31900 4148 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 3436 31480 3476 31520
rect 2668 31396 2708 31436
rect 1612 29968 1652 30008
rect 2572 29128 2612 29168
rect 1324 28960 1364 29000
rect 1324 28204 1364 28244
rect 1228 26776 1268 26816
rect 4012 31480 4052 31520
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4108 31312 4148 31352
rect 4972 32740 5012 32780
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 4780 32177 4820 32192
rect 4780 32152 4820 32177
rect 6508 34924 6548 34964
rect 6316 34000 6356 34040
rect 6412 33748 6452 33788
rect 7660 34924 7700 34964
rect 8812 35176 8852 35216
rect 8908 35092 8948 35132
rect 8812 34924 8852 34964
rect 8332 34588 8372 34628
rect 9196 35092 9236 35132
rect 9100 34588 9140 34628
rect 11884 35680 11924 35720
rect 10924 35176 10964 35216
rect 9676 34504 9716 34544
rect 10444 34504 10484 34544
rect 8332 34000 8372 34040
rect 6700 33916 6740 33956
rect 7468 33916 7508 33956
rect 6604 33664 6644 33704
rect 6412 33496 6452 33536
rect 6412 33328 6452 33368
rect 6124 32908 6164 32948
rect 5452 32824 5492 32864
rect 5356 32740 5396 32780
rect 4588 31480 4628 31520
rect 3724 30556 3764 30596
rect 4780 31480 4820 31520
rect 4972 31312 5012 31352
rect 6604 32824 6644 32864
rect 6508 32740 6548 32780
rect 5644 32656 5684 32696
rect 6316 32656 6356 32696
rect 8908 34000 8948 34040
rect 8620 33832 8660 33872
rect 6988 33748 7028 33788
rect 7180 33580 7220 33620
rect 6892 33160 6932 33200
rect 7084 32992 7124 33032
rect 6220 32152 6260 32192
rect 6700 32152 6740 32192
rect 6892 32824 6932 32864
rect 7084 32824 7124 32864
rect 6796 31480 6836 31520
rect 6892 31396 6932 31436
rect 4588 31144 4628 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3724 30304 3764 30344
rect 2764 29212 2804 29252
rect 3340 29884 3380 29924
rect 3628 29884 3668 29924
rect 3244 29212 3284 29252
rect 4108 29968 4148 30008
rect 3820 29800 3860 29840
rect 3532 29212 3572 29252
rect 3724 29128 3764 29168
rect 2956 29044 2996 29084
rect 3916 29128 3956 29168
rect 2764 28960 2804 29000
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3820 28456 3860 28496
rect 4684 30472 4724 30512
rect 4396 29968 4436 30008
rect 6124 30472 6164 30512
rect 5932 30304 5972 30344
rect 5548 29968 5588 30008
rect 5836 29968 5876 30008
rect 5068 29884 5108 29924
rect 4780 29800 4820 29840
rect 5164 29800 5204 29840
rect 5644 29800 5684 29840
rect 4588 29632 4628 29672
rect 4108 29380 4148 29420
rect 5260 29632 5300 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 5644 29380 5684 29420
rect 5356 29296 5396 29336
rect 5548 29296 5588 29336
rect 4204 29212 4244 29252
rect 5164 29212 5204 29252
rect 4684 29128 4724 29168
rect 4204 28456 4244 28496
rect 4876 28456 4916 28496
rect 4300 28288 4340 28328
rect 4108 28204 4148 28244
rect 3052 27700 3092 27740
rect 3340 27616 3380 27656
rect 2956 27364 2996 27404
rect 2764 27280 2804 27320
rect 3724 27616 3764 27656
rect 4780 28036 4820 28076
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 4204 27784 4244 27824
rect 4684 27784 4724 27824
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3628 27196 3668 27236
rect 3628 27028 3668 27068
rect 1228 26188 1268 26228
rect 3820 26776 3860 26816
rect 3628 26272 3668 26312
rect 4012 27448 4052 27488
rect 4108 27196 4148 27236
rect 4876 27784 4916 27824
rect 5740 29296 5780 29336
rect 6028 29296 6068 29336
rect 5836 29212 5876 29252
rect 6988 30640 7028 30680
rect 6604 30556 6644 30596
rect 6508 29632 6548 29672
rect 6316 29464 6356 29504
rect 9004 33832 9044 33872
rect 9388 34168 9428 34208
rect 10252 34336 10292 34376
rect 9580 33832 9620 33872
rect 11692 35092 11732 35132
rect 12076 35008 12116 35048
rect 13228 36436 13268 36476
rect 12940 35680 12980 35720
rect 12940 35260 12980 35300
rect 11596 34924 11636 34964
rect 10828 34336 10868 34376
rect 11212 34336 11252 34376
rect 11884 34588 11924 34628
rect 11692 34420 11732 34460
rect 11500 34252 11540 34292
rect 10636 34084 10676 34124
rect 7852 33328 7892 33368
rect 7564 32908 7604 32948
rect 7276 32740 7316 32780
rect 7660 32656 7700 32696
rect 8236 33160 8276 33200
rect 8140 32992 8180 33032
rect 8044 32824 8084 32864
rect 8236 32824 8276 32864
rect 7948 32656 7988 32696
rect 8140 32152 8180 32192
rect 8428 32740 8468 32780
rect 7180 30640 7220 30680
rect 7180 29632 7220 29672
rect 6220 29128 6260 29168
rect 7660 31480 7700 31520
rect 7468 30556 7508 30596
rect 8332 31480 8372 31520
rect 9196 33664 9236 33704
rect 9292 32908 9332 32948
rect 9868 33076 9908 33116
rect 9004 32824 9044 32864
rect 9676 32824 9716 32864
rect 8812 32740 8852 32780
rect 9676 31732 9716 31772
rect 8812 31480 8852 31520
rect 10540 33664 10580 33704
rect 9964 32824 10004 32864
rect 8716 31396 8756 31436
rect 8332 30976 8372 31016
rect 7564 30304 7604 30344
rect 7852 30220 7892 30260
rect 7564 29968 7604 30008
rect 7660 29800 7700 29840
rect 6124 29044 6164 29084
rect 5164 28288 5204 28328
rect 5068 27364 5108 27404
rect 6028 28120 6068 28160
rect 5356 28036 5396 28076
rect 5932 27616 5972 27656
rect 5164 27028 5204 27068
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 4588 26272 4628 26312
rect 4396 26188 4436 26228
rect 1036 25936 1076 25976
rect 1612 25936 1652 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 1132 24592 1172 24632
rect 3436 25348 3476 25388
rect 3532 25264 3572 25304
rect 2668 25180 2708 25220
rect 1228 23164 1268 23204
rect 2380 23836 2420 23876
rect 2284 23752 2324 23792
rect 2572 23752 2612 23792
rect 3628 25180 3668 25220
rect 2764 24592 2804 24632
rect 3532 24508 3572 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3532 23920 3572 23960
rect 4012 25684 4052 25724
rect 4012 25348 4052 25388
rect 4492 26104 4532 26144
rect 4780 26188 4820 26228
rect 5644 26692 5684 26732
rect 7276 29128 7316 29168
rect 7180 29044 7220 29084
rect 7372 29044 7412 29084
rect 5740 26272 5780 26312
rect 4396 25348 4436 25388
rect 4780 25264 4820 25304
rect 4492 25180 4532 25220
rect 4396 25096 4436 25136
rect 4204 24928 4244 24968
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4108 24508 4148 24548
rect 4492 24508 4532 24548
rect 4012 24004 4052 24044
rect 3820 23836 3860 23876
rect 3052 23752 3092 23792
rect 3148 23164 3188 23204
rect 652 22408 692 22448
rect 652 21568 692 21608
rect 268 20896 308 20936
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 1228 22828 1268 22868
rect 3628 23752 3668 23792
rect 3340 23248 3380 23288
rect 2476 22240 2516 22280
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3148 22240 3188 22280
rect 3628 22240 3668 22280
rect 5068 26104 5108 26144
rect 4972 25264 5012 25304
rect 5452 26104 5492 26144
rect 4876 24340 4916 24380
rect 4396 24004 4436 24044
rect 4204 23752 4244 23792
rect 4684 23836 4724 23876
rect 4780 23752 4820 23792
rect 5356 25180 5396 25220
rect 6700 28036 6740 28076
rect 7276 28288 7316 28328
rect 7468 28372 7508 28412
rect 7180 28204 7220 28244
rect 7372 28120 7412 28160
rect 7276 28036 7316 28076
rect 6796 27952 6836 27992
rect 6604 27784 6644 27824
rect 7084 27700 7124 27740
rect 6988 27196 7028 27236
rect 8140 29968 8180 30008
rect 7948 29296 7988 29336
rect 8044 29128 8084 29168
rect 7852 27952 7892 27992
rect 7756 27784 7796 27824
rect 7564 27700 7604 27740
rect 7660 27532 7700 27572
rect 6796 25684 6836 25724
rect 5356 24256 5396 24296
rect 5260 24004 5300 24044
rect 5836 24004 5876 24044
rect 5740 23920 5780 23960
rect 5644 23836 5684 23876
rect 4396 23584 4436 23624
rect 4588 23584 4628 23624
rect 3916 23500 3956 23540
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 4012 22912 4052 22952
rect 3916 22828 3956 22868
rect 2860 22156 2900 22196
rect 1804 21652 1844 21692
rect 2764 21652 2804 21692
rect 2668 21568 2708 21608
rect 2956 21652 2996 21692
rect 3916 21820 3956 21860
rect 3820 21568 3860 21608
rect 4204 23080 4244 23120
rect 4972 23584 5012 23624
rect 5164 23416 5204 23456
rect 4972 23164 5012 23204
rect 4492 22912 4532 22952
rect 4108 22156 4148 22196
rect 4108 21568 4148 21608
rect 4012 21484 4052 21524
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 5452 23080 5492 23120
rect 5548 22660 5588 22700
rect 6316 23920 6356 23960
rect 5932 23668 5972 23708
rect 6028 23248 6068 23288
rect 5740 23164 5780 23204
rect 6124 23164 6164 23204
rect 6316 22996 6356 23036
rect 4300 22240 4340 22280
rect 4876 22240 4916 22280
rect 5164 22156 5204 22196
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 5068 21820 5108 21860
rect 4492 21400 4532 21440
rect 5164 21736 5204 21776
rect 6796 24004 6836 24044
rect 6508 23248 6548 23288
rect 6700 23080 6740 23120
rect 6412 22408 6452 22448
rect 6508 22240 6548 22280
rect 6124 22156 6164 22196
rect 5836 21652 5876 21692
rect 5356 21484 5396 21524
rect 5068 21232 5108 21272
rect 1324 19048 1364 19088
rect 4204 20728 4244 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3724 19384 3764 19424
rect 4492 19384 4532 19424
rect 4204 19300 4244 19340
rect 3724 19132 3764 19172
rect 2572 18544 2612 18584
rect 2764 18544 2804 18584
rect 2956 18544 2996 18584
rect 3820 18544 3860 18584
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3628 17536 3668 17576
rect 1516 17200 1556 17240
rect 3532 17116 3572 17156
rect 3244 17032 3284 17072
rect 4492 19216 4532 19256
rect 5452 21400 5492 21440
rect 5260 20728 5300 20768
rect 5356 20056 5396 20096
rect 5548 20980 5588 21020
rect 5932 21484 5972 21524
rect 6604 22156 6644 22196
rect 6220 20980 6260 21020
rect 6508 20224 6548 20264
rect 5740 19888 5780 19928
rect 5836 19384 5876 19424
rect 6124 19216 6164 19256
rect 6796 21652 6836 21692
rect 7756 27448 7796 27488
rect 8716 31228 8756 31268
rect 8428 30472 8468 30512
rect 8428 29632 8468 29672
rect 8332 28876 8372 28916
rect 8236 28204 8276 28244
rect 8140 27616 8180 27656
rect 8044 27532 8084 27572
rect 7948 26440 7988 26480
rect 7852 26188 7892 26228
rect 7468 25348 7508 25388
rect 7852 25348 7892 25388
rect 6988 25180 7028 25220
rect 8236 25852 8276 25892
rect 8140 24760 8180 24800
rect 7468 24256 7508 24296
rect 7756 23920 7796 23960
rect 7180 23248 7220 23288
rect 7468 23164 7508 23204
rect 6988 23080 7028 23120
rect 7276 23080 7316 23120
rect 7084 22996 7124 23036
rect 6892 21568 6932 21608
rect 7756 22408 7796 22448
rect 7660 21568 7700 21608
rect 8044 24592 8084 24632
rect 8044 24256 8084 24296
rect 8428 27700 8468 27740
rect 8428 27196 8468 27236
rect 10060 31312 10100 31352
rect 9676 31228 9716 31268
rect 8812 30220 8852 30260
rect 8716 29968 8756 30008
rect 9676 30640 9716 30680
rect 9100 30052 9140 30092
rect 8716 29296 8756 29336
rect 8716 29128 8756 29168
rect 8620 29044 8660 29084
rect 9964 29884 10004 29924
rect 9100 29548 9140 29588
rect 10156 29128 10196 29168
rect 8716 28288 8756 28328
rect 8716 28120 8756 28160
rect 9292 28876 9332 28916
rect 10156 28288 10196 28328
rect 8908 27532 8948 27572
rect 8716 27448 8756 27488
rect 8620 27280 8660 27320
rect 10444 32824 10484 32864
rect 10828 32152 10868 32192
rect 10828 31732 10868 31772
rect 10444 31648 10484 31688
rect 11404 34168 11444 34208
rect 11212 33664 11252 33704
rect 11116 33076 11156 33116
rect 11116 32824 11156 32864
rect 11020 32152 11060 32192
rect 11020 31816 11060 31856
rect 12172 34420 12212 34460
rect 11980 34252 12020 34292
rect 12364 34168 12404 34208
rect 11692 34084 11732 34124
rect 11980 34084 12020 34124
rect 11788 33832 11828 33872
rect 11500 33328 11540 33368
rect 11212 31732 11252 31772
rect 11692 31900 11732 31940
rect 11692 31480 11732 31520
rect 10924 31312 10964 31352
rect 11020 30808 11060 30848
rect 10924 30640 10964 30680
rect 11116 30556 11156 30596
rect 10924 30388 10964 30428
rect 11500 30640 11540 30680
rect 11692 30640 11732 30680
rect 11404 30388 11444 30428
rect 11212 30304 11252 30344
rect 11116 30220 11156 30260
rect 11308 29968 11348 30008
rect 11308 29800 11348 29840
rect 11692 30304 11732 30344
rect 13132 34924 13172 34964
rect 13612 35260 13652 35300
rect 13228 34840 13268 34880
rect 13132 34588 13172 34628
rect 13228 34420 13268 34460
rect 12556 34252 12596 34292
rect 13036 34252 13076 34292
rect 12460 33832 12500 33872
rect 12364 31816 12404 31856
rect 12268 31732 12308 31772
rect 12172 31396 12212 31436
rect 11884 30808 11924 30848
rect 11884 30640 11924 30680
rect 11980 30472 12020 30512
rect 11884 30220 11924 30260
rect 11788 30136 11828 30176
rect 11788 29800 11828 29840
rect 12268 31312 12308 31352
rect 12172 30052 12212 30092
rect 12076 29800 12116 29840
rect 12268 29968 12308 30008
rect 13228 34000 13268 34040
rect 12940 33664 12980 33704
rect 12748 32908 12788 32948
rect 12652 32824 12692 32864
rect 12940 32656 12980 32696
rect 12460 31396 12500 31436
rect 12556 31228 12596 31268
rect 12556 29968 12596 30008
rect 12172 29128 12212 29168
rect 10348 28120 10388 28160
rect 8908 26944 8948 26984
rect 9292 26944 9332 26984
rect 9100 26440 9140 26480
rect 8524 26356 8564 26396
rect 9196 26272 9236 26312
rect 10060 26692 10100 26732
rect 9868 26272 9908 26312
rect 11404 27364 11444 27404
rect 11596 27364 11636 27404
rect 10540 26944 10580 26984
rect 10828 26776 10868 26816
rect 11020 26776 11060 26816
rect 10252 26104 10292 26144
rect 10924 26188 10964 26228
rect 9676 26020 9716 26060
rect 10156 26020 10196 26060
rect 9100 25264 9140 25304
rect 9292 24592 9332 24632
rect 8620 24004 8660 24044
rect 10060 25264 10100 25304
rect 11020 26020 11060 26060
rect 10444 25936 10484 25976
rect 10924 25936 10964 25976
rect 10060 24424 10100 24464
rect 10060 24004 10100 24044
rect 8620 23752 8660 23792
rect 8524 23668 8564 23708
rect 7948 22156 7988 22196
rect 8236 23164 8276 23204
rect 8332 23080 8372 23120
rect 8236 22996 8276 23036
rect 9772 23668 9812 23708
rect 10348 24844 10388 24884
rect 10252 24760 10292 24800
rect 11692 27196 11732 27236
rect 11308 26104 11348 26144
rect 11308 25348 11348 25388
rect 11116 25264 11156 25304
rect 11596 25264 11636 25304
rect 11308 25096 11348 25136
rect 11212 25012 11252 25052
rect 10828 24676 10868 24716
rect 10444 24424 10484 24464
rect 10156 23752 10196 23792
rect 10924 24592 10964 24632
rect 10732 24256 10772 24296
rect 11116 24004 11156 24044
rect 8620 23164 8660 23204
rect 9868 23164 9908 23204
rect 8716 22660 8756 22700
rect 8428 22576 8468 22616
rect 8140 22240 8180 22280
rect 8428 22156 8468 22196
rect 8140 21736 8180 21776
rect 9004 21736 9044 21776
rect 8044 21652 8084 21692
rect 6796 20224 6836 20264
rect 6988 19972 7028 20012
rect 7468 19972 7508 20012
rect 6796 19888 6836 19928
rect 8044 21400 8084 21440
rect 7948 20056 7988 20096
rect 7084 19888 7124 19928
rect 6892 19384 6932 19424
rect 4780 19132 4820 19172
rect 6028 19132 6068 19172
rect 4108 19048 4148 19088
rect 4204 18964 4244 19004
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4876 18544 4916 18584
rect 4396 17704 4436 17744
rect 4684 17872 4724 17912
rect 4012 17620 4052 17660
rect 3916 17452 3956 17492
rect 3820 17284 3860 17324
rect 3724 17200 3764 17240
rect 3340 16948 3380 16988
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4588 17536 4628 17576
rect 3820 16948 3860 16988
rect 4108 17116 4148 17156
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4972 17704 5012 17744
rect 4396 17200 4436 17240
rect 6316 18796 6356 18836
rect 7852 19132 7892 19172
rect 6988 18880 7028 18920
rect 7756 18880 7796 18920
rect 5164 17704 5204 17744
rect 5932 18124 5972 18164
rect 5260 17620 5300 17660
rect 5164 17536 5204 17576
rect 5068 17452 5108 17492
rect 4876 17200 4916 17240
rect 4204 17032 4244 17072
rect 4300 16864 4340 16904
rect 3628 16528 3668 16568
rect 4780 17032 4820 17072
rect 4684 16948 4724 16988
rect 4972 16864 5012 16904
rect 4684 16444 4724 16484
rect 844 15772 884 15812
rect 652 15688 692 15728
rect 940 15520 980 15560
rect 2860 16360 2900 16400
rect 3340 16360 3380 16400
rect 3628 16360 3668 16400
rect 4588 16360 4628 16400
rect 652 14848 692 14888
rect 1036 14092 1076 14132
rect 940 14008 980 14048
rect 3052 16192 3092 16232
rect 3148 16108 3188 16148
rect 3628 16108 3668 16148
rect 3244 15604 3284 15644
rect 4012 16192 4052 16232
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3628 15604 3668 15644
rect 3532 15520 3572 15560
rect 3340 15268 3380 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 2956 14848 2996 14888
rect 3436 14848 3476 14888
rect 2860 14680 2900 14720
rect 652 13168 692 13208
rect 2284 13168 2324 13208
rect 3244 14680 3284 14720
rect 3532 14680 3572 14720
rect 4012 15520 4052 15560
rect 4396 15604 4436 15644
rect 4492 15520 4532 15560
rect 3148 14092 3188 14132
rect 3724 14512 3764 14552
rect 4396 15100 4436 15140
rect 4012 14512 4052 14552
rect 3532 13840 3572 13880
rect 2860 12496 2900 12536
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 3628 12580 3668 12620
rect 3916 13840 3956 13880
rect 4300 14680 4340 14720
rect 4588 15352 4628 15392
rect 4684 15184 4724 15224
rect 4684 14932 4724 14972
rect 5164 16948 5204 16988
rect 5164 16780 5204 16820
rect 5356 17452 5396 17492
rect 6604 18124 6644 18164
rect 6700 17872 6740 17912
rect 5644 16780 5684 16820
rect 5452 16360 5492 16400
rect 5932 16444 5972 16484
rect 5644 16360 5684 16400
rect 5836 16192 5876 16232
rect 4972 15856 5012 15896
rect 5548 15856 5588 15896
rect 4972 15520 5012 15560
rect 5356 15520 5396 15560
rect 4876 15100 4916 15140
rect 4972 14932 5012 14972
rect 4780 14680 4820 14720
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4492 13168 4532 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 4204 12496 4244 12536
rect 5164 14512 5204 14552
rect 2956 12412 2996 12452
rect 3820 12412 3860 12452
rect 652 12328 692 12368
rect 4684 12496 4724 12536
rect 4972 12496 5012 12536
rect 5548 15184 5588 15224
rect 5452 15100 5492 15140
rect 5452 14596 5492 14636
rect 6124 15604 6164 15644
rect 6028 15184 6068 15224
rect 6412 16528 6452 16568
rect 6412 16192 6452 16232
rect 6508 16108 6548 16148
rect 6316 15520 6356 15560
rect 6604 15436 6644 15476
rect 7660 18796 7700 18836
rect 7948 18880 7988 18920
rect 9292 22660 9332 22700
rect 9964 23080 10004 23120
rect 11308 23752 11348 23792
rect 11404 23668 11444 23708
rect 11404 23332 11444 23372
rect 9388 22576 9428 22616
rect 9196 22240 9236 22280
rect 9388 22240 9428 22280
rect 10636 22660 10676 22700
rect 9772 22576 9812 22616
rect 8812 20560 8852 20600
rect 9292 20644 9332 20684
rect 10252 21652 10292 21692
rect 10348 21568 10388 21608
rect 11404 22492 11444 22532
rect 11020 22240 11060 22280
rect 10924 21736 10964 21776
rect 11596 21652 11636 21692
rect 11788 24592 11828 24632
rect 11980 27448 12020 27488
rect 11980 27028 12020 27068
rect 12268 27028 12308 27068
rect 12844 31480 12884 31520
rect 12748 31312 12788 31352
rect 13804 35092 13844 35132
rect 13708 35008 13748 35048
rect 13612 34252 13652 34292
rect 13612 34000 13652 34040
rect 13516 33076 13556 33116
rect 13996 35260 14036 35300
rect 14284 35176 14324 35216
rect 14572 35176 14612 35216
rect 14380 35092 14420 35132
rect 14092 34840 14132 34880
rect 14668 34840 14708 34880
rect 14860 34840 14900 34880
rect 14380 34756 14420 34796
rect 13900 34252 13940 34292
rect 13996 33664 14036 33704
rect 13804 33076 13844 33116
rect 13804 32824 13844 32864
rect 13996 32656 14036 32696
rect 13804 31900 13844 31940
rect 13420 31564 13460 31604
rect 13228 31480 13268 31520
rect 13708 31480 13748 31520
rect 13036 31396 13076 31436
rect 13324 31396 13364 31436
rect 13036 30976 13076 31016
rect 13612 31312 13652 31352
rect 13324 30808 13364 30848
rect 13132 30388 13172 30428
rect 13132 29884 13172 29924
rect 12844 29800 12884 29840
rect 13612 30976 13652 31016
rect 13516 30724 13556 30764
rect 13516 30304 13556 30344
rect 13420 30220 13460 30260
rect 13324 30136 13364 30176
rect 13612 30220 13652 30260
rect 13228 29632 13268 29672
rect 16300 35092 16340 35132
rect 16108 35008 16148 35048
rect 15436 34588 15476 34628
rect 14956 34504 14996 34544
rect 15820 34840 15860 34880
rect 14860 34252 14900 34292
rect 14764 34168 14804 34208
rect 14860 33412 14900 33452
rect 14380 32068 14420 32108
rect 13900 31228 13940 31268
rect 14092 30808 14132 30848
rect 13804 30640 13844 30680
rect 14188 30388 14228 30428
rect 13420 28456 13460 28496
rect 12748 28372 12788 28412
rect 13324 28372 13364 28412
rect 12844 27616 12884 27656
rect 13132 28288 13172 28328
rect 12652 27364 12692 27404
rect 12460 27196 12500 27236
rect 12460 26860 12500 26900
rect 12172 26776 12212 26816
rect 12556 26524 12596 26564
rect 13228 27196 13268 27236
rect 13036 26776 13076 26816
rect 12844 26692 12884 26732
rect 12652 26440 12692 26480
rect 12076 26104 12116 26144
rect 12268 25516 12308 25556
rect 12172 25096 12212 25136
rect 11980 24928 12020 24968
rect 11884 22492 11924 22532
rect 12364 25012 12404 25052
rect 12652 26104 12692 26144
rect 12556 25936 12596 25976
rect 12460 24928 12500 24968
rect 12076 23248 12116 23288
rect 12268 23584 12308 23624
rect 12844 25936 12884 25976
rect 13036 25852 13076 25892
rect 13036 25684 13076 25724
rect 12748 24592 12788 24632
rect 12460 23836 12500 23876
rect 12364 23332 12404 23372
rect 12940 25180 12980 25220
rect 12940 24340 12980 24380
rect 12844 23920 12884 23960
rect 12556 23752 12596 23792
rect 12940 23752 12980 23792
rect 12748 23584 12788 23624
rect 13132 25516 13172 25556
rect 13900 29884 13940 29924
rect 13996 29800 14036 29840
rect 13996 29128 14036 29168
rect 14764 32824 14804 32864
rect 15052 33076 15092 33116
rect 14956 32740 14996 32780
rect 14860 32656 14900 32696
rect 15244 33664 15284 33704
rect 15244 33412 15284 33452
rect 15340 33328 15380 33368
rect 15244 32824 15284 32864
rect 15628 34336 15668 34376
rect 15724 34252 15764 34292
rect 15436 32740 15476 32780
rect 15340 32152 15380 32192
rect 24460 36520 24500 36560
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 16492 35176 16532 35216
rect 18988 35848 19028 35888
rect 16780 35260 16820 35300
rect 16684 34924 16724 34964
rect 17164 35176 17204 35216
rect 17068 34840 17108 34880
rect 16972 34504 17012 34544
rect 16204 34336 16244 34376
rect 16588 34336 16628 34376
rect 16972 34336 17012 34376
rect 15916 33664 15956 33704
rect 18124 35176 18164 35216
rect 18316 35176 18356 35216
rect 17644 35092 17684 35132
rect 17452 35008 17492 35048
rect 17260 33748 17300 33788
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 18508 34588 18548 34628
rect 17740 34504 17780 34544
rect 18124 34420 18164 34460
rect 17932 33748 17972 33788
rect 16780 32908 16820 32948
rect 14764 31564 14804 31604
rect 14956 31480 14996 31520
rect 14476 30640 14516 30680
rect 14764 30220 14804 30260
rect 14668 29884 14708 29924
rect 14572 29800 14612 29840
rect 13900 28540 13940 28580
rect 14092 28540 14132 28580
rect 13804 28456 13844 28496
rect 13804 28288 13844 28328
rect 14092 28288 14132 28328
rect 14380 29212 14420 29252
rect 14284 29128 14324 29168
rect 15820 32068 15860 32108
rect 15916 31984 15956 32024
rect 15628 31480 15668 31520
rect 16108 32152 16148 32192
rect 15244 31312 15284 31352
rect 16012 31312 16052 31352
rect 16588 31984 16628 32024
rect 16492 31396 16532 31436
rect 16780 31648 16820 31688
rect 16684 31480 16724 31520
rect 16108 30724 16148 30764
rect 15820 29884 15860 29924
rect 15052 29800 15092 29840
rect 16300 30556 16340 30596
rect 16108 30388 16148 30428
rect 15052 29632 15092 29672
rect 14668 29128 14708 29168
rect 14476 28288 14516 28328
rect 13708 27616 13748 27656
rect 13612 27532 13652 27572
rect 14151 27616 14191 27656
rect 13900 27448 13940 27488
rect 13900 26860 13940 26900
rect 13324 25432 13364 25472
rect 13612 26104 13652 26144
rect 13612 25852 13652 25892
rect 13516 24844 13556 24884
rect 13420 24592 13460 24632
rect 14188 27196 14228 27236
rect 14284 27112 14324 27152
rect 14380 27028 14420 27068
rect 14380 26776 14420 26816
rect 13900 26608 13940 26648
rect 14284 26608 14324 26648
rect 14092 26440 14132 26480
rect 13900 25852 13940 25892
rect 13804 25432 13844 25472
rect 13804 25264 13844 25304
rect 13708 25180 13748 25220
rect 14188 26188 14228 26228
rect 14380 25936 14420 25976
rect 14284 25600 14324 25640
rect 14572 28120 14612 28160
rect 14764 27532 14804 27572
rect 14764 27364 14804 27404
rect 14668 27112 14708 27152
rect 14956 27616 14996 27656
rect 15340 29464 15380 29504
rect 16108 29212 16148 29252
rect 15436 29044 15476 29084
rect 16300 29128 16340 29168
rect 14860 27028 14900 27068
rect 14860 26776 14900 26816
rect 14668 26608 14708 26648
rect 14572 26524 14612 26564
rect 14668 26440 14708 26480
rect 14860 26608 14900 26648
rect 14860 26272 14900 26312
rect 15052 26692 15092 26732
rect 15052 26272 15092 26312
rect 15305 27364 15345 27404
rect 15244 27196 15284 27236
rect 15340 26776 15380 26816
rect 15244 26188 15284 26228
rect 14284 25432 14324 25472
rect 14764 25432 14804 25472
rect 14188 24928 14228 24968
rect 13708 24676 13748 24716
rect 13132 24340 13172 24380
rect 13900 24340 13940 24380
rect 13708 24004 13748 24044
rect 13612 23920 13652 23960
rect 12652 23248 12692 23288
rect 12556 23080 12596 23120
rect 12172 22660 12212 22700
rect 12364 22660 12404 22700
rect 12748 22660 12788 22700
rect 11884 21568 11924 21608
rect 9868 20728 9908 20768
rect 10348 20728 10388 20768
rect 9676 20644 9716 20684
rect 9004 20056 9044 20096
rect 9580 20560 9620 20600
rect 9292 20056 9332 20096
rect 10540 20560 10580 20600
rect 10156 19972 10196 20012
rect 9196 19888 9236 19928
rect 10348 19468 10388 19508
rect 8908 19300 8948 19340
rect 8332 19132 8372 19172
rect 6796 17032 6836 17072
rect 6796 16780 6836 16820
rect 6988 16360 7028 16400
rect 6988 16192 7028 16232
rect 7180 16192 7220 16232
rect 7852 17032 7892 17072
rect 7948 16780 7988 16820
rect 8140 17032 8180 17072
rect 10156 18880 10196 18920
rect 8428 18460 8468 18500
rect 8524 17536 8564 17576
rect 8428 16780 8468 16820
rect 8428 16444 8468 16484
rect 7852 16192 7892 16232
rect 7948 16108 7988 16148
rect 7852 15772 7892 15812
rect 7660 15692 7700 15728
rect 7660 15688 7700 15692
rect 8236 15688 8276 15728
rect 7852 15604 7892 15644
rect 8140 15604 8180 15644
rect 6412 15100 6452 15140
rect 5932 14848 5972 14888
rect 6220 14848 6260 14888
rect 6796 15184 6836 15224
rect 6604 14848 6644 14888
rect 5836 13840 5876 13880
rect 6028 13840 6068 13880
rect 5836 13168 5876 13208
rect 5836 12580 5876 12620
rect 5740 12496 5780 12536
rect 4492 12412 4532 12452
rect 5932 12496 5972 12536
rect 6892 15100 6932 15140
rect 7084 15016 7124 15056
rect 6508 13420 6548 13460
rect 6892 13420 6932 13460
rect 6796 13168 6836 13208
rect 8524 16192 8564 16232
rect 8716 17704 8756 17744
rect 10444 18796 10484 18836
rect 11500 20728 11540 20768
rect 10828 20644 10868 20684
rect 10828 20224 10868 20264
rect 11788 20224 11828 20264
rect 11308 20140 11348 20180
rect 10636 19468 10676 19508
rect 13612 23332 13652 23372
rect 13804 23332 13844 23372
rect 13516 23080 13556 23120
rect 12940 22324 12980 22364
rect 13420 22408 13460 22448
rect 13228 22324 13268 22364
rect 12940 21400 12980 21440
rect 13612 22660 13652 22700
rect 13708 22072 13748 22112
rect 14092 24592 14132 24632
rect 14476 25264 14516 25304
rect 14572 25132 14612 25136
rect 14572 25096 14612 25132
rect 14380 24676 14420 24716
rect 14188 24256 14228 24296
rect 14188 24088 14228 24128
rect 14092 23836 14132 23876
rect 13996 23668 14036 23708
rect 13996 23080 14036 23120
rect 13996 22408 14036 22448
rect 13900 21400 13940 21440
rect 13996 20812 14036 20852
rect 12940 20728 12980 20768
rect 12076 20056 12116 20096
rect 14284 23920 14324 23960
rect 14188 23584 14228 23624
rect 14284 22240 14324 22280
rect 14284 21568 14324 21608
rect 14476 24340 14516 24380
rect 14860 25264 14900 25304
rect 15052 25936 15092 25976
rect 16012 27616 16052 27656
rect 16012 27364 16052 27404
rect 17260 32908 17300 32948
rect 17644 31648 17684 31688
rect 17356 29884 17396 29924
rect 16588 28204 16628 28244
rect 16300 27616 16340 27656
rect 16492 27532 16532 27572
rect 16204 27196 16244 27236
rect 16780 27196 16820 27236
rect 17548 28204 17588 28244
rect 17452 27448 17492 27488
rect 17068 27196 17108 27236
rect 17356 27196 17396 27236
rect 16492 26692 16532 26732
rect 15628 26272 15668 26312
rect 15436 25516 15476 25556
rect 15244 25264 15284 25304
rect 15244 25096 15284 25136
rect 14860 24676 14900 24716
rect 14668 23920 14708 23960
rect 15052 24592 15092 24632
rect 16012 26356 16052 26396
rect 15916 26272 15956 26312
rect 16108 26104 16148 26144
rect 16108 25264 16148 25304
rect 16204 24844 16244 24884
rect 15244 24676 15284 24716
rect 14764 23836 14804 23876
rect 14668 23584 14708 23624
rect 14764 23500 14804 23540
rect 15052 24172 15092 24212
rect 15244 24088 15284 24128
rect 15340 24004 15380 24044
rect 15148 23836 15188 23876
rect 15052 23668 15092 23708
rect 15244 23584 15284 23624
rect 14956 23416 14996 23456
rect 15340 23416 15380 23456
rect 14860 23248 14900 23288
rect 15340 23164 15380 23204
rect 15148 22408 15188 22448
rect 15820 24592 15860 24632
rect 16012 24592 16052 24632
rect 16876 26440 16916 26480
rect 16588 25936 16628 25976
rect 17164 26440 17204 26480
rect 17260 26272 17300 26312
rect 17260 26020 17300 26060
rect 17740 31312 17780 31352
rect 18028 33664 18068 33704
rect 19564 35848 19604 35888
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 19276 34840 19316 34880
rect 18988 34351 19028 34376
rect 18988 34336 19028 34351
rect 19372 34504 19412 34544
rect 18892 34168 18932 34208
rect 18700 33748 18740 33788
rect 20044 34336 20084 34376
rect 19180 34168 19220 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 18124 32992 18164 33032
rect 18604 32908 18644 32948
rect 18892 33496 18932 33536
rect 18220 32824 18260 32864
rect 18124 32320 18164 32360
rect 19372 33748 19412 33788
rect 19660 33748 19700 33788
rect 19180 33664 19220 33704
rect 19180 33160 19220 33200
rect 19468 33328 19508 33368
rect 20332 33664 20372 33704
rect 21772 35344 21812 35384
rect 21196 35260 21236 35300
rect 23404 35260 23444 35300
rect 21196 34504 21236 34544
rect 21004 34336 21044 34376
rect 20044 33580 20084 33620
rect 19660 33076 19700 33116
rect 19372 32992 19412 33032
rect 19468 32824 19508 32864
rect 19756 32824 19796 32864
rect 20812 33580 20852 33620
rect 20332 33076 20372 33116
rect 20428 32824 20468 32864
rect 19372 32740 19412 32780
rect 18028 32152 18068 32192
rect 18412 32068 18452 32108
rect 17932 31984 17972 32024
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 18220 31312 18260 31352
rect 17836 30556 17876 30596
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 18700 30136 18740 30176
rect 18604 29968 18644 30008
rect 18796 29884 18836 29924
rect 18988 29884 19028 29924
rect 18700 29212 18740 29252
rect 18604 29128 18644 29168
rect 18892 29800 18932 29840
rect 20140 32740 20180 32780
rect 19564 32656 19604 32696
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 20044 32320 20084 32360
rect 19948 32152 19988 32192
rect 19372 31984 19412 32024
rect 19756 31480 19796 31520
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 19660 30640 19700 30680
rect 20332 31480 20372 31520
rect 20044 30640 20084 30680
rect 21292 34168 21332 34208
rect 21100 33664 21140 33704
rect 25900 36520 25940 36560
rect 25996 36436 26036 36476
rect 24076 35512 24116 35552
rect 25612 35512 25652 35552
rect 25804 35428 25844 35468
rect 25612 35344 25652 35384
rect 25420 34420 25460 34460
rect 22636 34336 22676 34376
rect 24556 34336 24596 34376
rect 23788 34168 23828 34208
rect 21580 33580 21620 33620
rect 21868 33664 21908 33704
rect 23596 33664 23636 33704
rect 24172 33664 24212 33704
rect 21484 33412 21524 33452
rect 21676 33412 21716 33452
rect 23212 33160 23252 33200
rect 21388 32992 21428 33032
rect 22156 32992 22196 33032
rect 21196 32320 21236 32360
rect 22540 32656 22580 32696
rect 21292 31984 21332 32024
rect 19468 29968 19508 30008
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 21196 30220 21236 30260
rect 21676 30220 21716 30260
rect 19660 29044 19700 29084
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 17932 28372 17972 28412
rect 18412 28288 18452 28328
rect 18988 28876 19028 28916
rect 18796 28204 18836 28244
rect 18700 28120 18740 28160
rect 20236 29128 20276 29168
rect 20140 28876 20180 28916
rect 20236 28792 20276 28832
rect 19756 28708 19796 28748
rect 19276 28456 19316 28496
rect 20812 29800 20852 29840
rect 20524 29296 20564 29336
rect 21100 29212 21140 29252
rect 22636 30304 22676 30344
rect 22348 30136 22388 30176
rect 23020 30052 23060 30092
rect 25036 34168 25076 34208
rect 25708 35092 25748 35132
rect 25516 34000 25556 34040
rect 25996 35344 26036 35384
rect 26092 35176 26132 35216
rect 25900 34336 25940 34376
rect 25996 34168 26036 34208
rect 26284 36688 26324 36728
rect 26380 35260 26420 35300
rect 27052 36436 27092 36476
rect 27628 37360 27668 37400
rect 27532 37192 27572 37232
rect 26860 35680 26900 35720
rect 28684 36688 28724 36728
rect 28972 36688 29012 36728
rect 29164 36100 29204 36140
rect 29452 36100 29492 36140
rect 28012 35680 28052 35720
rect 27724 35428 27764 35468
rect 26764 35176 26804 35216
rect 26476 35092 26516 35132
rect 26860 35092 26900 35132
rect 27052 35008 27092 35048
rect 26860 34504 26900 34544
rect 26284 34420 26324 34460
rect 27916 35008 27956 35048
rect 28300 35260 28340 35300
rect 28300 35008 28340 35048
rect 27532 34588 27572 34628
rect 28204 34588 28244 34628
rect 26188 34000 26228 34040
rect 26764 34000 26804 34040
rect 23692 33496 23732 33536
rect 24364 33496 24404 33536
rect 23788 33412 23828 33452
rect 28492 34420 28532 34460
rect 27916 34252 27956 34292
rect 26284 33412 26324 33452
rect 26956 33412 26996 33452
rect 25612 33160 25652 33200
rect 25612 32824 25652 32864
rect 23500 31564 23540 31604
rect 24844 32152 24884 32192
rect 24556 31480 24596 31520
rect 25228 31480 25268 31520
rect 24172 31144 24212 31184
rect 24748 31144 24788 31184
rect 25036 30808 25076 30848
rect 25420 30808 25460 30848
rect 24172 30640 24212 30680
rect 23884 30220 23924 30260
rect 25324 30136 25364 30176
rect 24364 30052 24404 30092
rect 21964 29296 22004 29336
rect 22924 29212 22964 29252
rect 21292 29044 21332 29084
rect 20428 28792 20468 28832
rect 20332 28624 20372 28664
rect 20716 28708 20756 28748
rect 19756 28288 19796 28328
rect 20236 28288 20276 28328
rect 20332 28204 20372 28244
rect 19276 28120 19316 28160
rect 20236 28120 20276 28160
rect 19180 28036 19220 28076
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 20524 28288 20564 28328
rect 21004 28204 21044 28244
rect 20716 28120 20756 28160
rect 19852 27700 19892 27740
rect 19564 27616 19604 27656
rect 18988 27364 19028 27404
rect 19372 27364 19412 27404
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 17740 27028 17780 27068
rect 18028 26944 18068 26984
rect 17548 26356 17588 26396
rect 18892 26692 18932 26732
rect 18700 26440 18740 26480
rect 18220 26188 18260 26228
rect 16684 25684 16724 25724
rect 16492 25348 16532 25388
rect 16972 25264 17012 25304
rect 16396 24760 16436 24800
rect 16396 24592 16436 24632
rect 15916 24424 15956 24464
rect 16684 24424 16724 24464
rect 15628 24088 15668 24128
rect 15532 23920 15572 23960
rect 16204 24004 16244 24044
rect 15724 23584 15764 23624
rect 15532 23416 15572 23456
rect 15628 23248 15668 23288
rect 16588 24004 16628 24044
rect 16396 23920 16436 23960
rect 16684 23836 16724 23876
rect 16780 23752 16820 23792
rect 17452 26020 17492 26060
rect 17452 25684 17492 25724
rect 17452 25348 17492 25388
rect 17740 26104 17780 26144
rect 18412 25936 18452 25976
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 17932 25348 17972 25388
rect 17548 25096 17588 25136
rect 17068 23920 17108 23960
rect 17356 23584 17396 23624
rect 16108 23416 16148 23456
rect 15436 22408 15476 22448
rect 15532 22240 15572 22280
rect 15724 23080 15764 23120
rect 16204 22240 16244 22280
rect 14668 20812 14708 20852
rect 12556 19972 12596 20012
rect 11308 19300 11348 19340
rect 10636 19216 10676 19256
rect 10828 19216 10868 19256
rect 10252 17704 10292 17744
rect 10540 18544 10580 18584
rect 10444 18460 10484 18500
rect 11788 19216 11828 19256
rect 11116 18628 11156 18668
rect 12076 19216 12116 19256
rect 12172 19048 12212 19088
rect 12268 18712 12308 18752
rect 11980 18628 12020 18668
rect 10636 18460 10676 18500
rect 11116 18460 11156 18500
rect 11212 18376 11252 18416
rect 10348 17536 10388 17576
rect 9388 17032 9428 17072
rect 8332 15520 8372 15560
rect 11308 17956 11348 17996
rect 11212 17536 11252 17576
rect 11596 18544 11636 18584
rect 13132 19048 13172 19088
rect 13324 18796 13364 18836
rect 11212 16360 11252 16400
rect 11692 16276 11732 16316
rect 8620 15688 8660 15728
rect 7948 15436 7988 15476
rect 8044 15016 8084 15056
rect 7948 14932 7988 14972
rect 7564 14176 7604 14216
rect 8524 15436 8564 15476
rect 8716 15520 8756 15560
rect 9100 15520 9140 15560
rect 8812 14848 8852 14888
rect 9100 14932 9140 14972
rect 9100 14680 9140 14720
rect 8140 14512 8180 14552
rect 8716 14176 8756 14216
rect 10540 15688 10580 15728
rect 9676 15520 9716 15560
rect 10156 15520 10196 15560
rect 10924 16192 10964 16232
rect 12268 17956 12308 17996
rect 12364 17704 12404 17744
rect 12940 18376 12980 18416
rect 12556 17704 12596 17744
rect 14476 19972 14516 20012
rect 13996 18460 14036 18500
rect 14188 18376 14228 18416
rect 13804 17704 13844 17744
rect 14188 17704 14228 17744
rect 12652 17620 12692 17660
rect 13612 17620 13652 17660
rect 14092 17620 14132 17660
rect 12940 16780 12980 16820
rect 12364 16192 12404 16232
rect 12748 16192 12788 16232
rect 9964 14932 10004 14972
rect 9580 14092 9620 14132
rect 7276 13420 7316 13460
rect 6412 12580 6452 12620
rect 7084 12496 7124 12536
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 6028 11656 6068 11696
rect 6988 12328 7028 12368
rect 8428 13252 8468 13292
rect 8620 12496 8660 12536
rect 8332 12412 8372 12452
rect 652 11488 692 11528
rect 7276 11404 7316 11444
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8044 11908 8084 11948
rect 8428 11908 8468 11948
rect 7660 11656 7700 11696
rect 7468 10984 7508 11024
rect 7276 10732 7316 10772
rect 7852 10732 7892 10772
rect 652 10648 692 10688
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 5548 10060 5588 10100
rect 652 9808 692 9848
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 7660 10144 7700 10184
rect 6988 10060 7028 10100
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 652 8968 692 9008
rect 3436 8800 3476 8840
rect 6124 8800 6164 8840
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 556 8128 596 8168
rect 4684 7960 4724 8000
rect 5932 8632 5972 8672
rect 4876 8044 4916 8084
rect 5164 7960 5204 8000
rect 5452 8044 5492 8084
rect 6220 8632 6260 8672
rect 2380 7708 2420 7748
rect 652 7288 692 7328
rect 3820 7708 3860 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4780 7456 4820 7496
rect 3628 7120 3668 7160
rect 4972 7792 5012 7832
rect 5356 7792 5396 7832
rect 5164 7456 5204 7496
rect 4972 7120 5012 7160
rect 5452 7372 5492 7412
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 652 6448 692 6488
rect 3724 6448 3764 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4876 6448 4916 6488
rect 4684 5776 4724 5816
rect 652 5608 692 5648
rect 4588 5608 4628 5648
rect 4396 5440 4436 5480
rect 4684 5440 4724 5480
rect 4204 5356 4244 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 4396 4936 4436 4976
rect 652 4768 692 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 3340 4180 3380 4220
rect 4492 4768 4532 4808
rect 4588 4348 4628 4388
rect 4684 4180 4724 4220
rect 5644 6364 5684 6404
rect 5548 5776 5588 5816
rect 5356 4768 5396 4808
rect 5932 7792 5972 7832
rect 6220 7876 6260 7916
rect 6700 8128 6740 8168
rect 5836 7540 5876 7580
rect 5836 7372 5876 7412
rect 6316 7792 6356 7832
rect 6220 7540 6260 7580
rect 6796 7540 6836 7580
rect 7948 9388 7988 9428
rect 7756 8212 7796 8252
rect 7372 7540 7412 7580
rect 6508 7120 6548 7160
rect 5836 6364 5876 6404
rect 5836 5692 5876 5732
rect 5740 5356 5780 5396
rect 6316 6784 6356 6824
rect 6220 6532 6260 6572
rect 6412 6475 6452 6488
rect 6412 6448 6452 6475
rect 7564 7960 7604 8000
rect 7660 7876 7700 7916
rect 7756 7708 7796 7748
rect 7660 7624 7700 7664
rect 7468 7456 7508 7496
rect 7468 7120 7508 7160
rect 7948 8632 7988 8672
rect 8428 11320 8468 11360
rect 8524 9976 8564 10016
rect 8140 9472 8180 9512
rect 8332 8212 8372 8252
rect 8236 8128 8276 8168
rect 8140 7372 8180 7412
rect 7756 6784 7796 6824
rect 7564 6364 7604 6404
rect 8428 7456 8468 7496
rect 7852 6448 7892 6488
rect 6028 6280 6068 6320
rect 7084 6280 7124 6320
rect 7660 6280 7700 6320
rect 5932 5020 5972 5060
rect 6220 5860 6260 5900
rect 6124 5608 6164 5648
rect 6124 5356 6164 5396
rect 6412 5440 6452 5480
rect 6220 4936 6260 4976
rect 5836 4180 5876 4220
rect 4588 4096 4628 4136
rect 4972 4096 5012 4136
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 652 3088 692 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 5836 2752 5876 2792
rect 652 2248 692 2288
rect 5452 2668 5492 2708
rect 6124 4180 6164 4220
rect 6316 4180 6356 4220
rect 6124 2668 6164 2708
rect 7372 6196 7412 6236
rect 7948 6196 7988 6236
rect 6796 5020 6836 5060
rect 7180 5440 7220 5480
rect 7468 5440 7508 5480
rect 6988 4180 7028 4220
rect 7180 5020 7220 5060
rect 6700 4096 6740 4136
rect 7084 4096 7124 4136
rect 6508 4012 6548 4052
rect 7372 4264 7412 4304
rect 7276 4096 7316 4136
rect 7948 5692 7988 5732
rect 8620 6952 8660 6992
rect 8428 6868 8468 6908
rect 10540 14008 10580 14048
rect 10828 14008 10868 14048
rect 11212 14008 11252 14048
rect 11212 13252 11252 13292
rect 8812 13168 8852 13208
rect 8812 12580 8852 12620
rect 9292 11908 9332 11948
rect 9292 10984 9332 11024
rect 9676 12412 9716 12452
rect 9580 12328 9620 12368
rect 8908 8464 8948 8504
rect 8908 7708 8948 7748
rect 8716 6784 8756 6824
rect 8332 6700 8372 6740
rect 8236 6280 8276 6320
rect 9484 10144 9524 10184
rect 9772 11236 9812 11276
rect 10060 11656 10100 11696
rect 9676 10144 9716 10184
rect 9388 9472 9428 9512
rect 9580 9472 9620 9512
rect 10156 10396 10196 10436
rect 9964 10312 10004 10352
rect 11788 14008 11828 14048
rect 11596 13840 11636 13880
rect 11980 13840 12020 13880
rect 11404 12580 11444 12620
rect 12268 13252 12308 13292
rect 11788 12244 11828 12284
rect 11980 11656 12020 11696
rect 10348 10984 10388 11024
rect 11020 10984 11060 11024
rect 10156 10060 10196 10100
rect 9100 9388 9140 9428
rect 9292 9388 9332 9428
rect 9964 9472 10004 9512
rect 10348 9976 10388 10016
rect 11692 11236 11732 11276
rect 11212 10732 11252 10772
rect 11308 10312 11348 10352
rect 10444 9472 10484 9512
rect 11500 10816 11540 10856
rect 11404 10060 11444 10100
rect 11308 9640 11348 9680
rect 9868 9388 9908 9428
rect 11212 9472 11252 9512
rect 11116 9388 11156 9428
rect 11020 9220 11060 9260
rect 9868 8884 9908 8924
rect 10348 8884 10388 8924
rect 10636 8800 10676 8840
rect 9388 8212 9428 8252
rect 9196 7960 9236 8000
rect 9196 7708 9236 7748
rect 9100 7372 9140 7412
rect 9868 7624 9908 7664
rect 9004 7120 9044 7160
rect 9100 6952 9140 6992
rect 8428 6616 8468 6656
rect 8524 6448 8564 6488
rect 8428 5608 8468 5648
rect 8812 6616 8852 6656
rect 9388 6784 9428 6824
rect 9292 6532 9332 6572
rect 9004 6448 9044 6488
rect 9772 6700 9812 6740
rect 9964 7540 10004 7580
rect 10732 8632 10772 8672
rect 10540 8464 10580 8504
rect 10252 7708 10292 7748
rect 10444 7708 10484 7748
rect 10732 7624 10772 7664
rect 10348 7540 10388 7580
rect 10636 7540 10676 7580
rect 10060 6784 10100 6824
rect 9964 6700 10004 6740
rect 9484 6616 9524 6656
rect 9868 6616 9908 6656
rect 9772 6532 9812 6572
rect 9484 6448 9524 6488
rect 8908 6280 8948 6320
rect 9196 6280 9236 6320
rect 9868 6280 9908 6320
rect 7756 5020 7796 5060
rect 7564 4348 7604 4388
rect 6892 2752 6932 2792
rect 7852 4264 7892 4304
rect 8524 4264 8564 4304
rect 7660 3760 7700 3800
rect 7948 3760 7988 3800
rect 7852 3340 7892 3380
rect 8140 4096 8180 4136
rect 8236 2752 8276 2792
rect 8044 2584 8084 2624
rect 8428 2584 8468 2624
rect 10060 5692 10100 5732
rect 9580 5104 9620 5144
rect 9676 5020 9716 5060
rect 9964 4936 10004 4976
rect 9388 4264 9428 4304
rect 10348 6616 10388 6656
rect 10348 6280 10388 6320
rect 10540 6448 10580 6488
rect 10924 7120 10964 7160
rect 11788 10060 11828 10100
rect 11692 9472 11732 9512
rect 12652 11908 12692 11948
rect 12460 11656 12500 11696
rect 12364 10732 12404 10772
rect 12556 10312 12596 10352
rect 12652 10228 12692 10268
rect 12076 9640 12116 9680
rect 11596 9388 11636 9428
rect 12652 9304 12692 9344
rect 11980 9220 12020 9260
rect 11692 8884 11732 8924
rect 13228 16192 13268 16232
rect 15148 20728 15188 20768
rect 15340 20644 15380 20684
rect 14860 19468 14900 19508
rect 15244 20308 15284 20348
rect 15148 19468 15188 19508
rect 14956 18712 14996 18752
rect 15052 18544 15092 18584
rect 14956 18460 14996 18500
rect 15436 20560 15476 20600
rect 15628 20728 15668 20768
rect 15436 20056 15476 20096
rect 15916 20644 15956 20684
rect 15820 20056 15860 20096
rect 15724 19384 15764 19424
rect 16972 23500 17012 23540
rect 17740 25264 17780 25304
rect 18028 25180 18068 25220
rect 18220 25180 18260 25220
rect 17836 25096 17876 25136
rect 17836 24592 17876 24632
rect 17644 24508 17684 24548
rect 17548 23836 17588 23876
rect 17740 23584 17780 23624
rect 17452 23080 17492 23120
rect 18508 25096 18548 25136
rect 19084 26692 19124 26732
rect 18796 26020 18836 26060
rect 18796 25348 18836 25388
rect 20236 27196 20276 27236
rect 19276 26776 19316 26816
rect 19660 26776 19700 26816
rect 19276 26440 19316 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 19372 26272 19412 26312
rect 19276 26188 19316 26228
rect 20620 27532 20660 27572
rect 19468 26104 19508 26144
rect 19372 26020 19412 26060
rect 19084 25684 19124 25724
rect 19372 25684 19412 25724
rect 19372 25348 19412 25388
rect 20332 26104 20372 26144
rect 21004 27448 21044 27488
rect 21196 27364 21236 27404
rect 20908 26188 20948 26228
rect 21100 26188 21140 26228
rect 20332 25852 20372 25892
rect 20524 25264 20564 25304
rect 19660 25096 19700 25136
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 19180 24004 19220 24044
rect 19084 23920 19124 23960
rect 16972 22492 17012 22532
rect 17644 22408 17684 22448
rect 16780 22072 16820 22112
rect 16876 21568 16916 21608
rect 17068 22072 17108 22112
rect 16684 20728 16724 20768
rect 17260 21652 17300 21692
rect 17836 21652 17876 21692
rect 17260 20812 17300 20852
rect 16876 20644 16916 20684
rect 16396 20560 16436 20600
rect 16300 20056 16340 20096
rect 16300 19468 16340 19508
rect 16300 19216 16340 19256
rect 15628 19048 15668 19088
rect 16684 20056 16724 20096
rect 19660 23836 19700 23876
rect 20044 23836 20084 23876
rect 19276 23752 19316 23792
rect 19756 23752 19796 23792
rect 19660 23584 19700 23624
rect 19276 23416 19316 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 18508 22408 18548 22448
rect 18124 22324 18164 22364
rect 18220 22240 18260 22280
rect 18028 22072 18068 22112
rect 18316 21568 18356 21608
rect 19180 22492 19220 22532
rect 19756 23248 19796 23288
rect 19372 23080 19412 23120
rect 18892 22156 18932 22196
rect 18700 21400 18740 21440
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 22732 28120 22772 28160
rect 21868 27448 21908 27488
rect 21964 26776 22004 26816
rect 21676 26440 21716 26480
rect 22060 26440 22100 26480
rect 26092 32992 26132 33032
rect 25996 32824 26036 32864
rect 26188 32908 26228 32948
rect 26860 32908 26900 32948
rect 25708 32740 25748 32780
rect 26380 32740 26420 32780
rect 25708 31312 25748 31352
rect 25996 32152 26036 32192
rect 26380 32152 26420 32192
rect 26188 31228 26228 31268
rect 26092 31060 26132 31100
rect 25708 30640 25748 30680
rect 25612 30388 25652 30428
rect 25516 29212 25556 29252
rect 25996 30220 26036 30260
rect 26380 31312 26420 31352
rect 26380 31144 26420 31184
rect 26860 31144 26900 31184
rect 26284 30136 26324 30176
rect 25804 29128 25844 29168
rect 26284 29128 26324 29168
rect 27436 33076 27476 33116
rect 27724 33664 27764 33704
rect 27628 33580 27668 33620
rect 27820 33580 27860 33620
rect 27532 32908 27572 32948
rect 27148 32488 27188 32528
rect 27052 31312 27092 31352
rect 26956 30640 26996 30680
rect 26476 30388 26516 30428
rect 26572 29716 26612 29756
rect 26572 29128 26612 29168
rect 26476 28876 26516 28916
rect 25324 28288 25364 28328
rect 23404 27700 23444 27740
rect 24268 27700 24308 27740
rect 24460 27700 24500 27740
rect 23212 27196 23252 27236
rect 23116 26440 23156 26480
rect 22732 26356 22772 26396
rect 21772 25852 21812 25892
rect 22348 26104 22388 26144
rect 22924 26104 22964 26144
rect 22828 26020 22868 26060
rect 22828 25348 22868 25388
rect 22060 25264 22100 25304
rect 22444 24592 22484 24632
rect 22252 24508 22292 24548
rect 20620 23836 20660 23876
rect 20620 23080 20660 23120
rect 19948 22240 19988 22280
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 20236 21400 20276 21440
rect 18988 20728 19028 20768
rect 18124 20644 18164 20684
rect 18892 20224 18932 20264
rect 17452 19468 17492 19508
rect 17932 19384 17972 19424
rect 18892 19972 18932 20012
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 17644 19048 17684 19088
rect 18028 19048 18068 19088
rect 15628 18544 15668 18584
rect 14668 17620 14708 17660
rect 14380 16864 14420 16904
rect 14572 16780 14612 16820
rect 15436 16948 15476 16988
rect 15244 16360 15284 16400
rect 15340 15856 15380 15896
rect 17740 17704 17780 17744
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 15916 17620 15956 17660
rect 16780 17620 16820 17660
rect 16684 17032 16724 17072
rect 15724 16192 15764 16232
rect 14188 15100 14228 15140
rect 15052 14848 15092 14888
rect 13420 14176 13460 14216
rect 13036 14092 13076 14132
rect 13324 14008 13364 14048
rect 12844 13840 12884 13880
rect 13036 13504 13076 13544
rect 13324 13168 13364 13208
rect 13132 13084 13172 13124
rect 13228 13000 13268 13040
rect 13516 14092 13556 14132
rect 12844 11656 12884 11696
rect 13900 14176 13940 14216
rect 13804 14092 13844 14132
rect 13804 13840 13844 13880
rect 13900 13756 13940 13796
rect 13996 13588 14036 13628
rect 14092 13504 14132 13544
rect 14380 13924 14420 13964
rect 14284 13840 14324 13880
rect 14188 13252 14228 13292
rect 15148 14680 15188 14720
rect 14572 13756 14612 13796
rect 14476 13504 14516 13544
rect 14380 13168 14420 13208
rect 14764 14008 14804 14048
rect 14956 14008 14996 14048
rect 15340 14512 15380 14552
rect 15244 13924 15284 13964
rect 15052 13840 15092 13880
rect 14860 13756 14900 13796
rect 14764 13588 14804 13628
rect 14668 13252 14708 13292
rect 13804 13000 13844 13040
rect 14284 13084 14324 13124
rect 14092 12832 14132 12872
rect 13996 12580 14036 12620
rect 14188 12496 14228 12536
rect 14476 13000 14516 13040
rect 14476 12748 14516 12788
rect 14380 12496 14420 12536
rect 13708 11908 13748 11948
rect 14380 12244 14420 12284
rect 14764 12916 14804 12956
rect 14956 12916 14996 12956
rect 14860 12748 14900 12788
rect 14956 12664 14996 12704
rect 15628 14176 15668 14216
rect 16012 15520 16052 15560
rect 15820 15436 15860 15476
rect 15916 14680 15956 14720
rect 15724 14008 15764 14048
rect 15532 13924 15572 13964
rect 15436 13336 15476 13376
rect 15244 13168 15284 13208
rect 15244 13000 15284 13040
rect 15148 12916 15188 12956
rect 15148 12748 15188 12788
rect 14668 12412 14708 12452
rect 14764 12328 14804 12368
rect 13996 11908 14036 11948
rect 13516 11488 13556 11528
rect 13900 11488 13940 11528
rect 13612 10816 13652 10856
rect 14572 11404 14612 11444
rect 15052 12496 15092 12536
rect 14956 12412 14996 12452
rect 15532 13168 15572 13208
rect 15820 13840 15860 13880
rect 15724 12916 15764 12956
rect 15628 12832 15668 12872
rect 15340 12664 15380 12704
rect 15724 12664 15764 12704
rect 15340 12496 15380 12536
rect 14956 11824 14996 11864
rect 14860 11656 14900 11696
rect 15340 11656 15380 11696
rect 15244 11488 15284 11528
rect 15148 11320 15188 11360
rect 15340 11320 15380 11360
rect 15052 11068 15092 11108
rect 13516 10396 13556 10436
rect 13420 9640 13460 9680
rect 12844 9304 12884 9344
rect 12268 8632 12308 8672
rect 12748 8632 12788 8672
rect 11212 7624 11252 7664
rect 11404 7120 11444 7160
rect 11596 6952 11636 6992
rect 11308 6868 11348 6908
rect 13516 9472 13556 9512
rect 14092 9976 14132 10016
rect 13900 9640 13940 9680
rect 13804 9556 13844 9596
rect 13420 9388 13460 9428
rect 13132 9304 13172 9344
rect 13996 9472 14036 9512
rect 15244 10900 15284 10940
rect 15052 10060 15092 10100
rect 15724 12496 15764 12536
rect 16300 15436 16340 15476
rect 16492 16360 16532 16400
rect 16492 16192 16532 16232
rect 16684 16192 16724 16232
rect 20812 20728 20852 20768
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 19660 20224 19700 20264
rect 19276 20056 19316 20096
rect 19372 19972 19412 20012
rect 19468 19888 19508 19928
rect 19276 19384 19316 19424
rect 21100 20560 21140 20600
rect 20908 20056 20948 20096
rect 19564 19300 19604 19340
rect 20716 19300 20756 19340
rect 19372 19216 19412 19256
rect 20812 19216 20852 19256
rect 21004 19216 21044 19256
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 21004 18880 21044 18920
rect 20908 18796 20948 18836
rect 20236 18544 20276 18584
rect 20140 17956 20180 17996
rect 18892 17620 18932 17660
rect 17932 17116 17972 17156
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 19372 17116 19412 17156
rect 18988 17032 19028 17072
rect 24268 27112 24308 27152
rect 24268 26944 24308 26984
rect 25132 27364 25172 27404
rect 24844 27280 24884 27320
rect 24748 27196 24788 27236
rect 24652 27112 24692 27152
rect 24748 27028 24788 27068
rect 24940 26944 24980 26984
rect 23884 26692 23924 26732
rect 24364 26692 24404 26732
rect 23308 26188 23348 26228
rect 23692 25516 23732 25556
rect 23596 25432 23636 25472
rect 24748 26608 24788 26648
rect 24940 26440 24980 26480
rect 26572 28624 26612 28664
rect 26764 28876 26804 28916
rect 26860 28624 26900 28664
rect 26668 28204 26708 28244
rect 26092 28036 26132 28076
rect 26284 28036 26324 28076
rect 26092 27616 26132 27656
rect 24556 26356 24596 26396
rect 25420 26356 25460 26396
rect 23788 24844 23828 24884
rect 23212 24088 23252 24128
rect 24268 26020 24308 26060
rect 25132 26104 25172 26144
rect 24844 25852 24884 25892
rect 25516 25516 25556 25556
rect 25900 26440 25940 26480
rect 27244 32320 27284 32360
rect 27340 31480 27380 31520
rect 27724 33076 27764 33116
rect 27820 32824 27860 32864
rect 27628 32656 27668 32696
rect 27820 32656 27860 32696
rect 27532 32488 27572 32528
rect 28588 34000 28628 34040
rect 28012 33664 28052 33704
rect 28588 33076 28628 33116
rect 28396 32992 28436 33032
rect 27916 32488 27956 32528
rect 28108 32656 28148 32696
rect 28012 32320 28052 32360
rect 27820 32152 27860 32192
rect 27628 31564 27668 31604
rect 27820 31480 27860 31520
rect 28012 31480 28052 31520
rect 28492 32824 28532 32864
rect 28684 32992 28724 33032
rect 27340 31144 27380 31184
rect 27916 31144 27956 31184
rect 27628 30808 27668 30848
rect 27724 30724 27764 30764
rect 27148 30304 27188 30344
rect 27244 29380 27284 29420
rect 27436 29296 27476 29336
rect 27244 29128 27284 29168
rect 28300 31312 28340 31352
rect 28396 31228 28436 31268
rect 27916 29716 27956 29756
rect 27628 29548 27668 29588
rect 27532 29128 27572 29168
rect 27436 29044 27476 29084
rect 27916 29212 27956 29252
rect 27916 28960 27956 29000
rect 28204 29380 28244 29420
rect 28108 29296 28148 29336
rect 28204 29212 28244 29252
rect 27724 28288 27764 28328
rect 26956 28204 26996 28244
rect 27724 27952 27764 27992
rect 26764 27616 26804 27656
rect 30796 36100 30836 36140
rect 31756 37360 31796 37400
rect 30988 36856 31028 36896
rect 31660 36856 31700 36896
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 32716 36772 32756 36812
rect 33292 36772 33332 36812
rect 31372 36520 31412 36560
rect 32044 36520 32084 36560
rect 30604 35680 30644 35720
rect 29740 35344 29780 35384
rect 30508 35344 30548 35384
rect 29836 35176 29876 35216
rect 30412 35176 30452 35216
rect 30124 35092 30164 35132
rect 29164 34588 29204 34628
rect 29452 34000 29492 34040
rect 29068 33916 29108 33956
rect 29644 35008 29684 35048
rect 29836 34420 29876 34460
rect 29932 34168 29972 34208
rect 30220 34504 30260 34544
rect 30028 33916 30068 33956
rect 29068 33496 29108 33536
rect 29164 32908 29204 32948
rect 29068 32824 29108 32864
rect 29356 32824 29396 32864
rect 28588 31480 28628 31520
rect 28588 30808 28628 30848
rect 28492 30388 28532 30428
rect 28396 30304 28436 30344
rect 28396 29128 28436 29168
rect 28780 29800 28820 29840
rect 29164 30304 29204 30344
rect 28684 29296 28724 29336
rect 28972 29296 29012 29336
rect 28684 29128 28724 29168
rect 28588 29044 28628 29084
rect 30892 35260 30932 35300
rect 30508 34840 30548 34880
rect 30412 34000 30452 34040
rect 30412 33580 30452 33620
rect 30316 33244 30356 33284
rect 30316 33076 30356 33116
rect 29548 32824 29588 32864
rect 30220 32824 30260 32864
rect 29548 30808 29588 30848
rect 29452 30220 29492 30260
rect 29260 29800 29300 29840
rect 30028 30640 30068 30680
rect 30316 30472 30356 30512
rect 29932 30388 29972 30428
rect 30892 34924 30932 34964
rect 30700 34420 30740 34460
rect 30988 34252 31028 34292
rect 30700 34168 30740 34208
rect 30604 33664 30644 33704
rect 30700 33076 30740 33116
rect 30508 32236 30548 32276
rect 30124 30220 30164 30260
rect 30124 29548 30164 29588
rect 29740 29296 29780 29336
rect 29932 29212 29972 29252
rect 30316 29296 30356 29336
rect 29260 29044 29300 29084
rect 30412 29128 30452 29168
rect 28588 28288 28628 28328
rect 29644 28456 29684 28496
rect 28876 28372 28916 28412
rect 28972 28204 29012 28244
rect 28012 27448 28052 27488
rect 27148 27364 27188 27404
rect 27724 27364 27764 27404
rect 26668 26524 26708 26564
rect 26380 26188 26420 26228
rect 25996 26104 26036 26144
rect 25804 25936 25844 25976
rect 26284 25852 26324 25892
rect 26956 25852 26996 25892
rect 26860 25432 26900 25472
rect 26380 25264 26420 25304
rect 25324 25180 25364 25220
rect 25132 24760 25172 24800
rect 25804 24760 25844 24800
rect 24556 24172 24596 24212
rect 22924 23752 22964 23792
rect 23308 23752 23348 23792
rect 22732 23668 22772 23708
rect 23500 23752 23540 23792
rect 23884 23752 23924 23792
rect 24076 23752 24116 23792
rect 24652 23752 24692 23792
rect 23212 23500 23252 23540
rect 23404 23668 23444 23708
rect 23404 23500 23444 23540
rect 23884 23080 23924 23120
rect 23308 22744 23348 22784
rect 23596 22744 23636 22784
rect 21292 21400 21332 21440
rect 22444 21400 22484 21440
rect 21292 20812 21332 20852
rect 22156 20812 22196 20852
rect 22348 20728 22388 20768
rect 21484 20560 21524 20600
rect 21676 20560 21716 20600
rect 21868 20140 21908 20180
rect 21772 19972 21812 20012
rect 22060 20140 22100 20180
rect 21964 20056 22004 20096
rect 21964 19888 22004 19928
rect 21868 19720 21908 19760
rect 21004 18544 21044 18584
rect 21196 18544 21236 18584
rect 20812 17704 20852 17744
rect 20812 17200 20852 17240
rect 18316 16948 18356 16988
rect 18796 16948 18836 16988
rect 17548 16864 17588 16904
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 17548 16192 17588 16232
rect 16780 15856 16820 15896
rect 16684 15520 16724 15560
rect 16972 15268 17012 15308
rect 16780 15184 16820 15224
rect 16396 15100 16436 15140
rect 18700 16192 18740 16232
rect 18508 15688 18548 15728
rect 18700 15520 18740 15560
rect 18892 16360 18932 16400
rect 20716 17032 20756 17072
rect 20908 17032 20948 17072
rect 21964 19468 22004 19508
rect 21868 18880 21908 18920
rect 21676 18544 21716 18584
rect 21868 18460 21908 18500
rect 21388 17956 21428 17996
rect 21484 17872 21524 17912
rect 19276 16360 19316 16400
rect 20140 16360 20180 16400
rect 20332 16360 20372 16400
rect 18988 16276 19028 16316
rect 19084 16192 19124 16232
rect 19180 16108 19220 16148
rect 19180 15520 19220 15560
rect 19660 16192 19700 16232
rect 19372 16108 19412 16148
rect 19852 16108 19892 16148
rect 20229 16192 20269 16232
rect 20332 16192 20372 16232
rect 19948 16024 19988 16064
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 19372 15688 19412 15728
rect 19564 15520 19604 15560
rect 20140 15940 20180 15980
rect 20524 16276 20564 16316
rect 20428 16108 20468 16148
rect 20716 16192 20756 16232
rect 20812 16024 20852 16064
rect 20620 15856 20660 15896
rect 20236 15688 20276 15728
rect 21196 16192 21236 16232
rect 21004 15856 21044 15896
rect 21292 15772 21332 15812
rect 22156 19384 22196 19424
rect 22444 20056 22484 20096
rect 22636 20560 22676 20600
rect 23116 22324 23156 22364
rect 23500 22492 23540 22532
rect 23788 22660 23828 22700
rect 23884 22576 23924 22616
rect 23692 22240 23732 22280
rect 23404 21400 23444 21440
rect 24844 23668 24884 23708
rect 24172 23584 24212 23624
rect 24076 22660 24116 22700
rect 24556 23332 24596 23372
rect 24460 23080 24500 23120
rect 24748 23080 24788 23120
rect 24556 22744 24596 22784
rect 24460 22492 24500 22532
rect 24556 22408 24596 22448
rect 24748 22828 24788 22868
rect 24364 22324 24404 22364
rect 24652 22156 24692 22196
rect 25036 23584 25076 23624
rect 25324 23752 25364 23792
rect 25036 23332 25076 23372
rect 25228 23332 25268 23372
rect 25804 24172 25844 24212
rect 25708 23752 25748 23792
rect 25420 23332 25460 23372
rect 25132 22996 25172 23036
rect 25324 22996 25364 23036
rect 25036 22912 25076 22952
rect 24748 22072 24788 22112
rect 24076 21568 24116 21608
rect 22540 19468 22580 19508
rect 22636 19384 22676 19424
rect 24364 21652 24404 21692
rect 26860 23920 26900 23960
rect 26668 23836 26708 23876
rect 25612 23164 25652 23204
rect 25900 22912 25940 22952
rect 25612 22660 25652 22700
rect 25132 22492 25172 22532
rect 25132 22324 25172 22364
rect 25036 22072 25076 22112
rect 25036 21652 25076 21692
rect 24460 21400 24500 21440
rect 22828 19300 22868 19340
rect 22540 19216 22580 19256
rect 23404 20056 23444 20096
rect 25036 21400 25076 21440
rect 25420 22240 25460 22280
rect 26092 23752 26132 23792
rect 26188 23584 26228 23624
rect 26092 23248 26132 23288
rect 26092 23080 26132 23120
rect 26284 23332 26324 23372
rect 26572 23668 26612 23708
rect 26476 23500 26516 23540
rect 26092 22660 26132 22700
rect 26284 22996 26324 23036
rect 26380 22828 26420 22868
rect 26764 23164 26804 23204
rect 26668 22912 26708 22952
rect 26572 22240 26612 22280
rect 26188 22156 26228 22196
rect 26476 22156 26516 22196
rect 25228 22072 25268 22112
rect 25996 22072 26036 22112
rect 25420 21988 25460 22028
rect 25324 21904 25364 21944
rect 25228 21652 25268 21692
rect 25900 21904 25940 21944
rect 25708 21736 25748 21776
rect 25612 21568 25652 21608
rect 25804 21568 25844 21608
rect 25708 21484 25748 21524
rect 25516 21400 25556 21440
rect 23500 19216 23540 19256
rect 22252 18880 22292 18920
rect 23308 18880 23348 18920
rect 22252 18544 22292 18584
rect 22348 18460 22388 18500
rect 23308 18712 23348 18752
rect 24076 18712 24116 18752
rect 22348 17956 22388 17996
rect 22252 17788 22292 17828
rect 21964 17200 22004 17240
rect 22636 18376 22676 18416
rect 22540 17788 22580 17828
rect 22444 17704 22484 17744
rect 22924 17704 22964 17744
rect 23308 18544 23348 18584
rect 23500 18544 23540 18584
rect 23500 18124 23540 18164
rect 23212 17704 23252 17744
rect 23116 17620 23156 17660
rect 23116 17452 23156 17492
rect 21868 17032 21908 17072
rect 21676 16780 21716 16820
rect 21772 16360 21812 16400
rect 21580 16024 21620 16064
rect 21772 15940 21812 15980
rect 21964 16360 22004 16400
rect 22636 17032 22676 17072
rect 22444 16276 22484 16316
rect 22348 16192 22388 16232
rect 22924 16192 22964 16232
rect 22636 16108 22676 16148
rect 22828 16108 22868 16148
rect 22540 16024 22580 16064
rect 23884 18544 23924 18584
rect 24076 18544 24116 18584
rect 23788 18040 23828 18080
rect 23692 17956 23732 17996
rect 24844 19888 24884 19928
rect 25036 19804 25076 19844
rect 24940 19300 24980 19340
rect 25228 20140 25268 20180
rect 25420 20140 25460 20180
rect 25228 19888 25268 19928
rect 24556 18544 24596 18584
rect 24172 18124 24212 18164
rect 23980 17872 24020 17912
rect 23596 17788 23636 17828
rect 23692 17704 23732 17744
rect 23596 17620 23636 17660
rect 23500 17536 23540 17576
rect 23404 17452 23444 17492
rect 23500 16948 23540 16988
rect 23212 16192 23252 16232
rect 23596 16276 23636 16316
rect 21484 15688 21524 15728
rect 21772 15688 21812 15728
rect 19372 15436 19412 15476
rect 18796 15352 18836 15392
rect 17836 15268 17876 15308
rect 17644 15016 17684 15056
rect 16876 14680 16916 14720
rect 16108 14008 16148 14048
rect 16972 14512 17012 14552
rect 16876 14092 16916 14132
rect 16396 13840 16436 13880
rect 16300 13756 16340 13796
rect 16300 13420 16340 13460
rect 15916 13336 15956 13376
rect 15916 13000 15956 13040
rect 16300 13168 16340 13208
rect 17068 14008 17108 14048
rect 17068 13420 17108 13460
rect 17260 14680 17300 14720
rect 17356 14512 17396 14552
rect 17260 14008 17300 14048
rect 18700 15184 18740 15224
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 17932 14848 17972 14888
rect 17836 14260 17876 14300
rect 17260 13168 17300 13208
rect 17164 13084 17204 13124
rect 16108 13000 16148 13040
rect 16492 13000 16532 13040
rect 16012 12748 16052 12788
rect 16204 12664 16244 12704
rect 15724 12244 15764 12284
rect 15724 11740 15764 11780
rect 15532 11656 15572 11696
rect 15628 11320 15668 11360
rect 15436 10900 15476 10940
rect 15916 11068 15956 11108
rect 15724 10984 15764 11024
rect 14668 9640 14708 9680
rect 14956 9640 14996 9680
rect 14284 9304 14324 9344
rect 13708 8884 13748 8924
rect 13420 8632 13460 8672
rect 13132 8128 13172 8168
rect 13036 7876 13076 7916
rect 13804 7876 13844 7916
rect 12844 7540 12884 7580
rect 14284 8632 14324 8672
rect 14284 8380 14324 8420
rect 14188 7876 14228 7916
rect 13996 7540 14036 7580
rect 14668 9388 14708 9428
rect 14572 9220 14612 9260
rect 14956 9472 14996 9512
rect 14860 9388 14900 9428
rect 15052 9136 15092 9176
rect 14860 8884 14900 8924
rect 14764 8800 14804 8840
rect 15244 9808 15284 9848
rect 16684 12496 16724 12536
rect 16588 12328 16628 12368
rect 16300 11656 16340 11696
rect 16588 11656 16628 11696
rect 17164 11824 17204 11864
rect 16972 11656 17012 11696
rect 16108 11488 16148 11528
rect 16300 11488 16340 11528
rect 16876 11488 16916 11528
rect 16396 11320 16436 11360
rect 16204 10984 16244 11024
rect 16108 10900 16148 10940
rect 15436 9724 15476 9764
rect 15340 9472 15380 9512
rect 15436 9388 15476 9428
rect 15532 8800 15572 8840
rect 15724 9808 15764 9848
rect 15916 9724 15956 9764
rect 15820 9640 15860 9680
rect 16108 10312 16148 10352
rect 17548 13252 17588 13292
rect 17740 14092 17780 14132
rect 18316 14680 18356 14720
rect 17932 13504 17972 13544
rect 18412 14512 18452 14552
rect 18892 14848 18932 14888
rect 18508 14260 18548 14300
rect 19660 15352 19700 15392
rect 19948 14848 19988 14888
rect 19852 14680 19892 14720
rect 20140 15520 20180 15560
rect 20620 15520 20660 15560
rect 20236 15268 20276 15308
rect 20236 15100 20276 15140
rect 20236 14764 20276 14804
rect 19660 14512 19700 14552
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 20140 14344 20180 14384
rect 18988 14092 19028 14132
rect 18892 14008 18932 14048
rect 18796 13840 18836 13880
rect 18988 13756 19028 13796
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 17452 13084 17492 13124
rect 17740 13168 17780 13208
rect 18028 13168 18068 13208
rect 18316 13168 18356 13208
rect 18604 13168 18644 13208
rect 17932 12748 17972 12788
rect 17836 12580 17876 12620
rect 17836 11908 17876 11948
rect 18508 12916 18548 12956
rect 18508 12580 18548 12620
rect 19468 14008 19508 14048
rect 19564 13924 19604 13964
rect 19084 13504 19124 13544
rect 19660 13504 19700 13544
rect 19948 14176 19988 14216
rect 19948 13924 19988 13964
rect 19276 13252 19316 13292
rect 19564 13252 19604 13292
rect 19084 13168 19124 13208
rect 19180 13084 19220 13124
rect 19084 12664 19124 12704
rect 19756 13168 19796 13208
rect 19564 13000 19604 13040
rect 19852 13000 19892 13040
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 19468 12664 19508 12704
rect 18796 12496 18836 12536
rect 18412 12412 18452 12452
rect 18988 12412 19028 12452
rect 18316 12328 18356 12368
rect 18796 12244 18836 12284
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 18988 12076 19028 12116
rect 18220 11740 18260 11780
rect 18377 11740 18417 11780
rect 18076 11572 18116 11612
rect 17932 11488 17972 11528
rect 17836 11404 17876 11444
rect 18892 11404 18932 11444
rect 17068 10816 17108 10856
rect 16204 9808 16244 9848
rect 16396 9808 16436 9848
rect 16012 9472 16052 9512
rect 15916 9304 15956 9344
rect 16204 9640 16244 9680
rect 16972 10060 17012 10100
rect 16780 9808 16820 9848
rect 16876 9724 16916 9764
rect 16588 9472 16628 9512
rect 15820 9220 15860 9260
rect 15724 8884 15764 8924
rect 15628 8632 15668 8672
rect 16108 9136 16148 9176
rect 14668 8464 14708 8504
rect 14764 8296 14804 8336
rect 16012 8464 16052 8504
rect 15340 7960 15380 8000
rect 14668 7876 14708 7916
rect 15532 7876 15572 7916
rect 15244 7540 15284 7580
rect 11884 7120 11924 7160
rect 12748 7120 12788 7160
rect 11884 6868 11924 6908
rect 11788 6700 11828 6740
rect 10444 5608 10484 5648
rect 10636 6196 10676 6236
rect 10732 5776 10772 5816
rect 10828 5692 10868 5732
rect 10732 5608 10772 5648
rect 10348 5020 10388 5060
rect 9196 3760 9236 3800
rect 9100 3592 9140 3632
rect 8716 3340 8756 3380
rect 9100 2752 9140 2792
rect 9388 3676 9428 3716
rect 9676 4096 9716 4136
rect 10252 4096 10292 4136
rect 10636 4264 10676 4304
rect 9964 4012 10004 4052
rect 9676 3928 9716 3968
rect 9580 3592 9620 3632
rect 9292 3424 9332 3464
rect 9484 3424 9524 3464
rect 8140 2416 8180 2456
rect 9292 2416 9332 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 9676 2416 9716 2456
rect 9484 1912 9524 1952
rect 844 1660 884 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 9964 1744 10004 1784
rect 9772 1240 9812 1280
rect 10156 1240 10196 1280
rect 11692 6112 11732 6152
rect 11116 6028 11156 6068
rect 11212 5944 11252 5984
rect 11596 5860 11636 5900
rect 11404 5692 11444 5732
rect 11308 5440 11348 5480
rect 11116 5356 11156 5396
rect 11404 5356 11444 5396
rect 11788 5860 11828 5900
rect 11692 5692 11732 5732
rect 12076 6448 12116 6488
rect 13228 7120 13268 7160
rect 11884 5692 11924 5732
rect 11596 5356 11636 5396
rect 11500 5272 11540 5312
rect 11692 5272 11732 5312
rect 11116 5020 11156 5060
rect 11500 5020 11540 5060
rect 11020 4936 11060 4976
rect 11308 4936 11348 4976
rect 11212 4348 11252 4388
rect 11020 4096 11060 4136
rect 10540 4012 10580 4052
rect 10636 3928 10676 3968
rect 10828 3760 10868 3800
rect 10444 3676 10484 3716
rect 11404 4264 11444 4304
rect 11788 5104 11828 5144
rect 11884 5020 11924 5060
rect 11692 4768 11732 4808
rect 11308 3760 11348 3800
rect 11404 3592 11444 3632
rect 11308 3424 11348 3464
rect 10732 1912 10772 1952
rect 12364 6028 12404 6068
rect 12940 6952 12980 6992
rect 12844 6448 12884 6488
rect 13036 6028 13076 6068
rect 12556 5860 12596 5900
rect 12268 5692 12308 5732
rect 12172 5608 12212 5648
rect 12748 5524 12788 5564
rect 12460 5440 12500 5480
rect 13132 5440 13172 5480
rect 13612 6952 13652 6992
rect 13612 6616 13652 6656
rect 13516 5944 13556 5984
rect 13804 6784 13844 6824
rect 13804 6280 13844 6320
rect 13420 5608 13460 5648
rect 14284 7120 14324 7160
rect 14193 6448 14233 6488
rect 14572 6700 14612 6740
rect 14476 6616 14516 6656
rect 14380 6448 14420 6488
rect 14668 6280 14708 6320
rect 15052 7120 15092 7160
rect 15052 6714 15092 6740
rect 15052 6700 15092 6714
rect 14764 6112 14804 6152
rect 13612 5524 13652 5564
rect 12364 4936 12404 4976
rect 11980 4600 12020 4640
rect 11884 4348 11924 4388
rect 11788 4096 11828 4136
rect 12940 4936 12980 4976
rect 13132 4936 13172 4976
rect 11884 3760 11924 3800
rect 11500 3172 11540 3212
rect 12460 4264 12500 4304
rect 12268 3424 12308 3464
rect 12076 3340 12116 3380
rect 12460 3172 12500 3212
rect 10540 1744 10580 1784
rect 13324 4600 13364 4640
rect 13804 5104 13844 5144
rect 14188 5440 14228 5480
rect 13996 5356 14036 5396
rect 14380 5776 14420 5816
rect 14860 5608 14900 5648
rect 14764 5356 14804 5396
rect 14284 5104 14324 5144
rect 14092 4936 14132 4976
rect 13996 4852 14036 4892
rect 14188 4684 14228 4724
rect 13420 4348 13460 4388
rect 14476 5020 14516 5060
rect 14572 4852 14612 4892
rect 15436 6784 15476 6824
rect 15340 6616 15380 6656
rect 15628 6616 15668 6656
rect 15724 6532 15764 6572
rect 15052 5608 15092 5648
rect 14956 5524 14996 5564
rect 15340 5356 15380 5396
rect 14956 5020 14996 5060
rect 14764 4768 14804 4808
rect 15148 4768 15188 4808
rect 14572 4264 14612 4304
rect 14380 4096 14420 4136
rect 14284 3928 14324 3968
rect 13420 3760 13460 3800
rect 14476 3592 14516 3632
rect 14764 4096 14804 4136
rect 14860 3676 14900 3716
rect 14764 3508 14804 3548
rect 15244 4264 15284 4304
rect 13132 3340 13172 3380
rect 15244 3340 15284 3380
rect 14092 2584 14132 2624
rect 15628 5776 15668 5816
rect 16492 9304 16532 9344
rect 16588 8800 16628 8840
rect 16780 8800 16820 8840
rect 16300 8632 16340 8672
rect 16492 7960 16532 8000
rect 16108 6784 16148 6824
rect 16300 6532 16340 6572
rect 16300 6280 16340 6320
rect 15724 5692 15764 5732
rect 15532 5440 15572 5480
rect 15532 5020 15572 5060
rect 15436 4768 15476 4808
rect 15436 3424 15476 3464
rect 15820 4768 15860 4808
rect 16396 5776 16436 5816
rect 16204 5440 16244 5480
rect 16108 5020 16148 5060
rect 16012 4936 16052 4976
rect 15916 3928 15956 3968
rect 15724 3760 15764 3800
rect 15820 3424 15860 3464
rect 15628 3256 15668 3296
rect 15724 3172 15764 3212
rect 15436 3004 15476 3044
rect 16108 4096 16148 4136
rect 16396 4936 16436 4976
rect 16972 9220 17012 9260
rect 17356 11068 17396 11108
rect 17452 10984 17492 11024
rect 17836 10984 17876 11024
rect 18316 10984 18356 11024
rect 17548 10900 17588 10940
rect 17356 10648 17396 10688
rect 19564 12580 19604 12620
rect 19852 12580 19892 12620
rect 19084 11992 19124 12032
rect 19468 12244 19508 12284
rect 19468 11824 19508 11864
rect 18508 10900 18548 10940
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 17548 10144 17588 10184
rect 17164 9304 17204 9344
rect 18892 10060 18932 10100
rect 19372 11740 19412 11780
rect 19180 11572 19220 11612
rect 19276 11488 19316 11528
rect 19756 12412 19796 12452
rect 19564 11656 19604 11696
rect 19756 11992 19796 12032
rect 19756 11824 19796 11864
rect 19660 11488 19700 11528
rect 20140 13168 20180 13208
rect 20140 12916 20180 12956
rect 20716 15436 20756 15476
rect 20812 15100 20852 15140
rect 20524 14512 20564 14552
rect 20620 14428 20660 14468
rect 20428 14008 20468 14048
rect 20428 13840 20468 13880
rect 20332 13168 20372 13208
rect 20524 13168 20564 13208
rect 20044 12496 20084 12536
rect 20236 12664 20276 12704
rect 20044 12244 20084 12284
rect 19948 11824 19988 11864
rect 19948 11656 19988 11696
rect 20201 11740 20241 11780
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 19084 10732 19124 10772
rect 18988 9976 19028 10016
rect 17548 9220 17588 9260
rect 16684 8380 16724 8420
rect 16972 7960 17012 8000
rect 17548 7120 17588 7160
rect 18028 7120 18068 7160
rect 17740 6700 17780 6740
rect 16876 6280 16916 6320
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 19852 10984 19892 11024
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 20332 11236 20372 11276
rect 20140 10732 20180 10772
rect 20332 10396 20372 10436
rect 20332 10228 20372 10268
rect 20044 9724 20084 9764
rect 20812 14008 20852 14048
rect 21484 15520 21524 15560
rect 21964 15520 22004 15560
rect 22252 15436 22292 15476
rect 22060 14848 22100 14888
rect 20908 13924 20948 13964
rect 21100 13168 21140 13208
rect 21292 14092 21332 14132
rect 21868 14680 21908 14720
rect 21676 14596 21716 14636
rect 21580 14512 21620 14552
rect 21676 14176 21716 14216
rect 21772 13924 21812 13964
rect 21614 13420 21654 13460
rect 21868 13420 21908 13460
rect 21484 13252 21524 13292
rect 20716 12664 20756 12704
rect 21196 12580 21236 12620
rect 20812 12496 20852 12536
rect 21484 13000 21524 13040
rect 21676 13000 21716 13040
rect 21580 12580 21620 12620
rect 20620 12076 20660 12116
rect 21868 12748 21908 12788
rect 21772 11656 21812 11696
rect 20620 11236 20660 11276
rect 20716 10732 20756 10772
rect 20812 10144 20852 10184
rect 20908 10060 20948 10100
rect 21388 10648 21428 10688
rect 22252 14176 22292 14216
rect 22156 14008 22196 14048
rect 22060 13420 22100 13460
rect 22060 13252 22100 13292
rect 22828 15772 22868 15812
rect 22732 15604 22772 15644
rect 22540 15520 22580 15560
rect 23020 15688 23060 15728
rect 22924 15520 22964 15560
rect 22444 15352 22484 15392
rect 23020 14596 23060 14636
rect 23020 14008 23060 14048
rect 22444 13168 22484 13208
rect 22252 11656 22292 11696
rect 22156 11068 22196 11108
rect 22060 10984 22100 11024
rect 21868 10732 21908 10772
rect 22540 12664 22580 12704
rect 23020 11656 23060 11696
rect 22540 11068 22580 11108
rect 22060 10396 22100 10436
rect 21484 10228 21524 10268
rect 21388 10060 21428 10100
rect 21676 8884 21716 8924
rect 20524 8716 20564 8756
rect 20332 8632 20372 8672
rect 19276 8380 19316 8420
rect 18796 7960 18836 8000
rect 19180 7960 19220 8000
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 18988 7120 19028 7160
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 20620 8296 20660 8336
rect 20524 7960 20564 8000
rect 21196 7960 21236 8000
rect 21484 7708 21524 7748
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 18124 6448 18164 6488
rect 19372 6448 19412 6488
rect 19564 6448 19604 6488
rect 18412 6280 18452 6320
rect 18124 6112 18164 6152
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 16300 4096 16340 4136
rect 17932 5608 17972 5648
rect 18124 5608 18164 5648
rect 17740 5020 17780 5060
rect 18028 4684 18068 4724
rect 16300 3424 16340 3464
rect 16108 3004 16148 3044
rect 16012 2752 16052 2792
rect 16012 2584 16052 2624
rect 16204 2752 16244 2792
rect 16588 3508 16628 3548
rect 16396 3340 16436 3380
rect 16492 3088 16532 3128
rect 16396 2836 16436 2876
rect 16300 2668 16340 2708
rect 18412 4768 18452 4808
rect 19180 5608 19220 5648
rect 20236 5608 20276 5648
rect 20332 5356 20372 5396
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 19372 4768 19412 4808
rect 18892 4684 18932 4724
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 19756 4096 19796 4136
rect 19852 4012 19892 4052
rect 19564 3928 19604 3968
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 21388 6952 21428 6992
rect 21772 6952 21812 6992
rect 21964 10144 22004 10184
rect 23692 16192 23732 16232
rect 23692 15940 23732 15980
rect 24268 17788 24308 17828
rect 24076 17536 24116 17576
rect 24076 17200 24116 17240
rect 23884 17032 23924 17072
rect 25516 19552 25556 19592
rect 25708 19888 25748 19928
rect 26572 21568 26612 21608
rect 26380 21400 26420 21440
rect 26092 20308 26132 20348
rect 26284 20224 26324 20264
rect 28492 28120 28532 28160
rect 28684 28120 28724 28160
rect 28684 27952 28724 27992
rect 28492 27616 28532 27656
rect 29068 27616 29108 27656
rect 29260 27616 29300 27656
rect 28588 27532 28628 27572
rect 28684 27448 28724 27488
rect 28492 27364 28532 27404
rect 27340 26524 27380 26564
rect 27628 26188 27668 26228
rect 27244 25852 27284 25892
rect 27724 26104 27764 26144
rect 27532 25768 27572 25808
rect 27532 25432 27572 25472
rect 27916 24592 27956 24632
rect 28396 26440 28436 26480
rect 28300 26104 28340 26144
rect 28108 24858 28148 24884
rect 28108 24844 28148 24858
rect 27244 23836 27284 23876
rect 27532 23836 27572 23876
rect 27724 23836 27764 23876
rect 27148 23668 27188 23708
rect 27340 23584 27380 23624
rect 27244 23332 27284 23372
rect 27628 23752 27668 23792
rect 27916 23752 27956 23792
rect 27724 23584 27764 23624
rect 27532 23416 27572 23456
rect 27436 23248 27476 23288
rect 27052 22828 27092 22868
rect 27052 22156 27092 22196
rect 26668 20224 26708 20264
rect 26380 20140 26420 20180
rect 27244 22240 27284 22280
rect 27820 23416 27860 23456
rect 27724 22744 27764 22784
rect 27532 22576 27572 22616
rect 27436 21736 27476 21776
rect 28396 26020 28436 26060
rect 29548 27651 29588 27656
rect 29548 27616 29588 27651
rect 29164 27364 29204 27404
rect 29740 27700 29780 27740
rect 28780 27028 28820 27068
rect 29644 26944 29684 26984
rect 28588 24592 28628 24632
rect 28300 24088 28340 24128
rect 28492 23752 28532 23792
rect 28972 26776 29012 26816
rect 29068 26524 29108 26564
rect 29548 26776 29588 26816
rect 29452 26440 29492 26480
rect 29740 26272 29780 26312
rect 29836 26104 29876 26144
rect 29548 25516 29588 25556
rect 29356 25432 29396 25472
rect 28876 24844 28916 24884
rect 30412 28288 30452 28328
rect 30892 33412 30932 33452
rect 30796 32908 30836 32948
rect 30604 30892 30644 30932
rect 30604 30724 30644 30764
rect 32044 35680 32084 35720
rect 31468 35092 31508 35132
rect 31276 35008 31316 35048
rect 31660 34672 31700 34712
rect 31756 34588 31796 34628
rect 31276 34420 31316 34460
rect 31084 33580 31124 33620
rect 31276 33412 31316 33452
rect 31468 33244 31508 33284
rect 31180 31312 31220 31352
rect 30892 31144 30932 31184
rect 32236 35176 32276 35216
rect 32236 34924 32276 34964
rect 32140 34672 32180 34712
rect 31948 34504 31988 34544
rect 31756 33916 31796 33956
rect 31852 33664 31892 33704
rect 32236 34336 32276 34376
rect 32140 33664 32180 33704
rect 31372 31144 31412 31184
rect 31276 30976 31316 31016
rect 30988 30892 31028 30932
rect 31084 30808 31124 30848
rect 31564 31144 31604 31184
rect 31756 31144 31796 31184
rect 31564 30976 31604 31016
rect 31180 30724 31220 30764
rect 30892 30472 30932 30512
rect 30700 29296 30740 29336
rect 30604 29128 30644 29168
rect 30700 28960 30740 29000
rect 30604 28876 30644 28916
rect 31372 30472 31412 30512
rect 30988 29800 31028 29840
rect 31084 29128 31124 29168
rect 30988 28960 31028 29000
rect 31084 28540 31124 28580
rect 30796 28456 30836 28496
rect 30412 27616 30452 27656
rect 30316 27028 30356 27068
rect 30316 26860 30356 26900
rect 30892 28288 30932 28328
rect 31372 28456 31412 28496
rect 31180 27868 31220 27908
rect 30700 27700 30740 27740
rect 30796 27280 30836 27320
rect 30700 27028 30740 27068
rect 31276 27784 31316 27824
rect 30988 27700 31028 27740
rect 31276 27448 31316 27488
rect 30988 27028 31028 27068
rect 30700 26776 30740 26816
rect 30700 26608 30740 26648
rect 30220 25432 30260 25472
rect 28876 23920 28916 23960
rect 28204 23668 28244 23708
rect 28300 23248 28340 23288
rect 28108 23164 28148 23204
rect 28588 23416 28628 23456
rect 28108 22996 28148 23036
rect 28780 23752 28820 23792
rect 28780 23248 28820 23288
rect 28684 22996 28724 23036
rect 28972 23836 29012 23876
rect 29164 23836 29204 23876
rect 28972 23584 29012 23624
rect 29452 23752 29492 23792
rect 29452 23584 29492 23624
rect 29260 23416 29300 23456
rect 29452 23416 29492 23456
rect 29068 23332 29108 23372
rect 29164 23164 29204 23204
rect 28972 23080 29012 23120
rect 29740 23248 29780 23288
rect 29548 23164 29588 23204
rect 30124 23080 30164 23120
rect 28876 22912 28916 22952
rect 28588 22828 28628 22868
rect 28588 22324 28628 22364
rect 27916 22156 27956 22196
rect 29164 22324 29204 22364
rect 28876 22240 28916 22280
rect 28780 22156 28820 22196
rect 30412 23080 30452 23120
rect 29932 22912 29972 22952
rect 29452 22072 29492 22112
rect 28588 21904 28628 21944
rect 27628 21568 27668 21608
rect 27532 21400 27572 21440
rect 27148 20308 27188 20348
rect 26092 19888 26132 19928
rect 26380 19972 26420 20012
rect 25996 19552 26036 19592
rect 25612 18880 25652 18920
rect 25899 18964 25939 19004
rect 24556 17704 24596 17744
rect 24364 17620 24404 17660
rect 24460 17452 24500 17492
rect 23980 16948 24020 16988
rect 23980 16444 24020 16484
rect 25516 18544 25556 18584
rect 25036 18376 25076 18416
rect 24652 17452 24692 17492
rect 24172 16696 24212 16736
rect 23308 15436 23348 15476
rect 23788 15184 23828 15224
rect 23212 14092 23252 14132
rect 23692 11656 23732 11696
rect 24940 17452 24980 17492
rect 24940 16528 24980 16568
rect 24748 16360 24788 16400
rect 24268 16192 24308 16232
rect 24172 15772 24212 15812
rect 24364 15940 24404 15980
rect 24556 16108 24596 16148
rect 24748 15940 24788 15980
rect 25420 17536 25460 17576
rect 25516 17368 25556 17408
rect 25228 17032 25268 17072
rect 25036 16192 25076 16232
rect 25036 15940 25076 15980
rect 24460 15856 24500 15896
rect 24844 15688 24884 15728
rect 24460 15436 24500 15476
rect 24748 15436 24788 15476
rect 24940 15520 24980 15560
rect 24172 15352 24212 15392
rect 24268 15100 24308 15140
rect 23980 14932 24020 14972
rect 23116 11236 23156 11276
rect 23020 10144 23060 10184
rect 23404 10228 23444 10268
rect 22444 10060 22484 10100
rect 23404 9472 23444 9512
rect 22828 9388 22868 9428
rect 22540 9052 22580 9092
rect 22732 8716 22772 8756
rect 22060 7960 22100 8000
rect 22540 7960 22580 8000
rect 22252 7540 22292 7580
rect 22252 7372 22292 7412
rect 22156 7288 22196 7328
rect 21580 6448 21620 6488
rect 20428 4684 20468 4724
rect 20044 4096 20084 4136
rect 20716 4096 20756 4136
rect 21868 5608 21908 5648
rect 21484 5356 21524 5396
rect 21484 4768 21524 4808
rect 20332 4012 20372 4052
rect 16684 3256 16724 3296
rect 16876 2836 16916 2876
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 16972 2668 17012 2708
rect 17836 2668 17876 2708
rect 18028 2668 18068 2708
rect 18700 2584 18740 2624
rect 19180 2584 19220 2624
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 20236 3172 20276 3212
rect 20716 3844 20756 3884
rect 21004 3760 21044 3800
rect 21292 3760 21332 3800
rect 21676 4096 21716 4136
rect 22636 7120 22676 7160
rect 22444 6448 22484 6488
rect 22252 6280 22292 6320
rect 22924 8464 22964 8504
rect 24172 11236 24212 11276
rect 24364 11068 24404 11108
rect 23788 10984 23828 11024
rect 23692 10228 23732 10268
rect 25804 18460 25844 18500
rect 25708 18376 25748 18416
rect 25708 17536 25748 17576
rect 25612 16696 25652 16736
rect 25324 16612 25364 16652
rect 25420 16444 25460 16484
rect 25132 15604 25172 15644
rect 24748 14932 24788 14972
rect 24844 13252 24884 13292
rect 24748 12328 24788 12368
rect 24748 10984 24788 11024
rect 24364 10144 24404 10184
rect 25132 13924 25172 13964
rect 25132 11068 25172 11108
rect 24844 10060 24884 10100
rect 23980 8800 24020 8840
rect 23404 8716 23444 8756
rect 23020 8380 23060 8420
rect 23116 7960 23156 8000
rect 23596 8464 23636 8504
rect 24172 9472 24212 9512
rect 24844 9556 24884 9596
rect 24556 9304 24596 9344
rect 24172 8968 24212 9008
rect 24076 8548 24116 8588
rect 23404 8128 23444 8168
rect 23020 7876 23060 7916
rect 23020 7708 23060 7748
rect 22924 7540 22964 7580
rect 23308 7876 23348 7916
rect 23500 7876 23540 7916
rect 23212 7540 23252 7580
rect 23465 7288 23505 7328
rect 23308 6952 23348 6992
rect 23116 6700 23156 6740
rect 22732 6532 22772 6572
rect 23212 6448 23252 6488
rect 22156 5608 22196 5648
rect 21964 4936 22004 4976
rect 22924 6280 22964 6320
rect 22348 5020 22388 5060
rect 22732 5020 22772 5060
rect 22156 4852 22196 4892
rect 22060 4768 22100 4808
rect 22156 4684 22196 4724
rect 22156 4096 22196 4136
rect 22060 3760 22100 3800
rect 20044 2080 20084 2120
rect 20812 2080 20852 2120
rect 21004 1912 21044 1952
rect 22060 2836 22100 2876
rect 21964 2668 22004 2708
rect 21868 2584 21908 2624
rect 23500 6952 23540 6992
rect 23404 6784 23444 6824
rect 24172 8128 24212 8168
rect 23692 7876 23732 7916
rect 23884 7540 23924 7580
rect 23788 7120 23828 7160
rect 24172 7960 24212 8000
rect 23980 7120 24020 7160
rect 24940 9304 24980 9344
rect 24652 8968 24692 9008
rect 24652 8800 24692 8840
rect 25324 15520 25364 15560
rect 25612 16360 25652 16400
rect 25708 15436 25748 15476
rect 25612 15352 25652 15392
rect 25612 15016 25652 15056
rect 26092 17956 26132 17996
rect 25996 17872 26036 17912
rect 25900 17536 25940 17576
rect 25900 17368 25940 17408
rect 26476 19804 26516 19844
rect 26956 20056 26996 20096
rect 26764 19720 26804 19760
rect 26668 19216 26708 19256
rect 27148 19048 27188 19088
rect 26764 18880 26804 18920
rect 26668 18712 26708 18752
rect 26668 18544 26708 18584
rect 26572 18460 26612 18500
rect 27148 17956 27188 17996
rect 27916 20056 27956 20096
rect 28012 19972 28052 20012
rect 28396 19888 28436 19928
rect 28300 19720 28340 19760
rect 26284 17872 26324 17912
rect 26188 17620 26228 17660
rect 26284 17452 26324 17492
rect 26764 17620 26804 17660
rect 26476 17536 26516 17576
rect 27244 17536 27284 17576
rect 26668 17284 26708 17324
rect 27052 17284 27092 17324
rect 26380 16444 26420 16484
rect 25900 15436 25940 15476
rect 25900 14764 25940 14804
rect 26572 16612 26612 16652
rect 26476 16360 26516 16400
rect 26956 16780 26996 16820
rect 26668 16276 26708 16316
rect 27148 17200 27188 17240
rect 27628 17536 27668 17576
rect 27724 17298 27764 17324
rect 27724 17284 27764 17298
rect 28108 18964 28148 19004
rect 30604 25852 30644 25892
rect 30604 25264 30644 25304
rect 30604 24592 30644 24632
rect 30988 26860 31028 26900
rect 30892 26776 30932 26816
rect 31084 26776 31124 26816
rect 31660 29800 31700 29840
rect 31756 29296 31796 29336
rect 31564 29128 31604 29168
rect 31756 29044 31796 29084
rect 32044 32152 32084 32192
rect 32140 32068 32180 32108
rect 35596 36520 35636 36560
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 32524 35260 32564 35300
rect 33196 35260 33236 35300
rect 32908 35176 32948 35216
rect 35212 35848 35252 35888
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 34732 35344 34772 35384
rect 34636 35260 34676 35300
rect 33964 35176 34004 35216
rect 33100 35092 33140 35132
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 32524 34588 32564 34628
rect 32428 34336 32468 34376
rect 32332 32824 32372 32864
rect 33772 34336 33812 34376
rect 33196 34000 33236 34040
rect 33772 34000 33812 34040
rect 32428 32320 32468 32360
rect 32332 32068 32372 32108
rect 31948 31480 31988 31520
rect 31948 30220 31988 30260
rect 31948 29800 31988 29840
rect 31948 29128 31988 29168
rect 31468 28288 31508 28328
rect 32428 31480 32468 31520
rect 32908 31480 32948 31520
rect 32236 31144 32276 31184
rect 32236 30220 32276 30260
rect 32428 30640 32468 30680
rect 34540 35176 34580 35216
rect 34348 35092 34388 35132
rect 34252 34840 34292 34880
rect 35116 35008 35156 35048
rect 35020 34336 35060 34376
rect 34348 34000 34388 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 34348 33664 34388 33704
rect 33676 33580 33716 33620
rect 33868 33580 33908 33620
rect 34252 33580 34292 33620
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 33484 32152 33524 32192
rect 33196 32068 33236 32108
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 32716 30220 32756 30260
rect 33004 30388 33044 30428
rect 32332 29380 32372 29420
rect 32908 29212 32948 29252
rect 33292 31312 33332 31352
rect 33580 31480 33620 31520
rect 33484 31396 33524 31436
rect 35404 35344 35444 35384
rect 35308 35260 35348 35300
rect 35404 35176 35444 35216
rect 35212 34084 35252 34124
rect 35788 35176 35828 35216
rect 36460 36520 36500 36560
rect 37612 36520 37652 36560
rect 36076 35848 36116 35888
rect 36076 35260 36116 35300
rect 35980 35176 36020 35216
rect 36460 35176 36500 35216
rect 36364 35008 36404 35048
rect 35788 34168 35828 34208
rect 35500 33916 35540 33956
rect 36364 33916 36404 33956
rect 36940 35092 36980 35132
rect 37612 35344 37652 35384
rect 39148 35428 39188 35468
rect 38284 35260 38324 35300
rect 38092 35176 38132 35216
rect 38668 35260 38708 35300
rect 39052 35260 39092 35300
rect 38476 34504 38516 34544
rect 37612 34420 37652 34460
rect 36940 34252 36980 34292
rect 36844 34168 36884 34208
rect 36460 33832 36500 33872
rect 36652 33664 36692 33704
rect 36556 33496 36596 33536
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 36076 32320 36116 32360
rect 34924 32152 34964 32192
rect 33964 31312 34004 31352
rect 33100 29800 33140 29840
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 33868 31144 33908 31184
rect 33868 30640 33908 30680
rect 33196 29296 33236 29336
rect 33580 29800 33620 29840
rect 34444 31480 34484 31520
rect 34252 30976 34292 31016
rect 35116 31312 35156 31352
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 34252 30640 34292 30680
rect 34444 30640 34484 30680
rect 35404 31144 35444 31184
rect 34348 30556 34388 30596
rect 34060 30052 34100 30092
rect 33964 29212 34004 29252
rect 33772 29128 33812 29168
rect 33676 29044 33716 29084
rect 34252 29128 34292 29168
rect 32428 28540 32468 28580
rect 32620 28540 32660 28580
rect 32140 27784 32180 27824
rect 31468 27448 31508 27488
rect 31372 27196 31412 27236
rect 31180 26356 31220 26396
rect 30988 25936 31028 25976
rect 30892 25600 30932 25640
rect 30796 25516 30836 25556
rect 31756 27616 31796 27656
rect 31756 27028 31796 27068
rect 31372 26860 31412 26900
rect 32140 26860 32180 26900
rect 31948 26776 31988 26816
rect 32236 26776 32276 26816
rect 31564 26440 31604 26480
rect 31756 26440 31796 26480
rect 33100 28960 33140 29000
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 34444 30388 34484 30428
rect 35308 30640 35348 30680
rect 35500 30556 35540 30596
rect 35116 30220 35156 30260
rect 34444 30136 34484 30176
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 35596 30220 35636 30260
rect 35980 30556 36020 30596
rect 36268 32908 36308 32948
rect 36268 32152 36308 32192
rect 36172 30472 36212 30512
rect 35884 30220 35924 30260
rect 35692 30052 35732 30092
rect 35788 29212 35828 29252
rect 35596 29044 35636 29084
rect 36268 30052 36308 30092
rect 35980 29884 36020 29924
rect 36652 30640 36692 30680
rect 36556 29884 36596 29924
rect 35980 29632 36020 29672
rect 36268 29800 36308 29840
rect 36460 29632 36500 29672
rect 36076 29044 36116 29084
rect 35212 28204 35252 28244
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 32812 27616 32852 27656
rect 33292 27616 33332 27656
rect 33964 27616 34004 27656
rect 32524 27196 32564 27236
rect 32428 26860 32468 26900
rect 33100 27448 33140 27488
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 32812 26776 32852 26816
rect 32524 26692 32564 26732
rect 32332 26272 32372 26312
rect 31372 26104 31412 26144
rect 31276 25516 31316 25556
rect 31180 25180 31220 25220
rect 30796 23752 30836 23792
rect 30700 23332 30740 23372
rect 30892 23332 30932 23372
rect 31660 25516 31700 25556
rect 33868 27196 33908 27236
rect 34156 25936 34196 25976
rect 32716 25852 32756 25892
rect 33580 25852 33620 25892
rect 32332 25768 32372 25808
rect 32524 25432 32564 25472
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 33868 25684 33908 25724
rect 32812 25432 32852 25472
rect 33004 25264 33044 25304
rect 32428 25180 32468 25220
rect 33292 25180 33332 25220
rect 34348 27616 34388 27656
rect 34444 26776 34484 26816
rect 35020 27616 35060 27656
rect 35212 27616 35252 27656
rect 34828 27448 34868 27488
rect 34348 25684 34388 25724
rect 34060 25264 34100 25304
rect 34348 25432 34388 25472
rect 34252 25264 34292 25304
rect 34156 25180 34196 25220
rect 34348 25180 34388 25220
rect 34156 25012 34196 25052
rect 33964 24592 34004 24632
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 31180 23164 31220 23204
rect 30796 23080 30836 23120
rect 31084 23080 31124 23120
rect 31468 23752 31508 23792
rect 31852 23164 31892 23204
rect 31756 23080 31796 23120
rect 31276 22996 31316 23036
rect 31180 22240 31220 22280
rect 34348 23836 34388 23876
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 35308 27532 35348 27572
rect 35692 27784 35732 27824
rect 36364 27700 36404 27740
rect 35596 27364 35636 27404
rect 35212 25936 35252 25976
rect 34540 25600 34580 25640
rect 34540 25432 34580 25472
rect 34924 25432 34964 25472
rect 35116 25432 35156 25472
rect 34828 25348 34868 25388
rect 34732 25180 34772 25220
rect 35020 25180 35060 25220
rect 34636 25096 34676 25136
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 35404 26608 35444 26648
rect 37324 34000 37364 34040
rect 37228 32908 37268 32948
rect 37516 33580 37556 33620
rect 38380 34000 38420 34040
rect 37612 32320 37652 32360
rect 40396 35428 40436 35468
rect 40300 35344 40340 35384
rect 38956 35092 38996 35132
rect 39052 34588 39092 34628
rect 39436 34672 39476 34712
rect 39532 34588 39572 34628
rect 40300 35092 40340 35132
rect 40684 35008 40724 35048
rect 39628 34504 39668 34544
rect 40108 34420 40148 34460
rect 39436 34252 39476 34292
rect 38572 34168 38612 34208
rect 38860 34168 38900 34208
rect 39052 34168 39092 34208
rect 39340 34168 39380 34208
rect 38860 33832 38900 33872
rect 38092 33580 38132 33620
rect 37900 33412 37940 33452
rect 37804 32320 37844 32360
rect 38284 33412 38324 33452
rect 38572 33664 38612 33704
rect 38956 33664 38996 33704
rect 39244 34000 39284 34040
rect 39916 34252 39956 34292
rect 40204 34336 40244 34376
rect 40972 35176 41012 35216
rect 40876 34588 40916 34628
rect 40588 34420 40628 34460
rect 40492 34336 40532 34376
rect 40780 34252 40820 34292
rect 40012 34168 40052 34208
rect 39532 33832 39572 33872
rect 40012 33748 40052 33788
rect 40108 33664 40148 33704
rect 39916 33496 39956 33536
rect 39148 32824 39188 32864
rect 38476 32152 38516 32192
rect 37036 30640 37076 30680
rect 37228 30640 37268 30680
rect 37708 30640 37748 30680
rect 37516 30220 37556 30260
rect 37132 30052 37172 30092
rect 37420 29884 37460 29924
rect 37324 29800 37364 29840
rect 37228 29128 37268 29168
rect 37132 29044 37172 29084
rect 37228 28876 37268 28916
rect 37708 30220 37748 30260
rect 37708 29632 37748 29672
rect 37228 28288 37268 28328
rect 38188 30640 38228 30680
rect 38380 30640 38420 30680
rect 39244 32152 39284 32192
rect 40300 32908 40340 32948
rect 40204 32488 40244 32528
rect 38668 30808 38708 30848
rect 40300 31144 40340 31184
rect 39244 30976 39284 31016
rect 38284 30304 38324 30344
rect 38380 29968 38420 30008
rect 38188 29212 38228 29252
rect 38764 30556 38804 30596
rect 38764 30304 38804 30344
rect 38476 29044 38516 29084
rect 38092 28624 38132 28664
rect 38380 28288 38420 28328
rect 39052 30640 39092 30680
rect 39532 30808 39572 30848
rect 39340 30556 39380 30596
rect 39148 30472 39188 30512
rect 40300 30472 40340 30512
rect 39052 29800 39092 29840
rect 39436 30220 39476 30260
rect 38956 29044 38996 29084
rect 39052 28624 39092 28664
rect 38860 28540 38900 28580
rect 39340 28540 39380 28580
rect 39820 29296 39860 29336
rect 40108 29044 40148 29084
rect 39436 28456 39476 28496
rect 38860 28288 38900 28328
rect 38380 27700 38420 27740
rect 36844 27028 36884 27068
rect 36268 26860 36308 26900
rect 35692 26776 35732 26816
rect 35980 26776 36020 26816
rect 36172 26776 36212 26816
rect 35884 26608 35924 26648
rect 36076 26608 36116 26648
rect 35500 25432 35540 25472
rect 35308 25348 35348 25388
rect 35212 25264 35252 25304
rect 35596 25180 35636 25220
rect 36076 25264 36116 25304
rect 34828 23584 34868 23624
rect 34252 22912 34292 22952
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 32908 22492 32948 22532
rect 30892 22072 30932 22112
rect 30988 21568 31028 21608
rect 28684 19300 28724 19340
rect 28780 18964 28820 19004
rect 28204 18880 28244 18920
rect 28588 18880 28628 18920
rect 28972 18880 29012 18920
rect 28396 18544 28436 18584
rect 29068 17956 29108 17996
rect 27916 17200 27956 17240
rect 27244 16948 27284 16988
rect 27148 16780 27188 16820
rect 27436 16780 27476 16820
rect 27244 16612 27284 16652
rect 27244 16360 27284 16400
rect 27052 16192 27092 16232
rect 26860 16024 26900 16064
rect 27244 15772 27284 15812
rect 26668 15688 26708 15728
rect 27244 15520 27284 15560
rect 27436 16360 27476 16400
rect 27628 16864 27668 16904
rect 29164 17872 29204 17912
rect 27820 16864 27860 16904
rect 27820 16444 27860 16484
rect 27532 16276 27572 16316
rect 28204 16444 28244 16484
rect 28108 16360 28148 16400
rect 28012 16192 28052 16232
rect 27436 16024 27476 16064
rect 27628 15940 27668 15980
rect 27724 15604 27764 15644
rect 26572 15184 26612 15224
rect 26284 15016 26324 15056
rect 26380 14764 26420 14804
rect 26860 14764 26900 14804
rect 25900 14596 25940 14636
rect 26092 14512 26132 14552
rect 26668 14512 26708 14552
rect 25516 14008 25556 14048
rect 27244 14260 27284 14300
rect 27052 14176 27092 14216
rect 26188 14092 26228 14132
rect 26284 14008 26324 14048
rect 26188 13924 26228 13964
rect 25708 13840 25748 13880
rect 25708 13252 25748 13292
rect 26092 13252 26132 13292
rect 25420 13168 25460 13208
rect 26476 13588 26516 13628
rect 26764 13504 26804 13544
rect 26476 13336 26516 13376
rect 26284 12664 26324 12704
rect 25900 12580 25940 12620
rect 26188 12496 26228 12536
rect 26764 13252 26804 13292
rect 26764 13084 26804 13124
rect 26764 12916 26804 12956
rect 26668 12748 26708 12788
rect 26572 12664 26612 12704
rect 26860 12832 26900 12872
rect 26092 12412 26132 12452
rect 25996 12328 26036 12368
rect 26284 12160 26324 12200
rect 26572 12328 26612 12368
rect 26380 11824 26420 11864
rect 25804 11572 25844 11612
rect 25612 11488 25652 11528
rect 26188 11656 26228 11696
rect 25804 11236 25844 11276
rect 25708 11152 25748 11192
rect 25420 10144 25460 10184
rect 25324 9976 25364 10016
rect 25228 9388 25268 9428
rect 25036 8800 25076 8840
rect 24748 8548 24788 8588
rect 25132 8548 25172 8588
rect 25036 8464 25076 8504
rect 24844 8380 24884 8420
rect 25036 8212 25076 8252
rect 25228 8464 25268 8504
rect 24713 7288 24753 7328
rect 24556 7204 24596 7244
rect 23884 7036 23924 7076
rect 23788 6952 23828 6992
rect 23692 6532 23732 6572
rect 23596 6448 23636 6488
rect 24268 6952 24308 6992
rect 23884 6616 23924 6656
rect 24076 6448 24116 6488
rect 23308 5608 23348 5648
rect 23212 5020 23252 5060
rect 23020 4936 23060 4976
rect 23692 4936 23732 4976
rect 23596 4852 23636 4892
rect 23788 4180 23828 4220
rect 23884 3928 23924 3968
rect 23596 3844 23636 3884
rect 23980 3172 24020 3212
rect 23980 2836 24020 2876
rect 23308 2668 23348 2708
rect 23596 2668 23636 2708
rect 23116 2584 23156 2624
rect 22252 1912 22292 1952
rect 22540 1912 22580 1952
rect 17452 1660 17492 1700
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 24268 6448 24308 6488
rect 25228 7960 25268 8000
rect 26092 11488 26132 11528
rect 26380 11656 26420 11696
rect 26764 12412 26804 12452
rect 26764 11824 26804 11864
rect 26668 11740 26708 11780
rect 27148 13840 27188 13880
rect 28108 15604 28148 15644
rect 28012 15520 28052 15560
rect 28204 15520 28244 15560
rect 28108 15184 28148 15224
rect 28775 17200 28815 17240
rect 28775 17032 28815 17072
rect 28972 17032 29012 17072
rect 28972 16780 29012 16820
rect 28876 16612 28916 16652
rect 29356 17956 29396 17996
rect 29260 17452 29300 17492
rect 29260 17284 29300 17324
rect 29164 17032 29204 17072
rect 29260 16780 29300 16820
rect 28684 16024 28724 16064
rect 29548 18628 29588 18668
rect 30316 20056 30356 20096
rect 29932 19888 29972 19928
rect 29836 18628 29876 18668
rect 29740 18544 29780 18584
rect 29452 17116 29492 17156
rect 29548 16948 29588 16988
rect 29452 16528 29492 16568
rect 29452 16360 29492 16400
rect 30796 19216 30836 19256
rect 30604 19048 30644 19088
rect 29932 16276 29972 16316
rect 29644 16108 29684 16148
rect 29068 16024 29108 16064
rect 29260 15940 29300 15980
rect 28780 15856 28820 15896
rect 30220 17536 30260 17576
rect 30220 17284 30260 17324
rect 31084 18544 31124 18584
rect 31660 19300 31700 19340
rect 31468 18964 31508 19004
rect 30604 17704 30644 17744
rect 30412 17032 30452 17072
rect 30220 16444 30260 16484
rect 30124 16192 30164 16232
rect 30508 16192 30548 16232
rect 29932 15940 29972 15980
rect 30604 15772 30644 15812
rect 29932 15688 29972 15728
rect 30508 15688 30548 15728
rect 28780 15436 28820 15476
rect 29548 15100 29588 15140
rect 28300 14764 28340 14804
rect 27916 14344 27956 14384
rect 28204 14344 28244 14384
rect 27532 13420 27572 13460
rect 28588 14680 28628 14720
rect 29740 14764 29780 14804
rect 28492 14260 28532 14300
rect 28588 14176 28628 14216
rect 28396 14092 28436 14132
rect 27340 12832 27380 12872
rect 28012 13168 28052 13208
rect 27820 12916 27860 12956
rect 27340 12664 27380 12704
rect 27724 12664 27764 12704
rect 26956 12160 26996 12200
rect 26956 11908 26996 11948
rect 27244 11992 27284 12032
rect 27148 11824 27188 11864
rect 26476 11152 26516 11192
rect 26668 11152 26708 11192
rect 26284 10984 26324 11024
rect 26476 10984 26516 11024
rect 27148 11656 27188 11696
rect 27628 12580 27668 12620
rect 27916 12832 27956 12872
rect 27532 12496 27572 12536
rect 27916 12496 27956 12536
rect 27436 12412 27476 12452
rect 28300 13672 28340 13712
rect 28204 13336 28244 13376
rect 28204 13084 28244 13124
rect 28972 14092 29012 14132
rect 29260 14344 29300 14384
rect 28876 13924 28916 13964
rect 28780 13840 28820 13880
rect 28588 13588 28628 13628
rect 28396 12916 28436 12956
rect 28684 13336 28724 13376
rect 28972 13840 29012 13880
rect 29164 13756 29204 13796
rect 29068 13588 29108 13628
rect 29452 14596 29492 14636
rect 29356 14092 29396 14132
rect 30988 17704 31028 17744
rect 30892 16108 30932 16148
rect 30700 15604 30740 15644
rect 30604 15184 30644 15224
rect 29836 14680 29876 14720
rect 29644 14596 29684 14636
rect 30028 14680 30068 14720
rect 29644 14176 29684 14216
rect 29932 14176 29972 14216
rect 29740 14008 29780 14048
rect 29836 13840 29876 13880
rect 29260 13420 29300 13460
rect 29260 13084 29300 13124
rect 30316 14596 30356 14636
rect 30220 13924 30260 13964
rect 30796 13756 30836 13796
rect 30412 13672 30452 13712
rect 30220 13336 30260 13376
rect 28972 13000 29012 13040
rect 28300 12328 28340 12368
rect 28492 12496 28532 12536
rect 29548 12916 29588 12956
rect 29068 12664 29108 12704
rect 29452 12664 29492 12704
rect 28972 12580 29012 12620
rect 28684 12412 28724 12452
rect 29164 12580 29204 12620
rect 29836 13168 29876 13208
rect 30028 13168 30068 13208
rect 29740 12916 29780 12956
rect 29356 12496 29396 12536
rect 29836 12496 29876 12536
rect 30796 13252 30836 13292
rect 30412 12916 30452 12956
rect 30700 13000 30740 13040
rect 30604 12832 30644 12872
rect 28492 12328 28532 12368
rect 29260 12328 29300 12368
rect 28108 12244 28148 12284
rect 28396 12244 28436 12284
rect 29068 11908 29108 11948
rect 29356 11740 29396 11780
rect 27436 11572 27476 11612
rect 29164 11488 29204 11528
rect 27340 11068 27380 11108
rect 27052 10984 27092 11024
rect 26668 10900 26708 10940
rect 26092 10732 26132 10772
rect 26380 10648 26420 10688
rect 26188 10480 26228 10520
rect 26284 10312 26324 10352
rect 26188 10144 26228 10184
rect 26956 10732 26996 10772
rect 27153 10312 27193 10352
rect 26284 9976 26324 10016
rect 25612 8548 25652 8588
rect 25612 8380 25652 8420
rect 25612 8212 25652 8252
rect 25900 8464 25940 8504
rect 25036 7876 25076 7916
rect 25324 7876 25364 7916
rect 25228 7708 25268 7748
rect 25767 7960 25807 8000
rect 26092 8632 26132 8672
rect 26188 8464 26228 8504
rect 25996 7960 26036 8000
rect 25516 7372 25556 7412
rect 25420 7288 25460 7328
rect 25036 7120 25076 7160
rect 25420 7120 25460 7160
rect 25228 7036 25268 7076
rect 25036 6868 25076 6908
rect 24940 6280 24980 6320
rect 25228 6448 25268 6488
rect 25420 6364 25460 6404
rect 24844 6112 24884 6152
rect 25132 6028 25172 6068
rect 24940 5776 24980 5816
rect 24268 5608 24308 5648
rect 24172 2752 24212 2792
rect 24844 4096 24884 4136
rect 25132 5608 25172 5648
rect 25324 5860 25364 5900
rect 25420 5608 25460 5648
rect 25324 5440 25364 5480
rect 25324 4600 25364 4640
rect 24556 2668 24596 2708
rect 23980 1996 24020 2036
rect 24460 2584 24500 2624
rect 25996 7288 26036 7328
rect 26764 9724 26804 9764
rect 26572 8632 26612 8672
rect 26380 8380 26420 8420
rect 26380 7288 26420 7328
rect 27052 10144 27092 10184
rect 29740 11908 29780 11948
rect 29644 11824 29684 11864
rect 29644 11488 29684 11528
rect 30220 12496 30260 12536
rect 30124 12412 30164 12452
rect 30412 12328 30452 12368
rect 30124 11824 30164 11864
rect 29356 11320 29396 11360
rect 30220 11572 30260 11612
rect 29260 11068 29300 11108
rect 28684 10816 28724 10856
rect 28876 10816 28916 10856
rect 29356 10984 29396 11024
rect 29260 10900 29300 10940
rect 29164 10480 29204 10520
rect 29644 10732 29684 10772
rect 29548 10480 29588 10520
rect 29836 10984 29876 11024
rect 30124 11152 30164 11192
rect 30124 10984 30164 11024
rect 30316 11152 30356 11192
rect 30028 10732 30068 10772
rect 27436 10144 27476 10184
rect 28204 10144 28244 10184
rect 27153 9976 27193 10016
rect 27340 9724 27380 9764
rect 27436 9640 27476 9680
rect 27820 9640 27860 9680
rect 28876 10060 28916 10100
rect 28588 9892 28628 9932
rect 27340 8884 27380 8924
rect 27340 8716 27380 8756
rect 27052 8632 27092 8672
rect 27244 8548 27284 8588
rect 27148 8464 27188 8504
rect 26668 7960 26708 8000
rect 26668 7792 26708 7832
rect 26572 7456 26612 7496
rect 26764 7624 26804 7664
rect 27724 8800 27764 8840
rect 27532 8380 27572 8420
rect 27244 7540 27284 7580
rect 27052 7456 27092 7496
rect 27153 7456 27193 7496
rect 26668 7120 26708 7160
rect 26668 6868 26708 6908
rect 25612 6112 25652 6152
rect 25612 5860 25652 5900
rect 25708 5776 25748 5816
rect 25612 5104 25652 5144
rect 25708 5020 25748 5060
rect 25996 6196 26036 6236
rect 25900 5104 25940 5144
rect 26188 6784 26228 6824
rect 26476 6784 26516 6824
rect 26572 6700 26612 6740
rect 26572 6532 26612 6572
rect 26860 7036 26900 7076
rect 26764 6616 26804 6656
rect 26284 6364 26324 6404
rect 25708 4096 25748 4136
rect 25612 4012 25652 4052
rect 25132 3676 25172 3716
rect 25516 3760 25556 3800
rect 25420 3340 25460 3380
rect 25804 3676 25844 3716
rect 25708 3340 25748 3380
rect 25228 2836 25268 2876
rect 25804 2836 25844 2876
rect 25420 2584 25460 2624
rect 26092 4936 26132 4976
rect 27207 7120 27247 7160
rect 27340 6784 27380 6824
rect 26668 6448 26708 6488
rect 26476 6280 26516 6320
rect 26668 6280 26708 6320
rect 26380 5104 26420 5144
rect 26284 5020 26324 5060
rect 27052 6448 27092 6488
rect 26956 6112 26996 6152
rect 26668 4936 26708 4976
rect 27052 5356 27092 5396
rect 27052 5104 27092 5144
rect 26188 4264 26228 4304
rect 26188 4096 26228 4136
rect 26092 4012 26132 4052
rect 25996 3928 26036 3968
rect 23980 1072 24020 1112
rect 25516 1072 25556 1112
rect 26668 4096 26708 4136
rect 26956 4936 26996 4976
rect 26572 3844 26612 3884
rect 26476 3760 26516 3800
rect 26860 3760 26900 3800
rect 26764 3676 26804 3716
rect 26380 3340 26420 3380
rect 26668 3424 26708 3464
rect 27628 5944 27668 5984
rect 27340 5356 27380 5396
rect 27340 5104 27380 5144
rect 27436 5020 27476 5060
rect 27340 4936 27380 4976
rect 27244 4852 27284 4892
rect 27148 4768 27188 4808
rect 27532 4936 27572 4976
rect 27628 4768 27668 4808
rect 27340 4096 27380 4136
rect 27244 3928 27284 3968
rect 27052 3172 27092 3212
rect 26572 2836 26612 2876
rect 26284 2584 26324 2624
rect 27244 2584 27284 2624
rect 27628 3760 27668 3800
rect 28300 9220 28340 9260
rect 28492 8800 28532 8840
rect 28396 8716 28436 8756
rect 27916 8632 27956 8672
rect 27916 8296 27956 8336
rect 28396 8296 28436 8336
rect 28876 9640 28916 9680
rect 28684 9472 28724 9512
rect 29164 10144 29204 10184
rect 29356 10144 29396 10184
rect 29452 9892 29492 9932
rect 28780 9304 28820 9344
rect 29068 9472 29108 9512
rect 29356 9472 29396 9512
rect 29644 10396 29684 10436
rect 30508 11152 30548 11192
rect 30700 10984 30740 11024
rect 30604 10900 30644 10940
rect 30124 10396 30164 10436
rect 29841 10144 29881 10184
rect 30412 10228 30452 10268
rect 30316 10060 30356 10100
rect 29740 9976 29780 10016
rect 29644 9724 29684 9764
rect 29644 9472 29684 9512
rect 29836 9892 29876 9932
rect 29548 9388 29588 9428
rect 29255 9304 29295 9344
rect 28972 9136 29012 9176
rect 29164 9136 29204 9176
rect 29068 8632 29108 8672
rect 30124 9724 30164 9764
rect 29932 9640 29972 9680
rect 29932 9472 29972 9512
rect 30604 10312 30644 10352
rect 30796 10228 30836 10268
rect 30316 9556 30356 9596
rect 30220 9052 30260 9092
rect 28876 8044 28916 8084
rect 28108 7792 28148 7832
rect 28012 7540 28052 7580
rect 28300 7960 28340 8000
rect 28492 7876 28532 7916
rect 29068 8212 29108 8252
rect 29836 8548 29876 8588
rect 29740 8296 29780 8336
rect 29260 7960 29300 8000
rect 28780 7792 28820 7832
rect 28780 7540 28820 7580
rect 28108 7120 28148 7160
rect 28204 6952 28244 6992
rect 28684 7456 28724 7496
rect 28492 6952 28532 6992
rect 28780 7204 28820 7244
rect 28684 7120 28724 7160
rect 29452 7708 29492 7748
rect 29356 7540 29396 7580
rect 28972 7456 29012 7496
rect 28876 7120 28916 7160
rect 29260 7288 29300 7328
rect 29836 7288 29876 7328
rect 29260 7120 29300 7160
rect 30028 8800 30068 8840
rect 30124 8548 30164 8588
rect 30220 8128 30260 8168
rect 30028 7792 30068 7832
rect 30281 7792 30321 7832
rect 29740 7120 29780 7160
rect 29452 7036 29492 7076
rect 29068 6532 29108 6572
rect 29452 6532 29492 6572
rect 28300 6364 28340 6404
rect 28204 6280 28244 6320
rect 27820 5440 27860 5480
rect 27916 5104 27956 5144
rect 27820 5020 27860 5060
rect 28780 6448 28820 6488
rect 28972 6364 29012 6404
rect 28684 5440 28724 5480
rect 28588 5104 28628 5144
rect 28204 4852 28244 4892
rect 28012 4768 28052 4808
rect 28204 4096 28244 4136
rect 27916 3928 27956 3968
rect 29164 6448 29204 6488
rect 29260 6196 29300 6236
rect 29740 6448 29780 6488
rect 29356 6028 29396 6068
rect 29068 4936 29108 4976
rect 29548 4600 29588 4640
rect 29740 4600 29780 4640
rect 28780 4096 28820 4136
rect 29260 4096 29300 4136
rect 28396 3844 28436 3884
rect 28300 3760 28340 3800
rect 29164 3760 29204 3800
rect 28492 3424 28532 3464
rect 28684 3424 28724 3464
rect 29740 4096 29780 4136
rect 28300 2836 28340 2876
rect 26668 1996 26708 2036
rect 30124 7120 30164 7160
rect 30220 7036 30260 7076
rect 30028 6196 30068 6236
rect 30220 5440 30260 5480
rect 30700 9556 30740 9596
rect 30508 9472 30548 9512
rect 30796 8716 30836 8756
rect 30700 8128 30740 8168
rect 30508 7960 30548 8000
rect 32332 20056 32372 20096
rect 31948 19804 31988 19844
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 33964 22492 34004 22532
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 35116 23332 35156 23372
rect 35884 24508 35924 24548
rect 36172 24508 36212 24548
rect 36652 26776 36692 26816
rect 37708 27196 37748 27236
rect 38188 27196 38228 27236
rect 36364 26608 36404 26648
rect 36460 25936 36500 25976
rect 36556 25768 36596 25808
rect 36652 25264 36692 25304
rect 36844 25936 36884 25976
rect 38284 26440 38324 26480
rect 36844 24256 36884 24296
rect 37324 24508 37364 24548
rect 35788 23752 35828 23792
rect 35788 23584 35828 23624
rect 35788 23416 35828 23456
rect 35692 23248 35732 23288
rect 35884 23164 35924 23204
rect 35308 23080 35348 23120
rect 35692 22996 35732 23036
rect 35020 22912 35060 22952
rect 35500 22828 35540 22868
rect 36748 23752 36788 23792
rect 36556 23248 36596 23288
rect 36460 23080 36500 23120
rect 37132 23332 37172 23372
rect 37228 23248 37268 23288
rect 36844 23080 36884 23120
rect 35980 22912 36020 22952
rect 37516 23752 37556 23792
rect 37708 23752 37748 23792
rect 37612 23584 37652 23624
rect 38764 27784 38804 27824
rect 38956 27784 38996 27824
rect 39148 27364 39188 27404
rect 39628 27364 39668 27404
rect 40012 28036 40052 28076
rect 39916 27616 39956 27656
rect 39820 27112 39860 27152
rect 38668 26944 38708 26984
rect 38476 26272 38516 26312
rect 38860 25684 38900 25724
rect 38476 25348 38516 25388
rect 40108 26776 40148 26816
rect 40300 26776 40340 26816
rect 39148 26188 39188 26228
rect 39340 26139 39380 26144
rect 39340 26104 39380 26139
rect 39820 26104 39860 26144
rect 40300 26104 40340 26144
rect 40492 32908 40532 32948
rect 40780 32824 40820 32864
rect 40588 32740 40628 32780
rect 40492 32236 40532 32276
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 41068 35092 41108 35132
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 41452 35092 41492 35132
rect 41260 35008 41300 35048
rect 41452 34588 41492 34628
rect 41164 34168 41204 34208
rect 41260 33748 41300 33788
rect 41068 32992 41108 33032
rect 41356 33160 41396 33200
rect 41452 32908 41492 32948
rect 41740 34168 41780 34208
rect 41836 33748 41876 33788
rect 41644 32740 41684 32780
rect 40972 32236 41012 32276
rect 41452 32152 41492 32192
rect 44428 35176 44468 35216
rect 45964 35176 46004 35216
rect 42892 34924 42932 34964
rect 42124 34420 42164 34460
rect 42220 34336 42260 34376
rect 42124 33748 42164 33788
rect 42220 33076 42260 33116
rect 42124 32992 42164 33032
rect 42028 32824 42068 32864
rect 42124 32656 42164 32696
rect 41932 32488 41972 32528
rect 42028 32404 42068 32444
rect 41932 32320 41972 32360
rect 41740 31144 41780 31184
rect 42508 31984 42548 32024
rect 40876 30220 40916 30260
rect 41260 30220 41300 30260
rect 41068 29716 41108 29756
rect 40876 29044 40916 29084
rect 41836 30220 41876 30260
rect 43756 34924 43796 34964
rect 43276 34672 43316 34712
rect 42892 34336 42932 34376
rect 42700 33580 42740 33620
rect 43372 34168 43412 34208
rect 43852 34168 43892 34208
rect 43084 33076 43124 33116
rect 42988 32992 43028 33032
rect 43084 32908 43124 32948
rect 42988 32824 43028 32864
rect 42700 32404 42740 32444
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 44140 33160 44180 33200
rect 44524 33160 44564 33200
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 43948 32824 43988 32864
rect 44716 32824 44756 32864
rect 43564 32740 43604 32780
rect 43276 32320 43316 32360
rect 43468 32236 43508 32276
rect 44140 32152 44180 32192
rect 43180 31984 43220 32024
rect 43084 31480 43124 31520
rect 42988 31396 43028 31436
rect 43372 31396 43412 31436
rect 43180 31312 43220 31352
rect 43084 31144 43124 31184
rect 43372 31144 43412 31184
rect 43180 30556 43220 30596
rect 42028 29968 42068 30008
rect 42316 29968 42356 30008
rect 42124 29800 42164 29840
rect 42988 29800 43028 29840
rect 41644 29716 41684 29756
rect 41836 29716 41876 29756
rect 41356 29632 41396 29672
rect 41260 29212 41300 29252
rect 40492 28288 40532 28328
rect 41644 29212 41684 29252
rect 43756 30976 43796 31016
rect 43564 30640 43604 30680
rect 43276 29716 43316 29756
rect 43468 29800 43508 29840
rect 42508 29632 42548 29672
rect 43372 29632 43412 29672
rect 43660 30388 43700 30428
rect 42892 29296 42932 29336
rect 41740 29044 41780 29084
rect 42220 28372 42260 28412
rect 40972 27700 41012 27740
rect 41740 27364 41780 27404
rect 42892 27952 42932 27992
rect 42892 27784 42932 27824
rect 44044 29212 44084 29252
rect 43276 29128 43316 29168
rect 43180 28456 43220 28496
rect 43084 28120 43124 28160
rect 43468 29044 43508 29084
rect 43372 28288 43412 28328
rect 43564 28372 43604 28412
rect 45964 32824 46004 32864
rect 46540 32656 46580 32696
rect 47020 32656 47060 32696
rect 45772 31900 45812 31940
rect 44620 31480 44660 31520
rect 45100 31480 45140 31520
rect 45676 31480 45716 31520
rect 44908 31312 44948 31352
rect 45100 31312 45140 31352
rect 44812 31228 44852 31268
rect 45580 31312 45620 31352
rect 45388 31228 45428 31268
rect 45868 31396 45908 31436
rect 46444 31396 46484 31436
rect 45676 31144 45716 31184
rect 45292 30976 45332 31016
rect 44812 30640 44852 30680
rect 45004 30640 45044 30680
rect 44908 30472 44948 30512
rect 44812 30388 44852 30428
rect 45100 29800 45140 29840
rect 46252 30640 46292 30680
rect 47116 32320 47156 32360
rect 47692 32320 47732 32360
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 47212 32152 47252 32192
rect 48076 32152 48116 32192
rect 47116 31900 47156 31940
rect 46924 31396 46964 31436
rect 46828 30724 46868 30764
rect 45292 30472 45332 30512
rect 45484 30388 45524 30428
rect 46444 30388 46484 30428
rect 43468 28120 43508 28160
rect 43660 28288 43700 28328
rect 45100 28372 45140 28412
rect 43372 27952 43412 27992
rect 41932 26776 41972 26816
rect 43180 27532 43220 27572
rect 42412 26776 42452 26816
rect 43084 26776 43124 26816
rect 40684 26440 40724 26480
rect 40876 26440 40916 26480
rect 41548 26440 41588 26480
rect 40588 26020 40628 26060
rect 39628 25768 39668 25808
rect 38956 25432 38996 25472
rect 40300 25432 40340 25472
rect 39916 25264 39956 25304
rect 40492 25264 40532 25304
rect 40780 26272 40820 26312
rect 40780 25852 40820 25892
rect 40684 25264 40724 25304
rect 38860 25180 38900 25220
rect 40012 25180 40052 25220
rect 38476 24676 38516 24716
rect 42220 26104 42260 26144
rect 41260 25516 41300 25556
rect 42892 26608 42932 26648
rect 42796 26104 42836 26144
rect 43276 26440 43316 26480
rect 43468 27364 43508 27404
rect 43372 26272 43412 26312
rect 43084 26104 43124 26144
rect 42508 25936 42548 25976
rect 41932 25348 41972 25388
rect 42316 25348 42356 25388
rect 41356 25264 41396 25304
rect 41740 25264 41780 25304
rect 40876 25180 40916 25220
rect 40972 24508 41012 24548
rect 38284 24256 38324 24296
rect 37900 23668 37940 23708
rect 37996 23500 38036 23540
rect 37420 23332 37460 23372
rect 37804 23332 37844 23372
rect 37804 23080 37844 23120
rect 37324 22996 37364 23036
rect 37996 22996 38036 23036
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 34348 21568 34388 21608
rect 36268 22156 36308 22196
rect 35692 22072 35732 22112
rect 33292 20896 33332 20936
rect 33292 20560 33332 20600
rect 33772 20560 33812 20600
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 34252 20224 34292 20264
rect 33100 19972 33140 20012
rect 33580 19972 33620 20012
rect 31852 18964 31892 19004
rect 31852 18796 31892 18836
rect 31564 18376 31604 18416
rect 31756 18376 31796 18416
rect 31756 17788 31796 17828
rect 31756 17368 31796 17408
rect 31660 16864 31700 16904
rect 31468 16360 31508 16400
rect 31372 15688 31412 15728
rect 32812 19216 32852 19256
rect 33004 19216 33044 19256
rect 32428 19132 32468 19172
rect 32044 18796 32084 18836
rect 32140 18040 32180 18080
rect 32044 17956 32084 17996
rect 32140 17872 32180 17912
rect 32044 17452 32084 17492
rect 31756 16360 31796 16400
rect 32332 17704 32372 17744
rect 32236 17452 32276 17492
rect 32044 16864 32084 16904
rect 32428 17200 32468 17240
rect 32428 17032 32468 17072
rect 31948 16696 31988 16736
rect 31948 16444 31988 16484
rect 31852 16192 31892 16232
rect 31660 15856 31700 15896
rect 31564 15772 31604 15812
rect 31564 15604 31604 15644
rect 31564 15268 31604 15308
rect 31468 14848 31508 14888
rect 31372 14680 31412 14720
rect 31660 14764 31700 14804
rect 31564 14512 31604 14552
rect 31468 13840 31508 13880
rect 31564 13336 31604 13376
rect 31372 13084 31412 13124
rect 31660 13084 31700 13124
rect 31468 12748 31508 12788
rect 31372 11656 31412 11696
rect 31852 15856 31892 15896
rect 32049 15520 32089 15560
rect 31948 15352 31988 15392
rect 31852 15268 31892 15308
rect 32332 16192 32372 16232
rect 32620 16780 32660 16820
rect 32423 15520 32463 15560
rect 33196 19804 33236 19844
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 33964 19552 34004 19592
rect 35116 19552 35156 19592
rect 33196 19048 33236 19088
rect 33676 18712 33716 18752
rect 33964 19216 34004 19256
rect 34060 19048 34100 19088
rect 33964 18964 34004 19004
rect 33868 18880 33908 18920
rect 33868 18544 33908 18584
rect 33580 18292 33620 18332
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 33388 17956 33428 17996
rect 33196 17788 33236 17828
rect 33100 17620 33140 17660
rect 34156 18964 34196 19004
rect 34252 18880 34292 18920
rect 34444 19216 34484 19256
rect 34348 18712 34388 18752
rect 34252 18460 34292 18500
rect 34156 17200 34196 17240
rect 33772 16780 33812 16820
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 32716 15856 32756 15896
rect 33100 16192 33140 16232
rect 33004 16108 33044 16148
rect 32908 16024 32948 16064
rect 33004 15856 33044 15896
rect 32908 15604 32948 15644
rect 32524 15268 32564 15308
rect 32428 15184 32468 15224
rect 32236 15016 32276 15056
rect 32140 14680 32180 14720
rect 33004 15184 33044 15224
rect 33100 15100 33140 15140
rect 32812 14764 32852 14804
rect 32524 14680 32564 14720
rect 32620 14428 32660 14468
rect 32812 14428 32852 14468
rect 32044 14344 32084 14384
rect 33004 14764 33044 14804
rect 32908 14176 32948 14216
rect 32332 14092 32372 14132
rect 31948 14008 31988 14048
rect 31756 12496 31796 12536
rect 32140 13840 32180 13880
rect 32236 13336 32276 13376
rect 32812 13336 32852 13376
rect 31852 12244 31892 12284
rect 32332 12244 32372 12284
rect 31756 11656 31796 11696
rect 32236 12160 32276 12200
rect 31852 11404 31892 11444
rect 31665 11236 31705 11276
rect 31564 11068 31604 11108
rect 31468 10984 31508 11024
rect 31372 10228 31412 10268
rect 31180 9892 31220 9932
rect 31468 8968 31508 9008
rect 33100 13252 33140 13292
rect 32524 12664 32564 12704
rect 33004 13168 33044 13208
rect 32908 12748 32948 12788
rect 32812 12580 32852 12620
rect 32716 11824 32756 11864
rect 32236 11068 32276 11108
rect 32044 10984 32084 11024
rect 33100 12664 33140 12704
rect 32716 11572 32756 11612
rect 34060 16444 34100 16484
rect 33292 16024 33332 16064
rect 33676 15604 33716 15644
rect 33772 15520 33812 15560
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 34060 15604 34100 15644
rect 34348 18208 34388 18248
rect 34348 17872 34388 17912
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 34540 18712 34580 18752
rect 35596 20224 35636 20264
rect 36940 21736 36980 21776
rect 35788 21568 35828 21608
rect 38188 23752 38228 23792
rect 38092 22660 38132 22700
rect 40492 24424 40532 24464
rect 41548 25180 41588 25220
rect 41452 24928 41492 24968
rect 41068 24256 41108 24296
rect 38956 23584 38996 23624
rect 38860 23332 38900 23372
rect 38572 22660 38612 22700
rect 37516 22240 37556 22280
rect 38764 22492 38804 22532
rect 37516 21736 37556 21776
rect 37324 21568 37364 21608
rect 37228 20980 37268 21020
rect 38668 22240 38708 22280
rect 35500 19552 35540 19592
rect 35404 19216 35444 19256
rect 35308 19048 35348 19088
rect 36364 19216 36404 19256
rect 34636 18292 34676 18332
rect 34924 18292 34964 18332
rect 34540 17872 34580 17912
rect 34732 17704 34772 17744
rect 35020 18208 35060 18248
rect 34636 17620 34676 17660
rect 35121 17788 35161 17828
rect 34444 17536 34484 17576
rect 34924 17536 34964 17576
rect 35121 17452 35161 17492
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 35116 17200 35156 17240
rect 35020 17116 35060 17156
rect 34348 16528 34388 16568
rect 34252 15940 34292 15980
rect 34636 16024 34676 16064
rect 34924 16024 34964 16064
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 34444 15772 34484 15812
rect 35020 15772 35060 15812
rect 34348 15688 34388 15728
rect 33868 14680 33908 14720
rect 33292 14344 33332 14384
rect 33676 14176 33716 14216
rect 33484 13840 33524 13880
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 33292 13168 33332 13208
rect 33388 13084 33428 13124
rect 33484 12664 33524 12704
rect 33196 12580 33236 12620
rect 33580 12580 33620 12620
rect 33292 12496 33332 12536
rect 34156 14680 34196 14720
rect 34156 13840 34196 13880
rect 34828 15688 34868 15728
rect 34636 15436 34676 15476
rect 34348 15184 34388 15224
rect 34444 14764 34484 14804
rect 34924 15520 34964 15560
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 34636 14176 34676 14216
rect 34348 14008 34388 14048
rect 35404 18544 35444 18584
rect 35596 18544 35636 18584
rect 35500 18040 35540 18080
rect 36076 18544 36116 18584
rect 35687 18292 35727 18332
rect 36076 17956 36116 17996
rect 35884 17872 35924 17912
rect 36172 17704 36212 17744
rect 36268 17620 36308 17660
rect 35692 17284 35732 17324
rect 35308 17116 35348 17156
rect 35596 15772 35636 15812
rect 35884 17284 35924 17324
rect 36308 17284 36348 17324
rect 36940 19216 36980 19256
rect 39340 22996 39380 23036
rect 40588 23500 40628 23540
rect 40012 22828 40052 22868
rect 39820 22660 39860 22700
rect 39052 22492 39092 22532
rect 38956 22240 38996 22280
rect 38956 21568 38996 21608
rect 39148 21568 39188 21608
rect 39052 20728 39092 20768
rect 38668 19888 38708 19928
rect 40204 22492 40244 22532
rect 39916 21316 39956 21356
rect 39916 20728 39956 20768
rect 40012 20056 40052 20096
rect 41068 23500 41108 23540
rect 41836 23752 41876 23792
rect 43180 25096 43220 25136
rect 43852 27700 43892 27740
rect 43948 27616 43988 27656
rect 43660 27532 43700 27572
rect 44524 28120 44564 28160
rect 45772 29800 45812 29840
rect 45964 29800 46004 29840
rect 45868 29632 45908 29672
rect 47500 31900 47540 31940
rect 47116 30640 47156 30680
rect 47884 31480 47924 31520
rect 48364 32152 48404 32192
rect 49804 32152 49844 32192
rect 48556 31900 48596 31940
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 48364 31480 48404 31520
rect 48268 31396 48308 31436
rect 47884 31228 47924 31268
rect 47692 30640 47732 30680
rect 47020 30388 47060 30428
rect 46924 29968 46964 30008
rect 46924 29716 46964 29756
rect 47308 29716 47348 29756
rect 47116 29632 47156 29672
rect 45004 27784 45044 27824
rect 45484 27784 45524 27824
rect 44428 27700 44468 27740
rect 44044 27280 44084 27320
rect 44140 26860 44180 26900
rect 45196 27616 45236 27656
rect 45100 27280 45140 27320
rect 44524 27028 44564 27068
rect 45004 26860 45044 26900
rect 43756 26608 43796 26648
rect 44332 26608 44372 26648
rect 43660 26272 43700 26312
rect 43468 25600 43508 25640
rect 43852 26272 43892 26312
rect 44236 26188 44276 26228
rect 44140 26104 44180 26144
rect 43852 25600 43892 25640
rect 45388 27616 45428 27656
rect 45388 27364 45428 27404
rect 45100 26356 45140 26396
rect 45292 26356 45332 26396
rect 44524 26272 44564 26312
rect 44428 26104 44468 26144
rect 44716 26104 44756 26144
rect 44908 26104 44948 26144
rect 44524 25600 44564 25640
rect 44140 25432 44180 25472
rect 44332 25432 44372 25472
rect 43852 25348 43892 25388
rect 44044 25096 44084 25136
rect 43948 24928 43988 24968
rect 44812 25432 44852 25472
rect 44620 25264 44660 25304
rect 45100 25348 45140 25388
rect 44716 25180 44756 25220
rect 44332 25096 44372 25136
rect 44236 24928 44276 24968
rect 43948 24676 43988 24716
rect 43372 23836 43412 23876
rect 44332 24844 44372 24884
rect 44524 24760 44564 24800
rect 44812 25012 44852 25052
rect 42988 23752 43028 23792
rect 40780 23416 40820 23456
rect 41740 23416 41780 23456
rect 40588 22828 40628 22868
rect 40396 22408 40436 22448
rect 40396 22156 40436 22196
rect 40300 21568 40340 21608
rect 40396 21400 40436 21440
rect 40492 21316 40532 21356
rect 41068 22744 41108 22784
rect 41932 23500 41972 23540
rect 41452 22996 41492 23036
rect 41356 22660 41396 22700
rect 40684 22492 40724 22532
rect 41164 21568 41204 21608
rect 43084 23248 43124 23288
rect 41548 22912 41588 22952
rect 42220 22912 42260 22952
rect 44044 23752 44084 23792
rect 43564 23080 43604 23120
rect 42700 22744 42740 22784
rect 42028 22660 42068 22700
rect 42316 22660 42356 22700
rect 41740 22576 41780 22616
rect 41644 22492 41684 22532
rect 42124 22492 42164 22532
rect 41548 22072 41588 22112
rect 41548 21568 41588 21608
rect 41452 21400 41492 21440
rect 40396 20056 40436 20096
rect 40300 19888 40340 19928
rect 37420 18628 37460 18668
rect 36556 17704 36596 17744
rect 37036 18040 37076 18080
rect 37324 18040 37364 18080
rect 37132 17956 37172 17996
rect 37228 17704 37268 17744
rect 36940 17620 36980 17660
rect 36844 17536 36884 17576
rect 36652 17452 36692 17492
rect 36460 17200 36500 17240
rect 36308 17116 36348 17156
rect 35788 16444 35828 16484
rect 35980 16444 36020 16484
rect 36556 16948 36596 16988
rect 36556 16780 36596 16820
rect 37228 17284 37268 17324
rect 37073 17116 37113 17156
rect 37804 18544 37844 18584
rect 37516 18208 37556 18248
rect 37420 17956 37460 17996
rect 37708 17872 37748 17912
rect 37516 17536 37556 17576
rect 37420 17452 37460 17492
rect 37324 17200 37364 17240
rect 37708 17536 37748 17576
rect 37900 18208 37940 18248
rect 37996 17704 38036 17744
rect 37324 16948 37364 16988
rect 36940 16612 36980 16652
rect 37420 16612 37460 16652
rect 36556 16444 36596 16484
rect 36748 16444 36788 16484
rect 37324 16444 37364 16484
rect 35980 16024 36020 16064
rect 35884 15772 35924 15812
rect 35596 15604 35636 15644
rect 35692 15520 35732 15560
rect 35404 15436 35444 15476
rect 35596 15352 35636 15392
rect 36268 16024 36308 16064
rect 36076 15688 36116 15728
rect 36172 15604 36212 15644
rect 36460 16192 36500 16232
rect 36652 16360 36692 16400
rect 37036 16360 37076 16400
rect 36556 15856 36596 15896
rect 36364 15772 36404 15812
rect 36076 15100 36116 15140
rect 36268 15352 36308 15392
rect 36364 15184 36404 15224
rect 36268 15100 36308 15140
rect 36556 15520 36596 15560
rect 36556 15268 36596 15308
rect 36844 15688 36884 15728
rect 37708 16864 37748 16904
rect 37612 16780 37652 16820
rect 37516 16528 37556 16568
rect 37516 16108 37556 16148
rect 37132 16024 37172 16064
rect 37324 15856 37364 15896
rect 37804 15856 37844 15896
rect 36940 15604 36980 15644
rect 37324 15604 37364 15644
rect 36748 15520 36788 15560
rect 39724 19216 39764 19256
rect 40684 19216 40724 19256
rect 38860 19048 38900 19088
rect 38764 17872 38804 17912
rect 38572 17704 38612 17744
rect 38572 17536 38612 17576
rect 38188 16864 38228 16904
rect 38092 16192 38132 16232
rect 37996 16060 38036 16064
rect 37996 16024 38036 16060
rect 38188 15940 38228 15980
rect 38092 15688 38132 15728
rect 36940 15436 36980 15476
rect 36844 15352 36884 15392
rect 37036 15352 37076 15392
rect 37132 14932 37172 14972
rect 37900 15520 37940 15560
rect 38188 15604 38228 15644
rect 37708 15436 37748 15476
rect 37612 15352 37652 15392
rect 37516 15184 37556 15224
rect 36268 14512 36308 14552
rect 36844 14512 36884 14552
rect 36076 14008 36116 14048
rect 36748 13756 36788 13796
rect 35212 13252 35252 13292
rect 34444 13168 34484 13208
rect 34060 12748 34100 12788
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 33196 11656 33236 11696
rect 33484 11908 33524 11948
rect 33580 11824 33620 11864
rect 33772 11824 33812 11864
rect 33100 11236 33140 11276
rect 32524 11068 32564 11108
rect 32716 11068 32756 11108
rect 32428 10984 32468 11024
rect 32524 10816 32564 10856
rect 32716 10564 32756 10604
rect 32812 10396 32852 10436
rect 32332 10312 32372 10352
rect 32236 10144 32276 10184
rect 32812 10228 32852 10268
rect 32332 9556 32372 9596
rect 31852 9472 31892 9512
rect 31564 8800 31604 8840
rect 31948 8968 31988 9008
rect 30892 7876 30932 7916
rect 30796 7624 30836 7664
rect 30604 7540 30644 7580
rect 31084 8464 31124 8504
rect 31468 8464 31508 8504
rect 31660 8632 31700 8672
rect 31660 8464 31700 8504
rect 31180 8044 31220 8084
rect 30988 7624 31028 7664
rect 31180 7876 31220 7916
rect 31948 8632 31988 8672
rect 31852 8380 31892 8420
rect 31852 8212 31892 8252
rect 31468 7960 31508 8000
rect 31372 7876 31412 7916
rect 31660 7792 31700 7832
rect 31564 7708 31604 7748
rect 31276 7372 31316 7412
rect 30892 7120 30932 7160
rect 31948 7960 31988 8000
rect 31756 7708 31796 7748
rect 31948 7708 31988 7748
rect 31756 7540 31796 7580
rect 31660 7204 31700 7244
rect 31564 6448 31604 6488
rect 31084 5860 31124 5900
rect 30892 5608 30932 5648
rect 31564 5608 31604 5648
rect 31852 6532 31892 6572
rect 30220 4852 30260 4892
rect 29356 3004 29396 3044
rect 29836 3004 29876 3044
rect 27724 1996 27764 2036
rect 28780 2584 28820 2624
rect 27532 1912 27572 1952
rect 28684 1912 28724 1952
rect 29452 2836 29492 2876
rect 29836 2836 29876 2876
rect 30508 4096 30548 4136
rect 31372 4096 31412 4136
rect 30412 3424 30452 3464
rect 33004 10816 33044 10856
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 33196 10312 33236 10352
rect 32908 10144 32948 10184
rect 33100 10144 33140 10184
rect 32620 10060 32660 10100
rect 33004 10060 33044 10100
rect 33004 9556 33044 9596
rect 32620 9472 32660 9512
rect 33100 9472 33140 9512
rect 32620 9136 32660 9176
rect 32428 8716 32468 8756
rect 32140 8464 32180 8504
rect 33004 9136 33044 9176
rect 32716 8632 32756 8672
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 33484 8800 33524 8840
rect 33196 8548 33236 8588
rect 32908 8464 32948 8504
rect 33100 8464 33140 8504
rect 33676 8669 33716 8672
rect 33676 8632 33716 8669
rect 32812 8380 32852 8420
rect 32620 8296 32660 8336
rect 32140 7876 32180 7916
rect 32428 7960 32468 8000
rect 32620 7876 32660 7916
rect 32620 7540 32660 7580
rect 32812 7540 32852 7580
rect 32332 7372 32372 7412
rect 32524 7372 32564 7412
rect 32044 7288 32084 7328
rect 32332 7120 32372 7160
rect 32044 6448 32084 6488
rect 32332 4096 32372 4136
rect 33484 8464 33524 8504
rect 33292 8212 33332 8252
rect 33484 7960 33524 8000
rect 33772 8044 33812 8084
rect 33772 7792 33812 7832
rect 33100 6868 33140 6908
rect 33676 7708 33716 7748
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 33484 7372 33524 7412
rect 33772 7372 33812 7412
rect 33964 11908 34004 11948
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 34540 12664 34580 12704
rect 35020 12580 35060 12620
rect 34732 11824 34772 11864
rect 35020 11824 35060 11864
rect 34252 11656 34292 11696
rect 33964 9388 34004 9428
rect 34348 11236 34388 11276
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 34348 10396 34388 10436
rect 34348 10228 34388 10268
rect 34732 10984 34772 11024
rect 34828 10816 34868 10856
rect 35020 10396 35060 10436
rect 35404 11320 35444 11360
rect 35404 11152 35444 11192
rect 35308 11068 35348 11108
rect 35500 10984 35540 11024
rect 35212 10732 35252 10772
rect 35500 10816 35540 10856
rect 35308 10228 35348 10268
rect 36268 12580 36308 12620
rect 35788 11320 35828 11360
rect 37324 14680 37364 14720
rect 37900 15184 37940 15224
rect 37612 14680 37652 14720
rect 38092 15100 38132 15140
rect 39436 17788 39476 17828
rect 38476 16780 38516 16820
rect 38380 16360 38420 16400
rect 38572 16192 38612 16232
rect 38380 15940 38420 15980
rect 38380 15268 38420 15308
rect 38188 14680 38228 14720
rect 37804 14008 37844 14048
rect 38092 13756 38132 13796
rect 38668 15856 38708 15896
rect 38668 15520 38708 15560
rect 38956 16192 38996 16232
rect 38668 15100 38708 15140
rect 38860 15100 38900 15140
rect 38764 13924 38804 13964
rect 38956 12664 38996 12704
rect 37612 12580 37652 12620
rect 39148 16024 39188 16064
rect 39244 15940 39284 15980
rect 39628 17032 39668 17072
rect 40012 19048 40052 19088
rect 40012 17704 40052 17744
rect 39916 17620 39956 17660
rect 42028 22240 42068 22280
rect 43180 22828 43220 22868
rect 42892 22660 42932 22700
rect 44908 24928 44948 24968
rect 45388 25516 45428 25556
rect 45100 24760 45140 24800
rect 45580 27532 45620 27572
rect 45580 27364 45620 27404
rect 45676 26188 45716 26228
rect 45676 25684 45716 25724
rect 46252 28120 46292 28160
rect 46156 27868 46196 27908
rect 45964 27616 46004 27656
rect 46540 28288 46580 28328
rect 47116 28876 47156 28916
rect 47020 28288 47060 28328
rect 46636 28204 46676 28244
rect 46828 28204 46868 28244
rect 46732 28120 46772 28160
rect 47788 30220 47828 30260
rect 47788 29968 47828 30008
rect 47788 28876 47828 28916
rect 47500 28456 47540 28496
rect 48268 30472 48308 30512
rect 48076 30220 48116 30260
rect 48268 30220 48308 30260
rect 48172 29716 48212 29756
rect 48076 29296 48116 29336
rect 47884 28288 47924 28328
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 49132 30724 49172 30764
rect 48460 30640 48500 30680
rect 48940 30472 48980 30512
rect 49996 30472 50036 30512
rect 48556 30388 48596 30428
rect 49612 30388 49652 30428
rect 48940 30304 48980 30344
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 48364 29800 48404 29840
rect 51244 30472 51284 30512
rect 50188 30304 50228 30344
rect 49420 29800 49460 29840
rect 50380 29800 50420 29840
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 49228 29296 49268 29336
rect 49036 29128 49076 29168
rect 50572 29128 50612 29168
rect 51628 30388 51668 30428
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 48940 28876 48980 28916
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 48268 28372 48308 28412
rect 48748 28288 48788 28328
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 47308 28120 47348 28160
rect 48652 28120 48692 28160
rect 47020 27868 47060 27908
rect 46444 27784 46484 27824
rect 46636 27784 46676 27824
rect 45964 27364 46004 27404
rect 46828 26776 46868 26816
rect 45868 25432 45908 25472
rect 45772 25264 45812 25304
rect 46156 25684 46196 25724
rect 45772 24928 45812 24968
rect 45676 24844 45716 24884
rect 44908 24592 44948 24632
rect 45004 24424 45044 24464
rect 44140 22996 44180 23036
rect 44428 22996 44468 23036
rect 43756 22912 43796 22952
rect 44620 23752 44660 23792
rect 44908 23752 44948 23792
rect 44812 23248 44852 23288
rect 44812 22912 44852 22952
rect 41932 22072 41972 22112
rect 43276 21400 43316 21440
rect 44524 21652 44564 21692
rect 44428 21568 44468 21608
rect 41644 20980 41684 21020
rect 44716 22324 44756 22364
rect 44716 21736 44756 21776
rect 45772 24676 45812 24716
rect 45676 24592 45716 24632
rect 45004 23248 45044 23288
rect 45004 22912 45044 22952
rect 46348 25852 46388 25892
rect 46252 25180 46292 25220
rect 46252 25012 46292 25052
rect 46732 25852 46772 25892
rect 46540 24928 46580 24968
rect 46348 24844 46388 24884
rect 46252 24760 46292 24800
rect 46540 24760 46580 24800
rect 46348 23500 46388 23540
rect 45772 23164 45812 23204
rect 45484 22576 45524 22616
rect 46156 23080 46196 23120
rect 46156 22660 46196 22700
rect 46540 22492 46580 22532
rect 46828 25432 46868 25472
rect 48652 27784 48692 27824
rect 47212 27700 47252 27740
rect 47116 27448 47156 27488
rect 47020 27364 47060 27404
rect 47596 27532 47636 27572
rect 47500 27448 47540 27488
rect 47692 27448 47732 27488
rect 47212 27280 47252 27320
rect 47308 26440 47348 26480
rect 48172 27616 48212 27656
rect 48268 27448 48308 27488
rect 48172 27280 48212 27320
rect 47980 27028 48020 27068
rect 47788 26692 47828 26732
rect 48172 26440 48212 26480
rect 47692 26356 47732 26396
rect 47212 26104 47252 26144
rect 47596 26104 47636 26144
rect 48076 26104 48116 26144
rect 48940 27616 48980 27656
rect 49228 27532 49268 27572
rect 48460 27448 48500 27488
rect 48748 27448 48788 27488
rect 49132 27448 49172 27488
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 48844 27028 48884 27068
rect 49036 27364 49076 27404
rect 48940 26860 48980 26900
rect 49996 28204 50036 28244
rect 49804 28120 49844 28160
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 49996 27784 50036 27824
rect 49612 26860 49652 26900
rect 50860 27784 50900 27824
rect 51628 28120 51668 28160
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 50668 27532 50708 27572
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 50188 26776 50228 26816
rect 50380 26776 50420 26816
rect 50860 26776 50900 26816
rect 49324 26692 49364 26732
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 49228 26272 49268 26312
rect 49804 26272 49844 26312
rect 48364 26104 48404 26144
rect 47500 25936 47540 25976
rect 47404 25012 47444 25052
rect 46924 24844 46964 24884
rect 48748 25936 48788 25976
rect 47500 24760 47540 24800
rect 47212 24592 47252 24632
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 47692 25180 47732 25220
rect 48460 25180 48500 25220
rect 48172 25012 48212 25052
rect 48268 24676 48308 24716
rect 49132 25936 49172 25976
rect 49036 25852 49076 25892
rect 48172 24508 48212 24548
rect 48940 24676 48980 24716
rect 48652 24508 48692 24548
rect 49900 26104 49940 26144
rect 50092 25852 50132 25892
rect 51628 26608 51668 26648
rect 52012 26608 52052 26648
rect 50956 26104 50996 26144
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 50764 26020 50804 26060
rect 51148 26020 51188 26060
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 48268 24172 48308 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 49516 23920 49556 23960
rect 47404 23164 47444 23204
rect 47020 22660 47060 22700
rect 46924 22408 46964 22448
rect 45388 21736 45428 21776
rect 47980 23080 48020 23120
rect 49132 23584 49172 23624
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 49132 23248 49172 23288
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 51820 24592 51860 24632
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 50764 23920 50804 23960
rect 49900 23080 49940 23120
rect 50668 23080 50708 23120
rect 51148 23584 51188 23624
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 47692 21652 47732 21692
rect 45484 21568 45524 21608
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 41068 17704 41108 17744
rect 40492 17032 40532 17072
rect 39820 16276 39860 16316
rect 39148 15184 39188 15224
rect 40300 16192 40340 16232
rect 40492 16192 40532 16232
rect 40108 16024 40148 16064
rect 40108 15604 40148 15644
rect 39820 15184 39860 15224
rect 39532 15100 39572 15140
rect 40972 16108 41012 16148
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 42316 16108 42356 16148
rect 41260 16024 41300 16064
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 40492 14932 40532 14972
rect 41548 14932 41588 14972
rect 39244 13924 39284 13964
rect 40396 14680 40436 14720
rect 39820 14008 39860 14048
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 39340 13336 39380 13376
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 36076 11572 36116 11612
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 37804 11572 37844 11612
rect 37516 11404 37556 11444
rect 37708 11404 37748 11444
rect 36076 11068 36116 11108
rect 35884 10732 35924 10772
rect 35692 10396 35732 10436
rect 35788 10228 35828 10268
rect 35020 9976 35060 10016
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 34252 9472 34292 9512
rect 34156 9220 34196 9260
rect 34444 9640 34484 9680
rect 34444 9388 34484 9428
rect 34545 9388 34585 9428
rect 34060 9052 34100 9092
rect 34348 9052 34388 9092
rect 34540 9052 34580 9092
rect 33964 8632 34004 8672
rect 34156 8716 34196 8756
rect 35212 9640 35252 9680
rect 35596 9976 35636 10016
rect 35212 9472 35252 9512
rect 36652 10144 36692 10184
rect 38092 10984 38132 11024
rect 38188 10312 38228 10352
rect 37900 10144 37940 10184
rect 35596 9304 35636 9344
rect 35404 9220 35444 9260
rect 34828 9052 34868 9092
rect 35116 9052 35156 9092
rect 34636 8884 34676 8924
rect 34252 8128 34292 8168
rect 34060 8044 34100 8084
rect 34828 8548 34868 8588
rect 35308 8632 35348 8672
rect 37324 9472 37364 9512
rect 36268 8716 36308 8756
rect 38764 11656 38804 11696
rect 39532 11656 39572 11696
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 38380 10144 38420 10184
rect 38668 10144 38708 10184
rect 38860 10060 38900 10100
rect 39820 10060 39860 10100
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 37996 9388 38036 9428
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 37996 8884 38036 8924
rect 39052 8884 39092 8924
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 35020 8296 35060 8336
rect 34348 7960 34388 8000
rect 34060 7708 34100 7748
rect 33964 7372 34004 7412
rect 33868 7120 33908 7160
rect 34348 7540 34388 7580
rect 33868 6448 33908 6488
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 33196 5608 33236 5648
rect 33484 5440 33524 5480
rect 35692 8128 35732 8168
rect 34924 7120 34964 7160
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 33964 5692 34004 5732
rect 34636 6448 34676 6488
rect 36652 8296 36692 8336
rect 36364 7792 36404 7832
rect 35212 7540 35252 7580
rect 34732 5692 34772 5732
rect 35020 5692 35060 5732
rect 35308 6616 35348 6656
rect 36748 7960 36788 8000
rect 37420 8044 37460 8084
rect 35788 7288 35828 7328
rect 36172 6616 36212 6656
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 37804 7960 37844 8000
rect 36940 7288 36980 7328
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 38092 7204 38132 7244
rect 38956 7204 38996 7244
rect 37228 7036 37268 7076
rect 37900 7036 37940 7076
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 34060 5524 34100 5564
rect 34636 5524 34676 5564
rect 35308 5608 35348 5648
rect 34444 5440 34484 5480
rect 34924 5440 34964 5480
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 30892 2584 30932 2624
rect 31852 2584 31892 2624
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 25612 904 25652 944
rect 25996 904 26036 944
rect 26476 904 26516 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37568 80 37588
rect 0 37528 268 37568
rect 308 37528 317 37568
rect 27427 37528 27436 37568
rect 27476 37528 27820 37568
rect 27860 37528 27869 37568
rect 0 37508 80 37528
rect 27619 37360 27628 37400
rect 27668 37360 31756 37400
rect 31796 37360 31805 37400
rect 26563 37192 26572 37232
rect 26612 37192 27532 37232
rect 27572 37192 27581 37232
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 30979 36856 30988 36896
rect 31028 36856 31660 36896
rect 31700 36856 31709 36896
rect 32707 36772 32716 36812
rect 32756 36772 33292 36812
rect 33332 36772 33341 36812
rect 0 36729 80 36748
rect 0 36728 125 36729
rect 0 36688 76 36728
rect 116 36688 125 36728
rect 26275 36688 26284 36728
rect 26324 36688 28684 36728
rect 28724 36688 28972 36728
rect 29012 36688 29021 36728
rect 0 36687 125 36688
rect 0 36668 80 36687
rect 13123 36520 13132 36560
rect 13172 36520 13900 36560
rect 13940 36520 13949 36560
rect 24451 36520 24460 36560
rect 24500 36520 25900 36560
rect 25940 36520 25949 36560
rect 31363 36520 31372 36560
rect 31412 36520 32044 36560
rect 32084 36520 35596 36560
rect 35636 36520 35645 36560
rect 36451 36520 36460 36560
rect 36500 36520 37612 36560
rect 37652 36520 37661 36560
rect 12643 36436 12652 36476
rect 12692 36436 13228 36476
rect 13268 36436 13277 36476
rect 25987 36436 25996 36476
rect 26036 36436 27052 36476
rect 27092 36436 27101 36476
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 29155 36100 29164 36140
rect 29204 36100 29452 36140
rect 29492 36100 30796 36140
rect 30836 36100 30845 36140
rect 0 35828 80 35908
rect 18979 35848 18988 35888
rect 19028 35848 19564 35888
rect 19604 35848 19613 35888
rect 35203 35848 35212 35888
rect 35252 35848 36076 35888
rect 36116 35848 36125 35888
rect 11875 35680 11884 35720
rect 11924 35680 12940 35720
rect 12980 35680 12989 35720
rect 26851 35680 26860 35720
rect 26900 35680 28012 35720
rect 28052 35680 28061 35720
rect 30595 35680 30604 35720
rect 30644 35680 32044 35720
rect 32084 35680 32093 35720
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 24067 35512 24076 35552
rect 24116 35512 25612 35552
rect 25652 35512 25661 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 25795 35428 25804 35468
rect 25844 35428 27724 35468
rect 27764 35428 27773 35468
rect 39139 35428 39148 35468
rect 39188 35428 40396 35468
rect 40436 35428 40445 35468
rect 21763 35344 21772 35384
rect 21812 35344 21821 35384
rect 25603 35344 25612 35384
rect 25652 35344 25996 35384
rect 26036 35344 26045 35384
rect 29731 35344 29740 35384
rect 29780 35344 30508 35384
rect 30548 35344 30557 35384
rect 34723 35344 34732 35384
rect 34772 35344 35404 35384
rect 35444 35344 35453 35384
rect 37603 35344 37612 35384
rect 37652 35344 40300 35384
rect 40340 35344 40349 35384
rect 21772 35300 21812 35344
rect 5923 35260 5932 35300
rect 5972 35260 6988 35300
rect 7028 35260 7037 35300
rect 12931 35260 12940 35300
rect 12980 35260 13612 35300
rect 13652 35260 13661 35300
rect 13987 35260 13996 35300
rect 14036 35260 16780 35300
rect 16820 35260 16829 35300
rect 21187 35260 21196 35300
rect 21236 35260 21812 35300
rect 23395 35260 23404 35300
rect 23444 35260 26380 35300
rect 26420 35260 26429 35300
rect 28291 35260 28300 35300
rect 28340 35260 30892 35300
rect 30932 35260 30941 35300
rect 32515 35260 32524 35300
rect 32564 35260 33196 35300
rect 33236 35260 33245 35300
rect 34627 35260 34636 35300
rect 34676 35260 35308 35300
rect 35348 35260 35357 35300
rect 36067 35260 36076 35300
rect 36116 35260 38284 35300
rect 38324 35260 38333 35300
rect 38659 35260 38668 35300
rect 38708 35260 39052 35300
rect 39092 35260 39101 35300
rect 4771 35176 4780 35216
rect 4820 35176 5356 35216
rect 5396 35176 5405 35216
rect 8803 35176 8812 35216
rect 8852 35176 10924 35216
rect 10964 35176 10973 35216
rect 14275 35176 14284 35216
rect 14324 35176 14333 35216
rect 14563 35176 14572 35216
rect 14612 35176 16492 35216
rect 16532 35176 16541 35216
rect 17155 35176 17164 35216
rect 17204 35176 18124 35216
rect 18164 35176 18316 35216
rect 18356 35176 18365 35216
rect 26083 35176 26092 35216
rect 26132 35176 26764 35216
rect 26804 35176 26813 35216
rect 29827 35176 29836 35216
rect 29876 35176 30412 35216
rect 30452 35176 30461 35216
rect 30508 35176 32236 35216
rect 32276 35176 32285 35216
rect 32899 35176 32908 35216
rect 32948 35176 33964 35216
rect 34004 35176 34540 35216
rect 34580 35176 34589 35216
rect 34636 35176 35404 35216
rect 35444 35176 35788 35216
rect 35828 35176 35837 35216
rect 35971 35176 35980 35216
rect 36020 35176 36460 35216
rect 36500 35176 36509 35216
rect 38083 35176 38092 35216
rect 38132 35176 40972 35216
rect 41012 35176 41021 35216
rect 44419 35176 44428 35216
rect 44468 35176 45964 35216
rect 46004 35176 46013 35216
rect 5443 35092 5452 35132
rect 5492 35092 6028 35132
rect 6068 35092 6077 35132
rect 8899 35092 8908 35132
rect 8948 35092 9196 35132
rect 9236 35092 9245 35132
rect 11683 35092 11692 35132
rect 11732 35092 13804 35132
rect 13844 35092 13853 35132
rect 0 34988 80 35068
rect 12067 35008 12076 35048
rect 12116 35008 13708 35048
rect 13748 35008 13757 35048
rect 14284 34964 14324 35176
rect 30508 35132 30548 35176
rect 34636 35132 34676 35176
rect 14371 35092 14380 35132
rect 14420 35092 16300 35132
rect 16340 35092 17644 35132
rect 17684 35092 17693 35132
rect 25699 35092 25708 35132
rect 25748 35092 26476 35132
rect 26516 35092 26860 35132
rect 26900 35092 28340 35132
rect 30115 35092 30124 35132
rect 30164 35092 30548 35132
rect 31459 35092 31468 35132
rect 31508 35092 33100 35132
rect 33140 35092 33149 35132
rect 34339 35092 34348 35132
rect 34388 35092 34676 35132
rect 35020 35092 36940 35132
rect 36980 35092 36989 35132
rect 38947 35092 38956 35132
rect 38996 35092 40300 35132
rect 40340 35092 41068 35132
rect 41108 35092 41452 35132
rect 41492 35092 41501 35132
rect 28300 35048 28340 35092
rect 35020 35048 35060 35092
rect 16099 35008 16108 35048
rect 16148 35008 17452 35048
rect 17492 35008 17501 35048
rect 27043 35008 27052 35048
rect 27092 35008 27916 35048
rect 27956 35008 27965 35048
rect 28291 35008 28300 35048
rect 28340 35008 29644 35048
rect 29684 35008 29693 35048
rect 31267 35008 31276 35048
rect 31316 35008 35060 35048
rect 35107 35008 35116 35048
rect 35156 35008 36364 35048
rect 36404 35008 36413 35048
rect 40675 35008 40684 35048
rect 40724 35008 41260 35048
rect 41300 35008 41309 35048
rect 6499 34924 6508 34964
rect 6548 34924 7660 34964
rect 7700 34924 8812 34964
rect 8852 34924 8861 34964
rect 11587 34924 11596 34964
rect 11636 34924 13132 34964
rect 13172 34924 13181 34964
rect 13228 34924 16684 34964
rect 16724 34924 16733 34964
rect 30883 34924 30892 34964
rect 30932 34924 32236 34964
rect 32276 34924 32285 34964
rect 42883 34924 42892 34964
rect 42932 34924 43756 34964
rect 43796 34924 43805 34964
rect 13132 34796 13172 34924
rect 13228 34880 13268 34924
rect 13219 34840 13228 34880
rect 13268 34840 13277 34880
rect 14083 34840 14092 34880
rect 14132 34840 14668 34880
rect 14708 34840 14717 34880
rect 14851 34840 14860 34880
rect 14900 34840 15820 34880
rect 15860 34840 17068 34880
rect 17108 34840 19276 34880
rect 19316 34840 19325 34880
rect 30499 34840 30508 34880
rect 30548 34840 34252 34880
rect 34292 34840 34301 34880
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 13132 34756 14380 34796
rect 14420 34756 14429 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 31651 34672 31660 34712
rect 31700 34672 32140 34712
rect 32180 34672 32189 34712
rect 39427 34672 39436 34712
rect 39476 34672 43276 34712
rect 43316 34672 43325 34712
rect 6019 34588 6028 34628
rect 6068 34588 8332 34628
rect 8372 34588 8381 34628
rect 9091 34588 9100 34628
rect 9140 34588 11884 34628
rect 11924 34588 11933 34628
rect 13123 34588 13132 34628
rect 13172 34588 15436 34628
rect 15476 34588 18508 34628
rect 18548 34588 18557 34628
rect 27523 34588 27532 34628
rect 27572 34588 28204 34628
rect 28244 34588 29164 34628
rect 29204 34588 29213 34628
rect 31747 34588 31756 34628
rect 31796 34588 32524 34628
rect 32564 34588 32573 34628
rect 39043 34588 39052 34628
rect 39092 34588 39532 34628
rect 39572 34588 39581 34628
rect 40867 34588 40876 34628
rect 40916 34588 41452 34628
rect 41492 34588 41501 34628
rect 9667 34504 9676 34544
rect 9716 34504 10444 34544
rect 10484 34504 10493 34544
rect 14947 34504 14956 34544
rect 14996 34504 16972 34544
rect 17012 34504 17021 34544
rect 17731 34504 17740 34544
rect 17780 34504 19372 34544
rect 19412 34504 21196 34544
rect 21236 34504 21245 34544
rect 26851 34504 26860 34544
rect 26900 34504 30220 34544
rect 30260 34504 31948 34544
rect 31988 34504 31997 34544
rect 38467 34504 38476 34544
rect 38516 34504 39628 34544
rect 39668 34504 39677 34544
rect 11683 34420 11692 34460
rect 11732 34420 12172 34460
rect 12212 34420 13228 34460
rect 13268 34420 13277 34460
rect 18115 34420 18124 34460
rect 18164 34420 19028 34460
rect 25411 34420 25420 34460
rect 25460 34420 26284 34460
rect 26324 34420 26333 34460
rect 28483 34420 28492 34460
rect 28532 34420 29836 34460
rect 29876 34420 30700 34460
rect 30740 34420 31276 34460
rect 31316 34420 32276 34460
rect 37603 34420 37612 34460
rect 37652 34420 39476 34460
rect 40099 34420 40108 34460
rect 40148 34420 40588 34460
rect 40628 34420 42124 34460
rect 42164 34420 42173 34460
rect 18988 34376 19028 34420
rect 32236 34376 32276 34420
rect 39436 34376 39476 34420
rect 3619 34336 3628 34376
rect 3668 34336 5644 34376
rect 5684 34336 5693 34376
rect 10243 34336 10252 34376
rect 10292 34336 10828 34376
rect 10868 34336 10877 34376
rect 11203 34336 11212 34376
rect 11252 34336 15628 34376
rect 15668 34336 15677 34376
rect 16195 34336 16204 34376
rect 16244 34336 16588 34376
rect 16628 34336 16972 34376
rect 17012 34336 17021 34376
rect 18979 34336 18988 34376
rect 19028 34336 19037 34376
rect 20035 34336 20044 34376
rect 20084 34336 21004 34376
rect 21044 34336 22636 34376
rect 22676 34336 24556 34376
rect 24596 34336 25900 34376
rect 25940 34336 25949 34376
rect 32227 34336 32236 34376
rect 32276 34336 32428 34376
rect 32468 34336 32477 34376
rect 33763 34336 33772 34376
rect 33812 34336 35020 34376
rect 35060 34336 35069 34376
rect 39436 34336 40204 34376
rect 40244 34336 40492 34376
rect 40532 34336 40541 34376
rect 42211 34336 42220 34376
rect 42260 34336 42892 34376
rect 42932 34336 42941 34376
rect 11491 34252 11500 34292
rect 11540 34252 11980 34292
rect 12020 34252 12556 34292
rect 12596 34252 13036 34292
rect 13076 34252 13085 34292
rect 13603 34252 13612 34292
rect 13652 34252 13900 34292
rect 13940 34252 13949 34292
rect 14851 34252 14860 34292
rect 14900 34252 15724 34292
rect 15764 34252 15773 34292
rect 27907 34252 27916 34292
rect 27956 34252 30988 34292
rect 31028 34252 31037 34292
rect 36931 34252 36940 34292
rect 36980 34252 39436 34292
rect 39476 34252 39485 34292
rect 39907 34252 39916 34292
rect 39956 34252 40780 34292
rect 40820 34252 40829 34292
rect 0 34148 80 34228
rect 9379 34168 9388 34208
rect 9428 34168 11404 34208
rect 11444 34168 11453 34208
rect 11980 34168 12364 34208
rect 12404 34168 14764 34208
rect 14804 34168 14813 34208
rect 18883 34168 18892 34208
rect 18932 34168 19180 34208
rect 19220 34168 19229 34208
rect 21283 34168 21292 34208
rect 21332 34168 23788 34208
rect 23828 34168 25036 34208
rect 25076 34168 25996 34208
rect 26036 34168 26045 34208
rect 29923 34168 29932 34208
rect 29972 34168 30700 34208
rect 30740 34168 30749 34208
rect 35779 34168 35788 34208
rect 35828 34168 36844 34208
rect 36884 34168 36893 34208
rect 38563 34168 38572 34208
rect 38612 34168 38860 34208
rect 38900 34168 39052 34208
rect 39092 34168 39340 34208
rect 39380 34168 40012 34208
rect 40052 34168 40061 34208
rect 41155 34168 41164 34208
rect 41204 34168 41740 34208
rect 41780 34168 41789 34208
rect 43363 34168 43372 34208
rect 43412 34168 43852 34208
rect 43892 34168 43901 34208
rect 11980 34124 12020 34168
rect 30700 34124 30740 34168
rect 4963 34084 4972 34124
rect 5012 34084 5836 34124
rect 5876 34084 5885 34124
rect 10627 34084 10636 34124
rect 10676 34084 11692 34124
rect 11732 34084 11741 34124
rect 11971 34084 11980 34124
rect 12020 34084 12029 34124
rect 30700 34084 35212 34124
rect 35252 34084 35261 34124
rect 28483 34040 28541 34041
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 4867 34000 4876 34040
rect 4916 34000 4925 34040
rect 5731 34000 5740 34040
rect 5780 34000 6316 34040
rect 6356 34000 6365 34040
rect 8323 34000 8332 34040
rect 8372 34000 8908 34040
rect 8948 34000 8957 34040
rect 13219 34000 13228 34040
rect 13268 34000 13612 34040
rect 13652 34000 13661 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 25507 34000 25516 34040
rect 25556 34000 26188 34040
rect 26228 34000 26764 34040
rect 26804 34000 26813 34040
rect 28483 34000 28492 34040
rect 28532 34000 28588 34040
rect 28628 34000 28637 34040
rect 29443 34000 29452 34040
rect 29492 34000 30412 34040
rect 30452 34000 30461 34040
rect 33187 34000 33196 34040
rect 33236 34000 33772 34040
rect 33812 34000 34348 34040
rect 34388 34000 34397 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 37315 34000 37324 34040
rect 37364 34000 38380 34040
rect 38420 34000 39244 34040
rect 39284 34000 39293 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 4876 33956 4916 34000
rect 28483 33999 28541 34000
rect 3235 33916 3244 33956
rect 3284 33916 6700 33956
rect 6740 33916 7468 33956
rect 7508 33916 7517 33956
rect 29059 33916 29068 33956
rect 29108 33916 30028 33956
rect 30068 33916 31756 33956
rect 31796 33916 31805 33956
rect 35491 33916 35500 33956
rect 35540 33916 36364 33956
rect 36404 33916 36413 33956
rect 5059 33832 5068 33872
rect 5108 33832 8620 33872
rect 8660 33832 9004 33872
rect 9044 33832 9580 33872
rect 9620 33832 9629 33872
rect 11779 33832 11788 33872
rect 11828 33832 12460 33872
rect 12500 33832 12509 33872
rect 36451 33832 36460 33872
rect 36500 33832 38860 33872
rect 38900 33832 39532 33872
rect 39572 33832 39581 33872
rect 5155 33748 5164 33788
rect 5204 33748 5972 33788
rect 6403 33748 6412 33788
rect 6452 33748 6988 33788
rect 7028 33748 7037 33788
rect 17251 33748 17260 33788
rect 17300 33748 17932 33788
rect 17972 33748 18700 33788
rect 18740 33748 19372 33788
rect 19412 33748 19660 33788
rect 19700 33748 19709 33788
rect 40003 33748 40012 33788
rect 40052 33748 41260 33788
rect 41300 33748 41836 33788
rect 41876 33748 42124 33788
rect 42164 33748 42173 33788
rect 5932 33704 5972 33748
rect 4675 33664 4684 33704
rect 4724 33664 5356 33704
rect 5396 33664 5405 33704
rect 5923 33664 5932 33704
rect 5972 33664 6604 33704
rect 6644 33664 9196 33704
rect 9236 33664 9245 33704
rect 10531 33664 10540 33704
rect 10580 33664 11212 33704
rect 11252 33664 12940 33704
rect 12980 33664 13996 33704
rect 14036 33664 14045 33704
rect 15235 33664 15244 33704
rect 15284 33664 15916 33704
rect 15956 33664 15965 33704
rect 18019 33664 18028 33704
rect 18068 33664 19180 33704
rect 19220 33664 19229 33704
rect 19276 33664 20332 33704
rect 20372 33664 20381 33704
rect 21091 33664 21100 33704
rect 21140 33664 21868 33704
rect 21908 33664 21917 33704
rect 23587 33664 23596 33704
rect 23636 33664 24172 33704
rect 24212 33664 24221 33704
rect 27715 33664 27724 33704
rect 27764 33664 28012 33704
rect 28052 33664 30604 33704
rect 30644 33664 30653 33704
rect 31843 33664 31852 33704
rect 31892 33664 32140 33704
rect 32180 33664 32189 33704
rect 34339 33664 34348 33704
rect 34388 33664 34397 33704
rect 36643 33664 36652 33704
rect 36692 33664 37820 33704
rect 38563 33664 38572 33704
rect 38612 33664 38956 33704
rect 38996 33664 40108 33704
rect 40148 33664 40157 33704
rect 19276 33620 19316 33664
rect 34348 33620 34388 33664
rect 37780 33620 37820 33664
rect 2755 33580 2764 33620
rect 2804 33580 4396 33620
rect 4436 33580 6028 33620
rect 6068 33580 7180 33620
rect 7220 33580 7229 33620
rect 18892 33580 19316 33620
rect 20035 33580 20044 33620
rect 20084 33580 20180 33620
rect 20803 33580 20812 33620
rect 20852 33580 21580 33620
rect 21620 33580 21629 33620
rect 27619 33580 27628 33620
rect 27668 33580 27820 33620
rect 27860 33580 29000 33620
rect 30403 33580 30412 33620
rect 30452 33580 31084 33620
rect 31124 33580 33676 33620
rect 33716 33580 33725 33620
rect 33859 33580 33868 33620
rect 33908 33580 34252 33620
rect 34292 33580 34301 33620
rect 34348 33580 37516 33620
rect 37556 33580 37565 33620
rect 37780 33580 38092 33620
rect 38132 33580 42700 33620
rect 42740 33580 42749 33620
rect 18892 33536 18932 33580
rect 4195 33496 4204 33536
rect 4244 33496 4972 33536
rect 5012 33496 6412 33536
rect 6452 33496 6461 33536
rect 18883 33496 18892 33536
rect 18932 33496 18941 33536
rect 20140 33452 20180 33580
rect 28960 33536 29000 33580
rect 23683 33496 23692 33536
rect 23732 33496 24364 33536
rect 24404 33496 24413 33536
rect 28960 33496 29068 33536
rect 29108 33496 29117 33536
rect 36547 33496 36556 33536
rect 36596 33496 39916 33536
rect 39956 33496 39965 33536
rect 14851 33412 14860 33452
rect 14900 33412 15244 33452
rect 15284 33412 15293 33452
rect 20140 33412 21484 33452
rect 21524 33412 21676 33452
rect 21716 33412 23788 33452
rect 23828 33412 23837 33452
rect 26275 33412 26284 33452
rect 26324 33412 26956 33452
rect 26996 33412 27005 33452
rect 30883 33412 30892 33452
rect 30932 33412 31276 33452
rect 31316 33412 31325 33452
rect 37891 33412 37900 33452
rect 37940 33412 38284 33452
rect 38324 33412 38333 33452
rect 0 33308 80 33388
rect 6403 33328 6412 33368
rect 6452 33328 7852 33368
rect 7892 33328 11500 33368
rect 11540 33328 11549 33368
rect 15331 33328 15340 33368
rect 15380 33328 19468 33368
rect 19508 33328 19517 33368
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 30307 33244 30316 33284
rect 30356 33244 31468 33284
rect 31508 33244 31517 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 6883 33160 6892 33200
rect 6932 33160 8236 33200
rect 8276 33160 8285 33200
rect 19171 33160 19180 33200
rect 19220 33160 23212 33200
rect 23252 33160 25612 33200
rect 25652 33160 25661 33200
rect 41347 33160 41356 33200
rect 41396 33160 44140 33200
rect 44180 33160 44524 33200
rect 44564 33160 44573 33200
rect 1315 33076 1324 33116
rect 1364 33076 4492 33116
rect 4532 33076 4541 33116
rect 4771 33076 4780 33116
rect 4820 33076 9868 33116
rect 9908 33076 9917 33116
rect 11107 33076 11116 33116
rect 11156 33076 13516 33116
rect 13556 33076 13565 33116
rect 13795 33076 13804 33116
rect 13844 33076 15052 33116
rect 15092 33076 15101 33116
rect 19651 33076 19660 33116
rect 19700 33076 20332 33116
rect 20372 33076 20381 33116
rect 27427 33076 27436 33116
rect 27476 33076 27724 33116
rect 27764 33076 28588 33116
rect 28628 33076 28637 33116
rect 30307 33076 30316 33116
rect 30356 33076 30700 33116
rect 30740 33076 30749 33116
rect 42211 33076 42220 33116
rect 42260 33076 43084 33116
rect 43124 33076 43133 33116
rect 2371 32992 2380 33032
rect 2420 32992 3724 33032
rect 3764 32992 3773 33032
rect 7075 32992 7084 33032
rect 7124 32992 8140 33032
rect 8180 32992 8189 33032
rect 18115 32992 18124 33032
rect 18164 32992 19372 33032
rect 19412 32992 19421 33032
rect 21379 32992 21388 33032
rect 21428 32992 22156 33032
rect 22196 32992 22205 33032
rect 26083 32992 26092 33032
rect 26132 32992 28396 33032
rect 28436 32992 28684 33032
rect 28724 32992 28733 33032
rect 41059 32992 41068 33032
rect 41108 32992 42124 33032
rect 42164 32992 42173 33032
rect 42979 32992 42988 33032
rect 43028 32992 43068 33032
rect 42988 32948 43028 32992
rect 1987 32908 1996 32948
rect 2036 32908 3052 32948
rect 3092 32908 3101 32948
rect 6115 32908 6124 32948
rect 6164 32908 7564 32948
rect 7604 32908 7613 32948
rect 9283 32908 9292 32948
rect 9332 32908 12748 32948
rect 12788 32908 12797 32948
rect 16771 32908 16780 32948
rect 16820 32908 17260 32948
rect 17300 32908 18604 32948
rect 18644 32908 18653 32948
rect 26179 32908 26188 32948
rect 26228 32908 26860 32948
rect 26900 32908 27532 32948
rect 27572 32908 29164 32948
rect 29204 32908 30796 32948
rect 30836 32908 30845 32948
rect 36259 32908 36268 32948
rect 36308 32908 37228 32948
rect 37268 32908 37820 32948
rect 40291 32908 40300 32948
rect 40340 32908 40492 32948
rect 40532 32908 40541 32948
rect 41443 32908 41452 32948
rect 41492 32908 43084 32948
rect 43124 32908 43133 32948
rect 37780 32864 37820 32908
rect 2179 32824 2188 32864
rect 2228 32824 2860 32864
rect 2900 32824 4012 32864
rect 4052 32824 4684 32864
rect 4724 32824 5452 32864
rect 5492 32824 6604 32864
rect 6644 32824 6892 32864
rect 6932 32824 6941 32864
rect 7075 32824 7084 32864
rect 7124 32824 8044 32864
rect 8084 32824 8093 32864
rect 8227 32824 8236 32864
rect 8276 32824 9004 32864
rect 9044 32824 9053 32864
rect 9667 32824 9676 32864
rect 9716 32824 9964 32864
rect 10004 32824 10444 32864
rect 10484 32824 11116 32864
rect 11156 32824 11165 32864
rect 12643 32824 12652 32864
rect 12692 32824 13804 32864
rect 13844 32824 13853 32864
rect 14755 32824 14764 32864
rect 14804 32824 15244 32864
rect 15284 32824 15293 32864
rect 18211 32824 18220 32864
rect 18260 32824 19468 32864
rect 19508 32824 19517 32864
rect 19747 32824 19756 32864
rect 19796 32824 20428 32864
rect 20468 32824 20477 32864
rect 25603 32824 25612 32864
rect 25652 32824 25996 32864
rect 26036 32824 26045 32864
rect 27811 32824 27820 32864
rect 27860 32824 27869 32864
rect 28483 32824 28492 32864
rect 28532 32824 29068 32864
rect 29108 32824 29117 32864
rect 29347 32824 29356 32864
rect 29396 32824 29548 32864
rect 29588 32824 29597 32864
rect 30211 32824 30220 32864
rect 30260 32824 32332 32864
rect 32372 32824 32381 32864
rect 37780 32824 39148 32864
rect 39188 32824 39197 32864
rect 40771 32824 40780 32864
rect 40820 32824 42028 32864
rect 42068 32824 42988 32864
rect 43028 32824 43948 32864
rect 43988 32824 44716 32864
rect 44756 32824 45964 32864
rect 46004 32824 46013 32864
rect 27820 32780 27860 32824
rect 2659 32740 2668 32780
rect 2708 32740 4204 32780
rect 4244 32740 4253 32780
rect 4963 32740 4972 32780
rect 5012 32740 5356 32780
rect 5396 32740 5405 32780
rect 6499 32740 6508 32780
rect 6548 32740 7276 32780
rect 7316 32740 7325 32780
rect 8419 32740 8428 32780
rect 8468 32740 8812 32780
rect 8852 32740 8861 32780
rect 14947 32740 14956 32780
rect 14996 32740 15436 32780
rect 15476 32740 15485 32780
rect 19363 32740 19372 32780
rect 19412 32740 20140 32780
rect 20180 32740 20189 32780
rect 25699 32740 25708 32780
rect 25748 32740 26380 32780
rect 26420 32740 26429 32780
rect 27628 32740 27860 32780
rect 40579 32740 40588 32780
rect 40628 32740 41644 32780
rect 41684 32740 41693 32780
rect 42124 32740 43564 32780
rect 43604 32740 43613 32780
rect 27628 32696 27668 32740
rect 42124 32696 42164 32740
rect 5635 32656 5644 32696
rect 5684 32656 6316 32696
rect 6356 32656 6365 32696
rect 7651 32656 7660 32696
rect 7700 32656 7948 32696
rect 7988 32656 7997 32696
rect 12931 32656 12940 32696
rect 12980 32656 13996 32696
rect 14036 32656 14860 32696
rect 14900 32656 14909 32696
rect 19555 32656 19564 32696
rect 19604 32656 22540 32696
rect 22580 32656 22589 32696
rect 27619 32656 27628 32696
rect 27668 32656 27677 32696
rect 27811 32656 27820 32696
rect 27860 32656 28108 32696
rect 28148 32656 28157 32696
rect 42115 32656 42124 32696
rect 42164 32656 42173 32696
rect 46531 32656 46540 32696
rect 46580 32656 47020 32696
rect 47060 32656 47069 32696
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 27139 32488 27148 32528
rect 27188 32488 27532 32528
rect 27572 32488 27916 32528
rect 27956 32488 27965 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 40195 32488 40204 32528
rect 40244 32488 41932 32528
rect 41972 32488 41981 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 42019 32404 42028 32444
rect 42068 32404 42700 32444
rect 42740 32404 42749 32444
rect 18115 32320 18124 32360
rect 18164 32320 20044 32360
rect 20084 32320 21196 32360
rect 21236 32320 21245 32360
rect 27235 32320 27244 32360
rect 27284 32320 28012 32360
rect 28052 32320 28061 32360
rect 32419 32320 32428 32360
rect 32468 32320 36076 32360
rect 36116 32320 36125 32360
rect 37603 32320 37612 32360
rect 37652 32320 37804 32360
rect 37844 32320 37853 32360
rect 41923 32320 41932 32360
rect 41972 32320 43276 32360
rect 43316 32320 43325 32360
rect 47107 32320 47116 32360
rect 47156 32320 47692 32360
rect 47732 32320 47741 32360
rect 30499 32236 30508 32276
rect 30548 32236 40492 32276
rect 40532 32236 40541 32276
rect 40963 32236 40972 32276
rect 41012 32236 43468 32276
rect 43508 32236 43517 32276
rect 4771 32192 4829 32193
rect 3715 32152 3724 32192
rect 3764 32152 4780 32192
rect 4820 32152 4829 32192
rect 6211 32152 6220 32192
rect 6260 32152 6700 32192
rect 6740 32152 6749 32192
rect 8131 32152 8140 32192
rect 8180 32152 10828 32192
rect 10868 32152 11020 32192
rect 11060 32152 11069 32192
rect 15331 32152 15340 32192
rect 15380 32152 16108 32192
rect 16148 32152 16157 32192
rect 18019 32152 18028 32192
rect 18068 32152 19948 32192
rect 19988 32152 20180 32192
rect 24835 32152 24844 32192
rect 24884 32152 25996 32192
rect 26036 32152 26045 32192
rect 26371 32152 26380 32192
rect 26420 32152 27820 32192
rect 27860 32152 27869 32192
rect 32035 32152 32044 32192
rect 32084 32152 33484 32192
rect 33524 32152 33533 32192
rect 34915 32152 34924 32192
rect 34964 32152 36268 32192
rect 36308 32152 36317 32192
rect 38467 32152 38476 32192
rect 38516 32152 39244 32192
rect 39284 32152 39293 32192
rect 41443 32152 41452 32192
rect 41492 32152 44140 32192
rect 44180 32152 44189 32192
rect 47203 32152 47212 32192
rect 47252 32152 48076 32192
rect 48116 32152 48125 32192
rect 48355 32152 48364 32192
rect 48404 32152 49804 32192
rect 49844 32152 49853 32192
rect 4771 32151 4829 32152
rect 14371 32068 14380 32108
rect 14420 32068 15820 32108
rect 15860 32068 18412 32108
rect 18452 32068 19412 32108
rect 19372 32024 19412 32068
rect 20140 32024 20180 32152
rect 32131 32068 32140 32108
rect 32180 32068 32332 32108
rect 32372 32068 33196 32108
rect 33236 32068 33245 32108
rect 15907 31984 15916 32024
rect 15956 31984 16588 32024
rect 16628 31984 17932 32024
rect 17972 31984 17981 32024
rect 19363 31984 19372 32024
rect 19412 31984 19421 32024
rect 20140 31984 21292 32024
rect 21332 31984 21341 32024
rect 42499 31984 42508 32024
rect 42548 31984 43180 32024
rect 43220 31984 43229 32024
rect 3523 31900 3532 31940
rect 3572 31900 4108 31940
rect 4148 31900 4157 31940
rect 11683 31900 11692 31940
rect 11732 31900 13804 31940
rect 13844 31900 13853 31940
rect 45763 31900 45772 31940
rect 45812 31900 47116 31940
rect 47156 31900 47165 31940
rect 47491 31900 47500 31940
rect 47540 31900 48556 31940
rect 48596 31900 48605 31940
rect 11011 31816 11020 31856
rect 11060 31816 12364 31856
rect 12404 31816 12413 31856
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 9667 31732 9676 31772
rect 9716 31732 10828 31772
rect 10868 31732 11212 31772
rect 11252 31732 11261 31772
rect 11320 31732 12268 31772
rect 12308 31732 12317 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31628 80 31708
rect 11320 31688 11360 31732
rect 10435 31648 10444 31688
rect 10484 31648 11360 31688
rect 16771 31648 16780 31688
rect 16820 31648 17644 31688
rect 17684 31648 17693 31688
rect 13123 31604 13181 31605
rect 13123 31564 13132 31604
rect 13172 31564 13420 31604
rect 13460 31564 14764 31604
rect 14804 31564 14813 31604
rect 23491 31564 23500 31604
rect 23540 31564 27628 31604
rect 27668 31564 27677 31604
rect 13123 31563 13181 31564
rect 2083 31480 2092 31520
rect 2132 31480 3436 31520
rect 3476 31480 3485 31520
rect 4003 31480 4012 31520
rect 4052 31480 4588 31520
rect 4628 31480 4637 31520
rect 4771 31480 4780 31520
rect 4820 31480 4829 31520
rect 6787 31480 6796 31520
rect 6836 31480 7660 31520
rect 7700 31480 7709 31520
rect 8323 31480 8332 31520
rect 8372 31480 8812 31520
rect 8852 31480 8861 31520
rect 11683 31480 11692 31520
rect 11732 31480 12844 31520
rect 12884 31480 12893 31520
rect 13219 31480 13228 31520
rect 13268 31480 13708 31520
rect 13748 31480 14956 31520
rect 14996 31480 15005 31520
rect 15619 31480 15628 31520
rect 15668 31480 16684 31520
rect 16724 31480 16733 31520
rect 19747 31480 19756 31520
rect 19796 31480 20332 31520
rect 20372 31480 20381 31520
rect 24547 31480 24556 31520
rect 24596 31480 25228 31520
rect 25268 31480 25277 31520
rect 27331 31480 27340 31520
rect 27380 31480 27820 31520
rect 27860 31480 27869 31520
rect 28003 31480 28012 31520
rect 28052 31480 28588 31520
rect 28628 31480 28637 31520
rect 31939 31480 31948 31520
rect 31988 31480 32428 31520
rect 32468 31480 32852 31520
rect 32899 31480 32908 31520
rect 32948 31480 33580 31520
rect 33620 31480 33629 31520
rect 34435 31480 34444 31520
rect 34484 31480 34493 31520
rect 43075 31480 43084 31520
rect 43124 31480 44620 31520
rect 44660 31480 44669 31520
rect 45091 31480 45100 31520
rect 45140 31480 45676 31520
rect 45716 31480 45725 31520
rect 47875 31480 47884 31520
rect 47924 31480 48364 31520
rect 48404 31480 48413 31520
rect 4780 31436 4820 31480
rect 32812 31436 32852 31480
rect 34444 31436 34484 31480
rect 2659 31396 2668 31436
rect 2708 31396 4820 31436
rect 6883 31396 6892 31436
rect 6932 31396 8716 31436
rect 8756 31396 8765 31436
rect 12163 31396 12172 31436
rect 12212 31396 12460 31436
rect 12500 31396 13036 31436
rect 13076 31396 13085 31436
rect 13315 31396 13324 31436
rect 13364 31396 16492 31436
rect 16532 31396 16541 31436
rect 32812 31396 33428 31436
rect 33475 31396 33484 31436
rect 33524 31396 34484 31436
rect 42979 31396 42988 31436
rect 43028 31396 43372 31436
rect 43412 31396 43421 31436
rect 44908 31396 45868 31436
rect 45908 31396 46444 31436
rect 46484 31396 46924 31436
rect 46964 31396 48268 31436
rect 48308 31396 48317 31436
rect 4099 31312 4108 31352
rect 4148 31312 4972 31352
rect 5012 31312 5021 31352
rect 1219 31144 1228 31184
rect 1268 31144 4588 31184
rect 4628 31144 4637 31184
rect 8332 31016 8372 31396
rect 33388 31352 33428 31396
rect 44908 31352 44948 31396
rect 10051 31312 10060 31352
rect 10100 31312 10924 31352
rect 10964 31312 10973 31352
rect 12259 31312 12268 31352
rect 12308 31312 12748 31352
rect 12788 31312 12797 31352
rect 13603 31312 13612 31352
rect 13652 31312 15244 31352
rect 15284 31312 15293 31352
rect 16003 31312 16012 31352
rect 16052 31312 17740 31352
rect 17780 31312 18220 31352
rect 18260 31312 18269 31352
rect 25699 31312 25708 31352
rect 25748 31312 26380 31352
rect 26420 31312 26429 31352
rect 27043 31312 27052 31352
rect 27092 31312 28300 31352
rect 28340 31312 28349 31352
rect 31171 31312 31180 31352
rect 31220 31312 33292 31352
rect 33332 31312 33341 31352
rect 33388 31312 33908 31352
rect 33955 31312 33964 31352
rect 34004 31312 35116 31352
rect 35156 31312 35165 31352
rect 43171 31312 43180 31352
rect 43220 31312 44908 31352
rect 44948 31312 44957 31352
rect 45091 31312 45100 31352
rect 45140 31312 45580 31352
rect 45620 31312 45629 31352
rect 8707 31228 8716 31268
rect 8756 31228 9676 31268
rect 9716 31228 9725 31268
rect 12547 31228 12556 31268
rect 12596 31228 13900 31268
rect 13940 31228 13949 31268
rect 26179 31228 26188 31268
rect 26228 31228 28396 31268
rect 28436 31228 28445 31268
rect 33868 31184 33908 31312
rect 44803 31228 44812 31268
rect 44852 31228 45388 31268
rect 45428 31228 45437 31268
rect 46600 31228 47884 31268
rect 47924 31228 47933 31268
rect 46600 31184 46640 31228
rect 24163 31144 24172 31184
rect 24212 31144 24748 31184
rect 24788 31144 26380 31184
rect 26420 31144 26429 31184
rect 26851 31144 26860 31184
rect 26900 31144 27340 31184
rect 27380 31144 27916 31184
rect 27956 31144 27965 31184
rect 30883 31144 30892 31184
rect 30932 31144 31372 31184
rect 31412 31144 31564 31184
rect 31604 31144 31613 31184
rect 31747 31144 31756 31184
rect 31796 31144 32236 31184
rect 32276 31144 32285 31184
rect 33859 31144 33868 31184
rect 33908 31144 35404 31184
rect 35444 31144 35453 31184
rect 40291 31144 40300 31184
rect 40340 31144 41740 31184
rect 41780 31144 43084 31184
rect 43124 31144 43133 31184
rect 43363 31144 43372 31184
rect 43412 31144 45676 31184
rect 45716 31144 46640 31184
rect 26860 31100 26900 31144
rect 26083 31060 26092 31100
rect 26132 31060 26900 31100
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 8323 30976 8332 31016
rect 8372 30976 8381 31016
rect 13027 30976 13036 31016
rect 13076 30976 13612 31016
rect 13652 30976 13661 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 31267 30976 31276 31016
rect 31316 30976 31564 31016
rect 31604 30976 34252 31016
rect 34292 30976 34301 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 39235 30976 39244 31016
rect 39284 30976 43756 31016
rect 43796 30976 45292 31016
rect 45332 30976 45341 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 30595 30892 30604 30932
rect 30644 30892 30988 30932
rect 31028 30892 31037 30932
rect 0 30788 80 30868
rect 11011 30808 11020 30848
rect 11060 30808 11884 30848
rect 11924 30808 12020 30848
rect 13315 30808 13324 30848
rect 13364 30808 14092 30848
rect 14132 30808 14141 30848
rect 25027 30808 25036 30848
rect 25076 30808 25420 30848
rect 25460 30808 27628 30848
rect 27668 30808 27677 30848
rect 28579 30808 28588 30848
rect 28628 30808 29000 30848
rect 29539 30808 29548 30848
rect 29588 30808 31084 30848
rect 31124 30808 31133 30848
rect 38659 30808 38668 30848
rect 38708 30808 39532 30848
rect 39572 30808 39581 30848
rect 6979 30640 6988 30680
rect 7028 30640 7180 30680
rect 7220 30640 7229 30680
rect 9667 30640 9676 30680
rect 9716 30640 9725 30680
rect 10915 30640 10924 30680
rect 10964 30640 11500 30680
rect 11540 30640 11549 30680
rect 11683 30640 11692 30680
rect 11732 30640 11884 30680
rect 11924 30640 11933 30680
rect 9676 30596 9716 30640
rect 3715 30556 3724 30596
rect 3764 30556 6604 30596
rect 6644 30556 7468 30596
rect 7508 30556 7517 30596
rect 9676 30556 11116 30596
rect 11156 30556 11165 30596
rect 4771 30512 4829 30513
rect 11980 30512 12020 30808
rect 28960 30764 29000 30808
rect 13507 30724 13516 30764
rect 13556 30724 16108 30764
rect 16148 30724 16157 30764
rect 25708 30724 27724 30764
rect 27764 30724 27773 30764
rect 28960 30724 30604 30764
rect 30644 30724 31180 30764
rect 31220 30724 31229 30764
rect 46819 30724 46828 30764
rect 46868 30724 49132 30764
rect 49172 30724 49181 30764
rect 25708 30680 25748 30724
rect 13795 30640 13804 30680
rect 13844 30640 14476 30680
rect 14516 30640 14525 30680
rect 19651 30640 19660 30680
rect 19700 30640 20044 30680
rect 20084 30640 20093 30680
rect 24163 30640 24172 30680
rect 24212 30640 25708 30680
rect 25748 30640 25757 30680
rect 26947 30640 26956 30680
rect 26996 30640 30028 30680
rect 30068 30640 32428 30680
rect 32468 30640 32477 30680
rect 33859 30640 33868 30680
rect 33908 30640 34252 30680
rect 34292 30640 34301 30680
rect 34435 30640 34444 30680
rect 34484 30640 35308 30680
rect 35348 30640 35357 30680
rect 36643 30640 36652 30680
rect 36692 30640 37036 30680
rect 37076 30640 37085 30680
rect 37219 30640 37228 30680
rect 37268 30640 37708 30680
rect 37748 30640 37757 30680
rect 38179 30640 38188 30680
rect 38228 30640 38237 30680
rect 38371 30640 38380 30680
rect 38420 30640 39052 30680
rect 39092 30640 39101 30680
rect 43555 30640 43564 30680
rect 43604 30640 44812 30680
rect 44852 30640 44861 30680
rect 44995 30640 45004 30680
rect 45044 30640 46252 30680
rect 46292 30640 47116 30680
rect 47156 30640 47165 30680
rect 47683 30640 47692 30680
rect 47732 30640 48460 30680
rect 48500 30640 48509 30680
rect 38188 30596 38228 30640
rect 45004 30596 45044 30640
rect 16291 30556 16300 30596
rect 16340 30556 17836 30596
rect 17876 30556 17885 30596
rect 34339 30556 34348 30596
rect 34388 30556 35500 30596
rect 35540 30556 35980 30596
rect 36020 30556 36029 30596
rect 38188 30556 38764 30596
rect 38804 30556 39340 30596
rect 39380 30556 43180 30596
rect 43220 30556 45044 30596
rect 4675 30472 4684 30512
rect 4724 30472 4780 30512
rect 4820 30472 4829 30512
rect 6115 30472 6124 30512
rect 6164 30472 8428 30512
rect 8468 30472 11924 30512
rect 11971 30472 11980 30512
rect 12020 30472 12029 30512
rect 30307 30472 30316 30512
rect 30356 30472 30892 30512
rect 30932 30472 30941 30512
rect 31363 30472 31372 30512
rect 31412 30472 36172 30512
rect 36212 30472 36221 30512
rect 39139 30472 39148 30512
rect 39188 30472 40300 30512
rect 40340 30472 40349 30512
rect 44899 30472 44908 30512
rect 44948 30472 45292 30512
rect 45332 30472 45341 30512
rect 48259 30472 48268 30512
rect 48308 30472 48940 30512
rect 48980 30472 48989 30512
rect 49987 30472 49996 30512
rect 50036 30472 51244 30512
rect 51284 30472 51293 30512
rect 4771 30471 4829 30472
rect 11884 30428 11924 30472
rect 10915 30388 10924 30428
rect 10964 30388 11404 30428
rect 11444 30388 11453 30428
rect 11884 30388 13132 30428
rect 13172 30388 14188 30428
rect 14228 30388 16108 30428
rect 16148 30388 16157 30428
rect 25603 30388 25612 30428
rect 25652 30388 26476 30428
rect 26516 30388 26525 30428
rect 28483 30388 28492 30428
rect 28532 30388 29932 30428
rect 29972 30388 29981 30428
rect 32995 30388 33004 30428
rect 33044 30388 34444 30428
rect 34484 30388 34493 30428
rect 43651 30388 43660 30428
rect 43700 30388 44812 30428
rect 44852 30388 44861 30428
rect 45475 30388 45484 30428
rect 45524 30388 46444 30428
rect 46484 30388 47020 30428
rect 47060 30388 47069 30428
rect 48268 30388 48556 30428
rect 48596 30388 48605 30428
rect 49603 30388 49612 30428
rect 49652 30388 51628 30428
rect 51668 30388 51677 30428
rect 3715 30304 3724 30344
rect 3764 30304 5932 30344
rect 5972 30304 7564 30344
rect 7604 30304 7613 30344
rect 11203 30304 11212 30344
rect 11252 30304 11692 30344
rect 11732 30304 11741 30344
rect 11788 30304 13516 30344
rect 13556 30304 13565 30344
rect 22627 30304 22636 30344
rect 22676 30304 27148 30344
rect 27188 30304 27197 30344
rect 28387 30304 28396 30344
rect 28436 30304 29164 30344
rect 29204 30304 29213 30344
rect 38275 30304 38284 30344
rect 38324 30304 38764 30344
rect 38804 30304 38813 30344
rect 11788 30260 11828 30304
rect 48268 30260 48308 30388
rect 48931 30304 48940 30344
rect 48980 30304 50188 30344
rect 50228 30304 50237 30344
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 7843 30220 7852 30260
rect 7892 30220 8812 30260
rect 8852 30220 8861 30260
rect 11107 30220 11116 30260
rect 11156 30220 11828 30260
rect 11875 30220 11884 30260
rect 11924 30220 13420 30260
rect 13460 30220 13469 30260
rect 13603 30220 13612 30260
rect 13652 30220 14764 30260
rect 14804 30220 14813 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 21187 30220 21196 30260
rect 21236 30220 21676 30260
rect 21716 30220 23884 30260
rect 23924 30220 25996 30260
rect 26036 30220 26045 30260
rect 28960 30220 29452 30260
rect 29492 30220 30124 30260
rect 30164 30220 31948 30260
rect 31988 30220 32236 30260
rect 32276 30220 32716 30260
rect 32756 30220 32765 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 35107 30220 35116 30260
rect 35156 30220 35596 30260
rect 35636 30220 35884 30260
rect 35924 30220 35933 30260
rect 37507 30220 37516 30260
rect 37556 30220 37708 30260
rect 37748 30220 39436 30260
rect 39476 30220 39485 30260
rect 40867 30220 40876 30260
rect 40916 30220 41260 30260
rect 41300 30220 41836 30260
rect 41876 30220 41885 30260
rect 47779 30220 47788 30260
rect 47828 30220 48076 30260
rect 48116 30220 48125 30260
rect 48259 30220 48268 30260
rect 48308 30220 48317 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 28960 30176 29000 30220
rect 11779 30136 11788 30176
rect 11828 30136 13324 30176
rect 13364 30136 13373 30176
rect 18691 30136 18700 30176
rect 18740 30136 22348 30176
rect 22388 30136 22397 30176
rect 25315 30136 25324 30176
rect 25364 30136 26284 30176
rect 26324 30136 29000 30176
rect 32716 30176 32756 30220
rect 32716 30136 34444 30176
rect 34484 30136 34493 30176
rect 9091 30052 9100 30092
rect 9140 30052 12172 30092
rect 12212 30052 23020 30092
rect 23060 30052 24364 30092
rect 24404 30052 24413 30092
rect 34051 30052 34060 30092
rect 34100 30052 35692 30092
rect 35732 30052 35741 30092
rect 36259 30052 36268 30092
rect 36308 30052 37132 30092
rect 37172 30052 37181 30092
rect 0 29948 80 30028
rect 1027 29968 1036 30008
rect 1076 29968 1612 30008
rect 1652 29968 1661 30008
rect 3340 29968 4108 30008
rect 4148 29968 4396 30008
rect 4436 29968 4445 30008
rect 5539 29968 5548 30008
rect 5588 29968 5597 30008
rect 5827 29968 5836 30008
rect 5876 29968 7564 30008
rect 7604 29968 8140 30008
rect 8180 29968 8716 30008
rect 8756 29968 8765 30008
rect 11299 29968 11308 30008
rect 11348 29968 12268 30008
rect 12308 29968 12556 30008
rect 12596 29968 12605 30008
rect 18595 29968 18604 30008
rect 18644 29968 19468 30008
rect 19508 29968 19517 30008
rect 38371 29968 38380 30008
rect 38420 29968 42028 30008
rect 42068 29968 42316 30008
rect 42356 29968 42365 30008
rect 46915 29968 46924 30008
rect 46964 29968 47788 30008
rect 47828 29968 47837 30008
rect 3340 29924 3380 29968
rect 5548 29924 5588 29968
rect 13123 29924 13181 29925
rect 3331 29884 3340 29924
rect 3380 29884 3389 29924
rect 3619 29884 3628 29924
rect 3668 29884 5068 29924
rect 5108 29884 5588 29924
rect 9955 29884 9964 29924
rect 10004 29884 13132 29924
rect 13172 29884 13900 29924
rect 13940 29884 13949 29924
rect 14659 29884 14668 29924
rect 14708 29884 15820 29924
rect 15860 29884 17356 29924
rect 17396 29884 17405 29924
rect 18787 29884 18796 29924
rect 18836 29884 18988 29924
rect 19028 29884 19037 29924
rect 35971 29884 35980 29924
rect 36020 29884 36556 29924
rect 36596 29884 37420 29924
rect 37460 29884 37469 29924
rect 13123 29883 13181 29884
rect 5635 29840 5693 29841
rect 18796 29840 18836 29884
rect 3811 29800 3820 29840
rect 3860 29800 4780 29840
rect 4820 29800 5164 29840
rect 5204 29800 5213 29840
rect 5550 29800 5644 29840
rect 5684 29800 5693 29840
rect 7651 29800 7660 29840
rect 7700 29800 11308 29840
rect 11348 29800 11357 29840
rect 11779 29800 11788 29840
rect 11828 29800 12076 29840
rect 12116 29800 12125 29840
rect 12835 29800 12844 29840
rect 12884 29800 13996 29840
rect 14036 29800 14045 29840
rect 14563 29800 14572 29840
rect 14612 29800 15052 29840
rect 15092 29800 18836 29840
rect 18883 29800 18892 29840
rect 18932 29800 20812 29840
rect 20852 29800 20861 29840
rect 28771 29800 28780 29840
rect 28820 29800 29260 29840
rect 29300 29800 29309 29840
rect 30979 29800 30988 29840
rect 31028 29800 31660 29840
rect 31700 29800 31948 29840
rect 31988 29800 31997 29840
rect 33091 29800 33100 29840
rect 33140 29800 33580 29840
rect 33620 29800 33629 29840
rect 36259 29800 36268 29840
rect 36308 29800 37324 29840
rect 37364 29800 37373 29840
rect 39043 29800 39052 29840
rect 39092 29800 42124 29840
rect 42164 29800 42988 29840
rect 43028 29800 43037 29840
rect 43459 29800 43468 29840
rect 43508 29800 45100 29840
rect 45140 29800 45772 29840
rect 45812 29800 45964 29840
rect 46004 29800 48364 29840
rect 48404 29800 49420 29840
rect 49460 29800 50380 29840
rect 50420 29800 50429 29840
rect 5635 29799 5693 29800
rect 26563 29716 26572 29756
rect 26612 29716 27916 29756
rect 27956 29716 27965 29756
rect 41059 29716 41068 29756
rect 41108 29716 41644 29756
rect 41684 29716 41693 29756
rect 41827 29716 41836 29756
rect 41876 29716 43276 29756
rect 43316 29716 46924 29756
rect 46964 29716 46973 29756
rect 47299 29716 47308 29756
rect 47348 29716 48172 29756
rect 48212 29716 48221 29756
rect 4579 29632 4588 29672
rect 4628 29632 4637 29672
rect 5251 29632 5260 29672
rect 5300 29632 6508 29672
rect 6548 29632 6557 29672
rect 7171 29632 7180 29672
rect 7220 29632 8428 29672
rect 8468 29632 8477 29672
rect 13219 29632 13228 29672
rect 13268 29632 15052 29672
rect 15092 29632 15101 29672
rect 35971 29632 35980 29672
rect 36020 29632 36460 29672
rect 36500 29632 36509 29672
rect 37699 29632 37708 29672
rect 37748 29632 41356 29672
rect 41396 29632 41405 29672
rect 42499 29632 42508 29672
rect 42548 29632 43372 29672
rect 43412 29632 43421 29672
rect 45859 29632 45868 29672
rect 45908 29632 47116 29672
rect 47156 29632 47165 29672
rect 4588 29588 4628 29632
rect 4588 29548 9100 29588
rect 9140 29548 9149 29588
rect 27619 29548 27628 29588
rect 27668 29548 30124 29588
rect 30164 29548 30173 29588
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 6307 29464 6316 29504
rect 6356 29464 15340 29504
rect 15380 29464 15389 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 4099 29380 4108 29420
rect 4148 29380 5644 29420
rect 5684 29380 5693 29420
rect 27235 29380 27244 29420
rect 27284 29380 28204 29420
rect 28244 29380 28253 29420
rect 29836 29380 32332 29420
rect 32372 29380 32381 29420
rect 5347 29296 5356 29336
rect 5396 29296 5548 29336
rect 5588 29296 5597 29336
rect 5731 29296 5740 29336
rect 5780 29296 6028 29336
rect 6068 29296 7948 29336
rect 7988 29296 8716 29336
rect 8756 29296 8765 29336
rect 20515 29296 20524 29336
rect 20564 29296 21964 29336
rect 22004 29296 22013 29336
rect 27427 29296 27436 29336
rect 27476 29296 28108 29336
rect 28148 29296 28684 29336
rect 28724 29296 28733 29336
rect 28963 29296 28972 29336
rect 29012 29296 29740 29336
rect 29780 29296 29789 29336
rect 29836 29252 29876 29380
rect 30307 29296 30316 29336
rect 30356 29296 30700 29336
rect 30740 29296 30749 29336
rect 31747 29296 31756 29336
rect 31796 29296 33196 29336
rect 33236 29296 33245 29336
rect 39811 29296 39820 29336
rect 39860 29296 42892 29336
rect 42932 29296 42941 29336
rect 48067 29296 48076 29336
rect 48116 29296 49228 29336
rect 49268 29296 49277 29336
rect 2755 29212 2764 29252
rect 2804 29212 3244 29252
rect 3284 29212 3293 29252
rect 3523 29212 3532 29252
rect 3572 29212 4204 29252
rect 4244 29212 4253 29252
rect 4300 29212 5164 29252
rect 5204 29212 5836 29252
rect 5876 29212 5885 29252
rect 14371 29212 14380 29252
rect 14420 29212 16108 29252
rect 16148 29212 18700 29252
rect 18740 29212 18749 29252
rect 21091 29212 21100 29252
rect 21140 29212 22924 29252
rect 22964 29212 22973 29252
rect 25507 29212 25516 29252
rect 25556 29212 27916 29252
rect 27956 29212 27965 29252
rect 28195 29212 28204 29252
rect 28244 29212 29876 29252
rect 29923 29212 29932 29252
rect 29972 29212 30740 29252
rect 32899 29212 32908 29252
rect 32948 29212 33964 29252
rect 34004 29212 35788 29252
rect 35828 29212 38188 29252
rect 38228 29212 38237 29252
rect 41251 29212 41260 29252
rect 41300 29212 41644 29252
rect 41684 29212 44044 29252
rect 44084 29212 44093 29252
rect 0 29108 80 29188
rect 4300 29168 4340 29212
rect 14083 29168 14141 29169
rect 20227 29168 20285 29169
rect 2563 29128 2572 29168
rect 2612 29128 3724 29168
rect 3764 29128 3773 29168
rect 3907 29128 3916 29168
rect 3956 29128 4340 29168
rect 4675 29128 4684 29168
rect 4724 29128 6220 29168
rect 6260 29128 6269 29168
rect 7267 29128 7276 29168
rect 7316 29128 8044 29168
rect 8084 29128 8093 29168
rect 8707 29128 8716 29168
rect 8756 29128 8765 29168
rect 10147 29128 10156 29168
rect 10196 29128 12172 29168
rect 12212 29128 12221 29168
rect 13987 29128 13996 29168
rect 14036 29128 14092 29168
rect 14132 29128 14141 29168
rect 14275 29128 14284 29168
rect 14324 29128 14668 29168
rect 14708 29128 14717 29168
rect 16291 29128 16300 29168
rect 16340 29128 18604 29168
rect 18644 29128 18653 29168
rect 20142 29128 20236 29168
rect 20276 29128 20285 29168
rect 25795 29128 25804 29168
rect 25844 29128 26284 29168
rect 26324 29128 26333 29168
rect 26563 29128 26572 29168
rect 26612 29128 27244 29168
rect 27284 29128 27293 29168
rect 27523 29128 27532 29168
rect 27572 29128 28396 29168
rect 28436 29128 28445 29168
rect 28675 29128 28684 29168
rect 28724 29128 29000 29168
rect 30403 29128 30412 29168
rect 30452 29128 30604 29168
rect 30644 29128 30653 29168
rect 3916 29084 3956 29128
rect 8716 29084 8756 29128
rect 14083 29127 14141 29128
rect 20227 29127 20285 29128
rect 26284 29084 26324 29128
rect 28960 29084 29000 29128
rect 30700 29084 30740 29212
rect 31075 29128 31084 29168
rect 31124 29128 31564 29168
rect 31604 29128 31613 29168
rect 31660 29128 31948 29168
rect 31988 29128 31997 29168
rect 33763 29128 33772 29168
rect 33812 29128 34252 29168
rect 34292 29128 34301 29168
rect 37219 29128 37228 29168
rect 37268 29128 43276 29168
rect 43316 29128 43325 29168
rect 49027 29128 49036 29168
rect 49076 29128 50572 29168
rect 50612 29128 50621 29168
rect 31660 29084 31700 29128
rect 2500 29044 2804 29084
rect 2947 29044 2956 29084
rect 2996 29044 3956 29084
rect 6115 29044 6124 29084
rect 6164 29044 7180 29084
rect 7220 29044 7229 29084
rect 7363 29044 7372 29084
rect 7412 29044 8620 29084
rect 8660 29044 8669 29084
rect 8716 29044 15436 29084
rect 15476 29044 15485 29084
rect 19651 29044 19660 29084
rect 19700 29044 21292 29084
rect 21332 29044 21341 29084
rect 26284 29044 27436 29084
rect 27476 29044 27485 29084
rect 27916 29044 28588 29084
rect 28628 29044 28637 29084
rect 28960 29044 29260 29084
rect 29300 29044 30644 29084
rect 2500 29000 2540 29044
rect 2764 29000 2804 29044
rect 27916 29000 27956 29044
rect 1315 28960 1324 29000
rect 1364 28960 2540 29000
rect 2724 28960 2764 29000
rect 2804 28960 2813 29000
rect 27876 28960 27916 29000
rect 27956 28960 27965 29000
rect 30604 28916 30644 29044
rect 30700 29044 31700 29084
rect 31747 29044 31756 29084
rect 31796 29044 33140 29084
rect 33667 29044 33676 29084
rect 33716 29044 35596 29084
rect 35636 29044 36076 29084
rect 36116 29044 37132 29084
rect 37172 29044 37181 29084
rect 37228 29044 38476 29084
rect 38516 29044 38956 29084
rect 38996 29044 39005 29084
rect 40099 29044 40108 29084
rect 40148 29044 40876 29084
rect 40916 29044 40925 29084
rect 41731 29044 41740 29084
rect 41780 29044 43468 29084
rect 43508 29044 43517 29084
rect 30700 29000 30740 29044
rect 33100 29000 33140 29044
rect 30691 28960 30700 29000
rect 30740 28960 30749 29000
rect 30796 28960 30988 29000
rect 31028 28960 31037 29000
rect 33091 28960 33100 29000
rect 33140 28960 33149 29000
rect 30796 28916 30836 28960
rect 37228 28916 37268 29044
rect 8323 28876 8332 28916
rect 8372 28876 9292 28916
rect 9332 28876 9341 28916
rect 18979 28876 18988 28916
rect 19028 28876 20140 28916
rect 20180 28876 20189 28916
rect 26467 28876 26476 28916
rect 26516 28876 26764 28916
rect 26804 28876 26813 28916
rect 30595 28876 30604 28916
rect 30644 28876 30836 28916
rect 37219 28876 37228 28916
rect 37268 28876 37277 28916
rect 47107 28876 47116 28916
rect 47156 28876 47788 28916
rect 47828 28876 48940 28916
rect 48980 28876 48989 28916
rect 20227 28792 20236 28832
rect 20276 28792 20428 28832
rect 20468 28792 20477 28832
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 19747 28708 19756 28748
rect 19796 28708 20716 28748
rect 20756 28708 20765 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 20140 28624 20332 28664
rect 20372 28624 20381 28664
rect 26563 28624 26572 28664
rect 26612 28624 26860 28664
rect 26900 28624 26909 28664
rect 38083 28624 38092 28664
rect 38132 28624 39052 28664
rect 39092 28624 39101 28664
rect 20140 28580 20180 28624
rect 13891 28540 13900 28580
rect 13940 28540 14092 28580
rect 14132 28540 14141 28580
rect 20044 28540 20180 28580
rect 31075 28540 31084 28580
rect 31124 28540 32428 28580
rect 32468 28540 32620 28580
rect 32660 28540 32669 28580
rect 38851 28540 38860 28580
rect 38900 28540 39340 28580
rect 39380 28540 39389 28580
rect 20044 28496 20084 28540
rect 3811 28456 3820 28496
rect 3860 28456 4204 28496
rect 4244 28456 4876 28496
rect 4916 28456 4925 28496
rect 13411 28456 13420 28496
rect 13460 28456 13804 28496
rect 13844 28456 13853 28496
rect 19267 28456 19276 28496
rect 19316 28456 20084 28496
rect 28960 28456 29644 28496
rect 29684 28456 29693 28496
rect 30787 28456 30796 28496
rect 30836 28456 31372 28496
rect 31412 28456 31421 28496
rect 39427 28456 39436 28496
rect 39476 28456 39485 28496
rect 43171 28456 43180 28496
rect 43220 28456 47500 28496
rect 47540 28456 47549 28496
rect 28960 28412 29000 28456
rect 4300 28372 7468 28412
rect 7508 28372 7517 28412
rect 12739 28372 12748 28412
rect 12788 28372 13324 28412
rect 13364 28372 17932 28412
rect 17972 28372 28876 28412
rect 28916 28372 29000 28412
rect 39436 28412 39476 28456
rect 39436 28372 42220 28412
rect 42260 28372 43564 28412
rect 43604 28372 43613 28412
rect 45091 28372 45100 28412
rect 45140 28372 48268 28412
rect 48308 28372 48317 28412
rect 0 28268 80 28348
rect 4300 28328 4340 28372
rect 5635 28328 5693 28329
rect 20227 28328 20285 28329
rect 4291 28288 4300 28328
rect 4340 28288 4349 28328
rect 5155 28288 5164 28328
rect 5204 28288 5644 28328
rect 5684 28288 5693 28328
rect 7267 28288 7276 28328
rect 7316 28288 8716 28328
rect 8756 28288 8765 28328
rect 10147 28288 10156 28328
rect 10196 28288 13132 28328
rect 13172 28288 13181 28328
rect 13795 28288 13804 28328
rect 13844 28288 13853 28328
rect 14083 28288 14092 28328
rect 14132 28288 14476 28328
rect 14516 28288 14525 28328
rect 18403 28288 18412 28328
rect 18452 28288 19756 28328
rect 19796 28288 19805 28328
rect 20142 28288 20236 28328
rect 20276 28288 20524 28328
rect 20564 28288 20573 28328
rect 25315 28288 25324 28328
rect 25364 28288 27724 28328
rect 27764 28288 27773 28328
rect 28579 28288 28588 28328
rect 28628 28288 30412 28328
rect 30452 28288 30461 28328
rect 30883 28288 30892 28328
rect 30932 28288 31468 28328
rect 31508 28288 31517 28328
rect 37219 28288 37228 28328
rect 37268 28288 38380 28328
rect 38420 28288 38860 28328
rect 38900 28288 38909 28328
rect 40483 28288 40492 28328
rect 40532 28288 43372 28328
rect 43412 28288 43421 28328
rect 43651 28288 43660 28328
rect 43700 28288 43709 28328
rect 46531 28288 46540 28328
rect 46580 28288 47020 28328
rect 47060 28288 47069 28328
rect 47875 28288 47884 28328
rect 47924 28288 48748 28328
rect 48788 28288 48797 28328
rect 5635 28287 5693 28288
rect 13804 28244 13844 28288
rect 20227 28287 20285 28288
rect 43660 28244 43700 28288
rect 1315 28204 1324 28244
rect 1364 28204 4108 28244
rect 4148 28204 4157 28244
rect 7171 28204 7180 28244
rect 7220 28204 8236 28244
rect 8276 28204 8285 28244
rect 13804 28204 16588 28244
rect 16628 28204 17548 28244
rect 17588 28204 18796 28244
rect 18836 28204 18845 28244
rect 20323 28204 20332 28244
rect 20372 28204 21004 28244
rect 21044 28204 21053 28244
rect 26659 28204 26668 28244
rect 26708 28204 26956 28244
rect 26996 28204 27005 28244
rect 28492 28204 28972 28244
rect 29012 28204 29021 28244
rect 32740 28204 35212 28244
rect 35252 28204 35261 28244
rect 43660 28204 46636 28244
rect 46676 28204 46685 28244
rect 46819 28204 46828 28244
rect 46868 28204 49996 28244
rect 50036 28204 50045 28244
rect 20611 28160 20669 28161
rect 28492 28160 28532 28204
rect 32740 28160 32780 28204
rect 6019 28120 6028 28160
rect 6068 28120 7372 28160
rect 7412 28120 7421 28160
rect 8707 28120 8716 28160
rect 8756 28120 10348 28160
rect 10388 28120 14572 28160
rect 14612 28120 14621 28160
rect 18691 28120 18700 28160
rect 18740 28120 19276 28160
rect 19316 28120 20236 28160
rect 20276 28120 20285 28160
rect 20592 28120 20620 28160
rect 20660 28120 20716 28160
rect 20756 28120 22732 28160
rect 22772 28120 22781 28160
rect 28483 28120 28492 28160
rect 28532 28120 28541 28160
rect 28675 28120 28684 28160
rect 28724 28120 32780 28160
rect 43075 28120 43084 28160
rect 43124 28120 43468 28160
rect 43508 28120 43517 28160
rect 44515 28120 44524 28160
rect 44564 28120 46252 28160
rect 46292 28120 46732 28160
rect 46772 28120 46781 28160
rect 47299 28120 47308 28160
rect 47348 28120 48652 28160
rect 48692 28120 48701 28160
rect 49795 28120 49804 28160
rect 49844 28120 51628 28160
rect 51668 28120 51677 28160
rect 14572 28076 14612 28120
rect 20611 28119 20669 28120
rect 4771 28036 4780 28076
rect 4820 28036 5356 28076
rect 5396 28036 6700 28076
rect 6740 28036 7276 28076
rect 7316 28036 7325 28076
rect 14572 28036 19180 28076
rect 19220 28036 19229 28076
rect 26083 28036 26092 28076
rect 26132 28036 26284 28076
rect 26324 28036 40012 28076
rect 40052 28036 40061 28076
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 6787 27952 6796 27992
rect 6836 27952 7852 27992
rect 7892 27952 7901 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 27715 27952 27724 27992
rect 27764 27952 28684 27992
rect 28724 27952 28733 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 42883 27952 42892 27992
rect 42932 27952 43372 27992
rect 43412 27952 43421 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 31171 27908 31229 27909
rect 31086 27868 31180 27908
rect 31220 27868 31229 27908
rect 46147 27868 46156 27908
rect 46196 27868 47020 27908
rect 47060 27868 47069 27908
rect 31171 27867 31229 27868
rect 4195 27784 4204 27824
rect 4244 27784 4253 27824
rect 4675 27784 4684 27824
rect 4724 27784 4876 27824
rect 4916 27784 6604 27824
rect 6644 27784 6653 27824
rect 7747 27784 7756 27824
rect 7796 27784 7805 27824
rect 31267 27784 31276 27824
rect 31316 27784 32140 27824
rect 32180 27784 32189 27824
rect 35683 27784 35692 27824
rect 35732 27784 38764 27824
rect 38804 27784 38956 27824
rect 38996 27784 39005 27824
rect 42883 27784 42892 27824
rect 42932 27784 45004 27824
rect 45044 27784 45053 27824
rect 45475 27784 45484 27824
rect 45524 27784 46444 27824
rect 46484 27784 46493 27824
rect 46627 27784 46636 27824
rect 46676 27784 48652 27824
rect 48692 27784 48701 27824
rect 49987 27784 49996 27824
rect 50036 27784 50860 27824
rect 50900 27784 50909 27824
rect 4204 27740 4244 27784
rect 7756 27740 7796 27784
rect 3043 27700 3052 27740
rect 3092 27700 4244 27740
rect 7075 27700 7084 27740
rect 7124 27700 7564 27740
rect 7604 27700 7613 27740
rect 7756 27700 8428 27740
rect 8468 27700 8477 27740
rect 19843 27700 19852 27740
rect 19892 27700 23404 27740
rect 23444 27700 24268 27740
rect 24308 27700 24317 27740
rect 24451 27700 24460 27740
rect 24500 27700 29740 27740
rect 29780 27700 29789 27740
rect 29836 27700 30700 27740
rect 30740 27700 30988 27740
rect 31028 27700 31037 27740
rect 36355 27700 36364 27740
rect 36404 27700 38380 27740
rect 38420 27700 38429 27740
rect 40963 27700 40972 27740
rect 41012 27700 43796 27740
rect 43843 27700 43852 27740
rect 43892 27700 44428 27740
rect 44468 27700 44477 27740
rect 45196 27700 47212 27740
rect 47252 27700 47261 27740
rect 3331 27616 3340 27656
rect 3380 27616 3724 27656
rect 3764 27616 3773 27656
rect 0 27428 80 27508
rect 4012 27488 4052 27700
rect 28483 27656 28541 27657
rect 29836 27656 29876 27700
rect 43756 27656 43796 27700
rect 45196 27656 45236 27700
rect 5923 27616 5932 27656
rect 5972 27616 8140 27656
rect 8180 27616 8189 27656
rect 12835 27616 12844 27656
rect 12884 27616 13708 27656
rect 13748 27616 13757 27656
rect 14142 27616 14151 27656
rect 14191 27616 14956 27656
rect 14996 27616 15005 27656
rect 16003 27616 16012 27656
rect 16052 27616 16061 27656
rect 16291 27616 16300 27656
rect 16340 27616 19564 27656
rect 19604 27616 19613 27656
rect 26083 27616 26092 27656
rect 26132 27616 26764 27656
rect 26804 27616 26813 27656
rect 28398 27616 28492 27656
rect 28532 27616 28541 27656
rect 29059 27616 29068 27656
rect 29108 27616 29117 27656
rect 29251 27616 29260 27656
rect 29300 27616 29548 27656
rect 29588 27616 29876 27656
rect 30403 27616 30412 27656
rect 30452 27616 31756 27656
rect 31796 27616 31805 27656
rect 32803 27616 32812 27656
rect 32852 27616 33292 27656
rect 33332 27616 33341 27656
rect 33955 27616 33964 27656
rect 34004 27616 34348 27656
rect 34388 27616 34397 27656
rect 35011 27616 35020 27656
rect 35060 27616 35212 27656
rect 35252 27616 39916 27656
rect 39956 27616 39965 27656
rect 43756 27616 43948 27656
rect 43988 27616 43997 27656
rect 45187 27616 45196 27656
rect 45236 27616 45245 27656
rect 45379 27616 45388 27656
rect 45428 27616 45964 27656
rect 46004 27616 46013 27656
rect 48163 27616 48172 27656
rect 48212 27616 48940 27656
rect 48980 27616 48989 27656
rect 16012 27572 16052 27616
rect 28483 27615 28541 27616
rect 20611 27572 20669 27573
rect 28579 27572 28637 27573
rect 7651 27532 7660 27572
rect 7700 27532 8044 27572
rect 8084 27532 8908 27572
rect 8948 27532 8957 27572
rect 13603 27532 13612 27572
rect 13652 27532 14764 27572
rect 14804 27532 14813 27572
rect 16012 27532 16492 27572
rect 16532 27532 16541 27572
rect 20526 27532 20620 27572
rect 20660 27532 20669 27572
rect 28494 27532 28588 27572
rect 28628 27532 28637 27572
rect 29068 27572 29108 27616
rect 29068 27532 35308 27572
rect 35348 27532 35357 27572
rect 43171 27532 43180 27572
rect 43220 27532 43660 27572
rect 43700 27532 43709 27572
rect 45571 27532 45580 27572
rect 45620 27532 45629 27572
rect 47587 27532 47596 27572
rect 47636 27532 49228 27572
rect 49268 27532 50668 27572
rect 50708 27532 50717 27572
rect 20611 27531 20669 27532
rect 28579 27531 28637 27532
rect 45580 27488 45620 27532
rect 4003 27448 4012 27488
rect 4052 27448 4061 27488
rect 7747 27448 7756 27488
rect 7796 27448 8716 27488
rect 8756 27448 11444 27488
rect 11971 27448 11980 27488
rect 12020 27448 13900 27488
rect 13940 27448 13949 27488
rect 13996 27448 17452 27488
rect 17492 27448 17501 27488
rect 20995 27448 21004 27488
rect 21044 27448 21868 27488
rect 21908 27448 21917 27488
rect 28003 27448 28012 27488
rect 28052 27448 28684 27488
rect 28724 27448 31276 27488
rect 31316 27448 31468 27488
rect 31508 27448 31517 27488
rect 33091 27448 33100 27488
rect 33140 27448 34828 27488
rect 34868 27448 34877 27488
rect 45388 27448 45620 27488
rect 46600 27448 47116 27488
rect 47156 27448 47500 27488
rect 47540 27448 47549 27488
rect 47683 27448 47692 27488
rect 47732 27448 48268 27488
rect 48308 27448 48317 27488
rect 48451 27448 48460 27488
rect 48500 27448 48748 27488
rect 48788 27448 49132 27488
rect 49172 27448 49181 27488
rect 11404 27404 11444 27448
rect 13996 27404 14036 27448
rect 45388 27404 45428 27448
rect 2947 27364 2956 27404
rect 2996 27364 5068 27404
rect 5108 27364 5117 27404
rect 11395 27364 11404 27404
rect 11444 27364 11596 27404
rect 11636 27364 11645 27404
rect 12643 27364 12652 27404
rect 12692 27364 14036 27404
rect 14755 27364 14764 27404
rect 14804 27364 14813 27404
rect 15296 27364 15305 27404
rect 15345 27364 16012 27404
rect 16052 27364 16061 27404
rect 18979 27364 18988 27404
rect 19028 27364 19372 27404
rect 19412 27364 21196 27404
rect 21236 27364 21245 27404
rect 25123 27364 25132 27404
rect 25172 27364 27148 27404
rect 27188 27364 27197 27404
rect 27715 27364 27724 27404
rect 27764 27364 28492 27404
rect 28532 27364 29164 27404
rect 29204 27364 29213 27404
rect 35587 27364 35596 27404
rect 35636 27364 39148 27404
rect 39188 27364 39628 27404
rect 39668 27364 39677 27404
rect 41731 27364 41740 27404
rect 41780 27364 43468 27404
rect 43508 27364 43517 27404
rect 45379 27364 45388 27404
rect 45428 27364 45437 27404
rect 45571 27364 45580 27404
rect 45620 27364 45964 27404
rect 46004 27364 46013 27404
rect 14764 27320 14804 27364
rect 46600 27320 46640 27448
rect 47011 27364 47020 27404
rect 47060 27364 49036 27404
rect 49076 27364 49085 27404
rect 2755 27280 2764 27320
rect 2804 27280 8620 27320
rect 8660 27280 8669 27320
rect 14764 27280 24844 27320
rect 24884 27280 24893 27320
rect 30787 27280 30796 27320
rect 30836 27280 44044 27320
rect 44084 27280 44093 27320
rect 45091 27280 45100 27320
rect 45140 27280 46640 27320
rect 47203 27280 47212 27320
rect 47252 27280 48172 27320
rect 48212 27280 48221 27320
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 3619 27196 3628 27236
rect 3668 27196 4108 27236
rect 4148 27196 4157 27236
rect 6979 27196 6988 27236
rect 7028 27196 8428 27236
rect 8468 27196 11692 27236
rect 11732 27196 11741 27236
rect 12451 27196 12460 27236
rect 12500 27196 13228 27236
rect 13268 27196 14188 27236
rect 14228 27196 15244 27236
rect 15284 27196 16204 27236
rect 16244 27196 16780 27236
rect 16820 27196 17068 27236
rect 17108 27196 17356 27236
rect 17396 27196 17405 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 20227 27196 20236 27236
rect 20276 27196 23212 27236
rect 23252 27196 23261 27236
rect 24268 27196 24748 27236
rect 24788 27196 24797 27236
rect 31363 27196 31372 27236
rect 31412 27196 32524 27236
rect 32564 27196 32573 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 33859 27196 33868 27236
rect 33908 27196 37708 27236
rect 37748 27196 38188 27236
rect 38228 27196 38237 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 24268 27152 24308 27196
rect 14275 27112 14284 27152
rect 14324 27112 14668 27152
rect 14708 27112 24268 27152
rect 24308 27112 24317 27152
rect 24643 27112 24652 27152
rect 24692 27112 39820 27152
rect 39860 27112 39869 27152
rect 3619 27028 3628 27068
rect 3668 27028 5164 27068
rect 5204 27028 5213 27068
rect 11971 27028 11980 27068
rect 12020 27028 12268 27068
rect 12308 27028 12317 27068
rect 14371 27028 14380 27068
rect 14420 27028 14860 27068
rect 14900 27028 14909 27068
rect 17731 27028 17740 27068
rect 17780 27028 24748 27068
rect 24788 27028 24797 27068
rect 28771 27028 28780 27068
rect 28820 27028 30316 27068
rect 30356 27028 30365 27068
rect 30691 27028 30700 27068
rect 30740 27028 30988 27068
rect 31028 27028 31037 27068
rect 31747 27028 31756 27068
rect 31796 27028 36844 27068
rect 36884 27028 36893 27068
rect 44515 27028 44524 27068
rect 44564 27028 47980 27068
rect 48020 27028 48844 27068
rect 48884 27028 48893 27068
rect 8899 26944 8908 26984
rect 8948 26944 9292 26984
rect 9332 26944 9341 26984
rect 10531 26944 10540 26984
rect 10580 26944 18028 26984
rect 18068 26944 18077 26984
rect 24259 26944 24268 26984
rect 24308 26944 24940 26984
rect 24980 26944 24989 26984
rect 29635 26944 29644 26984
rect 29684 26944 38668 26984
rect 38708 26944 38717 26984
rect 11320 26860 12460 26900
rect 12500 26860 12509 26900
rect 13891 26860 13900 26900
rect 13940 26860 30316 26900
rect 30356 26860 30365 26900
rect 30979 26860 30988 26900
rect 31028 26860 31372 26900
rect 31412 26860 31421 26900
rect 32131 26860 32140 26900
rect 32180 26860 32428 26900
rect 32468 26860 32477 26900
rect 36076 26860 36268 26900
rect 36308 26860 36317 26900
rect 44131 26860 44140 26900
rect 44180 26860 45004 26900
rect 45044 26860 45053 26900
rect 48931 26860 48940 26900
rect 48980 26860 49612 26900
rect 49652 26860 49661 26900
rect 11320 26816 11360 26860
rect 1219 26776 1228 26816
rect 1268 26776 3820 26816
rect 3860 26776 3869 26816
rect 10819 26776 10828 26816
rect 10868 26776 10877 26816
rect 11011 26776 11020 26816
rect 11060 26776 11360 26816
rect 12163 26776 12172 26816
rect 12212 26776 12221 26816
rect 13027 26776 13036 26816
rect 13076 26776 14380 26816
rect 14420 26776 14860 26816
rect 14900 26776 14909 26816
rect 15331 26776 15340 26816
rect 15380 26776 19276 26816
rect 19316 26776 19325 26816
rect 19651 26776 19660 26816
rect 19700 26776 21964 26816
rect 22004 26776 22013 26816
rect 28963 26776 28972 26816
rect 29012 26776 29548 26816
rect 29588 26776 29597 26816
rect 30691 26776 30700 26816
rect 30740 26776 30892 26816
rect 30932 26776 30941 26816
rect 31075 26776 31084 26816
rect 31124 26776 31948 26816
rect 31988 26776 31997 26816
rect 32227 26776 32236 26816
rect 32276 26776 32812 26816
rect 32852 26776 32861 26816
rect 34435 26776 34444 26816
rect 34484 26776 35692 26816
rect 35732 26776 35980 26816
rect 36020 26776 36029 26816
rect 10828 26732 10868 26776
rect 12172 26732 12212 26776
rect 19660 26732 19700 26776
rect 36076 26732 36116 26860
rect 36163 26776 36172 26816
rect 36212 26776 36652 26816
rect 36692 26776 36701 26816
rect 40099 26776 40108 26816
rect 40148 26776 40300 26816
rect 40340 26776 41932 26816
rect 41972 26776 42412 26816
rect 42452 26776 42461 26816
rect 43075 26776 43084 26816
rect 43124 26776 46828 26816
rect 46868 26776 50188 26816
rect 50228 26776 50380 26816
rect 50420 26776 50860 26816
rect 50900 26776 50909 26816
rect 5635 26692 5644 26732
rect 5684 26692 10060 26732
rect 10100 26692 12212 26732
rect 12835 26692 12844 26732
rect 12884 26692 15052 26732
rect 15092 26692 16492 26732
rect 16532 26692 16541 26732
rect 18883 26692 18892 26732
rect 18932 26692 19084 26732
rect 19124 26692 19700 26732
rect 23875 26692 23884 26732
rect 23924 26692 24364 26732
rect 24404 26692 24413 26732
rect 32515 26692 32524 26732
rect 32564 26692 36116 26732
rect 47779 26692 47788 26732
rect 47828 26692 49324 26732
rect 49364 26692 49373 26732
rect 0 26588 80 26668
rect 13891 26608 13900 26648
rect 13940 26608 14284 26648
rect 14324 26608 14333 26648
rect 14659 26608 14668 26648
rect 14708 26608 14860 26648
rect 14900 26608 14909 26648
rect 24739 26608 24748 26648
rect 24788 26608 30700 26648
rect 30740 26608 30749 26648
rect 35395 26608 35404 26648
rect 35444 26608 35884 26648
rect 35924 26608 35933 26648
rect 36067 26608 36076 26648
rect 36116 26608 36364 26648
rect 36404 26608 36413 26648
rect 42883 26608 42892 26648
rect 42932 26608 43756 26648
rect 43796 26608 44332 26648
rect 44372 26608 44381 26648
rect 51619 26608 51628 26648
rect 51668 26608 52012 26648
rect 52052 26608 52061 26648
rect 12547 26524 12556 26564
rect 12596 26524 14572 26564
rect 14612 26524 14621 26564
rect 26659 26524 26668 26564
rect 26708 26524 27340 26564
rect 27380 26524 29068 26564
rect 29108 26524 29117 26564
rect 13027 26480 13085 26481
rect 14083 26480 14141 26481
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 7939 26440 7948 26480
rect 7988 26440 9100 26480
rect 9140 26440 9149 26480
rect 12643 26440 12652 26480
rect 12692 26440 13036 26480
rect 13076 26440 13085 26480
rect 13998 26440 14092 26480
rect 14132 26440 14141 26480
rect 14659 26440 14668 26480
rect 14708 26440 16876 26480
rect 16916 26440 16925 26480
rect 17155 26440 17164 26480
rect 17204 26440 18700 26480
rect 18740 26440 19276 26480
rect 19316 26440 19325 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 21667 26440 21676 26480
rect 21716 26440 22060 26480
rect 22100 26440 23116 26480
rect 23156 26440 23165 26480
rect 24931 26440 24940 26480
rect 24980 26440 25900 26480
rect 25940 26440 25949 26480
rect 28387 26440 28396 26480
rect 28436 26440 29452 26480
rect 29492 26440 31564 26480
rect 31604 26440 31756 26480
rect 31796 26440 31805 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 38275 26440 38284 26480
rect 38324 26440 40684 26480
rect 40724 26440 40733 26480
rect 40867 26440 40876 26480
rect 40916 26440 41548 26480
rect 41588 26440 41597 26480
rect 43267 26440 43276 26480
rect 43316 26440 43892 26480
rect 47299 26440 47308 26480
rect 47348 26440 48172 26480
rect 48212 26440 48221 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 13027 26439 13085 26440
rect 14083 26439 14141 26440
rect 31171 26396 31229 26397
rect 8515 26356 8524 26396
rect 8564 26356 16012 26396
rect 16052 26356 16061 26396
rect 16108 26356 17548 26396
rect 17588 26356 22732 26396
rect 22772 26356 22781 26396
rect 24547 26356 24556 26396
rect 24596 26356 25420 26396
rect 25460 26356 25469 26396
rect 31086 26356 31180 26396
rect 31220 26356 31229 26396
rect 16108 26312 16148 26356
rect 31171 26355 31229 26356
rect 19171 26312 19229 26313
rect 43852 26312 43892 26440
rect 47587 26396 47645 26397
rect 45091 26356 45100 26396
rect 45140 26356 45292 26396
rect 45332 26356 47596 26396
rect 47636 26356 47692 26396
rect 47732 26356 47741 26396
rect 47587 26355 47645 26356
rect 3619 26272 3628 26312
rect 3668 26272 4532 26312
rect 4579 26272 4588 26312
rect 4628 26272 5740 26312
rect 5780 26272 5789 26312
rect 9187 26272 9196 26312
rect 9236 26272 9868 26312
rect 9908 26272 9917 26312
rect 14851 26272 14860 26312
rect 14900 26272 14940 26312
rect 15043 26272 15052 26312
rect 15092 26272 15628 26312
rect 15668 26272 15916 26312
rect 15956 26272 16148 26312
rect 17251 26272 17260 26312
rect 17300 26272 18260 26312
rect 4492 26228 4532 26272
rect 14860 26228 14900 26272
rect 18220 26228 18260 26272
rect 19171 26272 19180 26312
rect 19220 26272 19372 26312
rect 19412 26272 19421 26312
rect 29731 26272 29740 26312
rect 29780 26272 32332 26312
rect 32372 26272 32381 26312
rect 38467 26272 38476 26312
rect 38516 26272 40780 26312
rect 40820 26272 40829 26312
rect 43363 26272 43372 26312
rect 43412 26272 43660 26312
rect 43700 26272 43709 26312
rect 43843 26272 43852 26312
rect 43892 26272 44372 26312
rect 44515 26272 44524 26312
rect 44564 26272 49228 26312
rect 49268 26272 49804 26312
rect 49844 26272 49853 26312
rect 19171 26271 19229 26272
rect 39139 26228 39197 26229
rect 44332 26228 44372 26272
rect 1219 26188 1228 26228
rect 1268 26188 4396 26228
rect 4436 26188 4445 26228
rect 4492 26188 4780 26228
rect 4820 26188 7852 26228
rect 7892 26188 7901 26228
rect 10915 26188 10924 26228
rect 10964 26188 12116 26228
rect 12076 26144 12116 26188
rect 12652 26188 14188 26228
rect 14228 26188 15244 26228
rect 15284 26188 15293 26228
rect 18211 26188 18220 26228
rect 18260 26188 18269 26228
rect 19267 26188 19276 26228
rect 19316 26188 20908 26228
rect 20948 26188 20957 26228
rect 21091 26188 21100 26228
rect 21140 26188 23308 26228
rect 23348 26188 23357 26228
rect 26371 26188 26380 26228
rect 26420 26188 27628 26228
rect 27668 26188 27677 26228
rect 39054 26188 39148 26228
rect 39188 26188 39197 26228
rect 12652 26144 12692 26188
rect 39139 26187 39197 26188
rect 39820 26188 44236 26228
rect 44276 26188 44285 26228
rect 44332 26188 45676 26228
rect 45716 26188 48116 26228
rect 25987 26144 26045 26145
rect 29827 26144 29885 26145
rect 39820 26144 39860 26188
rect 47587 26144 47645 26145
rect 48076 26144 48116 26188
rect 4483 26104 4492 26144
rect 4532 26104 5068 26144
rect 5108 26104 5452 26144
rect 5492 26104 5501 26144
rect 10156 26104 10252 26144
rect 10292 26104 11308 26144
rect 11348 26104 11357 26144
rect 12067 26104 12076 26144
rect 12116 26104 12652 26144
rect 12692 26104 12701 26144
rect 13603 26104 13612 26144
rect 13652 26104 13661 26144
rect 16099 26104 16108 26144
rect 16148 26104 17740 26144
rect 17780 26104 17789 26144
rect 19459 26104 19468 26144
rect 19508 26104 20332 26144
rect 20372 26104 20381 26144
rect 22339 26104 22348 26144
rect 22388 26104 22924 26144
rect 22964 26104 22973 26144
rect 25123 26104 25132 26144
rect 25172 26104 25181 26144
rect 25902 26104 25996 26144
rect 26036 26104 26045 26144
rect 27715 26104 27724 26144
rect 27764 26104 28300 26144
rect 28340 26104 28349 26144
rect 29742 26104 29836 26144
rect 29876 26104 29885 26144
rect 31363 26104 31372 26144
rect 31412 26104 39340 26144
rect 39380 26104 39389 26144
rect 39811 26104 39820 26144
rect 39860 26104 39869 26144
rect 40291 26104 40300 26144
rect 40340 26104 42220 26144
rect 42260 26104 42269 26144
rect 42787 26104 42796 26144
rect 42836 26104 43084 26144
rect 43124 26104 43133 26144
rect 44131 26104 44140 26144
rect 44180 26104 44428 26144
rect 44468 26104 44716 26144
rect 44756 26104 44765 26144
rect 44899 26104 44908 26144
rect 44948 26104 47212 26144
rect 47252 26104 47261 26144
rect 47502 26104 47596 26144
rect 47636 26104 47645 26144
rect 48067 26104 48076 26144
rect 48116 26104 48125 26144
rect 48355 26104 48364 26144
rect 48404 26104 49900 26144
rect 49940 26104 50956 26144
rect 50996 26104 51005 26144
rect 10156 26060 10196 26104
rect 13612 26060 13652 26104
rect 25132 26060 25172 26104
rect 25987 26103 26045 26104
rect 29827 26103 29885 26104
rect 39340 26060 39380 26104
rect 47587 26103 47645 26104
rect 9667 26020 9676 26060
rect 9716 26020 10156 26060
rect 10196 26020 10205 26060
rect 11011 26020 11020 26060
rect 11060 26020 13652 26060
rect 17251 26020 17260 26060
rect 17300 26020 17452 26060
rect 17492 26020 17501 26060
rect 18787 26020 18796 26060
rect 18836 26020 19372 26060
rect 19412 26020 19421 26060
rect 22819 26020 22828 26060
rect 22868 26020 24268 26060
rect 24308 26020 24317 26060
rect 25132 26020 28396 26060
rect 28436 26020 28445 26060
rect 39340 26020 40588 26060
rect 40628 26020 40637 26060
rect 47500 26020 50764 26060
rect 50804 26020 51148 26060
rect 51188 26020 51197 26060
rect 47500 25976 47540 26020
rect 1027 25936 1036 25976
rect 1076 25936 1612 25976
rect 1652 25936 1661 25976
rect 10435 25936 10444 25976
rect 10484 25936 10924 25976
rect 10964 25936 10973 25976
rect 11320 25936 12556 25976
rect 12596 25936 12605 25976
rect 12835 25936 12844 25976
rect 12884 25936 14380 25976
rect 14420 25936 14429 25976
rect 15043 25936 15052 25976
rect 15092 25936 16588 25976
rect 16628 25936 16637 25976
rect 18403 25936 18412 25976
rect 18452 25936 25804 25976
rect 25844 25936 25853 25976
rect 30979 25936 30988 25976
rect 31028 25936 34100 25976
rect 34147 25936 34156 25976
rect 34196 25936 35212 25976
rect 35252 25936 35261 25976
rect 36451 25936 36460 25976
rect 36500 25936 36844 25976
rect 36884 25936 36893 25976
rect 42499 25936 42508 25976
rect 42548 25936 47500 25976
rect 47540 25936 47549 25976
rect 48739 25936 48748 25976
rect 48788 25936 49132 25976
rect 49172 25936 49181 25976
rect 11320 25892 11360 25936
rect 30595 25892 30653 25893
rect 34060 25892 34100 25936
rect 8227 25852 8236 25892
rect 8276 25852 11360 25892
rect 13027 25852 13036 25892
rect 13076 25852 13612 25892
rect 13652 25852 13661 25892
rect 13891 25852 13900 25892
rect 13940 25852 20180 25892
rect 20323 25852 20332 25892
rect 20372 25852 21772 25892
rect 21812 25852 21821 25892
rect 24835 25852 24844 25892
rect 24884 25852 26284 25892
rect 26324 25852 26333 25892
rect 26947 25852 26956 25892
rect 26996 25852 27244 25892
rect 27284 25852 27293 25892
rect 30510 25852 30604 25892
rect 30644 25852 30653 25892
rect 32707 25852 32716 25892
rect 32756 25852 33580 25892
rect 33620 25852 33629 25892
rect 34060 25852 40780 25892
rect 40820 25852 40829 25892
rect 46339 25852 46348 25892
rect 46388 25852 46732 25892
rect 46772 25852 46781 25892
rect 49027 25852 49036 25892
rect 49076 25852 50092 25892
rect 50132 25852 50141 25892
rect 0 25748 80 25828
rect 20140 25808 20180 25852
rect 30595 25851 30653 25852
rect 20140 25768 27532 25808
rect 27572 25768 27581 25808
rect 32323 25768 32332 25808
rect 32372 25768 36556 25808
rect 36596 25768 39628 25808
rect 39668 25768 39677 25808
rect 13027 25724 13085 25725
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 4003 25684 4012 25724
rect 4052 25684 6796 25724
rect 6836 25684 6845 25724
rect 12942 25684 13036 25724
rect 13076 25684 13085 25724
rect 16675 25684 16684 25724
rect 16724 25684 17452 25724
rect 17492 25684 17501 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 19075 25684 19084 25724
rect 19124 25684 19372 25724
rect 19412 25684 19421 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 33859 25684 33868 25724
rect 33908 25684 34348 25724
rect 34388 25684 34397 25724
rect 34732 25684 38860 25724
rect 38900 25684 38909 25724
rect 45667 25684 45676 25724
rect 45716 25684 46156 25724
rect 46196 25684 46205 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 13027 25683 13085 25684
rect 14275 25600 14284 25640
rect 14324 25600 30892 25640
rect 30932 25600 30941 25640
rect 31660 25600 34540 25640
rect 34580 25600 34589 25640
rect 25507 25556 25565 25557
rect 31660 25556 31700 25600
rect 34732 25556 34772 25684
rect 43459 25600 43468 25640
rect 43508 25600 43852 25640
rect 43892 25600 44524 25640
rect 44564 25600 44573 25640
rect 41251 25556 41309 25557
rect 12259 25516 12268 25556
rect 12308 25516 13132 25556
rect 13172 25516 13181 25556
rect 15427 25516 15436 25556
rect 15476 25516 23692 25556
rect 23732 25516 23741 25556
rect 25422 25516 25516 25556
rect 25556 25516 25565 25556
rect 25507 25515 25565 25516
rect 28960 25516 29548 25556
rect 29588 25516 29597 25556
rect 30787 25516 30796 25556
rect 30836 25516 31276 25556
rect 31316 25516 31660 25556
rect 31700 25516 31709 25556
rect 31756 25516 34772 25556
rect 41166 25516 41260 25556
rect 41300 25516 41309 25556
rect 28960 25472 29000 25516
rect 31756 25472 31796 25516
rect 41251 25515 41309 25516
rect 41356 25516 45388 25556
rect 45428 25516 45437 25556
rect 41356 25472 41396 25516
rect 13315 25432 13324 25472
rect 13364 25432 13804 25472
rect 13844 25432 13853 25472
rect 14275 25432 14284 25472
rect 14324 25432 14764 25472
rect 14804 25432 14813 25472
rect 23587 25432 23596 25472
rect 23636 25432 26860 25472
rect 26900 25432 27532 25472
rect 27572 25432 29000 25472
rect 29347 25432 29356 25472
rect 29396 25432 30220 25472
rect 30260 25432 31796 25472
rect 32515 25432 32524 25472
rect 32564 25432 32573 25472
rect 32803 25432 32812 25472
rect 32852 25432 34348 25472
rect 34388 25432 34397 25472
rect 34531 25432 34540 25472
rect 34580 25432 34924 25472
rect 34964 25432 35116 25472
rect 35156 25432 35500 25472
rect 35540 25432 35549 25472
rect 38947 25432 38956 25472
rect 38996 25432 39005 25472
rect 40291 25432 40300 25472
rect 40340 25432 41396 25472
rect 42316 25432 44140 25472
rect 44180 25432 44189 25472
rect 44323 25432 44332 25472
rect 44372 25432 44812 25472
rect 44852 25432 44861 25472
rect 45859 25432 45868 25472
rect 45908 25432 46828 25472
rect 46868 25432 46877 25472
rect 32524 25388 32564 25432
rect 38956 25388 38996 25432
rect 42316 25388 42356 25432
rect 3427 25348 3436 25388
rect 3476 25348 4012 25388
rect 4052 25348 4061 25388
rect 4387 25348 4396 25388
rect 4436 25348 7468 25388
rect 7508 25348 7852 25388
rect 7892 25348 11308 25388
rect 11348 25348 11357 25388
rect 16483 25348 16492 25388
rect 16532 25348 17452 25388
rect 17492 25348 17932 25388
rect 17972 25348 17981 25388
rect 18787 25348 18796 25388
rect 18836 25348 19372 25388
rect 19412 25348 19421 25388
rect 20140 25348 22828 25388
rect 22868 25348 22877 25388
rect 32524 25348 32948 25388
rect 34819 25348 34828 25388
rect 34868 25348 35308 25388
rect 35348 25348 38476 25388
rect 38516 25348 38996 25388
rect 41560 25348 41932 25388
rect 41972 25348 42316 25388
rect 42356 25348 42365 25388
rect 43843 25348 43852 25388
rect 43892 25348 45100 25388
rect 45140 25348 45149 25388
rect 20140 25304 20180 25348
rect 3523 25264 3532 25304
rect 3572 25264 4780 25304
rect 4820 25264 4972 25304
rect 5012 25264 5021 25304
rect 9091 25264 9100 25304
rect 9140 25264 10060 25304
rect 10100 25264 10109 25304
rect 11107 25264 11116 25304
rect 11156 25264 11596 25304
rect 11636 25264 11645 25304
rect 13795 25264 13804 25304
rect 13844 25264 14476 25304
rect 14516 25264 14525 25304
rect 14851 25264 14860 25304
rect 14900 25264 15244 25304
rect 15284 25264 15293 25304
rect 16099 25264 16108 25304
rect 16148 25264 16972 25304
rect 17012 25264 17740 25304
rect 17780 25264 20180 25304
rect 20515 25264 20524 25304
rect 20564 25264 22060 25304
rect 22100 25264 22109 25304
rect 26371 25264 26380 25304
rect 26420 25264 30604 25304
rect 30644 25264 30653 25304
rect 32908 25220 32948 25348
rect 41560 25304 41600 25348
rect 32995 25264 33004 25304
rect 33044 25264 34060 25304
rect 34100 25264 34109 25304
rect 34243 25264 34252 25304
rect 34292 25264 35212 25304
rect 35252 25264 35261 25304
rect 36067 25264 36076 25304
rect 36116 25264 36652 25304
rect 36692 25264 36701 25304
rect 39907 25264 39916 25304
rect 39956 25264 40492 25304
rect 40532 25264 40541 25304
rect 40675 25264 40684 25304
rect 40724 25264 41356 25304
rect 41396 25264 41600 25304
rect 41731 25264 41740 25304
rect 41780 25264 44564 25304
rect 44611 25264 44620 25304
rect 44660 25264 45772 25304
rect 45812 25264 45821 25304
rect 2659 25180 2668 25220
rect 2708 25180 3628 25220
rect 3668 25180 4492 25220
rect 4532 25180 5356 25220
rect 5396 25180 5405 25220
rect 6979 25180 6988 25220
rect 7028 25180 12940 25220
rect 12980 25180 13708 25220
rect 13748 25180 18028 25220
rect 18068 25180 18077 25220
rect 18211 25180 18220 25220
rect 18260 25180 25324 25220
rect 25364 25180 25373 25220
rect 31171 25180 31180 25220
rect 31220 25180 32428 25220
rect 32468 25180 32852 25220
rect 32908 25180 33292 25220
rect 33332 25180 33341 25220
rect 33388 25180 34156 25220
rect 34196 25180 34205 25220
rect 34339 25180 34348 25220
rect 34388 25180 34732 25220
rect 34772 25180 34781 25220
rect 35011 25180 35020 25220
rect 35060 25180 35596 25220
rect 35636 25180 35645 25220
rect 38851 25180 38860 25220
rect 38900 25180 40012 25220
rect 40052 25180 40876 25220
rect 40916 25180 40925 25220
rect 41539 25180 41548 25220
rect 41588 25180 44468 25220
rect 32812 25136 32852 25180
rect 33388 25136 33428 25180
rect 4204 25096 4396 25136
rect 4436 25096 4445 25136
rect 11299 25096 11308 25136
rect 11348 25096 12172 25136
rect 12212 25096 12221 25136
rect 14563 25096 14572 25136
rect 14612 25096 15244 25136
rect 15284 25096 17548 25136
rect 17588 25096 17836 25136
rect 17876 25096 17885 25136
rect 18499 25096 18508 25136
rect 18548 25096 19660 25136
rect 19700 25096 19709 25136
rect 32812 25096 33428 25136
rect 34156 25096 34636 25136
rect 34676 25096 34685 25136
rect 43171 25096 43180 25136
rect 43220 25096 44044 25136
rect 44084 25096 44332 25136
rect 44372 25096 44381 25136
rect 0 24908 80 24988
rect 4204 24968 4244 25096
rect 34156 25052 34196 25096
rect 11203 25012 11212 25052
rect 11252 25012 12364 25052
rect 12404 25012 12413 25052
rect 34147 25012 34156 25052
rect 34196 25012 34205 25052
rect 44428 24968 44468 25180
rect 44524 25052 44564 25264
rect 44707 25180 44716 25220
rect 44756 25180 46252 25220
rect 46292 25180 46301 25220
rect 47683 25180 47692 25220
rect 47732 25180 48460 25220
rect 48500 25180 48509 25220
rect 44524 25012 44812 25052
rect 44852 25012 44861 25052
rect 46243 25012 46252 25052
rect 46292 25012 47404 25052
rect 47444 25012 48172 25052
rect 48212 25012 48221 25052
rect 4195 24928 4204 24968
rect 4244 24928 4253 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 11971 24928 11980 24968
rect 12020 24928 12460 24968
rect 12500 24928 14188 24968
rect 14228 24928 14237 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 41443 24928 41452 24968
rect 41492 24928 43948 24968
rect 43988 24928 44236 24968
rect 44276 24928 44285 24968
rect 44428 24928 44908 24968
rect 44948 24928 44957 24968
rect 45763 24928 45772 24968
rect 45812 24928 46540 24968
rect 46580 24928 46589 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 10339 24844 10348 24884
rect 10388 24844 13516 24884
rect 13556 24844 13565 24884
rect 16195 24844 16204 24884
rect 16244 24844 23788 24884
rect 23828 24844 23837 24884
rect 28099 24844 28108 24884
rect 28148 24844 28876 24884
rect 28916 24844 28925 24884
rect 44323 24844 44332 24884
rect 44372 24844 45676 24884
rect 45716 24844 46292 24884
rect 46339 24844 46348 24884
rect 46388 24844 46924 24884
rect 46964 24844 46973 24884
rect 46252 24800 46292 24844
rect 8131 24760 8140 24800
rect 8180 24760 10252 24800
rect 10292 24760 10301 24800
rect 16387 24760 16396 24800
rect 16436 24760 20180 24800
rect 25123 24760 25132 24800
rect 25172 24760 25804 24800
rect 25844 24760 25853 24800
rect 44515 24760 44524 24800
rect 44564 24760 45100 24800
rect 45140 24760 45149 24800
rect 46243 24760 46252 24800
rect 46292 24760 46301 24800
rect 46531 24760 46540 24800
rect 46580 24760 47500 24800
rect 47540 24760 47549 24800
rect 20140 24716 20180 24760
rect 10819 24676 10828 24716
rect 10868 24676 11828 24716
rect 13699 24676 13708 24716
rect 13748 24676 14380 24716
rect 14420 24676 14429 24716
rect 14851 24676 14860 24716
rect 14900 24676 15244 24716
rect 15284 24676 15293 24716
rect 20140 24676 27956 24716
rect 11788 24632 11828 24676
rect 27916 24632 27956 24676
rect 34060 24676 38476 24716
rect 38516 24676 38525 24716
rect 43939 24676 43948 24716
rect 43988 24676 45772 24716
rect 45812 24676 45821 24716
rect 48259 24676 48268 24716
rect 48308 24676 48940 24716
rect 48980 24676 48989 24716
rect 1123 24592 1132 24632
rect 1172 24592 2764 24632
rect 2804 24592 2813 24632
rect 8035 24592 8044 24632
rect 8084 24592 9292 24632
rect 9332 24592 9341 24632
rect 10915 24592 10924 24632
rect 10964 24592 11360 24632
rect 11779 24592 11788 24632
rect 11828 24592 11837 24632
rect 12739 24592 12748 24632
rect 12788 24592 13420 24632
rect 13460 24592 13469 24632
rect 14083 24592 14092 24632
rect 14132 24592 14141 24632
rect 15043 24592 15052 24632
rect 15092 24592 15820 24632
rect 15860 24592 15869 24632
rect 16003 24592 16012 24632
rect 16052 24592 16396 24632
rect 16436 24592 16445 24632
rect 17827 24592 17836 24632
rect 17876 24592 22444 24632
rect 22484 24592 22493 24632
rect 27907 24592 27916 24632
rect 27956 24592 27965 24632
rect 28579 24592 28588 24632
rect 28628 24592 29000 24632
rect 30595 24592 30604 24632
rect 30644 24592 33964 24632
rect 34004 24592 34013 24632
rect 11320 24548 11360 24592
rect 14092 24548 14132 24592
rect 19171 24548 19229 24549
rect 28960 24548 29000 24592
rect 34060 24548 34100 24676
rect 44899 24592 44908 24632
rect 44948 24592 45676 24632
rect 45716 24592 45725 24632
rect 46600 24592 47212 24632
rect 47252 24592 51820 24632
rect 51860 24592 51869 24632
rect 46600 24548 46640 24592
rect 3523 24508 3532 24548
rect 3572 24508 4108 24548
rect 4148 24508 4492 24548
rect 4532 24508 4541 24548
rect 11320 24508 14132 24548
rect 14476 24508 17644 24548
rect 17684 24508 17693 24548
rect 19171 24508 19180 24548
rect 19220 24508 22252 24548
rect 22292 24508 22301 24548
rect 28960 24508 34100 24548
rect 35875 24508 35884 24548
rect 35924 24508 36172 24548
rect 36212 24508 37324 24548
rect 37364 24508 37373 24548
rect 40963 24508 40972 24548
rect 41012 24508 46640 24548
rect 48163 24508 48172 24548
rect 48212 24508 48652 24548
rect 48692 24508 48701 24548
rect 14476 24464 14516 24508
rect 19171 24507 19229 24508
rect 10051 24424 10060 24464
rect 10100 24424 10444 24464
rect 10484 24424 10493 24464
rect 11320 24424 14516 24464
rect 15907 24424 15916 24464
rect 15956 24424 16684 24464
rect 16724 24424 16733 24464
rect 40483 24424 40492 24464
rect 40532 24424 45004 24464
rect 45044 24424 45053 24464
rect 11320 24380 11360 24424
rect 4867 24340 4876 24380
rect 4916 24340 11360 24380
rect 12931 24340 12940 24380
rect 12980 24340 13132 24380
rect 13172 24340 13181 24380
rect 13891 24340 13900 24380
rect 13940 24340 14476 24380
rect 14516 24340 14525 24380
rect 5347 24256 5356 24296
rect 5396 24256 7468 24296
rect 7508 24256 8044 24296
rect 8084 24256 8093 24296
rect 10723 24256 10732 24296
rect 10772 24256 12500 24296
rect 14179 24256 14188 24296
rect 14228 24256 15092 24296
rect 36835 24256 36844 24296
rect 36884 24256 38284 24296
rect 38324 24256 38333 24296
rect 41059 24256 41068 24296
rect 41108 24256 41600 24296
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 0 24068 80 24148
rect 12460 24044 12500 24256
rect 15052 24212 15092 24256
rect 24451 24212 24509 24213
rect 41560 24212 41600 24256
rect 15043 24172 15052 24212
rect 15092 24172 15101 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 24432 24172 24460 24212
rect 24500 24172 24556 24212
rect 24596 24172 25804 24212
rect 25844 24172 25853 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 41560 24172 48268 24212
rect 48308 24172 48317 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 24451 24171 24509 24172
rect 14179 24088 14188 24128
rect 14228 24088 15244 24128
rect 15284 24088 15628 24128
rect 15668 24088 15677 24128
rect 23203 24088 23212 24128
rect 23252 24088 23261 24128
rect 28291 24088 28300 24128
rect 28340 24088 28349 24128
rect 19171 24044 19229 24045
rect 4003 24004 4012 24044
rect 4052 24004 4396 24044
rect 4436 24004 5260 24044
rect 5300 24004 5836 24044
rect 5876 24004 5885 24044
rect 6787 24004 6796 24044
rect 6836 24004 8620 24044
rect 8660 24004 8669 24044
rect 10051 24004 10060 24044
rect 10100 24004 11116 24044
rect 11156 24004 11165 24044
rect 12460 24004 13708 24044
rect 13748 24004 15340 24044
rect 15380 24004 16204 24044
rect 16244 24004 16588 24044
rect 16628 24004 16637 24044
rect 19086 24004 19180 24044
rect 19220 24004 19229 24044
rect 3523 23920 3532 23960
rect 3572 23920 5740 23960
rect 5780 23920 5789 23960
rect 6307 23920 6316 23960
rect 6356 23920 7756 23960
rect 7796 23920 7805 23960
rect 3532 23876 3572 23920
rect 12460 23876 12500 24004
rect 19171 24003 19229 24004
rect 23212 23960 23252 24088
rect 28300 23960 28340 24088
rect 12835 23920 12844 23960
rect 12884 23920 13612 23960
rect 13652 23920 14284 23960
rect 14324 23920 14333 23960
rect 14659 23920 14668 23960
rect 14708 23920 15532 23960
rect 15572 23920 15581 23960
rect 16387 23920 16396 23960
rect 16436 23920 17068 23960
rect 17108 23920 17117 23960
rect 19075 23920 19084 23960
rect 19124 23920 19796 23960
rect 23212 23920 23540 23960
rect 26851 23920 26860 23960
rect 26900 23920 28876 23960
rect 28916 23920 28925 23960
rect 49507 23920 49516 23960
rect 49556 23920 50764 23960
rect 50804 23920 50813 23960
rect 2371 23836 2380 23876
rect 2420 23836 3572 23876
rect 3811 23836 3820 23876
rect 3860 23836 4684 23876
rect 4724 23836 5644 23876
rect 5684 23836 5693 23876
rect 12451 23836 12460 23876
rect 12500 23836 12509 23876
rect 14083 23836 14092 23876
rect 14132 23836 14764 23876
rect 14804 23836 14813 23876
rect 15139 23836 15148 23876
rect 15188 23836 15197 23876
rect 16675 23836 16684 23876
rect 16724 23836 17548 23876
rect 17588 23836 19660 23876
rect 19700 23836 19709 23876
rect 15148 23792 15188 23836
rect 19756 23792 19796 23920
rect 23500 23876 23540 23920
rect 20035 23836 20044 23876
rect 20084 23836 20620 23876
rect 20660 23836 20669 23876
rect 23500 23836 25172 23876
rect 26659 23836 26668 23876
rect 26708 23836 27244 23876
rect 27284 23836 27532 23876
rect 27572 23836 27581 23876
rect 27715 23836 27724 23876
rect 27764 23836 28972 23876
rect 29012 23836 29021 23876
rect 29155 23836 29164 23876
rect 29204 23836 30836 23876
rect 34339 23836 34348 23876
rect 34388 23836 43372 23876
rect 43412 23836 43421 23876
rect 23500 23792 23540 23836
rect 2275 23752 2284 23792
rect 2324 23752 2572 23792
rect 2612 23752 2621 23792
rect 3043 23752 3052 23792
rect 3092 23752 3101 23792
rect 3619 23752 3628 23792
rect 3668 23752 4204 23792
rect 4244 23752 4780 23792
rect 4820 23752 4829 23792
rect 8611 23752 8620 23792
rect 8660 23752 10156 23792
rect 10196 23752 11308 23792
rect 11348 23752 11357 23792
rect 12547 23752 12556 23792
rect 12596 23752 12940 23792
rect 12980 23752 12989 23792
rect 15148 23752 16780 23792
rect 16820 23752 19276 23792
rect 19316 23752 19325 23792
rect 19747 23752 19756 23792
rect 19796 23752 19805 23792
rect 22915 23752 22924 23792
rect 22964 23752 23308 23792
rect 23348 23752 23357 23792
rect 23491 23752 23500 23792
rect 23540 23752 23549 23792
rect 23875 23752 23884 23792
rect 23924 23752 23933 23792
rect 24067 23752 24076 23792
rect 24116 23752 24652 23792
rect 24692 23752 24701 23792
rect 3052 23708 3092 23752
rect 23884 23708 23924 23752
rect 3052 23668 5932 23708
rect 5972 23668 5981 23708
rect 8515 23668 8524 23708
rect 8564 23668 9772 23708
rect 9812 23668 11404 23708
rect 11444 23668 11453 23708
rect 13987 23668 13996 23708
rect 14036 23668 15052 23708
rect 15092 23668 15101 23708
rect 22723 23668 22732 23708
rect 22772 23668 23404 23708
rect 23444 23668 23453 23708
rect 23884 23668 24844 23708
rect 24884 23668 24893 23708
rect 25132 23624 25172 23836
rect 25315 23792 25373 23793
rect 25699 23792 25757 23793
rect 25230 23752 25324 23792
rect 25364 23752 25373 23792
rect 25614 23752 25708 23792
rect 25748 23752 25757 23792
rect 26083 23752 26092 23792
rect 26132 23752 27628 23792
rect 27668 23752 27677 23792
rect 27907 23752 27916 23792
rect 27956 23752 28492 23792
rect 28532 23752 28541 23792
rect 28771 23752 28780 23792
rect 28820 23752 29452 23792
rect 29492 23752 29501 23792
rect 25315 23751 25373 23752
rect 25699 23751 25757 23752
rect 25708 23708 25748 23751
rect 25708 23668 26572 23708
rect 26612 23668 26621 23708
rect 27139 23668 27148 23708
rect 27188 23668 28204 23708
rect 28244 23668 28253 23708
rect 27724 23624 27764 23668
rect 3916 23584 4396 23624
rect 4436 23584 4445 23624
rect 4579 23584 4588 23624
rect 4628 23584 4972 23624
rect 5012 23584 5021 23624
rect 12259 23584 12268 23624
rect 12308 23584 12748 23624
rect 12788 23584 12797 23624
rect 14179 23584 14188 23624
rect 14228 23584 14668 23624
rect 14708 23584 14717 23624
rect 15235 23584 15244 23624
rect 15284 23584 15724 23624
rect 15764 23584 15773 23624
rect 17347 23584 17356 23624
rect 17396 23584 17740 23624
rect 17780 23584 17789 23624
rect 19651 23584 19660 23624
rect 19700 23584 19988 23624
rect 24163 23584 24172 23624
rect 24212 23584 25036 23624
rect 25076 23584 25085 23624
rect 25132 23584 26036 23624
rect 26179 23584 26188 23624
rect 26228 23584 27340 23624
rect 27380 23584 27389 23624
rect 27715 23584 27724 23624
rect 27764 23584 27773 23624
rect 28963 23584 28972 23624
rect 29012 23584 29452 23624
rect 29492 23584 29501 23624
rect 3916 23540 3956 23584
rect 3907 23500 3916 23540
rect 3956 23500 3965 23540
rect 14755 23500 14764 23540
rect 14804 23500 16972 23540
rect 17012 23500 17021 23540
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 5155 23416 5164 23456
rect 5204 23416 14956 23456
rect 14996 23416 15005 23456
rect 15331 23416 15340 23456
rect 15380 23416 15532 23456
rect 15572 23416 15581 23456
rect 16099 23416 16108 23456
rect 16148 23416 19276 23456
rect 19316 23416 19325 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 19948 23372 19988 23584
rect 24355 23540 24413 23541
rect 25996 23540 26036 23584
rect 23203 23500 23212 23540
rect 23252 23500 23404 23540
rect 23444 23500 24364 23540
rect 24404 23500 25940 23540
rect 25996 23500 26476 23540
rect 26516 23500 26525 23540
rect 27340 23500 29396 23540
rect 24355 23499 24413 23500
rect 25900 23456 25940 23500
rect 27340 23456 27380 23500
rect 25900 23416 27380 23456
rect 27523 23416 27532 23456
rect 27572 23416 27820 23456
rect 27860 23416 28588 23456
rect 28628 23416 29260 23456
rect 29300 23416 29309 23456
rect 28195 23372 28253 23373
rect 29356 23372 29396 23500
rect 29548 23456 29588 23836
rect 30796 23792 30836 23836
rect 30787 23752 30796 23792
rect 30836 23752 31468 23792
rect 31508 23752 31517 23792
rect 35779 23752 35788 23792
rect 35828 23752 36748 23792
rect 36788 23752 37516 23792
rect 37556 23752 37565 23792
rect 37699 23752 37708 23792
rect 37748 23752 38188 23792
rect 38228 23752 38237 23792
rect 41827 23752 41836 23792
rect 41876 23752 42988 23792
rect 43028 23752 44044 23792
rect 44084 23752 44620 23792
rect 44660 23752 44908 23792
rect 44948 23752 44957 23792
rect 37516 23708 37556 23752
rect 37516 23668 37900 23708
rect 37940 23668 37949 23708
rect 34819 23584 34828 23624
rect 34868 23584 35788 23624
rect 35828 23584 35837 23624
rect 37603 23584 37612 23624
rect 37652 23584 38956 23624
rect 38996 23584 39005 23624
rect 49123 23584 49132 23624
rect 49172 23584 51148 23624
rect 51188 23584 51197 23624
rect 37987 23500 37996 23540
rect 38036 23500 40588 23540
rect 40628 23500 41068 23540
rect 41108 23500 41117 23540
rect 41923 23500 41932 23540
rect 41972 23500 46348 23540
rect 46388 23500 46397 23540
rect 29443 23416 29452 23456
rect 29492 23416 29588 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 35779 23416 35788 23456
rect 35828 23416 40780 23456
rect 40820 23416 41740 23456
rect 41780 23416 41789 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 11395 23332 11404 23372
rect 11444 23332 12364 23372
rect 12404 23332 12413 23372
rect 13603 23332 13612 23372
rect 13652 23332 13804 23372
rect 13844 23332 13853 23372
rect 19756 23332 19988 23372
rect 24547 23332 24556 23372
rect 24596 23332 25036 23372
rect 25076 23332 25085 23372
rect 25219 23332 25228 23372
rect 25268 23332 25277 23372
rect 25411 23332 25420 23372
rect 25460 23332 26284 23372
rect 26324 23332 26333 23372
rect 27235 23332 27244 23372
rect 27284 23332 28204 23372
rect 28244 23332 28253 23372
rect 0 23228 80 23308
rect 19756 23288 19796 23332
rect 25123 23288 25181 23289
rect 25228 23288 25268 23332
rect 28195 23331 28253 23332
rect 28300 23332 29068 23372
rect 29108 23332 29117 23372
rect 29356 23332 30700 23372
rect 30740 23332 30892 23372
rect 30932 23332 30941 23372
rect 35107 23332 35116 23372
rect 35156 23332 37132 23372
rect 37172 23332 37181 23372
rect 37411 23332 37420 23372
rect 37460 23332 37804 23372
rect 37844 23332 38860 23372
rect 38900 23332 38909 23372
rect 3331 23248 3340 23288
rect 3380 23248 6028 23288
rect 6068 23248 6077 23288
rect 6499 23248 6508 23288
rect 6548 23248 7180 23288
rect 7220 23248 7229 23288
rect 12067 23248 12076 23288
rect 12116 23248 12652 23288
rect 12692 23248 12701 23288
rect 14851 23248 14860 23288
rect 14900 23248 15628 23288
rect 15668 23248 15677 23288
rect 19747 23248 19756 23288
rect 19796 23248 19805 23288
rect 25123 23248 25132 23288
rect 25172 23248 25268 23288
rect 25411 23288 25469 23289
rect 28300 23288 28340 23332
rect 25411 23248 25420 23288
rect 25460 23248 26092 23288
rect 26132 23248 26141 23288
rect 27427 23248 27436 23288
rect 27476 23248 28300 23288
rect 28340 23248 28349 23288
rect 28771 23248 28780 23288
rect 28820 23248 29740 23288
rect 29780 23248 29789 23288
rect 35683 23248 35692 23288
rect 35732 23248 36556 23288
rect 36596 23248 36605 23288
rect 37219 23248 37228 23288
rect 37268 23248 43084 23288
rect 43124 23248 43133 23288
rect 44803 23248 44812 23288
rect 44852 23248 45004 23288
rect 45044 23248 49132 23288
rect 49172 23248 49181 23288
rect 25123 23247 25181 23248
rect 25411 23247 25469 23248
rect 1219 23164 1228 23204
rect 1268 23164 3148 23204
rect 3188 23164 3197 23204
rect 4963 23164 4972 23204
rect 5012 23164 5740 23204
rect 5780 23164 5789 23204
rect 6115 23164 6124 23204
rect 6164 23164 7468 23204
rect 7508 23164 7517 23204
rect 8227 23164 8236 23204
rect 8276 23164 8620 23204
rect 8660 23164 9868 23204
rect 9908 23164 9917 23204
rect 11320 23164 15340 23204
rect 15380 23164 15389 23204
rect 23884 23164 25612 23204
rect 25652 23164 26764 23204
rect 26804 23164 26813 23204
rect 28099 23164 28108 23204
rect 28148 23164 29164 23204
rect 29204 23164 29548 23204
rect 29588 23164 29597 23204
rect 31171 23164 31180 23204
rect 31220 23164 31852 23204
rect 31892 23164 31901 23204
rect 35875 23164 35884 23204
rect 35924 23164 36884 23204
rect 45763 23164 45772 23204
rect 45812 23164 47404 23204
rect 47444 23164 47453 23204
rect 11320 23120 11360 23164
rect 23884 23120 23924 23164
rect 24451 23120 24509 23121
rect 36844 23120 36884 23164
rect 4195 23080 4204 23120
rect 4244 23080 5452 23120
rect 5492 23080 5501 23120
rect 6691 23080 6700 23120
rect 6740 23080 6988 23120
rect 7028 23080 7037 23120
rect 7267 23080 7276 23120
rect 7316 23080 8332 23120
rect 8372 23080 8381 23120
rect 9955 23080 9964 23120
rect 10004 23080 11360 23120
rect 12547 23080 12556 23120
rect 12596 23080 13516 23120
rect 13556 23080 13565 23120
rect 13987 23080 13996 23120
rect 14036 23080 15724 23120
rect 15764 23080 15773 23120
rect 17443 23080 17452 23120
rect 17492 23080 19372 23120
rect 19412 23080 20620 23120
rect 20660 23080 20669 23120
rect 23875 23080 23884 23120
rect 23924 23080 23933 23120
rect 24366 23080 24460 23120
rect 24500 23080 24509 23120
rect 24739 23080 24748 23120
rect 24788 23080 26092 23120
rect 26132 23080 26141 23120
rect 28108 23080 28972 23120
rect 29012 23080 29021 23120
rect 30115 23080 30124 23120
rect 30164 23080 30412 23120
rect 30452 23080 30796 23120
rect 30836 23080 30845 23120
rect 31075 23080 31084 23120
rect 31124 23080 31756 23120
rect 31796 23080 31805 23120
rect 35299 23080 35308 23120
rect 35348 23080 36460 23120
rect 36500 23080 36509 23120
rect 36835 23080 36844 23120
rect 36884 23080 37804 23120
rect 37844 23080 37853 23120
rect 43555 23080 43564 23120
rect 43604 23080 46156 23120
rect 46196 23080 47980 23120
rect 48020 23080 49900 23120
rect 49940 23080 50668 23120
rect 50708 23080 50717 23120
rect 24451 23079 24509 23080
rect 6307 22996 6316 23036
rect 6356 22996 7084 23036
rect 7124 22996 8236 23036
rect 8276 22996 8285 23036
rect 24460 22952 24500 23079
rect 25123 23036 25181 23037
rect 28108 23036 28148 23080
rect 25038 22996 25132 23036
rect 25172 22996 25181 23036
rect 25315 22996 25324 23036
rect 25364 22996 26284 23036
rect 26324 22996 26333 23036
rect 28099 22996 28108 23036
rect 28148 22996 28157 23036
rect 28675 22996 28684 23036
rect 28724 22996 31276 23036
rect 31316 22996 31325 23036
rect 35683 22996 35692 23036
rect 35732 22996 37324 23036
rect 37364 22996 37996 23036
rect 38036 22996 39340 23036
rect 39380 22996 39389 23036
rect 41443 22996 41452 23036
rect 41492 22996 44140 23036
rect 44180 22996 44428 23036
rect 44468 22996 44477 23036
rect 25123 22995 25181 22996
rect 28684 22952 28724 22996
rect 4003 22912 4012 22952
rect 4052 22912 4492 22952
rect 4532 22912 4541 22952
rect 24460 22912 25036 22952
rect 25076 22912 25085 22952
rect 25891 22912 25900 22952
rect 25940 22912 26668 22952
rect 26708 22912 28724 22952
rect 28867 22912 28876 22952
rect 28916 22912 29932 22952
rect 29972 22912 29981 22952
rect 34243 22912 34252 22952
rect 34292 22912 35020 22952
rect 35060 22912 35980 22952
rect 36020 22912 36029 22952
rect 41539 22912 41548 22952
rect 41588 22912 42220 22952
rect 42260 22912 42269 22952
rect 43747 22912 43756 22952
rect 43796 22912 44812 22952
rect 44852 22912 45004 22952
rect 45044 22912 45053 22952
rect 24460 22868 24500 22912
rect 35491 22868 35549 22869
rect 1219 22828 1228 22868
rect 1268 22828 3916 22868
rect 3956 22828 3965 22868
rect 23308 22828 24500 22868
rect 24739 22828 24748 22868
rect 24788 22828 26380 22868
rect 26420 22828 27052 22868
rect 27092 22828 28588 22868
rect 28628 22828 28637 22868
rect 35406 22828 35500 22868
rect 35540 22828 35549 22868
rect 40003 22828 40012 22868
rect 40052 22828 40588 22868
rect 40628 22828 43180 22868
rect 43220 22828 43229 22868
rect 23308 22784 23348 22828
rect 35491 22827 35549 22828
rect 24739 22784 24797 22785
rect 23299 22744 23308 22784
rect 23348 22744 23357 22784
rect 23587 22744 23596 22784
rect 23636 22744 24556 22784
rect 24596 22744 24605 22784
rect 24739 22744 24748 22784
rect 24788 22744 27724 22784
rect 27764 22744 27773 22784
rect 41059 22744 41068 22784
rect 41108 22744 42700 22784
rect 42740 22744 42749 22784
rect 24739 22743 24797 22744
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 5539 22660 5548 22700
rect 5588 22660 8716 22700
rect 8756 22660 9292 22700
rect 9332 22660 9341 22700
rect 10627 22660 10636 22700
rect 10676 22660 12172 22700
rect 12212 22660 12364 22700
rect 12404 22660 12413 22700
rect 12739 22660 12748 22700
rect 12788 22660 13612 22700
rect 13652 22660 13661 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 23779 22660 23788 22700
rect 23828 22660 24076 22700
rect 24116 22660 24125 22700
rect 25603 22660 25612 22700
rect 25652 22660 26092 22700
rect 26132 22660 26141 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 38083 22660 38092 22700
rect 38132 22660 38572 22700
rect 38612 22660 39820 22700
rect 39860 22660 41300 22700
rect 41347 22660 41356 22700
rect 41396 22660 42028 22700
rect 42068 22660 42077 22700
rect 42307 22660 42316 22700
rect 42356 22660 42892 22700
rect 42932 22660 42941 22700
rect 46147 22660 46156 22700
rect 46196 22660 47020 22700
rect 47060 22660 47069 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 25315 22616 25373 22617
rect 8419 22576 8428 22616
rect 8468 22576 9388 22616
rect 9428 22576 9772 22616
rect 9812 22576 9821 22616
rect 23875 22576 23884 22616
rect 23924 22576 25324 22616
rect 25364 22576 25373 22616
rect 25315 22575 25373 22576
rect 25507 22616 25565 22617
rect 41260 22616 41300 22660
rect 25507 22576 25516 22616
rect 25556 22576 27532 22616
rect 27572 22576 27581 22616
rect 41260 22576 41600 22616
rect 41731 22576 41740 22616
rect 41780 22576 45484 22616
rect 45524 22576 45533 22616
rect 25507 22575 25565 22576
rect 41560 22532 41600 22576
rect 11395 22492 11404 22532
rect 11444 22492 11884 22532
rect 11924 22492 11933 22532
rect 16963 22492 16972 22532
rect 17012 22492 19180 22532
rect 19220 22492 19229 22532
rect 23491 22492 23500 22532
rect 23540 22492 24460 22532
rect 24500 22492 25132 22532
rect 25172 22492 25181 22532
rect 32899 22492 32908 22532
rect 32948 22492 33964 22532
rect 34004 22492 34013 22532
rect 38755 22492 38764 22532
rect 38804 22492 39052 22532
rect 39092 22492 40204 22532
rect 40244 22492 40684 22532
rect 40724 22492 40733 22532
rect 41560 22492 41644 22532
rect 41684 22492 41693 22532
rect 42115 22492 42124 22532
rect 42164 22492 46540 22532
rect 46580 22492 46589 22532
rect 0 22448 80 22468
rect 24739 22448 24797 22449
rect 0 22408 652 22448
rect 692 22408 701 22448
rect 6403 22408 6412 22448
rect 6452 22408 7756 22448
rect 7796 22408 7805 22448
rect 13411 22408 13420 22448
rect 13460 22408 13996 22448
rect 14036 22408 14045 22448
rect 15139 22408 15148 22448
rect 15188 22408 15436 22448
rect 15476 22408 15485 22448
rect 17635 22408 17644 22448
rect 17684 22408 18508 22448
rect 18548 22408 18557 22448
rect 24547 22408 24556 22448
rect 24596 22408 24748 22448
rect 24788 22408 24797 22448
rect 40387 22408 40396 22448
rect 40436 22408 46924 22448
rect 46964 22408 46973 22448
rect 0 22388 80 22408
rect 24739 22407 24797 22408
rect 44716 22364 44756 22408
rect 12931 22324 12940 22364
rect 12980 22324 13228 22364
rect 13268 22324 18124 22364
rect 18164 22324 18173 22364
rect 23107 22324 23116 22364
rect 23156 22324 24364 22364
rect 24404 22324 25132 22364
rect 25172 22324 25181 22364
rect 28579 22324 28588 22364
rect 28628 22324 29164 22364
rect 29204 22324 29213 22364
rect 44707 22324 44716 22364
rect 44756 22324 44765 22364
rect 2467 22240 2476 22280
rect 2516 22240 3148 22280
rect 3188 22240 3197 22280
rect 3619 22240 3628 22280
rect 3668 22240 4300 22280
rect 4340 22240 4876 22280
rect 4916 22240 4925 22280
rect 6499 22240 6508 22280
rect 6548 22240 8140 22280
rect 8180 22240 8189 22280
rect 9187 22240 9196 22280
rect 9236 22240 9388 22280
rect 9428 22240 11020 22280
rect 11060 22240 11069 22280
rect 14275 22240 14284 22280
rect 14324 22240 15532 22280
rect 15572 22240 16204 22280
rect 16244 22240 16253 22280
rect 18211 22240 18220 22280
rect 18260 22240 19948 22280
rect 19988 22240 19997 22280
rect 23683 22240 23692 22280
rect 23732 22240 25420 22280
rect 25460 22240 25469 22280
rect 26563 22240 26572 22280
rect 26612 22240 27244 22280
rect 27284 22240 27293 22280
rect 28867 22240 28876 22280
rect 28916 22240 31180 22280
rect 31220 22240 31229 22280
rect 37507 22240 37516 22280
rect 37556 22240 38668 22280
rect 38708 22240 38717 22280
rect 38947 22240 38956 22280
rect 38996 22240 42028 22280
rect 42068 22240 42077 22280
rect 2851 22156 2860 22196
rect 2900 22156 4108 22196
rect 4148 22156 5164 22196
rect 5204 22156 5213 22196
rect 6115 22156 6124 22196
rect 6164 22156 6604 22196
rect 6644 22156 7948 22196
rect 7988 22156 8428 22196
rect 8468 22156 8477 22196
rect 16780 22156 18892 22196
rect 18932 22156 18941 22196
rect 24643 22156 24652 22196
rect 24692 22156 26188 22196
rect 26228 22156 26237 22196
rect 26467 22156 26476 22196
rect 26516 22156 27052 22196
rect 27092 22156 27916 22196
rect 27956 22156 28780 22196
rect 28820 22156 28829 22196
rect 36259 22156 36268 22196
rect 36308 22156 40396 22196
rect 40436 22156 40445 22196
rect 16780 22112 16820 22156
rect 13699 22072 13708 22112
rect 13748 22072 16780 22112
rect 16820 22072 16829 22112
rect 17059 22072 17068 22112
rect 17108 22072 18028 22112
rect 18068 22072 18077 22112
rect 24739 22072 24748 22112
rect 24788 22072 25036 22112
rect 25076 22072 25085 22112
rect 25219 22072 25228 22112
rect 25268 22072 25996 22112
rect 26036 22072 26045 22112
rect 29443 22072 29452 22112
rect 29492 22072 30892 22112
rect 30932 22072 35692 22112
rect 35732 22072 35741 22112
rect 41539 22072 41548 22112
rect 41588 22072 41932 22112
rect 41972 22072 41981 22112
rect 25699 22028 25757 22029
rect 25411 21988 25420 22028
rect 25460 21988 25708 22028
rect 25748 21988 25757 22028
rect 25699 21987 25757 21988
rect 25411 21944 25469 21945
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 25315 21904 25324 21944
rect 25364 21904 25420 21944
rect 25460 21904 25469 21944
rect 25891 21904 25900 21944
rect 25940 21904 28588 21944
rect 28628 21904 28637 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 25411 21903 25469 21904
rect 3907 21820 3916 21860
rect 3956 21820 5068 21860
rect 5108 21820 5117 21860
rect 5155 21736 5164 21776
rect 5204 21736 6836 21776
rect 8131 21736 8140 21776
rect 8180 21736 9004 21776
rect 9044 21736 10924 21776
rect 10964 21736 10973 21776
rect 25699 21736 25708 21776
rect 25748 21736 27436 21776
rect 27476 21736 27485 21776
rect 36931 21736 36940 21776
rect 36980 21736 37516 21776
rect 37556 21736 37565 21776
rect 44707 21736 44716 21776
rect 44756 21736 45388 21776
rect 45428 21736 45437 21776
rect 6796 21692 6836 21736
rect 24355 21692 24413 21693
rect 1795 21652 1804 21692
rect 1844 21652 2764 21692
rect 2804 21652 2813 21692
rect 2947 21652 2956 21692
rect 2996 21652 5836 21692
rect 5876 21652 5885 21692
rect 6787 21652 6796 21692
rect 6836 21652 8044 21692
rect 8084 21652 8093 21692
rect 10243 21652 10252 21692
rect 10292 21652 11596 21692
rect 11636 21652 11645 21692
rect 17251 21652 17260 21692
rect 17300 21652 17836 21692
rect 17876 21652 17885 21692
rect 24270 21652 24364 21692
rect 24404 21652 24413 21692
rect 25027 21652 25036 21692
rect 25076 21652 25228 21692
rect 25268 21652 25277 21692
rect 44515 21652 44524 21692
rect 44564 21652 47692 21692
rect 47732 21652 47741 21692
rect 24355 21651 24413 21652
rect 0 21608 80 21628
rect 35203 21608 35261 21609
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 2659 21568 2668 21608
rect 2708 21568 3820 21608
rect 3860 21568 3869 21608
rect 4099 21568 4108 21608
rect 4148 21568 6892 21608
rect 6932 21568 7660 21608
rect 7700 21568 7709 21608
rect 10339 21568 10348 21608
rect 10388 21568 11884 21608
rect 11924 21568 14284 21608
rect 14324 21568 14333 21608
rect 16867 21568 16876 21608
rect 16916 21568 18316 21608
rect 18356 21568 18365 21608
rect 24067 21568 24076 21608
rect 24116 21568 25612 21608
rect 25652 21568 25661 21608
rect 25795 21568 25804 21608
rect 25844 21568 26572 21608
rect 26612 21568 26621 21608
rect 27619 21568 27628 21608
rect 27668 21568 30988 21608
rect 31028 21568 31037 21608
rect 34339 21568 34348 21608
rect 34388 21568 35212 21608
rect 35252 21568 35788 21608
rect 35828 21568 35837 21608
rect 37315 21568 37324 21608
rect 37364 21568 38956 21608
rect 38996 21568 39005 21608
rect 39139 21568 39148 21608
rect 39188 21568 40300 21608
rect 40340 21568 40349 21608
rect 41155 21568 41164 21608
rect 41204 21568 41548 21608
rect 41588 21568 41597 21608
rect 44419 21568 44428 21608
rect 44468 21568 45484 21608
rect 45524 21568 45533 21608
rect 0 21548 80 21568
rect 35203 21567 35261 21568
rect 4003 21484 4012 21524
rect 4052 21484 5356 21524
rect 5396 21484 5932 21524
rect 5972 21484 5981 21524
rect 24460 21484 25708 21524
rect 25748 21484 25757 21524
rect 24460 21440 24500 21484
rect 4483 21400 4492 21440
rect 4532 21400 5108 21440
rect 5443 21400 5452 21440
rect 5492 21400 8044 21440
rect 8084 21400 8093 21440
rect 12931 21400 12940 21440
rect 12980 21400 13900 21440
rect 13940 21400 13949 21440
rect 18691 21400 18700 21440
rect 18740 21400 20236 21440
rect 20276 21400 21292 21440
rect 21332 21400 22444 21440
rect 22484 21400 23404 21440
rect 23444 21400 23453 21440
rect 24451 21400 24460 21440
rect 24500 21400 24509 21440
rect 25027 21400 25036 21440
rect 25076 21400 25516 21440
rect 25556 21400 25565 21440
rect 26371 21400 26380 21440
rect 26420 21400 27532 21440
rect 27572 21400 27581 21440
rect 40387 21400 40396 21440
rect 40436 21400 41452 21440
rect 41492 21400 43276 21440
rect 43316 21400 43325 21440
rect 5068 21272 5108 21400
rect 39907 21316 39916 21356
rect 39956 21316 40492 21356
rect 40532 21316 40541 21356
rect 5059 21232 5068 21272
rect 5108 21232 5117 21272
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 5539 20980 5548 21020
rect 5588 20980 6220 21020
rect 6260 20980 6269 21020
rect 37219 20980 37228 21020
rect 37268 20980 41644 21020
rect 41684 20980 41693 21020
rect 259 20896 268 20936
rect 308 20896 33292 20936
rect 33332 20896 33341 20936
rect 13987 20812 13996 20852
rect 14036 20812 14668 20852
rect 14708 20812 17260 20852
rect 17300 20812 17309 20852
rect 21283 20812 21292 20852
rect 21332 20812 22156 20852
rect 22196 20812 22205 20852
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 4195 20728 4204 20768
rect 4244 20728 5260 20768
rect 5300 20728 5309 20768
rect 9859 20728 9868 20768
rect 9908 20728 10348 20768
rect 10388 20728 10397 20768
rect 11491 20728 11500 20768
rect 11540 20728 12940 20768
rect 12980 20728 12989 20768
rect 15139 20728 15148 20768
rect 15188 20728 15628 20768
rect 15668 20728 15677 20768
rect 16675 20728 16684 20768
rect 16724 20728 18988 20768
rect 19028 20728 19037 20768
rect 20803 20728 20812 20768
rect 20852 20728 22348 20768
rect 22388 20728 22397 20768
rect 39043 20728 39052 20768
rect 39092 20728 39916 20768
rect 39956 20728 39965 20768
rect 0 20708 80 20728
rect 9283 20644 9292 20684
rect 9332 20644 9676 20684
rect 9716 20644 10828 20684
rect 10868 20644 10877 20684
rect 15331 20644 15340 20684
rect 15380 20644 15916 20684
rect 15956 20644 16876 20684
rect 16916 20644 16925 20684
rect 18115 20644 18124 20684
rect 18164 20644 29000 20684
rect 28960 20600 29000 20644
rect 8803 20560 8812 20600
rect 8852 20560 9580 20600
rect 9620 20560 10540 20600
rect 10580 20560 10589 20600
rect 15427 20560 15436 20600
rect 15476 20560 16396 20600
rect 16436 20560 16445 20600
rect 21091 20560 21100 20600
rect 21140 20560 21484 20600
rect 21524 20560 21533 20600
rect 21667 20560 21676 20600
rect 21716 20560 22636 20600
rect 22676 20560 22685 20600
rect 28960 20560 33292 20600
rect 33332 20560 33772 20600
rect 33812 20560 33821 20600
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 15148 20308 15244 20348
rect 15284 20308 15293 20348
rect 26083 20308 26092 20348
rect 26132 20308 27148 20348
rect 27188 20308 27197 20348
rect 6499 20224 6508 20264
rect 6548 20224 6796 20264
rect 6836 20224 6845 20264
rect 10819 20224 10828 20264
rect 10868 20224 11788 20264
rect 11828 20224 11837 20264
rect 11280 20140 11308 20180
rect 11348 20140 11444 20180
rect 11404 20096 11444 20140
rect 15148 20096 15188 20308
rect 18883 20224 18892 20264
rect 18932 20224 19660 20264
rect 19700 20224 19709 20264
rect 26275 20224 26284 20264
rect 26324 20224 26668 20264
rect 26708 20224 26717 20264
rect 34243 20224 34252 20264
rect 34292 20224 35596 20264
rect 35636 20224 35645 20264
rect 21859 20140 21868 20180
rect 21908 20140 22060 20180
rect 22100 20140 22109 20180
rect 25219 20140 25228 20180
rect 25268 20140 25420 20180
rect 25460 20140 26380 20180
rect 26420 20140 26429 20180
rect 16675 20096 16733 20097
rect 31939 20096 31997 20097
rect 5347 20056 5356 20096
rect 5396 20056 7948 20096
rect 7988 20056 7997 20096
rect 8995 20056 9004 20096
rect 9044 20056 9292 20096
rect 9332 20056 9341 20096
rect 11404 20056 12076 20096
rect 12116 20056 12125 20096
rect 15148 20056 15436 20096
rect 15476 20056 15485 20096
rect 15811 20056 15820 20096
rect 15860 20056 16300 20096
rect 16340 20056 16349 20096
rect 16590 20056 16684 20096
rect 16724 20056 16733 20096
rect 19267 20056 19276 20096
rect 19316 20056 20908 20096
rect 20948 20056 20957 20096
rect 21955 20056 21964 20096
rect 22004 20056 22444 20096
rect 22484 20056 22493 20096
rect 23395 20056 23404 20096
rect 23444 20056 26956 20096
rect 26996 20056 27005 20096
rect 27907 20056 27916 20096
rect 27956 20056 30316 20096
rect 30356 20056 30365 20096
rect 31939 20056 31948 20096
rect 31988 20056 32332 20096
rect 32372 20056 32381 20096
rect 40003 20056 40012 20096
rect 40052 20056 40396 20096
rect 40436 20056 40445 20096
rect 9004 20012 9044 20056
rect 16675 20055 16733 20056
rect 31939 20055 31997 20056
rect 16684 20012 16724 20055
rect 6979 19972 6988 20012
rect 7028 19972 7468 20012
rect 7508 19972 9044 20012
rect 10147 19972 10156 20012
rect 10196 19972 12556 20012
rect 12596 19972 14476 20012
rect 14516 19972 16724 20012
rect 18883 19972 18892 20012
rect 18932 19972 19372 20012
rect 19412 19972 21772 20012
rect 21812 19972 21821 20012
rect 26371 19972 26380 20012
rect 26420 19972 28012 20012
rect 28052 19972 28061 20012
rect 33091 19972 33100 20012
rect 33140 19972 33580 20012
rect 33620 19972 33629 20012
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 5731 19888 5740 19928
rect 5780 19888 6796 19928
rect 6836 19888 6845 19928
rect 7075 19888 7084 19928
rect 7124 19888 9196 19928
rect 9236 19888 9245 19928
rect 19459 19888 19468 19928
rect 19508 19888 21964 19928
rect 22004 19888 22013 19928
rect 24835 19888 24844 19928
rect 24884 19888 25228 19928
rect 25268 19888 25277 19928
rect 25699 19888 25708 19928
rect 25748 19888 26092 19928
rect 26132 19888 26141 19928
rect 28387 19888 28396 19928
rect 28436 19888 29932 19928
rect 29972 19888 29981 19928
rect 38659 19888 38668 19928
rect 38708 19888 40300 19928
rect 40340 19888 40349 19928
rect 0 19868 80 19888
rect 25027 19804 25036 19844
rect 25076 19804 26476 19844
rect 26516 19804 26525 19844
rect 31939 19804 31948 19844
rect 31988 19804 33196 19844
rect 33236 19804 33245 19844
rect 21859 19720 21868 19760
rect 21908 19720 26764 19760
rect 26804 19720 28300 19760
rect 28340 19720 28349 19760
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 25507 19552 25516 19592
rect 25556 19552 25996 19592
rect 26036 19552 26045 19592
rect 33955 19552 33964 19592
rect 34004 19552 35116 19592
rect 35156 19552 35500 19592
rect 35540 19552 35549 19592
rect 10339 19468 10348 19508
rect 10388 19468 10636 19508
rect 10676 19468 10685 19508
rect 14851 19468 14860 19508
rect 14900 19468 15148 19508
rect 15188 19468 15197 19508
rect 16291 19468 16300 19508
rect 16340 19468 17452 19508
rect 17492 19468 17501 19508
rect 21955 19468 21964 19508
rect 22004 19468 22540 19508
rect 22580 19468 22589 19508
rect 3715 19384 3724 19424
rect 3764 19384 4492 19424
rect 4532 19384 4541 19424
rect 5827 19384 5836 19424
rect 5876 19384 6892 19424
rect 6932 19384 6941 19424
rect 15715 19384 15724 19424
rect 15764 19384 15773 19424
rect 17923 19384 17932 19424
rect 17972 19384 19276 19424
rect 19316 19384 19325 19424
rect 22147 19384 22156 19424
rect 22196 19384 22636 19424
rect 22676 19384 22685 19424
rect 4195 19340 4253 19341
rect 4110 19300 4204 19340
rect 4244 19300 4253 19340
rect 8899 19300 8908 19340
rect 8948 19300 11308 19340
rect 11348 19300 11357 19340
rect 4195 19299 4253 19300
rect 3724 19216 4492 19256
rect 4532 19216 4541 19256
rect 6115 19216 6124 19256
rect 6164 19216 10636 19256
rect 10676 19216 10828 19256
rect 10868 19216 10877 19256
rect 11779 19216 11788 19256
rect 11828 19216 12076 19256
rect 12116 19216 12125 19256
rect 3724 19172 3764 19216
rect 3715 19132 3724 19172
rect 3764 19132 3773 19172
rect 4204 19132 4780 19172
rect 4820 19132 6028 19172
rect 6068 19132 7852 19172
rect 7892 19132 8332 19172
rect 8372 19132 8381 19172
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 1315 19048 1324 19088
rect 1364 19048 4108 19088
rect 4148 19048 4157 19088
rect 0 19028 80 19048
rect 4204 19004 4244 19132
rect 15724 19088 15764 19384
rect 28579 19340 28637 19341
rect 19555 19300 19564 19340
rect 19604 19300 20716 19340
rect 20756 19300 22828 19340
rect 22868 19300 22877 19340
rect 24931 19300 24940 19340
rect 24980 19300 28588 19340
rect 28628 19300 28684 19340
rect 28724 19300 31660 19340
rect 31700 19300 31709 19340
rect 28579 19299 28637 19300
rect 26659 19256 26717 19257
rect 16291 19216 16300 19256
rect 16340 19216 19372 19256
rect 19412 19216 19421 19256
rect 20803 19216 20812 19256
rect 20852 19216 21004 19256
rect 21044 19216 21053 19256
rect 22531 19216 22540 19256
rect 22580 19216 23500 19256
rect 23540 19216 23549 19256
rect 26574 19216 26668 19256
rect 26708 19216 26717 19256
rect 30787 19216 30796 19256
rect 30836 19216 32812 19256
rect 32852 19216 33004 19256
rect 33044 19216 33053 19256
rect 33955 19216 33964 19256
rect 34004 19216 34444 19256
rect 34484 19216 34493 19256
rect 35395 19216 35404 19256
rect 35444 19216 36364 19256
rect 36404 19216 36940 19256
rect 36980 19216 36989 19256
rect 39715 19216 39724 19256
rect 39764 19216 40684 19256
rect 40724 19216 40733 19256
rect 26659 19215 26717 19216
rect 32419 19172 32477 19173
rect 32334 19132 32428 19172
rect 32468 19132 32477 19172
rect 32419 19131 32477 19132
rect 18691 19088 18749 19089
rect 34243 19088 34301 19089
rect 12163 19048 12172 19088
rect 12212 19048 13132 19088
rect 13172 19048 13181 19088
rect 15619 19048 15628 19088
rect 15668 19048 17644 19088
rect 17684 19048 17693 19088
rect 18019 19048 18028 19088
rect 18068 19048 18700 19088
rect 18740 19048 27148 19088
rect 27188 19048 30604 19088
rect 30644 19048 30653 19088
rect 33187 19048 33196 19088
rect 33236 19048 34060 19088
rect 34100 19048 34109 19088
rect 34243 19048 34252 19088
rect 34292 19048 35308 19088
rect 35348 19048 35357 19088
rect 38851 19048 38860 19088
rect 38900 19048 40012 19088
rect 40052 19048 40061 19088
rect 18691 19047 18749 19048
rect 34243 19047 34301 19048
rect 25699 19004 25757 19005
rect 4195 18964 4204 19004
rect 4244 18964 4253 19004
rect 25699 18964 25708 19004
rect 25748 18964 25899 19004
rect 25939 18964 25948 19004
rect 28099 18964 28108 19004
rect 28148 18964 28780 19004
rect 28820 18964 31468 19004
rect 31508 18964 31852 19004
rect 31892 18964 31901 19004
rect 33955 18964 33964 19004
rect 34004 18964 34156 19004
rect 34196 18964 34205 19004
rect 25699 18963 25757 18964
rect 23107 18920 23165 18921
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 6979 18880 6988 18920
rect 7028 18880 7756 18920
rect 7796 18880 7948 18920
rect 7988 18880 10156 18920
rect 10196 18880 10205 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 20995 18880 21004 18920
rect 21044 18880 21868 18920
rect 21908 18880 21917 18920
rect 22243 18880 22252 18920
rect 22292 18880 22301 18920
rect 23107 18880 23116 18920
rect 23156 18880 23308 18920
rect 23348 18880 23357 18920
rect 25603 18880 25612 18920
rect 25652 18880 26764 18920
rect 26804 18880 28204 18920
rect 28244 18880 28253 18920
rect 28579 18880 28588 18920
rect 28628 18880 28972 18920
rect 29012 18880 29021 18920
rect 33859 18880 33868 18920
rect 33908 18880 34252 18920
rect 34292 18880 34301 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 22252 18836 22292 18880
rect 23107 18879 23165 18880
rect 6307 18796 6316 18836
rect 6356 18796 7660 18836
rect 7700 18796 7709 18836
rect 10435 18796 10444 18836
rect 10484 18796 13324 18836
rect 13364 18796 13373 18836
rect 20899 18796 20908 18836
rect 20948 18796 26708 18836
rect 31843 18796 31852 18836
rect 31892 18796 32044 18836
rect 32084 18796 32093 18836
rect 26668 18752 26708 18796
rect 12259 18712 12268 18752
rect 12308 18712 14956 18752
rect 14996 18712 15005 18752
rect 23299 18712 23308 18752
rect 23348 18712 24076 18752
rect 24116 18712 24125 18752
rect 26659 18712 26668 18752
rect 26708 18712 26717 18752
rect 33667 18712 33676 18752
rect 33716 18712 33725 18752
rect 34339 18712 34348 18752
rect 34388 18712 34540 18752
rect 34580 18712 34589 18752
rect 33676 18668 33716 18712
rect 11107 18628 11116 18668
rect 11156 18628 11980 18668
rect 12020 18628 12029 18668
rect 29539 18628 29548 18668
rect 29588 18628 29836 18668
rect 29876 18628 29885 18668
rect 33676 18628 37420 18668
rect 37460 18628 37469 18668
rect 35596 18584 35636 18628
rect 2563 18544 2572 18584
rect 2612 18544 2764 18584
rect 2804 18544 2956 18584
rect 2996 18544 3005 18584
rect 3811 18544 3820 18584
rect 3860 18544 4876 18584
rect 4916 18544 4925 18584
rect 10531 18544 10540 18584
rect 10580 18544 11596 18584
rect 11636 18544 11645 18584
rect 15043 18544 15052 18584
rect 15092 18544 15628 18584
rect 15668 18544 15677 18584
rect 20227 18544 20236 18584
rect 20276 18544 21004 18584
rect 21044 18544 21053 18584
rect 21187 18544 21196 18584
rect 21236 18544 21676 18584
rect 21716 18544 21725 18584
rect 22243 18544 22252 18584
rect 22292 18544 23308 18584
rect 23348 18544 23357 18584
rect 23491 18544 23500 18584
rect 23540 18544 23884 18584
rect 23924 18544 24076 18584
rect 24116 18544 24556 18584
rect 24596 18544 24605 18584
rect 25507 18544 25516 18584
rect 25556 18544 26668 18584
rect 26708 18544 26717 18584
rect 28387 18544 28396 18584
rect 28436 18544 29740 18584
rect 29780 18544 31084 18584
rect 31124 18544 31133 18584
rect 33859 18544 33868 18584
rect 33908 18544 35404 18584
rect 35444 18544 35453 18584
rect 35587 18544 35596 18584
rect 35636 18544 35645 18584
rect 36067 18544 36076 18584
rect 36116 18544 37804 18584
rect 37844 18544 37853 18584
rect 34243 18500 34301 18501
rect 8419 18460 8428 18500
rect 8468 18460 10444 18500
rect 10484 18460 10636 18500
rect 10676 18460 11116 18500
rect 11156 18460 11165 18500
rect 11320 18460 13996 18500
rect 14036 18460 14956 18500
rect 14996 18460 15005 18500
rect 21859 18460 21868 18500
rect 21908 18460 22348 18500
rect 22388 18460 22397 18500
rect 25795 18460 25804 18500
rect 25844 18460 26572 18500
rect 26612 18460 26621 18500
rect 34158 18460 34252 18500
rect 34292 18460 34301 18500
rect 11320 18416 11360 18460
rect 34243 18459 34301 18460
rect 11203 18376 11212 18416
rect 11252 18376 11360 18416
rect 12931 18376 12940 18416
rect 12980 18376 14188 18416
rect 14228 18376 14237 18416
rect 22627 18376 22636 18416
rect 22676 18376 25036 18416
rect 25076 18376 25708 18416
rect 25748 18376 31564 18416
rect 31604 18376 31756 18416
rect 31796 18376 31805 18416
rect 33571 18292 33580 18332
rect 33620 18292 34636 18332
rect 34676 18292 34685 18332
rect 34915 18292 34924 18332
rect 34964 18292 35687 18332
rect 35727 18292 35736 18332
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 34339 18208 34348 18248
rect 34388 18208 35020 18248
rect 35060 18208 37516 18248
rect 37556 18208 37900 18248
rect 37940 18208 37949 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 5923 18124 5932 18164
rect 5972 18124 6604 18164
rect 6644 18124 6653 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 23491 18124 23500 18164
rect 23540 18124 24172 18164
rect 24212 18124 24221 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 23779 18080 23837 18081
rect 23694 18040 23788 18080
rect 23828 18040 23837 18080
rect 23779 18039 23837 18040
rect 24067 17996 24125 17997
rect 11299 17956 11308 17996
rect 11348 17956 12268 17996
rect 12308 17956 12317 17996
rect 20131 17956 20140 17996
rect 20180 17956 21388 17996
rect 21428 17956 22348 17996
rect 22388 17956 22397 17996
rect 23683 17956 23692 17996
rect 23732 17956 24076 17996
rect 24116 17956 24125 17996
rect 24067 17955 24125 17956
rect 4675 17872 4684 17912
rect 4724 17872 6700 17912
rect 6740 17872 6749 17912
rect 21475 17872 21484 17912
rect 21524 17872 23980 17912
rect 24020 17872 24029 17912
rect 24172 17828 24212 18124
rect 32131 18040 32140 18080
rect 32180 18040 35500 18080
rect 35540 18040 37036 18080
rect 37076 18040 37324 18080
rect 37364 18040 37373 18080
rect 26083 17956 26092 17996
rect 26132 17956 27148 17996
rect 27188 17956 27197 17996
rect 29059 17956 29068 17996
rect 29108 17956 29356 17996
rect 29396 17956 29405 17996
rect 32035 17956 32044 17996
rect 32084 17956 33388 17996
rect 33428 17956 36076 17996
rect 36116 17956 36125 17996
rect 37123 17956 37132 17996
rect 37172 17956 37420 17996
rect 37460 17956 37469 17996
rect 25987 17872 25996 17912
rect 26036 17872 26284 17912
rect 26324 17872 26333 17912
rect 29155 17872 29164 17912
rect 29204 17872 32140 17912
rect 32180 17872 32189 17912
rect 34339 17872 34348 17912
rect 34388 17872 34540 17912
rect 34580 17872 35884 17912
rect 35924 17872 35933 17912
rect 37699 17872 37708 17912
rect 37748 17872 38764 17912
rect 38804 17872 38813 17912
rect 22243 17788 22252 17828
rect 22292 17788 22540 17828
rect 22580 17788 22589 17828
rect 23212 17788 23596 17828
rect 23636 17788 23645 17828
rect 24172 17788 24268 17828
rect 24308 17788 24317 17828
rect 31747 17788 31756 17828
rect 31796 17788 33196 17828
rect 33236 17788 35121 17828
rect 35161 17788 35170 17828
rect 37780 17788 39436 17828
rect 39476 17788 39485 17828
rect 23212 17744 23252 17788
rect 34435 17744 34493 17745
rect 37780 17744 37820 17788
rect 4387 17704 4396 17744
rect 4436 17704 4972 17744
rect 5012 17704 5164 17744
rect 5204 17704 5213 17744
rect 8707 17704 8716 17744
rect 8756 17704 10252 17744
rect 10292 17704 10301 17744
rect 12355 17704 12364 17744
rect 12404 17704 12556 17744
rect 12596 17704 12605 17744
rect 13795 17704 13804 17744
rect 13844 17704 14188 17744
rect 14228 17704 14237 17744
rect 17731 17704 17740 17744
rect 17780 17704 20812 17744
rect 20852 17704 20861 17744
rect 22435 17704 22444 17744
rect 22484 17704 22924 17744
rect 22964 17704 22973 17744
rect 23203 17704 23212 17744
rect 23252 17704 23261 17744
rect 23683 17704 23692 17744
rect 23732 17704 24556 17744
rect 24596 17704 24605 17744
rect 30595 17704 30604 17744
rect 30644 17704 30988 17744
rect 31028 17704 32332 17744
rect 32372 17704 32381 17744
rect 34435 17704 34444 17744
rect 34484 17704 34732 17744
rect 34772 17704 34781 17744
rect 36163 17704 36172 17744
rect 36212 17704 36556 17744
rect 36596 17704 36605 17744
rect 37219 17704 37228 17744
rect 37268 17704 37820 17744
rect 37987 17704 37996 17744
rect 38036 17704 38572 17744
rect 38612 17704 40012 17744
rect 40052 17704 41068 17744
rect 41108 17704 41117 17744
rect 34435 17703 34493 17704
rect 23107 17660 23165 17661
rect 26179 17660 26237 17661
rect 4003 17620 4012 17660
rect 4052 17620 5260 17660
rect 5300 17620 5309 17660
rect 11320 17620 12652 17660
rect 12692 17620 12701 17660
rect 13603 17620 13612 17660
rect 13652 17620 14092 17660
rect 14132 17620 14668 17660
rect 14708 17620 15916 17660
rect 15956 17620 15965 17660
rect 16771 17620 16780 17660
rect 16820 17620 18892 17660
rect 18932 17620 18941 17660
rect 23022 17620 23116 17660
rect 23156 17620 23165 17660
rect 23587 17620 23596 17660
rect 23636 17620 24364 17660
rect 24404 17620 24413 17660
rect 26094 17620 26188 17660
rect 26228 17620 26237 17660
rect 26755 17620 26764 17660
rect 26804 17620 33100 17660
rect 33140 17620 33149 17660
rect 34348 17620 34636 17660
rect 34676 17620 36268 17660
rect 36308 17620 36884 17660
rect 36931 17620 36940 17660
rect 36980 17620 37748 17660
rect 4195 17576 4253 17577
rect 11320 17576 11360 17620
rect 23107 17619 23165 17620
rect 26179 17619 26237 17620
rect 23779 17576 23837 17577
rect 34348 17576 34388 17620
rect 36844 17576 36884 17620
rect 37708 17576 37748 17620
rect 38572 17620 39916 17660
rect 39956 17620 39965 17660
rect 38572 17576 38612 17620
rect 3619 17536 3628 17576
rect 3668 17536 4204 17576
rect 4244 17536 4253 17576
rect 4579 17536 4588 17576
rect 4628 17536 5164 17576
rect 5204 17536 5213 17576
rect 8515 17536 8524 17576
rect 8564 17536 10348 17576
rect 10388 17536 11212 17576
rect 11252 17536 11360 17576
rect 23491 17536 23500 17576
rect 23540 17536 23788 17576
rect 23828 17536 23837 17576
rect 24067 17536 24076 17576
rect 24116 17536 25420 17576
rect 25460 17536 25469 17576
rect 25699 17536 25708 17576
rect 25748 17536 25900 17576
rect 25940 17536 26476 17576
rect 26516 17536 26525 17576
rect 27235 17536 27244 17576
rect 27284 17536 27628 17576
rect 27668 17536 27677 17576
rect 30211 17536 30220 17576
rect 30260 17536 34388 17576
rect 34435 17536 34444 17576
rect 34484 17536 34924 17576
rect 34964 17536 34973 17576
rect 36835 17536 36844 17576
rect 36884 17536 37516 17576
rect 37556 17536 37565 17576
rect 37699 17536 37708 17576
rect 37748 17536 37757 17576
rect 38563 17536 38572 17576
rect 38612 17536 38621 17576
rect 4195 17535 4253 17536
rect 23779 17535 23837 17536
rect 3907 17452 3916 17492
rect 3956 17452 5068 17492
rect 5108 17452 5356 17492
rect 5396 17452 5405 17492
rect 23107 17452 23116 17492
rect 23156 17452 23404 17492
rect 23444 17452 24460 17492
rect 24500 17452 24509 17492
rect 24643 17452 24652 17492
rect 24692 17452 24940 17492
rect 24980 17452 24989 17492
rect 26275 17452 26284 17492
rect 26324 17452 29260 17492
rect 29300 17452 32044 17492
rect 32084 17452 32236 17492
rect 32276 17452 32285 17492
rect 35112 17452 35121 17492
rect 35161 17452 35300 17492
rect 36643 17452 36652 17492
rect 36692 17452 37420 17492
rect 37460 17452 37469 17492
rect 0 17408 80 17428
rect 31756 17408 31796 17452
rect 35260 17408 35300 17452
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 25507 17368 25516 17408
rect 25556 17368 25900 17408
rect 25940 17368 29000 17408
rect 31747 17368 31756 17408
rect 31796 17368 31836 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 35260 17368 36308 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 28960 17324 29000 17368
rect 3811 17284 3820 17324
rect 3860 17284 3869 17324
rect 26659 17284 26668 17324
rect 26708 17284 27052 17324
rect 27092 17284 27724 17324
rect 27764 17284 27773 17324
rect 28960 17284 29260 17324
rect 29300 17284 30220 17324
rect 30260 17284 30269 17324
rect 35683 17284 35692 17324
rect 35732 17284 35884 17324
rect 35924 17284 35933 17324
rect 36268 17284 36308 17368
rect 36547 17324 36605 17325
rect 36348 17284 36357 17324
rect 36547 17284 36556 17324
rect 36596 17284 37228 17324
rect 37268 17284 37277 17324
rect 1507 17200 1516 17240
rect 1556 17200 3724 17240
rect 3764 17200 3773 17240
rect 3820 17156 3860 17284
rect 36547 17283 36605 17284
rect 24067 17240 24125 17241
rect 37315 17240 37373 17241
rect 4387 17200 4396 17240
rect 4436 17200 4876 17240
rect 4916 17200 4925 17240
rect 20803 17200 20812 17240
rect 20852 17200 21964 17240
rect 22004 17200 22013 17240
rect 23982 17200 24076 17240
rect 24116 17200 24125 17240
rect 27139 17200 27148 17240
rect 27188 17200 27916 17240
rect 27956 17200 27965 17240
rect 28766 17200 28775 17240
rect 28815 17200 32428 17240
rect 32468 17200 32477 17240
rect 34147 17200 34156 17240
rect 34196 17200 35116 17240
rect 35156 17200 36460 17240
rect 36500 17200 36509 17240
rect 37230 17200 37324 17240
rect 37364 17200 37373 17240
rect 24067 17199 24125 17200
rect 3523 17116 3532 17156
rect 3572 17116 4108 17156
rect 4148 17116 4157 17156
rect 17923 17116 17932 17156
rect 17972 17116 19372 17156
rect 19412 17116 19421 17156
rect 29068 17116 29452 17156
rect 29492 17116 29501 17156
rect 29068 17072 29108 17116
rect 3235 17032 3244 17072
rect 3284 17032 4204 17072
rect 4244 17032 4780 17072
rect 4820 17032 4829 17072
rect 6787 17032 6796 17072
rect 6836 17032 7852 17072
rect 7892 17032 7901 17072
rect 8131 17032 8140 17072
rect 8180 17032 9388 17072
rect 9428 17032 9437 17072
rect 16675 17032 16684 17072
rect 16724 17032 18988 17072
rect 19028 17032 19037 17072
rect 20707 17032 20716 17072
rect 20756 17032 20908 17072
rect 20948 17032 21868 17072
rect 21908 17032 21917 17072
rect 22627 17032 22636 17072
rect 22676 17032 23884 17072
rect 23924 17032 23933 17072
rect 25219 17032 25228 17072
rect 25268 17032 28775 17072
rect 28815 17032 28824 17072
rect 28963 17032 28972 17072
rect 29012 17032 29108 17072
rect 29155 17032 29164 17072
rect 29204 17032 30412 17072
rect 30452 17032 30461 17072
rect 3331 16948 3340 16988
rect 3380 16948 3820 16988
rect 3860 16948 3869 16988
rect 4675 16948 4684 16988
rect 4724 16948 5164 16988
rect 5204 16948 5213 16988
rect 15427 16948 15436 16988
rect 15476 16948 18316 16988
rect 18356 16948 18796 16988
rect 18836 16948 18845 16988
rect 23491 16948 23500 16988
rect 23540 16948 23980 16988
rect 24020 16948 24029 16988
rect 27235 16948 27244 16988
rect 27284 16948 29548 16988
rect 29588 16948 29597 16988
rect 32044 16904 32084 17200
rect 37315 17199 37373 17200
rect 35011 17116 35020 17156
rect 35060 17116 35308 17156
rect 35348 17116 35357 17156
rect 36299 17116 36308 17156
rect 36348 17116 37073 17156
rect 37113 17116 37122 17156
rect 32419 17032 32428 17072
rect 32468 17032 39628 17072
rect 39668 17032 40492 17072
rect 40532 17032 40541 17072
rect 36547 16948 36556 16988
rect 36596 16948 37324 16988
rect 37364 16948 37373 16988
rect 4291 16864 4300 16904
rect 4340 16864 4972 16904
rect 5012 16864 5021 16904
rect 14371 16864 14380 16904
rect 14420 16864 17548 16904
rect 17588 16864 17597 16904
rect 27619 16864 27628 16904
rect 27668 16864 27820 16904
rect 27860 16864 27869 16904
rect 31651 16864 31660 16904
rect 31700 16864 31709 16904
rect 32035 16864 32044 16904
rect 32084 16864 32093 16904
rect 37699 16864 37708 16904
rect 37748 16864 38188 16904
rect 38228 16864 38237 16904
rect 21571 16820 21629 16821
rect 31660 16820 31700 16864
rect 5155 16780 5164 16820
rect 5204 16780 5644 16820
rect 5684 16780 5693 16820
rect 6787 16780 6796 16820
rect 6836 16780 7948 16820
rect 7988 16780 8428 16820
rect 8468 16780 8477 16820
rect 12931 16780 12940 16820
rect 12980 16780 14572 16820
rect 14612 16780 14621 16820
rect 21571 16780 21580 16820
rect 21620 16780 21676 16820
rect 21716 16780 21725 16820
rect 26947 16780 26956 16820
rect 26996 16780 27148 16820
rect 27188 16780 27436 16820
rect 27476 16780 27485 16820
rect 28963 16780 28972 16820
rect 29012 16780 29260 16820
rect 29300 16780 29309 16820
rect 31660 16780 32620 16820
rect 32660 16780 33772 16820
rect 33812 16780 36556 16820
rect 36596 16780 36605 16820
rect 37603 16780 37612 16820
rect 37652 16780 38476 16820
rect 38516 16780 38525 16820
rect 21571 16779 21629 16780
rect 32035 16736 32093 16737
rect 24163 16696 24172 16736
rect 24212 16696 25612 16736
rect 25652 16696 25661 16736
rect 31939 16696 31948 16736
rect 31988 16696 32044 16736
rect 32084 16696 32093 16736
rect 32035 16695 32093 16696
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 25315 16612 25324 16652
rect 25364 16612 26572 16652
rect 26612 16612 27244 16652
rect 27284 16612 27293 16652
rect 28867 16612 28876 16652
rect 28916 16612 33236 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 36931 16612 36940 16652
rect 36980 16612 37420 16652
rect 37460 16612 37469 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 33196 16568 33236 16612
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 3619 16528 3628 16568
rect 3668 16528 6412 16568
rect 6452 16528 6461 16568
rect 24931 16528 24940 16568
rect 24980 16528 29452 16568
rect 29492 16528 31988 16568
rect 33196 16528 34348 16568
rect 34388 16528 34397 16568
rect 37507 16528 37516 16568
rect 37556 16528 40436 16568
rect 0 16508 80 16528
rect 18979 16484 19037 16485
rect 31555 16484 31613 16485
rect 31948 16484 31988 16528
rect 36547 16484 36605 16485
rect 4675 16444 4684 16484
rect 4724 16444 5684 16484
rect 5923 16444 5932 16484
rect 5972 16444 8428 16484
rect 8468 16444 8477 16484
rect 18979 16444 18988 16484
rect 19028 16444 20372 16484
rect 23971 16444 23980 16484
rect 24020 16444 25420 16484
rect 25460 16444 26380 16484
rect 26420 16444 26429 16484
rect 27811 16444 27820 16484
rect 27860 16444 28204 16484
rect 28244 16444 28253 16484
rect 30211 16444 30220 16484
rect 30260 16444 31564 16484
rect 31604 16444 31613 16484
rect 31939 16444 31948 16484
rect 31988 16444 34060 16484
rect 34100 16444 34109 16484
rect 35779 16444 35788 16484
rect 35828 16444 35980 16484
rect 36020 16444 36029 16484
rect 36462 16444 36556 16484
rect 36596 16444 36605 16484
rect 36739 16444 36748 16484
rect 36788 16444 37324 16484
rect 37364 16444 39572 16484
rect 5644 16400 5684 16444
rect 18979 16443 19037 16444
rect 20332 16400 20372 16444
rect 31555 16443 31613 16444
rect 36547 16443 36605 16444
rect 32419 16400 32477 16401
rect 39532 16400 39572 16444
rect 40396 16400 40436 16528
rect 2851 16360 2860 16400
rect 2900 16360 3340 16400
rect 3380 16360 3628 16400
rect 3668 16360 3677 16400
rect 4579 16360 4588 16400
rect 4628 16360 5452 16400
rect 5492 16360 5501 16400
rect 5635 16360 5644 16400
rect 5684 16360 6988 16400
rect 7028 16360 7037 16400
rect 11203 16360 11212 16400
rect 11252 16360 11732 16400
rect 15235 16360 15244 16400
rect 15284 16360 16492 16400
rect 16532 16360 16541 16400
rect 18883 16360 18892 16400
rect 18932 16360 19276 16400
rect 19316 16360 20140 16400
rect 20180 16360 20189 16400
rect 20323 16360 20332 16400
rect 20372 16360 20381 16400
rect 21763 16360 21772 16400
rect 21812 16360 21964 16400
rect 22004 16360 24748 16400
rect 24788 16360 24797 16400
rect 25603 16360 25612 16400
rect 25652 16360 26476 16400
rect 26516 16360 26525 16400
rect 27235 16360 27244 16400
rect 27284 16360 27436 16400
rect 27476 16360 27485 16400
rect 28099 16360 28108 16400
rect 28148 16360 29452 16400
rect 29492 16360 29501 16400
rect 31459 16360 31468 16400
rect 31508 16360 31756 16400
rect 31796 16360 31805 16400
rect 32419 16360 32428 16400
rect 32468 16360 36652 16400
rect 36692 16360 36701 16400
rect 37027 16360 37036 16400
rect 37076 16360 38380 16400
rect 38420 16360 38429 16400
rect 39532 16360 40340 16400
rect 40396 16360 40532 16400
rect 11692 16316 11732 16360
rect 32419 16359 32477 16360
rect 11683 16276 11692 16316
rect 11732 16276 11741 16316
rect 18979 16276 18988 16316
rect 19028 16276 20372 16316
rect 20515 16276 20524 16316
rect 20564 16276 21236 16316
rect 22435 16276 22444 16316
rect 22484 16276 23596 16316
rect 23636 16276 23645 16316
rect 23692 16276 26668 16316
rect 26708 16276 26717 16316
rect 27523 16276 27532 16316
rect 27572 16276 29932 16316
rect 29972 16276 29981 16316
rect 35404 16276 39820 16316
rect 39860 16276 39869 16316
rect 20131 16232 20189 16233
rect 20332 16232 20372 16276
rect 21196 16233 21236 16276
rect 21187 16232 21245 16233
rect 23692 16232 23732 16276
rect 24259 16232 24317 16233
rect 3043 16192 3052 16232
rect 3092 16192 4012 16232
rect 4052 16192 4061 16232
rect 5827 16192 5836 16232
rect 5876 16192 6412 16232
rect 6452 16192 6988 16232
rect 7028 16192 7037 16232
rect 7171 16192 7180 16232
rect 7220 16192 7852 16232
rect 7892 16192 7901 16232
rect 8515 16192 8524 16232
rect 8564 16192 8573 16232
rect 10915 16192 10924 16232
rect 10964 16192 12364 16232
rect 12404 16192 12413 16232
rect 12739 16192 12748 16232
rect 12788 16192 13228 16232
rect 13268 16192 13277 16232
rect 15715 16192 15724 16232
rect 15764 16192 16492 16232
rect 16532 16192 16541 16232
rect 16675 16192 16684 16232
rect 16724 16192 17548 16232
rect 17588 16192 17597 16232
rect 18691 16192 18700 16232
rect 18740 16192 19084 16232
rect 19124 16192 19660 16232
rect 19700 16192 19709 16232
rect 20131 16192 20140 16232
rect 20180 16192 20229 16232
rect 20269 16192 20278 16232
rect 20323 16192 20332 16232
rect 20372 16192 20716 16232
rect 20756 16192 20765 16232
rect 21102 16192 21196 16232
rect 21236 16192 21245 16232
rect 22339 16192 22348 16232
rect 22388 16192 22924 16232
rect 22964 16192 22973 16232
rect 23203 16192 23212 16232
rect 23252 16192 23692 16232
rect 23732 16192 23741 16232
rect 24174 16192 24268 16232
rect 24308 16192 25036 16232
rect 25076 16192 25085 16232
rect 27043 16192 27052 16232
rect 27092 16192 28012 16232
rect 28052 16192 28061 16232
rect 30115 16192 30124 16232
rect 30164 16192 30508 16232
rect 30548 16192 31852 16232
rect 31892 16192 31901 16232
rect 32323 16192 32332 16232
rect 32372 16192 33100 16232
rect 33140 16192 33149 16232
rect 8524 16148 8564 16192
rect 20131 16191 20189 16192
rect 21187 16191 21245 16192
rect 24259 16191 24317 16192
rect 3139 16108 3148 16148
rect 3188 16108 3628 16148
rect 3668 16108 3677 16148
rect 6499 16108 6508 16148
rect 6548 16108 7948 16148
rect 7988 16108 8564 16148
rect 19171 16108 19180 16148
rect 19220 16108 19372 16148
rect 19412 16108 19421 16148
rect 19843 16108 19852 16148
rect 19892 16108 20428 16148
rect 20468 16108 20477 16148
rect 22627 16108 22636 16148
rect 22676 16108 22828 16148
rect 22868 16108 24556 16148
rect 24596 16108 24605 16148
rect 27436 16064 27476 16192
rect 35404 16148 35444 16276
rect 40300 16232 40340 16360
rect 40492 16232 40532 16360
rect 36451 16192 36460 16232
rect 36500 16192 37820 16232
rect 38083 16192 38092 16232
rect 38132 16192 38572 16232
rect 38612 16192 38956 16232
rect 38996 16192 39005 16232
rect 40291 16192 40300 16232
rect 40340 16192 40349 16232
rect 40483 16192 40492 16232
rect 40532 16192 40541 16232
rect 29616 16108 29644 16148
rect 29684 16108 30892 16148
rect 30932 16108 30941 16148
rect 32995 16108 33004 16148
rect 33044 16108 35444 16148
rect 37315 16148 37373 16149
rect 37780 16148 37820 16192
rect 37315 16108 37324 16148
rect 37364 16108 37516 16148
rect 37556 16108 37565 16148
rect 37780 16108 40972 16148
rect 41012 16108 42316 16148
rect 42356 16108 42365 16148
rect 19939 16024 19948 16064
rect 19988 16024 20812 16064
rect 20852 16024 21580 16064
rect 21620 16024 21908 16064
rect 22531 16024 22540 16064
rect 22580 16024 26860 16064
rect 26900 16024 26909 16064
rect 27427 16024 27436 16064
rect 27476 16024 27485 16064
rect 28675 16024 28684 16064
rect 28724 16024 29068 16064
rect 29108 16024 29117 16064
rect 21868 15980 21908 16024
rect 26860 15980 26900 16024
rect 20131 15940 20140 15980
rect 20180 15940 21772 15980
rect 21812 15940 21821 15980
rect 21868 15940 23692 15980
rect 23732 15940 23741 15980
rect 24355 15940 24364 15980
rect 24404 15940 24748 15980
rect 24788 15940 25036 15980
rect 25076 15940 25085 15980
rect 26860 15940 27628 15980
rect 27668 15940 29260 15980
rect 29300 15940 29309 15980
rect 15427 15896 15485 15897
rect 24451 15896 24509 15897
rect 29740 15896 29780 16108
rect 37315 16107 37373 16108
rect 32419 16064 32477 16065
rect 37699 16064 37757 16065
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 4963 15856 4972 15896
rect 5012 15856 5548 15896
rect 5588 15856 5597 15896
rect 15331 15856 15340 15896
rect 15380 15856 15436 15896
rect 15476 15856 16780 15896
rect 16820 15856 16829 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 20611 15856 20620 15896
rect 20660 15856 21004 15896
rect 21044 15856 21053 15896
rect 24366 15856 24460 15896
rect 24500 15856 28780 15896
rect 28820 15856 28829 15896
rect 28876 15856 29780 15896
rect 29836 16024 32428 16064
rect 32468 16024 32477 16064
rect 32899 16024 32908 16064
rect 32948 16024 33292 16064
rect 33332 16024 33341 16064
rect 34627 16024 34636 16064
rect 34676 16024 34924 16064
rect 34964 16024 34973 16064
rect 35971 16024 35980 16064
rect 36020 16024 36268 16064
rect 36308 16024 36317 16064
rect 37123 16024 37132 16064
rect 37172 16024 37708 16064
rect 37748 16024 37996 16064
rect 38036 16024 39148 16064
rect 39188 16024 39197 16064
rect 40099 16024 40108 16064
rect 40148 16024 41260 16064
rect 41300 16024 41309 16064
rect 15427 15855 15485 15856
rect 24451 15855 24509 15856
rect 20227 15812 20285 15813
rect 28876 15812 28916 15856
rect 29836 15812 29876 16024
rect 32419 16023 32477 16024
rect 34636 15980 34676 16024
rect 37699 16023 37757 16024
rect 29923 15940 29932 15980
rect 29972 15940 34252 15980
rect 34292 15940 34676 15980
rect 38179 15940 38188 15980
rect 38228 15940 38380 15980
rect 38420 15940 39244 15980
rect 39284 15940 39293 15980
rect 31651 15856 31660 15896
rect 31700 15856 31852 15896
rect 31892 15856 31901 15896
rect 32707 15856 32716 15896
rect 32756 15856 33004 15896
rect 33044 15856 33053 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 36547 15856 36556 15896
rect 36596 15856 37324 15896
rect 37364 15856 37373 15896
rect 37795 15856 37804 15896
rect 37844 15856 38668 15896
rect 38708 15856 38717 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 835 15772 844 15812
rect 884 15772 7316 15812
rect 7843 15772 7852 15812
rect 7892 15772 9140 15812
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 0 15668 80 15688
rect 7276 15644 7316 15772
rect 7651 15688 7660 15728
rect 7700 15688 8236 15728
rect 8276 15688 8620 15728
rect 8660 15688 8669 15728
rect 9100 15644 9140 15772
rect 20140 15772 20236 15812
rect 20276 15772 21292 15812
rect 21332 15772 22828 15812
rect 22868 15772 22877 15812
rect 22924 15772 24172 15812
rect 24212 15772 24221 15812
rect 27235 15772 27244 15812
rect 27284 15772 28916 15812
rect 28960 15772 29876 15812
rect 30595 15772 30604 15812
rect 30644 15772 31564 15812
rect 31604 15772 31613 15812
rect 34435 15772 34444 15812
rect 34484 15772 35020 15812
rect 35060 15772 35596 15812
rect 35636 15772 35884 15812
rect 35924 15772 36364 15812
rect 36404 15772 36980 15812
rect 20140 15728 20180 15772
rect 20227 15771 20285 15772
rect 21667 15728 21725 15729
rect 22924 15728 22964 15772
rect 28960 15728 29000 15772
rect 36940 15728 36980 15772
rect 10531 15688 10540 15728
rect 10580 15688 10589 15728
rect 18499 15688 18508 15728
rect 18548 15688 19372 15728
rect 19412 15688 20180 15728
rect 20227 15688 20236 15728
rect 20276 15688 20285 15728
rect 21475 15688 21484 15728
rect 21524 15688 21533 15728
rect 21648 15688 21676 15728
rect 21716 15688 21772 15728
rect 21812 15688 22964 15728
rect 23011 15688 23020 15728
rect 23060 15688 24844 15728
rect 24884 15688 24893 15728
rect 26659 15688 26668 15728
rect 26708 15688 29000 15728
rect 29923 15688 29932 15728
rect 29972 15688 30508 15728
rect 30548 15688 31372 15728
rect 31412 15688 31421 15728
rect 34339 15688 34348 15728
rect 34388 15688 34828 15728
rect 34868 15688 34877 15728
rect 36067 15688 36076 15728
rect 36116 15688 36844 15728
rect 36884 15688 36893 15728
rect 36940 15688 38092 15728
rect 38132 15688 38141 15728
rect 10540 15644 10580 15688
rect 3235 15604 3244 15644
rect 3284 15604 3628 15644
rect 3668 15604 4052 15644
rect 4387 15604 4396 15644
rect 4436 15604 6124 15644
rect 6164 15604 6173 15644
rect 7276 15604 7852 15644
rect 7892 15604 8140 15644
rect 8180 15604 8189 15644
rect 9100 15604 10580 15644
rect 4012 15560 4052 15604
rect 9100 15560 9140 15604
rect 931 15520 940 15560
rect 980 15520 3532 15560
rect 3572 15520 3581 15560
rect 4003 15520 4012 15560
rect 4052 15520 4492 15560
rect 4532 15520 4972 15560
rect 5012 15520 5021 15560
rect 5347 15520 5356 15560
rect 5396 15520 6316 15560
rect 6356 15520 6365 15560
rect 8323 15520 8332 15560
rect 8372 15520 8716 15560
rect 8756 15520 8765 15560
rect 9091 15520 9100 15560
rect 9140 15520 9149 15560
rect 9667 15520 9676 15560
rect 9716 15520 10156 15560
rect 10196 15520 10205 15560
rect 16003 15520 16012 15560
rect 16052 15520 16684 15560
rect 16724 15520 16733 15560
rect 18691 15520 18700 15560
rect 18740 15520 19180 15560
rect 19220 15520 19564 15560
rect 19604 15520 20140 15560
rect 20180 15520 20189 15560
rect 20236 15476 20276 15688
rect 21484 15644 21524 15688
rect 21667 15687 21725 15688
rect 31555 15644 31613 15645
rect 37123 15644 37181 15645
rect 21484 15604 22732 15644
rect 22772 15604 25132 15644
rect 25172 15604 25181 15644
rect 27715 15604 27724 15644
rect 27764 15604 28108 15644
rect 28148 15604 28157 15644
rect 28960 15604 30700 15644
rect 30740 15604 30749 15644
rect 31470 15604 31564 15644
rect 31604 15604 32908 15644
rect 32948 15604 32957 15644
rect 33667 15604 33676 15644
rect 33716 15604 34060 15644
rect 34100 15604 35596 15644
rect 35636 15604 36172 15644
rect 36212 15604 36884 15644
rect 36931 15604 36940 15644
rect 36980 15604 37132 15644
rect 37172 15604 37181 15644
rect 37315 15604 37324 15644
rect 37364 15604 37373 15644
rect 37780 15604 38188 15644
rect 38228 15604 40108 15644
rect 40148 15604 40157 15644
rect 27715 15560 27773 15561
rect 28960 15560 29000 15604
rect 31555 15603 31613 15604
rect 20611 15520 20620 15560
rect 20660 15520 21484 15560
rect 21524 15520 21964 15560
rect 22004 15520 22013 15560
rect 22531 15520 22540 15560
rect 22580 15520 22924 15560
rect 22964 15520 22973 15560
rect 24931 15520 24940 15560
rect 24980 15520 25324 15560
rect 25364 15520 25373 15560
rect 25420 15520 27244 15560
rect 27284 15520 27293 15560
rect 27715 15520 27724 15560
rect 27764 15520 28012 15560
rect 28052 15520 28061 15560
rect 28195 15520 28204 15560
rect 28244 15520 29000 15560
rect 32040 15520 32049 15560
rect 32089 15520 32423 15560
rect 32463 15520 32472 15560
rect 33763 15520 33772 15560
rect 33812 15520 34924 15560
rect 34964 15520 34973 15560
rect 35683 15520 35692 15560
rect 35732 15520 36556 15560
rect 36596 15520 36605 15560
rect 36739 15520 36748 15560
rect 36788 15520 36797 15560
rect 25420 15476 25460 15520
rect 27715 15519 27773 15520
rect 36748 15476 36788 15520
rect 6595 15436 6604 15476
rect 6644 15436 6653 15476
rect 7939 15436 7948 15476
rect 7988 15436 8524 15476
rect 8564 15436 8573 15476
rect 15811 15436 15820 15476
rect 15860 15436 16300 15476
rect 16340 15436 16349 15476
rect 19363 15436 19372 15476
rect 19412 15436 20716 15476
rect 20756 15436 20765 15476
rect 22243 15436 22252 15476
rect 22292 15436 23308 15476
rect 23348 15436 23357 15476
rect 24451 15436 24460 15476
rect 24500 15436 24748 15476
rect 24788 15436 25460 15476
rect 25699 15436 25708 15476
rect 25748 15436 25900 15476
rect 25940 15436 25949 15476
rect 28771 15436 28780 15476
rect 28820 15436 32468 15476
rect 34627 15436 34636 15476
rect 34676 15436 35404 15476
rect 35444 15436 36788 15476
rect 6604 15392 6644 15436
rect 4579 15352 4588 15392
rect 4628 15352 6644 15392
rect 18787 15352 18796 15392
rect 18836 15352 19660 15392
rect 19700 15352 19709 15392
rect 3331 15268 3340 15308
rect 3380 15268 4436 15308
rect 4396 15140 4436 15268
rect 6604 15224 6644 15352
rect 22252 15308 22292 15436
rect 32035 15392 32093 15393
rect 22435 15352 22444 15392
rect 22484 15352 24172 15392
rect 24212 15352 25612 15392
rect 25652 15352 25661 15392
rect 31939 15352 31948 15392
rect 31988 15352 32044 15392
rect 32084 15352 32093 15392
rect 32035 15351 32093 15352
rect 16963 15268 16972 15308
rect 17012 15268 17836 15308
rect 17876 15268 17885 15308
rect 20227 15268 20236 15308
rect 20276 15268 22292 15308
rect 31555 15268 31564 15308
rect 31604 15268 31852 15308
rect 31892 15268 31901 15308
rect 32428 15224 32468 15436
rect 36844 15392 36884 15604
rect 37123 15603 37181 15604
rect 37324 15560 37364 15604
rect 37780 15560 37820 15604
rect 37324 15520 37820 15560
rect 37891 15520 37900 15560
rect 37940 15520 38668 15560
rect 38708 15520 38717 15560
rect 37699 15476 37757 15477
rect 36931 15436 36940 15476
rect 36980 15436 37556 15476
rect 37614 15436 37708 15476
rect 37748 15436 37757 15476
rect 37516 15392 37556 15436
rect 37699 15435 37757 15436
rect 35587 15352 35596 15392
rect 35636 15352 36268 15392
rect 36308 15352 36317 15392
rect 36835 15352 36844 15392
rect 36884 15352 36893 15392
rect 37027 15352 37036 15392
rect 37076 15352 37085 15392
rect 37516 15352 37612 15392
rect 37652 15352 37661 15392
rect 32515 15308 32573 15309
rect 37036 15308 37076 15352
rect 32515 15268 32524 15308
rect 32564 15268 36500 15308
rect 36547 15268 36556 15308
rect 36596 15268 36605 15308
rect 37036 15268 38380 15308
rect 38420 15268 38429 15308
rect 32515 15267 32573 15268
rect 4675 15184 4684 15224
rect 4724 15184 5396 15224
rect 5539 15184 5548 15224
rect 5588 15184 6028 15224
rect 6068 15184 6077 15224
rect 6604 15184 6796 15224
rect 6836 15184 6845 15224
rect 16771 15184 16780 15224
rect 16820 15184 18700 15224
rect 18740 15184 18749 15224
rect 23779 15184 23788 15224
rect 23828 15184 26572 15224
rect 26612 15184 28108 15224
rect 28148 15184 30604 15224
rect 30644 15184 30653 15224
rect 32419 15184 32428 15224
rect 32468 15184 33004 15224
rect 33044 15184 33053 15224
rect 33100 15184 34348 15224
rect 34388 15184 36364 15224
rect 36404 15184 36413 15224
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 4387 15100 4396 15140
rect 4436 15100 4876 15140
rect 4916 15100 4925 15140
rect 5356 15056 5396 15184
rect 20803 15140 20861 15141
rect 24259 15140 24317 15141
rect 25699 15140 25757 15141
rect 33100 15140 33140 15184
rect 5443 15100 5452 15140
rect 5492 15100 6412 15140
rect 6452 15100 6892 15140
rect 6932 15100 6941 15140
rect 14179 15100 14188 15140
rect 14228 15100 16396 15140
rect 16436 15100 16445 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 20227 15100 20236 15140
rect 20276 15100 20285 15140
rect 20718 15100 20812 15140
rect 20852 15100 20861 15140
rect 24174 15100 24268 15140
rect 24308 15100 25708 15140
rect 25748 15100 25757 15140
rect 29539 15100 29548 15140
rect 29588 15100 33100 15140
rect 33140 15100 33149 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 36067 15100 36076 15140
rect 36116 15100 36268 15140
rect 36308 15100 36317 15140
rect 5923 15056 5981 15057
rect 17635 15056 17693 15057
rect 20131 15056 20189 15057
rect 5356 15016 5932 15056
rect 5972 15016 7084 15056
rect 7124 15016 8044 15056
rect 8084 15016 8093 15056
rect 17550 15016 17644 15056
rect 17684 15016 20140 15056
rect 20180 15016 20189 15056
rect 5923 15015 5981 15016
rect 17635 15015 17693 15016
rect 20131 15015 20189 15016
rect 18787 14972 18845 14973
rect 20236 14972 20276 15100
rect 20803 15099 20861 15100
rect 24259 15099 24317 15100
rect 25699 15099 25757 15100
rect 27715 15056 27773 15057
rect 36460 15056 36500 15268
rect 36556 15224 36596 15268
rect 36556 15184 37516 15224
rect 37556 15184 37565 15224
rect 37780 15184 37900 15224
rect 37940 15184 38900 15224
rect 39139 15184 39148 15224
rect 39188 15184 39820 15224
rect 39860 15184 39869 15224
rect 37780 15140 37820 15184
rect 38860 15140 38900 15184
rect 36940 15100 37820 15140
rect 38083 15100 38092 15140
rect 38132 15100 38668 15140
rect 38708 15100 38717 15140
rect 38851 15100 38860 15140
rect 38900 15100 39532 15140
rect 39572 15100 39581 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 36940 15056 36980 15100
rect 25603 15016 25612 15056
rect 25652 15016 26284 15056
rect 26324 15016 27724 15056
rect 27764 15016 27773 15056
rect 32227 15016 32236 15056
rect 32276 15016 32285 15056
rect 36460 15016 36980 15056
rect 27715 15015 27773 15016
rect 31939 14972 31997 14973
rect 4675 14932 4684 14972
rect 4724 14932 4972 14972
rect 5012 14932 7948 14972
rect 7988 14932 7997 14972
rect 9091 14932 9100 14972
rect 9140 14932 9964 14972
rect 10004 14932 10013 14972
rect 18787 14932 18796 14972
rect 18836 14932 20276 14972
rect 23971 14932 23980 14972
rect 24020 14932 24748 14972
rect 24788 14932 31948 14972
rect 31988 14932 31997 14972
rect 18787 14931 18845 14932
rect 31939 14931 31997 14932
rect 0 14888 80 14908
rect 19939 14888 19997 14889
rect 32236 14888 32276 15016
rect 37123 14972 37181 14973
rect 37038 14932 37132 14972
rect 37172 14932 37181 14972
rect 40483 14932 40492 14972
rect 40532 14932 41548 14972
rect 41588 14932 41597 14972
rect 37123 14931 37181 14932
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 2947 14848 2956 14888
rect 2996 14848 3436 14888
rect 3476 14848 5932 14888
rect 5972 14848 5981 14888
rect 6211 14848 6220 14888
rect 6260 14848 6604 14888
rect 6644 14848 6653 14888
rect 8803 14848 8812 14888
rect 8852 14848 9140 14888
rect 15043 14848 15052 14888
rect 15092 14848 17932 14888
rect 17972 14848 17981 14888
rect 18883 14848 18892 14888
rect 18932 14848 19948 14888
rect 19988 14848 22060 14888
rect 22100 14848 22109 14888
rect 31459 14848 31468 14888
rect 31508 14848 32276 14888
rect 0 14828 80 14848
rect 9100 14720 9140 14848
rect 19939 14847 19997 14848
rect 20227 14804 20285 14805
rect 20227 14764 20236 14804
rect 20276 14764 20370 14804
rect 25891 14764 25900 14804
rect 25940 14764 26380 14804
rect 26420 14764 26860 14804
rect 26900 14764 28300 14804
rect 28340 14764 29740 14804
rect 29780 14764 29789 14804
rect 31651 14764 31660 14804
rect 31700 14764 32812 14804
rect 32852 14764 32861 14804
rect 32995 14764 33004 14804
rect 33044 14764 34444 14804
rect 34484 14764 34493 14804
rect 20227 14763 20285 14764
rect 2851 14680 2860 14720
rect 2900 14680 3244 14720
rect 3284 14680 3293 14720
rect 3523 14680 3532 14720
rect 3572 14680 4300 14720
rect 4340 14680 4780 14720
rect 4820 14680 4829 14720
rect 9091 14680 9100 14720
rect 9140 14680 9149 14720
rect 15139 14680 15148 14720
rect 15188 14680 15916 14720
rect 15956 14680 16876 14720
rect 16916 14680 16925 14720
rect 17251 14680 17260 14720
rect 17300 14680 18316 14720
rect 18356 14680 18365 14720
rect 19843 14680 19852 14720
rect 19892 14680 21868 14720
rect 21908 14680 21917 14720
rect 28579 14680 28588 14720
rect 28628 14680 29000 14720
rect 29827 14680 29836 14720
rect 29876 14680 30028 14720
rect 30068 14680 30077 14720
rect 31363 14680 31372 14720
rect 31412 14680 32140 14720
rect 32180 14680 32189 14720
rect 32515 14680 32524 14720
rect 32564 14680 33868 14720
rect 33908 14680 34156 14720
rect 34196 14680 34205 14720
rect 37315 14680 37324 14720
rect 37364 14680 37612 14720
rect 37652 14680 37661 14720
rect 38179 14680 38188 14720
rect 38228 14680 40396 14720
rect 40436 14680 40445 14720
rect 21667 14636 21725 14637
rect 28960 14636 29000 14680
rect 4012 14596 5452 14636
rect 5492 14596 5501 14636
rect 21582 14596 21676 14636
rect 21716 14596 21725 14636
rect 23011 14596 23020 14636
rect 23060 14596 25900 14636
rect 25940 14596 25949 14636
rect 28960 14596 29452 14636
rect 29492 14596 29501 14636
rect 29635 14596 29644 14636
rect 29684 14596 30316 14636
rect 30356 14596 30365 14636
rect 4012 14552 4052 14596
rect 21667 14595 21725 14596
rect 32035 14552 32093 14553
rect 32611 14552 32669 14553
rect 3715 14512 3724 14552
rect 3764 14512 4012 14552
rect 4052 14512 4061 14552
rect 5155 14512 5164 14552
rect 5204 14512 8140 14552
rect 8180 14512 8189 14552
rect 15331 14512 15340 14552
rect 15380 14512 16972 14552
rect 17012 14512 17356 14552
rect 17396 14512 18412 14552
rect 18452 14512 18461 14552
rect 19651 14512 19660 14552
rect 19700 14512 19709 14552
rect 20515 14512 20524 14552
rect 20564 14512 21580 14552
rect 21620 14512 21629 14552
rect 26083 14512 26092 14552
rect 26132 14512 26668 14552
rect 26708 14512 31564 14552
rect 31604 14512 31613 14552
rect 32035 14512 32044 14552
rect 32084 14512 32620 14552
rect 32660 14512 36268 14552
rect 36308 14512 36844 14552
rect 36884 14512 36893 14552
rect 19660 14468 19700 14512
rect 32035 14511 32093 14512
rect 32611 14511 32669 14512
rect 19660 14428 20620 14468
rect 20660 14428 20669 14468
rect 32611 14428 32620 14468
rect 32660 14428 32812 14468
rect 32852 14428 32861 14468
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 20131 14344 20140 14384
rect 20180 14344 20189 14384
rect 27907 14344 27916 14384
rect 27956 14344 28204 14384
rect 28244 14344 29260 14384
rect 29300 14344 29309 14384
rect 32035 14344 32044 14384
rect 32084 14344 33292 14384
rect 33332 14344 33341 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 17827 14260 17836 14300
rect 17876 14260 18508 14300
rect 18548 14260 18557 14300
rect 18787 14216 18845 14217
rect 20035 14216 20093 14217
rect 7555 14176 7564 14216
rect 7604 14176 8716 14216
rect 8756 14176 8765 14216
rect 13411 14176 13420 14216
rect 13460 14176 13900 14216
rect 13940 14176 15628 14216
rect 15668 14176 18796 14216
rect 18836 14176 18845 14216
rect 19939 14176 19948 14216
rect 19988 14176 20044 14216
rect 20084 14176 20093 14216
rect 18787 14175 18845 14176
rect 20035 14175 20093 14176
rect 19171 14132 19229 14133
rect 20140 14132 20180 14344
rect 27235 14260 27244 14300
rect 27284 14260 28492 14300
rect 28532 14260 28541 14300
rect 29923 14216 29981 14217
rect 21667 14176 21676 14216
rect 21716 14176 22252 14216
rect 22292 14176 22301 14216
rect 27043 14176 27052 14216
rect 27092 14176 27101 14216
rect 28579 14176 28588 14216
rect 28628 14176 29644 14216
rect 29684 14176 29693 14216
rect 29838 14176 29932 14216
rect 29972 14176 29981 14216
rect 32899 14176 32908 14216
rect 32948 14176 33676 14216
rect 33716 14176 34636 14216
rect 34676 14176 34685 14216
rect 26179 14132 26237 14133
rect 1027 14092 1036 14132
rect 1076 14092 3148 14132
rect 3188 14092 3197 14132
rect 9571 14092 9580 14132
rect 9620 14092 13036 14132
rect 13076 14092 13085 14132
rect 13507 14092 13516 14132
rect 13556 14092 13804 14132
rect 13844 14092 15764 14132
rect 16867 14092 16876 14132
rect 16916 14092 17740 14132
rect 17780 14092 18988 14132
rect 19028 14092 19037 14132
rect 19171 14092 19180 14132
rect 19220 14092 21292 14132
rect 21332 14092 23212 14132
rect 23252 14092 23261 14132
rect 26094 14092 26188 14132
rect 26228 14092 26237 14132
rect 0 14048 80 14068
rect 14947 14048 15005 14049
rect 15724 14048 15764 14092
rect 18988 14048 19028 14092
rect 19171 14091 19229 14092
rect 26179 14091 26237 14092
rect 27052 14048 27092 14176
rect 29923 14175 29981 14176
rect 28387 14092 28396 14132
rect 28436 14092 28972 14132
rect 29012 14092 29021 14132
rect 29347 14092 29356 14132
rect 29396 14092 32332 14132
rect 32372 14092 32381 14132
rect 31939 14048 31997 14049
rect 0 14008 940 14048
rect 980 14008 989 14048
rect 10531 14008 10540 14048
rect 10580 14008 10828 14048
rect 10868 14008 11212 14048
rect 11252 14008 11788 14048
rect 11828 14008 11837 14048
rect 13315 14008 13324 14048
rect 13364 14008 14764 14048
rect 14804 14008 14813 14048
rect 14947 14008 14956 14048
rect 14996 14008 15090 14048
rect 15715 14008 15724 14048
rect 15764 14008 16108 14048
rect 16148 14008 16157 14048
rect 17059 14008 17068 14048
rect 17108 14008 17260 14048
rect 17300 14008 17309 14048
rect 18883 14008 18892 14048
rect 18932 14008 18941 14048
rect 18988 14008 19468 14048
rect 19508 14008 20428 14048
rect 20468 14008 20812 14048
rect 20852 14008 20861 14048
rect 22147 14008 22156 14048
rect 22196 14008 23020 14048
rect 23060 14008 23069 14048
rect 25507 14008 25516 14048
rect 25556 14008 26284 14048
rect 26324 14008 26333 14048
rect 27052 14008 29740 14048
rect 29780 14008 29789 14048
rect 31854 14008 31948 14048
rect 31988 14008 31997 14048
rect 34339 14008 34348 14048
rect 34388 14008 36076 14048
rect 36116 14008 36125 14048
rect 37795 14008 37804 14048
rect 37844 14008 39820 14048
rect 39860 14008 39869 14048
rect 0 13988 80 14008
rect 14947 14007 15005 14008
rect 15235 13964 15293 13965
rect 18892 13964 18932 14008
rect 31939 14007 31997 14008
rect 19939 13964 19997 13965
rect 28195 13964 28253 13965
rect 14188 13924 14380 13964
rect 14420 13924 14429 13964
rect 15150 13924 15244 13964
rect 15284 13924 15293 13964
rect 15523 13924 15532 13964
rect 15572 13924 18740 13964
rect 18892 13924 19564 13964
rect 19604 13924 19613 13964
rect 19854 13924 19948 13964
rect 19988 13924 19997 13964
rect 20899 13924 20908 13964
rect 20948 13924 21772 13964
rect 21812 13924 25132 13964
rect 25172 13924 25181 13964
rect 26179 13924 26188 13964
rect 26228 13924 28204 13964
rect 28244 13924 28253 13964
rect 28867 13924 28876 13964
rect 28916 13924 30220 13964
rect 30260 13924 30269 13964
rect 38755 13924 38764 13964
rect 38804 13924 39244 13964
rect 39284 13924 39293 13964
rect 14188 13880 14228 13924
rect 15235 13923 15293 13924
rect 3523 13840 3532 13880
rect 3572 13840 3916 13880
rect 3956 13840 3965 13880
rect 5827 13840 5836 13880
rect 5876 13840 6028 13880
rect 6068 13840 6077 13880
rect 11587 13840 11596 13880
rect 11636 13840 11980 13880
rect 12020 13840 12844 13880
rect 12884 13840 12893 13880
rect 13795 13840 13804 13880
rect 13844 13840 14228 13880
rect 14275 13840 14284 13880
rect 14324 13840 15052 13880
rect 15092 13840 15101 13880
rect 15811 13840 15820 13880
rect 15860 13840 16396 13880
rect 16436 13840 16445 13880
rect 18700 13796 18740 13924
rect 19939 13923 19997 13924
rect 28195 13923 28253 13924
rect 19948 13880 19988 13923
rect 18787 13840 18796 13880
rect 18836 13840 19988 13880
rect 20035 13880 20093 13881
rect 20035 13840 20044 13880
rect 20084 13840 20428 13880
rect 20468 13840 20477 13880
rect 25699 13840 25708 13880
rect 25748 13840 27148 13880
rect 27188 13840 27197 13880
rect 28771 13840 28780 13880
rect 28820 13840 28972 13880
rect 29012 13840 29836 13880
rect 29876 13840 29885 13880
rect 31459 13840 31468 13880
rect 31508 13840 32140 13880
rect 32180 13840 32189 13880
rect 33475 13840 33484 13880
rect 33524 13840 34156 13880
rect 34196 13840 34205 13880
rect 20035 13839 20093 13840
rect 28963 13796 29021 13797
rect 13891 13756 13900 13796
rect 13940 13756 14572 13796
rect 14612 13756 14860 13796
rect 14900 13756 16300 13796
rect 16340 13756 16349 13796
rect 18700 13756 18988 13796
rect 19028 13756 19037 13796
rect 28963 13756 28972 13796
rect 29012 13756 29164 13796
rect 29204 13756 30796 13796
rect 30836 13756 30845 13796
rect 36739 13756 36748 13796
rect 36788 13756 38092 13796
rect 38132 13756 38141 13796
rect 28963 13755 29021 13756
rect 28291 13672 28300 13712
rect 28340 13672 30412 13712
rect 30452 13672 30461 13712
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 13987 13588 13996 13628
rect 14036 13588 14764 13628
rect 14804 13588 14813 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 26467 13588 26476 13628
rect 26516 13588 28588 13628
rect 28628 13588 29068 13628
rect 29108 13588 29117 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 18019 13544 18077 13545
rect 26755 13544 26813 13545
rect 13027 13504 13036 13544
rect 13076 13504 14092 13544
rect 14132 13504 14476 13544
rect 14516 13504 14525 13544
rect 17923 13504 17932 13544
rect 17972 13504 18028 13544
rect 18068 13504 18077 13544
rect 19075 13504 19084 13544
rect 19124 13504 19660 13544
rect 19700 13504 19709 13544
rect 26670 13504 26764 13544
rect 26804 13504 26813 13544
rect 18019 13503 18077 13504
rect 26755 13503 26813 13504
rect 21571 13460 21629 13461
rect 6499 13420 6508 13460
rect 6548 13420 6892 13460
rect 6932 13420 7276 13460
rect 7316 13420 7325 13460
rect 16291 13420 16300 13460
rect 16340 13420 17068 13460
rect 17108 13420 17117 13460
rect 17164 13420 20180 13460
rect 15331 13376 15389 13377
rect 17164 13376 17204 13420
rect 19171 13376 19229 13377
rect 15331 13336 15340 13376
rect 15380 13336 15436 13376
rect 15476 13336 15916 13376
rect 15956 13336 17204 13376
rect 17260 13336 19180 13376
rect 19220 13336 19229 13376
rect 20140 13376 20180 13420
rect 21571 13420 21580 13460
rect 21654 13420 21715 13460
rect 21859 13420 21868 13460
rect 21908 13420 22060 13460
rect 22100 13420 22109 13460
rect 27523 13420 27532 13460
rect 27572 13420 29260 13460
rect 29300 13420 29309 13460
rect 21571 13419 21629 13420
rect 28003 13376 28061 13377
rect 20140 13336 26476 13376
rect 26516 13336 26525 13376
rect 28003 13336 28012 13376
rect 28052 13336 28204 13376
rect 28244 13336 28253 13376
rect 28675 13336 28684 13376
rect 28724 13336 30220 13376
rect 30260 13336 30269 13376
rect 31555 13336 31564 13376
rect 31604 13336 32236 13376
rect 32276 13336 32285 13376
rect 32803 13336 32812 13376
rect 32852 13336 39340 13376
rect 39380 13336 39389 13376
rect 15331 13335 15389 13336
rect 17260 13292 17300 13336
rect 19171 13335 19229 13336
rect 28003 13335 28061 13336
rect 20035 13292 20093 13293
rect 8419 13252 8428 13292
rect 8468 13252 11212 13292
rect 11252 13252 11261 13292
rect 12259 13252 12268 13292
rect 12308 13252 14188 13292
rect 14228 13252 14668 13292
rect 14708 13252 14717 13292
rect 15244 13252 17300 13292
rect 17539 13252 17548 13292
rect 17588 13252 19276 13292
rect 19316 13252 19325 13292
rect 19555 13252 19564 13292
rect 19604 13252 20044 13292
rect 20084 13252 21484 13292
rect 21524 13252 22060 13292
rect 22100 13252 22109 13292
rect 24835 13252 24844 13292
rect 24884 13252 25708 13292
rect 25748 13252 26092 13292
rect 26132 13252 26764 13292
rect 26804 13252 29876 13292
rect 30787 13252 30796 13292
rect 30836 13252 33100 13292
rect 33140 13252 35212 13292
rect 35252 13252 35261 13292
rect 0 13208 80 13228
rect 15244 13208 15284 13252
rect 17260 13208 17300 13252
rect 20035 13251 20093 13252
rect 17731 13208 17789 13209
rect 18019 13208 18077 13209
rect 28003 13208 28061 13209
rect 29836 13208 29876 13252
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 2275 13168 2284 13208
rect 2324 13168 4492 13208
rect 4532 13168 5836 13208
rect 5876 13168 5885 13208
rect 6787 13168 6796 13208
rect 6836 13168 8812 13208
rect 8852 13168 8861 13208
rect 13315 13168 13324 13208
rect 13364 13168 14380 13208
rect 14420 13168 14429 13208
rect 15235 13168 15244 13208
rect 15284 13168 15293 13208
rect 15523 13168 15532 13208
rect 15572 13168 16300 13208
rect 16340 13168 16349 13208
rect 17251 13168 17260 13208
rect 17300 13168 17309 13208
rect 17646 13168 17740 13208
rect 17780 13168 17789 13208
rect 17934 13168 18028 13208
rect 18068 13168 18316 13208
rect 18356 13168 18365 13208
rect 18595 13168 18604 13208
rect 18644 13168 19084 13208
rect 19124 13168 19133 13208
rect 19747 13168 19756 13208
rect 19796 13168 20140 13208
rect 20180 13168 20189 13208
rect 20323 13168 20332 13208
rect 20372 13168 20524 13208
rect 20564 13168 21100 13208
rect 21140 13168 21149 13208
rect 22435 13168 22444 13208
rect 22484 13168 22493 13208
rect 25411 13168 25420 13208
rect 25460 13168 25469 13208
rect 27918 13168 28012 13208
rect 28052 13168 28061 13208
rect 29827 13168 29836 13208
rect 29876 13168 29885 13208
rect 30019 13168 30028 13208
rect 30068 13168 30108 13208
rect 32995 13168 33004 13208
rect 33044 13168 33292 13208
rect 33332 13168 34444 13208
rect 34484 13168 34493 13208
rect 0 13148 80 13168
rect 17731 13167 17789 13168
rect 18019 13167 18077 13168
rect 22444 13124 22484 13168
rect 13123 13084 13132 13124
rect 13172 13084 14284 13124
rect 14324 13084 14333 13124
rect 17155 13084 17164 13124
rect 17204 13084 17452 13124
rect 17492 13084 17501 13124
rect 19171 13084 19180 13124
rect 19220 13084 22484 13124
rect 25420 13124 25460 13168
rect 28003 13167 28061 13168
rect 28195 13124 28253 13125
rect 30028 13124 30068 13168
rect 25420 13084 26764 13124
rect 26804 13084 26813 13124
rect 28110 13084 28204 13124
rect 28244 13084 29260 13124
rect 29300 13084 31372 13124
rect 31412 13084 31421 13124
rect 31651 13084 31660 13124
rect 31700 13084 33388 13124
rect 33428 13084 33437 13124
rect 28195 13083 28253 13084
rect 19843 13040 19901 13041
rect 13219 13000 13228 13040
rect 13268 13000 13804 13040
rect 13844 13000 13853 13040
rect 14467 13000 14476 13040
rect 14516 13000 15244 13040
rect 15284 13000 15293 13040
rect 15907 13000 15916 13040
rect 15956 13000 16108 13040
rect 16148 13000 16492 13040
rect 16532 13000 19564 13040
rect 19604 13000 19613 13040
rect 19758 13000 19852 13040
rect 19892 13000 19901 13040
rect 21475 13000 21484 13040
rect 21524 13000 21676 13040
rect 21716 13000 21725 13040
rect 28963 13000 28972 13040
rect 29012 13000 30700 13040
rect 30740 13000 30749 13040
rect 13804 12956 13844 13000
rect 19843 12999 19901 13000
rect 14947 12956 15005 12957
rect 15715 12956 15773 12957
rect 29731 12956 29789 12957
rect 13804 12916 14764 12956
rect 14804 12916 14813 12956
rect 14947 12916 14956 12956
rect 14996 12916 15090 12956
rect 15139 12916 15148 12956
rect 15188 12916 15197 12956
rect 15630 12916 15724 12956
rect 15764 12916 15773 12956
rect 18499 12916 18508 12956
rect 18548 12916 20140 12956
rect 20180 12916 20189 12956
rect 26755 12916 26764 12956
rect 26804 12916 27820 12956
rect 27860 12916 27869 12956
rect 28387 12916 28396 12956
rect 28436 12916 29548 12956
rect 29588 12916 29597 12956
rect 29646 12916 29740 12956
rect 29780 12916 29789 12956
rect 30403 12916 30412 12956
rect 30452 12916 32948 12956
rect 14947 12915 15005 12916
rect 15148 12872 15188 12916
rect 15715 12915 15773 12916
rect 15619 12872 15677 12873
rect 28963 12872 29021 12873
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 14083 12832 14092 12872
rect 14132 12832 15188 12872
rect 15534 12832 15628 12872
rect 15668 12832 15677 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 26851 12832 26860 12872
rect 26900 12832 26909 12872
rect 27331 12832 27340 12872
rect 27380 12832 27389 12872
rect 27907 12832 27916 12872
rect 27956 12832 28972 12872
rect 29012 12832 29021 12872
rect 29548 12872 29588 12916
rect 29731 12915 29789 12916
rect 29548 12832 30604 12872
rect 30644 12832 30653 12872
rect 15619 12831 15677 12832
rect 26659 12788 26717 12789
rect 14467 12748 14476 12788
rect 14516 12748 14860 12788
rect 14900 12748 14909 12788
rect 15139 12748 15148 12788
rect 15188 12748 16012 12788
rect 16052 12748 16061 12788
rect 17923 12748 17932 12788
rect 17972 12748 21868 12788
rect 21908 12748 21917 12788
rect 26574 12748 26668 12788
rect 26708 12748 26717 12788
rect 14947 12664 14956 12704
rect 14996 12664 15340 12704
rect 15380 12664 15389 12704
rect 15715 12664 15724 12704
rect 15764 12664 16204 12704
rect 16244 12664 16253 12704
rect 19075 12664 19084 12704
rect 19124 12664 19468 12704
rect 19508 12664 19517 12704
rect 19564 12620 19604 12748
rect 26659 12747 26717 12748
rect 20227 12664 20236 12704
rect 20276 12664 20716 12704
rect 20756 12664 20765 12704
rect 20812 12664 22540 12704
rect 22580 12664 22589 12704
rect 26275 12664 26284 12704
rect 26324 12664 26572 12704
rect 26612 12664 26621 12704
rect 20812 12620 20852 12664
rect 26860 12620 26900 12832
rect 27340 12788 27380 12832
rect 28963 12831 29021 12832
rect 32908 12788 32948 12916
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 27340 12748 31468 12788
rect 31508 12748 31517 12788
rect 32899 12748 32908 12788
rect 32948 12748 34060 12788
rect 34100 12748 34109 12788
rect 27331 12664 27340 12704
rect 27380 12664 27724 12704
rect 27764 12664 27773 12704
rect 29059 12664 29068 12704
rect 29108 12664 29452 12704
rect 29492 12664 29501 12704
rect 32515 12664 32524 12704
rect 32564 12664 33100 12704
rect 33140 12664 33149 12704
rect 33475 12664 33484 12704
rect 33524 12664 34540 12704
rect 34580 12664 38956 12704
rect 38996 12664 39005 12704
rect 3619 12580 3628 12620
rect 3668 12580 4724 12620
rect 5827 12580 5836 12620
rect 5876 12580 6412 12620
rect 6452 12580 6461 12620
rect 8803 12580 8812 12620
rect 8852 12580 11404 12620
rect 11444 12580 11453 12620
rect 13987 12580 13996 12620
rect 14036 12580 17836 12620
rect 17876 12580 17885 12620
rect 18499 12580 18508 12620
rect 18548 12580 18557 12620
rect 19555 12580 19564 12620
rect 19604 12580 19613 12620
rect 19843 12580 19852 12620
rect 19892 12580 20852 12620
rect 21187 12580 21196 12620
rect 21236 12580 21580 12620
rect 21620 12580 21629 12620
rect 25891 12580 25900 12620
rect 25940 12580 27628 12620
rect 27668 12580 27677 12620
rect 28963 12580 28972 12620
rect 29012 12580 29164 12620
rect 29204 12580 32812 12620
rect 32852 12580 32861 12620
rect 33187 12580 33196 12620
rect 33236 12580 33580 12620
rect 33620 12580 35020 12620
rect 35060 12580 35069 12620
rect 36259 12580 36268 12620
rect 36308 12580 37612 12620
rect 37652 12580 37661 12620
rect 4684 12536 4724 12580
rect 5923 12536 5981 12537
rect 18508 12536 18548 12580
rect 20803 12536 20861 12537
rect 2851 12496 2860 12536
rect 2900 12496 4204 12536
rect 4244 12496 4253 12536
rect 4675 12496 4684 12536
rect 4724 12496 4733 12536
rect 4963 12496 4972 12536
rect 5012 12496 5740 12536
rect 5780 12496 5789 12536
rect 5923 12496 5932 12536
rect 5972 12496 6066 12536
rect 7075 12496 7084 12536
rect 7124 12496 8620 12536
rect 8660 12496 8669 12536
rect 14179 12496 14188 12536
rect 14228 12496 14380 12536
rect 14420 12496 15052 12536
rect 15092 12496 15340 12536
rect 15380 12496 15389 12536
rect 15715 12496 15724 12536
rect 15764 12496 16684 12536
rect 16724 12496 16733 12536
rect 16780 12496 18548 12536
rect 18787 12496 18796 12536
rect 18836 12496 20044 12536
rect 20084 12496 20093 12536
rect 20718 12496 20812 12536
rect 20852 12496 20861 12536
rect 26179 12496 26188 12536
rect 26228 12496 26804 12536
rect 27523 12496 27532 12536
rect 27572 12496 27916 12536
rect 27956 12496 27965 12536
rect 28483 12496 28492 12536
rect 28532 12496 28541 12536
rect 29347 12496 29356 12536
rect 29396 12496 29836 12536
rect 29876 12496 30220 12536
rect 30260 12496 30269 12536
rect 31747 12496 31756 12536
rect 31796 12496 33292 12536
rect 33332 12496 33341 12536
rect 4972 12452 5012 12496
rect 5923 12495 5981 12496
rect 15715 12452 15773 12453
rect 16780 12452 16820 12496
rect 20803 12495 20861 12496
rect 18787 12452 18845 12453
rect 2947 12412 2956 12452
rect 2996 12412 3820 12452
rect 3860 12412 3869 12452
rect 4483 12412 4492 12452
rect 4532 12412 5012 12452
rect 8323 12412 8332 12452
rect 8372 12412 9676 12452
rect 9716 12412 9725 12452
rect 14659 12412 14668 12452
rect 14708 12412 14956 12452
rect 14996 12412 15005 12452
rect 15715 12412 15724 12452
rect 15764 12412 16820 12452
rect 18403 12412 18412 12452
rect 18452 12412 18796 12452
rect 18836 12412 18845 12452
rect 15715 12411 15773 12412
rect 18787 12411 18845 12412
rect 18979 12452 19037 12453
rect 19747 12452 19805 12453
rect 18979 12412 18988 12452
rect 19028 12412 19122 12452
rect 19662 12412 19756 12452
rect 19796 12412 19805 12452
rect 18979 12411 19037 12412
rect 19747 12411 19805 12412
rect 25987 12452 26045 12453
rect 26764 12452 26804 12496
rect 28492 12452 28532 12496
rect 25987 12412 25996 12452
rect 26036 12412 26092 12452
rect 26132 12412 26141 12452
rect 26755 12412 26764 12452
rect 26804 12412 26813 12452
rect 26860 12412 27284 12452
rect 27427 12412 27436 12452
rect 27476 12412 28532 12452
rect 28675 12412 28684 12452
rect 28724 12412 30124 12452
rect 30164 12412 30173 12452
rect 25987 12411 26045 12412
rect 0 12368 80 12388
rect 15619 12368 15677 12369
rect 26860 12368 26900 12412
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 6979 12328 6988 12368
rect 7028 12328 9580 12368
rect 9620 12328 9629 12368
rect 14755 12328 14764 12368
rect 14804 12328 15628 12368
rect 15668 12328 16588 12368
rect 16628 12328 16637 12368
rect 18307 12328 18316 12368
rect 18356 12328 24748 12368
rect 24788 12328 24797 12368
rect 25987 12328 25996 12368
rect 26036 12328 26572 12368
rect 26612 12328 26900 12368
rect 27244 12368 27284 12412
rect 27244 12328 28300 12368
rect 28340 12328 28349 12368
rect 28483 12328 28492 12368
rect 28532 12328 29260 12368
rect 29300 12328 30412 12368
rect 30452 12328 30461 12368
rect 0 12308 80 12328
rect 15619 12327 15677 12328
rect 11779 12284 11837 12285
rect 14947 12284 15005 12285
rect 18883 12284 18941 12285
rect 19747 12284 19805 12285
rect 20035 12284 20093 12285
rect 11694 12244 11788 12284
rect 11828 12244 11837 12284
rect 14371 12244 14380 12284
rect 14420 12244 14956 12284
rect 14996 12244 15724 12284
rect 15764 12244 15773 12284
rect 18787 12244 18796 12284
rect 18836 12244 18892 12284
rect 18932 12244 18941 12284
rect 19459 12244 19468 12284
rect 19508 12244 19756 12284
rect 19796 12244 19892 12284
rect 19950 12244 20044 12284
rect 20084 12244 20093 12284
rect 24748 12284 24788 12328
rect 24748 12244 28108 12284
rect 28148 12244 28396 12284
rect 28436 12244 28445 12284
rect 31843 12244 31852 12284
rect 31892 12244 32332 12284
rect 32372 12244 32381 12284
rect 11779 12243 11837 12244
rect 14947 12243 15005 12244
rect 18883 12243 18941 12244
rect 19747 12243 19805 12244
rect 19852 12200 19892 12244
rect 20035 12243 20093 12244
rect 34435 12200 34493 12201
rect 19852 12160 24692 12200
rect 26275 12160 26284 12200
rect 26324 12160 26956 12200
rect 26996 12160 32236 12200
rect 32276 12160 34444 12200
rect 34484 12160 34493 12200
rect 19939 12116 19997 12117
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 18979 12076 18988 12116
rect 19028 12076 19948 12116
rect 19988 12076 19997 12116
rect 19939 12075 19997 12076
rect 20131 12116 20189 12117
rect 20131 12076 20140 12116
rect 20180 12076 20620 12116
rect 20660 12076 20669 12116
rect 20131 12075 20189 12076
rect 19075 11992 19084 12032
rect 19124 11992 19756 12032
rect 19796 11992 19805 12032
rect 24652 11948 24692 12160
rect 34435 12159 34493 12160
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 26659 12032 26717 12033
rect 26659 11992 26668 12032
rect 26708 11992 27244 12032
rect 27284 11992 27293 12032
rect 26659 11991 26717 11992
rect 26755 11948 26813 11949
rect 8035 11908 8044 11948
rect 8084 11908 8428 11948
rect 8468 11908 9292 11948
rect 9332 11908 9341 11948
rect 12643 11908 12652 11948
rect 12692 11908 13708 11948
rect 13748 11908 13757 11948
rect 13987 11908 13996 11948
rect 14036 11908 17836 11948
rect 17876 11908 17885 11948
rect 24652 11908 26764 11948
rect 26804 11908 26956 11948
rect 26996 11908 27005 11948
rect 29059 11908 29068 11948
rect 29108 11908 29740 11948
rect 29780 11908 29789 11948
rect 33475 11908 33484 11948
rect 33524 11908 33964 11948
rect 34004 11908 34013 11948
rect 26755 11907 26813 11908
rect 17923 11864 17981 11865
rect 35011 11864 35069 11865
rect 14947 11824 14956 11864
rect 14996 11824 15860 11864
rect 17155 11824 17164 11864
rect 17204 11824 17932 11864
rect 17972 11824 17981 11864
rect 15820 11780 15860 11824
rect 17923 11823 17981 11824
rect 18220 11824 19468 11864
rect 19508 11824 19517 11864
rect 19747 11824 19756 11864
rect 19796 11824 19948 11864
rect 19988 11824 19997 11864
rect 26371 11824 26380 11864
rect 26420 11824 26460 11864
rect 26755 11824 26764 11864
rect 26804 11824 27148 11864
rect 27188 11824 27197 11864
rect 29635 11824 29644 11864
rect 29684 11824 30124 11864
rect 30164 11824 30173 11864
rect 32707 11824 32716 11864
rect 32756 11824 33580 11864
rect 33620 11824 33629 11864
rect 33763 11824 33772 11864
rect 33812 11824 34732 11864
rect 34772 11824 34781 11864
rect 34926 11824 35020 11864
rect 35060 11824 35069 11864
rect 18220 11780 18260 11824
rect 21571 11780 21629 11781
rect 26380 11780 26420 11824
rect 35011 11823 35069 11824
rect 29731 11780 29789 11781
rect 15340 11740 15724 11780
rect 15764 11740 15773 11780
rect 15820 11740 18220 11780
rect 18260 11740 18269 11780
rect 18321 11740 18377 11780
rect 18417 11740 19372 11780
rect 19412 11740 20201 11780
rect 20241 11740 21580 11780
rect 21620 11740 21629 11780
rect 15340 11696 15380 11740
rect 18321 11696 18361 11740
rect 21571 11739 21629 11740
rect 26188 11740 26668 11780
rect 26708 11740 26717 11780
rect 29347 11740 29356 11780
rect 29396 11740 29740 11780
rect 29780 11740 33236 11780
rect 26083 11696 26141 11697
rect 26188 11696 26228 11740
rect 29731 11739 29789 11740
rect 33196 11696 33236 11740
rect 6019 11656 6028 11696
rect 6068 11656 7660 11696
rect 7700 11656 7709 11696
rect 10051 11656 10060 11696
rect 10100 11656 11980 11696
rect 12020 11656 12029 11696
rect 12451 11656 12460 11696
rect 12500 11656 12844 11696
rect 12884 11656 12893 11696
rect 14851 11656 14860 11696
rect 14900 11656 15340 11696
rect 15380 11656 15389 11696
rect 15523 11656 15532 11696
rect 15572 11656 16300 11696
rect 16340 11656 16588 11696
rect 16628 11656 16637 11696
rect 16963 11656 16972 11696
rect 17012 11656 18361 11696
rect 19180 11656 19564 11696
rect 19604 11656 19948 11696
rect 19988 11656 19997 11696
rect 21763 11656 21772 11696
rect 21812 11656 22252 11696
rect 22292 11656 22301 11696
rect 23011 11656 23020 11696
rect 23060 11656 23692 11696
rect 23732 11656 23741 11696
rect 26083 11656 26092 11696
rect 26132 11656 26188 11696
rect 26228 11656 26237 11696
rect 26371 11656 26380 11696
rect 26420 11656 27148 11696
rect 27188 11656 27197 11696
rect 31363 11656 31372 11696
rect 31412 11656 31756 11696
rect 31796 11656 31805 11696
rect 33187 11656 33196 11696
rect 33236 11656 34252 11696
rect 34292 11656 38764 11696
rect 38804 11656 39532 11696
rect 39572 11656 39581 11696
rect 17923 11612 17981 11613
rect 19180 11612 19220 11656
rect 26083 11655 26141 11656
rect 17923 11572 17932 11612
rect 17972 11572 18076 11612
rect 18116 11572 19180 11612
rect 19220 11572 19229 11612
rect 25795 11572 25804 11612
rect 25844 11572 27436 11612
rect 27476 11572 27485 11612
rect 30211 11572 30220 11612
rect 30260 11572 32716 11612
rect 32756 11572 36076 11612
rect 36116 11572 37804 11612
rect 37844 11572 37853 11612
rect 17923 11571 17981 11572
rect 0 11528 80 11548
rect 15235 11528 15293 11529
rect 16099 11528 16157 11529
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 13507 11488 13516 11528
rect 13556 11488 13900 11528
rect 13940 11488 13949 11528
rect 15150 11488 15244 11528
rect 15284 11488 15293 11528
rect 16014 11488 16108 11528
rect 16148 11488 16157 11528
rect 16291 11488 16300 11528
rect 16340 11488 16876 11528
rect 16916 11488 16925 11528
rect 17923 11488 17932 11528
rect 17972 11488 19276 11528
rect 19316 11488 19325 11528
rect 19651 11488 19660 11528
rect 19700 11488 19709 11528
rect 25603 11488 25612 11528
rect 25652 11488 26092 11528
rect 26132 11488 26141 11528
rect 29155 11488 29164 11528
rect 29204 11488 29644 11528
rect 29684 11488 29693 11528
rect 0 11468 80 11488
rect 15235 11487 15293 11488
rect 16099 11487 16157 11488
rect 15427 11444 15485 11445
rect 19660 11444 19700 11488
rect 7267 11404 7276 11444
rect 7316 11404 8468 11444
rect 14563 11404 14572 11444
rect 14612 11404 15140 11444
rect 8428 11360 8468 11404
rect 15100 11360 15140 11404
rect 15427 11404 15436 11444
rect 15476 11404 15668 11444
rect 17827 11404 17836 11444
rect 17876 11404 18892 11444
rect 18932 11404 19700 11444
rect 31843 11404 31852 11444
rect 31892 11404 37516 11444
rect 37556 11404 37708 11444
rect 37748 11404 37757 11444
rect 15427 11403 15485 11404
rect 15331 11360 15389 11361
rect 15628 11360 15668 11404
rect 16387 11360 16445 11361
rect 29923 11360 29981 11361
rect 35788 11360 35828 11404
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 8388 11320 8428 11360
rect 8468 11320 8477 11360
rect 15100 11320 15148 11360
rect 15188 11320 15197 11360
rect 15331 11320 15340 11360
rect 15380 11320 15474 11360
rect 15588 11320 15628 11360
rect 15668 11320 15677 11360
rect 16302 11320 16396 11360
rect 16436 11320 16445 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 29347 11320 29356 11360
rect 29396 11320 29932 11360
rect 29972 11320 29981 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 35395 11320 35404 11360
rect 35444 11320 35453 11360
rect 35748 11320 35788 11360
rect 35828 11320 35837 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 15331 11319 15389 11320
rect 16387 11319 16445 11320
rect 29923 11319 29981 11320
rect 35404 11276 35444 11320
rect 9763 11236 9772 11276
rect 9812 11236 11540 11276
rect 11683 11236 11692 11276
rect 11732 11236 20332 11276
rect 20372 11236 20381 11276
rect 20611 11236 20620 11276
rect 20660 11236 23116 11276
rect 23156 11236 24172 11276
rect 24212 11236 24221 11276
rect 25795 11236 25804 11276
rect 25844 11236 31665 11276
rect 31705 11236 31714 11276
rect 33091 11236 33100 11276
rect 33140 11236 34348 11276
rect 34388 11236 35444 11276
rect 7459 10984 7468 11024
rect 7508 10984 9292 11024
rect 9332 10984 9341 11024
rect 10339 10984 10348 11024
rect 10388 10984 11020 11024
rect 11060 10984 11069 11024
rect 11500 10856 11540 11236
rect 25987 11192 26045 11193
rect 35011 11192 35069 11193
rect 25699 11152 25708 11192
rect 25748 11152 25996 11192
rect 26036 11152 26476 11192
rect 26516 11152 26525 11192
rect 26659 11152 26668 11192
rect 26708 11152 30124 11192
rect 30164 11152 30316 11192
rect 30356 11152 30508 11192
rect 30548 11152 30557 11192
rect 35011 11152 35020 11192
rect 35060 11152 35404 11192
rect 35444 11152 35453 11192
rect 25987 11151 26045 11152
rect 35011 11151 35069 11152
rect 15715 11108 15773 11109
rect 15043 11068 15052 11108
rect 15092 11068 15724 11108
rect 15764 11068 15916 11108
rect 15956 11068 17356 11108
rect 17396 11068 17405 11108
rect 22147 11068 22156 11108
rect 22196 11068 22540 11108
rect 22580 11068 22589 11108
rect 24355 11068 24364 11108
rect 24404 11068 25132 11108
rect 25172 11068 25181 11108
rect 26284 11068 27340 11108
rect 27380 11068 27389 11108
rect 29251 11068 29260 11108
rect 29300 11068 29309 11108
rect 30700 11068 31564 11108
rect 31604 11068 32236 11108
rect 32276 11068 32524 11108
rect 32564 11068 32716 11108
rect 32756 11068 32765 11108
rect 35299 11068 35308 11108
rect 35348 11068 36076 11108
rect 36116 11068 36125 11108
rect 15715 11067 15773 11068
rect 26284 11024 26324 11068
rect 29260 11024 29300 11068
rect 30700 11024 30740 11068
rect 32515 11024 32573 11025
rect 15715 10984 15724 11024
rect 15764 10984 16204 11024
rect 16244 10984 16253 11024
rect 17443 10984 17452 11024
rect 17492 10984 17836 11024
rect 17876 10984 17885 11024
rect 18307 10984 18316 11024
rect 18356 10984 19852 11024
rect 19892 10984 19901 11024
rect 22051 10984 22060 11024
rect 22100 10984 23788 11024
rect 23828 10984 24748 11024
rect 24788 10984 24797 11024
rect 26275 10984 26284 11024
rect 26324 10984 26333 11024
rect 26467 10984 26476 11024
rect 26516 10984 27052 11024
rect 27092 10984 27101 11024
rect 29260 10984 29356 11024
rect 29396 10984 29405 11024
rect 29827 10984 29836 11024
rect 29876 10984 30124 11024
rect 30164 10984 30173 11024
rect 30691 10984 30700 11024
rect 30740 10984 30749 11024
rect 31459 10984 31468 11024
rect 31508 10984 32044 11024
rect 32084 10984 32093 11024
rect 32419 10984 32428 11024
rect 32468 10984 32524 11024
rect 32564 10984 32573 11024
rect 34723 10984 34732 11024
rect 34772 10984 35500 11024
rect 35540 10984 38092 11024
rect 38132 10984 38141 11024
rect 32515 10983 32573 10984
rect 15907 10940 15965 10941
rect 18691 10940 18749 10941
rect 26659 10940 26717 10941
rect 15235 10900 15244 10940
rect 15284 10900 15436 10940
rect 15476 10900 15916 10940
rect 15956 10900 16108 10940
rect 16148 10900 16157 10940
rect 17539 10900 17548 10940
rect 17588 10900 18508 10940
rect 18548 10900 18700 10940
rect 18740 10900 18749 10940
rect 26574 10900 26668 10940
rect 26708 10900 26717 10940
rect 29251 10900 29260 10940
rect 29300 10900 30604 10940
rect 30644 10900 30653 10940
rect 15907 10899 15965 10900
rect 18691 10899 18749 10900
rect 26659 10899 26717 10900
rect 17731 10856 17789 10857
rect 11491 10816 11500 10856
rect 11540 10816 11549 10856
rect 13603 10816 13612 10856
rect 13652 10816 17068 10856
rect 17108 10816 17740 10856
rect 17780 10816 28684 10856
rect 28724 10816 28733 10856
rect 28867 10816 28876 10856
rect 28916 10816 32524 10856
rect 32564 10816 33004 10856
rect 33044 10816 33053 10856
rect 34819 10816 34828 10856
rect 34868 10816 35500 10856
rect 35540 10816 35549 10856
rect 17731 10815 17789 10816
rect 7267 10732 7276 10772
rect 7316 10732 7852 10772
rect 7892 10732 7901 10772
rect 11203 10732 11212 10772
rect 11252 10732 12364 10772
rect 12404 10732 12413 10772
rect 19075 10732 19084 10772
rect 19124 10732 20140 10772
rect 20180 10732 20189 10772
rect 20707 10732 20716 10772
rect 20756 10732 21868 10772
rect 21908 10732 21917 10772
rect 26083 10732 26092 10772
rect 26132 10732 26956 10772
rect 26996 10732 27005 10772
rect 29635 10732 29644 10772
rect 29684 10732 30028 10772
rect 30068 10732 30077 10772
rect 35203 10732 35212 10772
rect 35252 10732 35884 10772
rect 35924 10732 35933 10772
rect 0 10688 80 10708
rect 26380 10688 26420 10732
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 17347 10648 17356 10688
rect 17396 10648 21388 10688
rect 21428 10648 21437 10688
rect 26371 10648 26380 10688
rect 26420 10648 26460 10688
rect 0 10628 80 10648
rect 33091 10604 33149 10605
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 32707 10564 32716 10604
rect 32756 10564 33100 10604
rect 33140 10564 33149 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 33091 10563 33149 10564
rect 20140 10480 26188 10520
rect 26228 10480 26237 10520
rect 29155 10480 29164 10520
rect 29204 10480 29548 10520
rect 29588 10480 29597 10520
rect 10147 10396 10156 10436
rect 10196 10396 13516 10436
rect 13556 10396 13565 10436
rect 16099 10352 16157 10353
rect 9955 10312 9964 10352
rect 10004 10312 11308 10352
rect 11348 10312 12556 10352
rect 12596 10312 12605 10352
rect 16014 10312 16108 10352
rect 16148 10312 16157 10352
rect 16099 10311 16157 10312
rect 20140 10268 20180 10480
rect 20323 10396 20332 10436
rect 20372 10396 22060 10436
rect 22100 10396 22109 10436
rect 29260 10396 29644 10436
rect 29684 10396 30124 10436
rect 30164 10396 30173 10436
rect 32803 10396 32812 10436
rect 32852 10396 34348 10436
rect 34388 10396 34397 10436
rect 35011 10396 35020 10436
rect 35060 10396 35692 10436
rect 35732 10396 35741 10436
rect 26275 10312 26284 10352
rect 26324 10312 27153 10352
rect 27193 10312 27202 10352
rect 29260 10268 29300 10396
rect 12643 10228 12652 10268
rect 12692 10228 20180 10268
rect 20323 10228 20332 10268
rect 20372 10228 21484 10268
rect 21524 10228 21533 10268
rect 23395 10228 23404 10268
rect 23444 10228 23692 10268
rect 23732 10228 23741 10268
rect 27436 10228 29300 10268
rect 29356 10312 30604 10352
rect 30644 10312 30653 10352
rect 32323 10312 32332 10352
rect 32372 10312 33196 10352
rect 33236 10312 33245 10352
rect 37780 10312 38188 10352
rect 38228 10312 38237 10352
rect 27436 10184 27476 10228
rect 29356 10184 29396 10312
rect 32515 10268 32573 10269
rect 37780 10268 37820 10312
rect 30403 10228 30412 10268
rect 30452 10228 30796 10268
rect 30836 10228 31372 10268
rect 31412 10228 32524 10268
rect 32564 10228 32812 10268
rect 32852 10228 32861 10268
rect 34339 10228 34348 10268
rect 34388 10228 35308 10268
rect 35348 10228 35788 10268
rect 35828 10228 37820 10268
rect 32515 10227 32573 10228
rect 7651 10144 7660 10184
rect 7700 10144 9484 10184
rect 9524 10144 9533 10184
rect 9667 10144 9676 10184
rect 9716 10144 17548 10184
rect 17588 10144 17597 10184
rect 20803 10144 20812 10184
rect 20852 10144 21964 10184
rect 22004 10144 23020 10184
rect 23060 10144 23069 10184
rect 24355 10144 24364 10184
rect 24404 10144 25420 10184
rect 25460 10144 25469 10184
rect 26179 10144 26188 10184
rect 26228 10144 27052 10184
rect 27092 10144 27436 10184
rect 27476 10144 27485 10184
rect 28195 10144 28204 10184
rect 28244 10144 29164 10184
rect 29204 10144 29213 10184
rect 29347 10144 29356 10184
rect 29396 10144 29405 10184
rect 29832 10144 29841 10184
rect 29881 10144 32180 10184
rect 32227 10144 32236 10184
rect 32276 10144 32908 10184
rect 32948 10144 32957 10184
rect 33091 10144 33100 10184
rect 33140 10144 33149 10184
rect 36643 10144 36652 10184
rect 36692 10144 37900 10184
rect 37940 10144 38380 10184
rect 38420 10144 38668 10184
rect 38708 10144 38717 10184
rect 32140 10100 32180 10144
rect 33100 10100 33140 10144
rect 5539 10060 5548 10100
rect 5588 10060 6988 10100
rect 7028 10060 7037 10100
rect 10147 10060 10156 10100
rect 10196 10060 11404 10100
rect 11444 10060 11453 10100
rect 11779 10060 11788 10100
rect 11828 10060 15052 10100
rect 15092 10060 15101 10100
rect 16963 10060 16972 10100
rect 17012 10060 18892 10100
rect 18932 10060 18941 10100
rect 20899 10060 20908 10100
rect 20948 10060 21388 10100
rect 21428 10060 22444 10100
rect 22484 10060 22493 10100
rect 24835 10060 24844 10100
rect 24884 10060 28876 10100
rect 28916 10060 28925 10100
rect 29740 10060 30316 10100
rect 30356 10060 30365 10100
rect 32140 10060 32620 10100
rect 32660 10060 33004 10100
rect 33044 10060 33053 10100
rect 33100 10060 38860 10100
rect 38900 10060 39820 10100
rect 39860 10060 39869 10100
rect 29740 10016 29780 10060
rect 8515 9976 8524 10016
rect 8564 9976 10348 10016
rect 10388 9976 10397 10016
rect 14083 9976 14092 10016
rect 14132 9976 18988 10016
rect 19028 9976 19037 10016
rect 25315 9976 25324 10016
rect 25364 9976 26284 10016
rect 26324 9976 26333 10016
rect 27144 9976 27153 10016
rect 27193 9976 29684 10016
rect 29731 9976 29740 10016
rect 29780 9976 29789 10016
rect 35011 9976 35020 10016
rect 35060 9976 35596 10016
rect 35636 9976 35645 10016
rect 18019 9932 18077 9933
rect 29644 9932 29684 9976
rect 15244 9892 18028 9932
rect 18068 9892 18077 9932
rect 28579 9892 28588 9932
rect 28628 9892 29452 9932
rect 29492 9892 29501 9932
rect 29644 9892 29836 9932
rect 29876 9892 31180 9932
rect 31220 9892 31229 9932
rect 0 9848 80 9868
rect 15244 9848 15284 9892
rect 18019 9891 18077 9892
rect 15715 9848 15773 9849
rect 16195 9848 16253 9849
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 15235 9808 15244 9848
rect 15284 9808 15293 9848
rect 15630 9808 15724 9848
rect 15764 9808 15773 9848
rect 16110 9808 16204 9848
rect 16244 9808 16253 9848
rect 16387 9808 16396 9848
rect 16436 9808 16780 9848
rect 16820 9808 16829 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 0 9788 80 9808
rect 15715 9807 15773 9808
rect 16195 9807 16253 9808
rect 15427 9724 15436 9764
rect 15476 9724 15916 9764
rect 15956 9724 16876 9764
rect 16916 9724 16925 9764
rect 20035 9724 20044 9764
rect 20084 9724 20180 9764
rect 26755 9724 26764 9764
rect 26804 9724 27340 9764
rect 27380 9724 27389 9764
rect 29635 9724 29644 9764
rect 29684 9724 30124 9764
rect 30164 9724 30173 9764
rect 14947 9680 15005 9681
rect 11299 9640 11308 9680
rect 11348 9640 12076 9680
rect 12116 9640 12125 9680
rect 13411 9640 13420 9680
rect 13460 9640 13900 9680
rect 13940 9640 14668 9680
rect 14708 9640 14717 9680
rect 14862 9640 14956 9680
rect 14996 9640 15005 9680
rect 15811 9640 15820 9680
rect 15860 9640 16204 9680
rect 16244 9640 16253 9680
rect 14947 9639 15005 9640
rect 9580 9556 13804 9596
rect 13844 9556 13853 9596
rect 9580 9512 9620 9556
rect 8131 9472 8140 9512
rect 8180 9472 9388 9512
rect 9428 9472 9437 9512
rect 9571 9472 9580 9512
rect 9620 9472 9629 9512
rect 9955 9472 9964 9512
rect 10004 9472 10444 9512
rect 10484 9472 10493 9512
rect 11203 9472 11212 9512
rect 11252 9472 11692 9512
rect 11732 9472 11741 9512
rect 13507 9472 13516 9512
rect 13556 9472 13996 9512
rect 14036 9472 14045 9512
rect 14947 9472 14956 9512
rect 14996 9472 15340 9512
rect 15380 9472 15389 9512
rect 16003 9472 16012 9512
rect 16052 9472 16588 9512
rect 16628 9472 16637 9512
rect 20140 9428 20180 9724
rect 27427 9640 27436 9680
rect 27476 9640 27820 9680
rect 27860 9640 28876 9680
rect 28916 9640 29932 9680
rect 29972 9640 29981 9680
rect 34435 9640 34444 9680
rect 34484 9640 35212 9680
rect 35252 9640 35261 9680
rect 34819 9596 34877 9597
rect 24835 9556 24844 9596
rect 24884 9556 29684 9596
rect 30307 9556 30316 9596
rect 30356 9556 30700 9596
rect 30740 9556 32332 9596
rect 32372 9556 33004 9596
rect 33044 9556 34828 9596
rect 34868 9556 34877 9596
rect 29644 9512 29684 9556
rect 34819 9555 34877 9556
rect 31843 9512 31901 9513
rect 32611 9512 32669 9513
rect 33091 9512 33149 9513
rect 23395 9472 23404 9512
rect 23444 9472 24172 9512
rect 24212 9472 24221 9512
rect 28675 9472 28684 9512
rect 28724 9472 29068 9512
rect 29108 9472 29356 9512
rect 29396 9472 29405 9512
rect 29635 9472 29644 9512
rect 29684 9472 29693 9512
rect 29923 9472 29932 9512
rect 29972 9472 30508 9512
rect 30548 9472 30557 9512
rect 31758 9472 31852 9512
rect 31892 9472 31901 9512
rect 32526 9472 32620 9512
rect 32660 9472 32669 9512
rect 33006 9472 33100 9512
rect 33140 9472 33149 9512
rect 34243 9472 34252 9512
rect 34292 9472 35212 9512
rect 35252 9472 37324 9512
rect 37364 9472 37373 9512
rect 31843 9471 31901 9472
rect 32611 9471 32669 9472
rect 33091 9471 33149 9472
rect 34819 9428 34877 9429
rect 7939 9388 7948 9428
rect 7988 9388 9100 9428
rect 9140 9388 9149 9428
rect 9283 9388 9292 9428
rect 9332 9388 9868 9428
rect 9908 9388 9917 9428
rect 11107 9388 11116 9428
rect 11156 9388 11596 9428
rect 11636 9388 13420 9428
rect 13460 9388 13469 9428
rect 14659 9388 14668 9428
rect 14708 9388 14860 9428
rect 14900 9388 15436 9428
rect 15476 9388 15485 9428
rect 16012 9388 22828 9428
rect 22868 9388 22877 9428
rect 25219 9388 25228 9428
rect 25268 9388 25277 9428
rect 28780 9388 29548 9428
rect 29588 9388 29597 9428
rect 33955 9388 33964 9428
rect 34004 9388 34444 9428
rect 34484 9388 34493 9428
rect 34536 9388 34545 9428
rect 34585 9388 34594 9428
rect 34819 9388 34828 9428
rect 34868 9388 37996 9428
rect 38036 9388 38045 9428
rect 15907 9344 15965 9345
rect 12643 9304 12652 9344
rect 12692 9304 12844 9344
rect 12884 9304 12893 9344
rect 13123 9304 13132 9344
rect 13172 9304 14284 9344
rect 14324 9304 14333 9344
rect 15822 9304 15916 9344
rect 15956 9304 15965 9344
rect 15907 9303 15965 9304
rect 11011 9220 11020 9260
rect 11060 9220 11980 9260
rect 12020 9220 12029 9260
rect 14563 9220 14572 9260
rect 14612 9220 15820 9260
rect 15860 9220 15869 9260
rect 16012 9176 16052 9388
rect 25228 9344 25268 9388
rect 28780 9344 28820 9388
rect 33859 9344 33917 9345
rect 34540 9344 34580 9388
rect 34819 9387 34877 9388
rect 16483 9304 16492 9344
rect 16532 9304 17164 9344
rect 17204 9304 17213 9344
rect 24547 9304 24556 9344
rect 24596 9304 24940 9344
rect 24980 9304 25268 9344
rect 28771 9304 28780 9344
rect 28820 9304 28829 9344
rect 28960 9304 29255 9344
rect 29295 9304 29304 9344
rect 33859 9304 33868 9344
rect 33908 9304 35596 9344
rect 35636 9304 35645 9344
rect 28960 9260 29000 9304
rect 33859 9303 33917 9304
rect 16963 9220 16972 9260
rect 17012 9220 17548 9260
rect 17588 9220 17597 9260
rect 28291 9220 28300 9260
rect 28340 9220 29000 9260
rect 34147 9220 34156 9260
rect 34196 9220 35404 9260
rect 35444 9220 35453 9260
rect 16195 9176 16253 9177
rect 15043 9136 15052 9176
rect 15092 9136 16052 9176
rect 16099 9136 16108 9176
rect 16148 9136 16204 9176
rect 16244 9136 16253 9176
rect 28963 9136 28972 9176
rect 29012 9136 29164 9176
rect 29204 9136 32620 9176
rect 32660 9136 33004 9176
rect 33044 9136 33053 9176
rect 16195 9135 16253 9136
rect 34051 9092 34109 9093
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 22531 9052 22540 9092
rect 22580 9052 30220 9092
rect 30260 9052 30269 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 33966 9052 34060 9092
rect 34100 9052 34109 9092
rect 34339 9052 34348 9092
rect 34388 9052 34397 9092
rect 34531 9052 34540 9092
rect 34580 9052 34828 9092
rect 34868 9052 35116 9092
rect 35156 9052 35165 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 34051 9051 34109 9052
rect 0 9008 80 9028
rect 34348 9008 34388 9052
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 24163 8968 24172 9008
rect 24212 8968 24652 9008
rect 24692 8968 24701 9008
rect 31459 8968 31468 9008
rect 31508 8968 31948 9008
rect 31988 8968 31997 9008
rect 33580 8968 34388 9008
rect 0 8948 80 8968
rect 9859 8884 9868 8924
rect 9908 8884 10348 8924
rect 10388 8884 11692 8924
rect 11732 8884 11741 8924
rect 13699 8884 13708 8924
rect 13748 8884 14860 8924
rect 14900 8884 14909 8924
rect 15715 8884 15724 8924
rect 15764 8884 16820 8924
rect 21667 8884 21676 8924
rect 21716 8884 27340 8924
rect 27380 8884 27389 8924
rect 16780 8840 16820 8884
rect 18787 8840 18845 8841
rect 25027 8840 25085 8841
rect 27715 8840 27773 8841
rect 31939 8840 31997 8841
rect 33580 8840 33620 8968
rect 34060 8884 34636 8924
rect 34676 8884 34685 8924
rect 37987 8884 37996 8924
rect 38036 8884 39052 8924
rect 39092 8884 39101 8924
rect 3427 8800 3436 8840
rect 3476 8800 6124 8840
rect 6164 8800 6173 8840
rect 10627 8800 10636 8840
rect 10676 8800 14764 8840
rect 14804 8800 14813 8840
rect 15523 8800 15532 8840
rect 15572 8800 16588 8840
rect 16628 8800 16637 8840
rect 16771 8800 16780 8840
rect 16820 8800 18796 8840
rect 18836 8800 18845 8840
rect 23971 8800 23980 8840
rect 24020 8800 24652 8840
rect 24692 8800 24701 8840
rect 24942 8800 25036 8840
rect 25076 8800 25085 8840
rect 27630 8800 27724 8840
rect 27764 8800 27773 8840
rect 28483 8800 28492 8840
rect 28532 8800 30028 8840
rect 30068 8800 30077 8840
rect 31555 8800 31564 8840
rect 31604 8800 31948 8840
rect 31988 8800 31997 8840
rect 33475 8800 33484 8840
rect 33524 8800 33620 8840
rect 33859 8840 33917 8841
rect 33859 8800 33868 8840
rect 33908 8800 33917 8840
rect 18787 8799 18845 8800
rect 25027 8799 25085 8800
rect 27715 8799 27773 8800
rect 31939 8799 31997 8800
rect 33859 8799 33917 8800
rect 20515 8716 20524 8756
rect 20564 8716 22732 8756
rect 22772 8716 23404 8756
rect 23444 8716 23453 8756
rect 27331 8716 27340 8756
rect 27380 8716 28396 8756
rect 28436 8716 28445 8756
rect 30787 8716 30796 8756
rect 30836 8716 32428 8756
rect 32468 8716 32477 8756
rect 33868 8672 33908 8799
rect 34060 8672 34100 8884
rect 34147 8716 34156 8756
rect 34196 8716 36268 8756
rect 36308 8716 36317 8756
rect 5923 8632 5932 8672
rect 5972 8632 6220 8672
rect 6260 8632 6269 8672
rect 7939 8632 7948 8672
rect 7988 8632 10732 8672
rect 10772 8632 12268 8672
rect 12308 8632 12317 8672
rect 12739 8632 12748 8672
rect 12788 8632 13420 8672
rect 13460 8632 14284 8672
rect 14324 8632 14333 8672
rect 15619 8632 15628 8672
rect 15668 8632 16300 8672
rect 16340 8632 16349 8672
rect 20323 8632 20332 8672
rect 20372 8632 26092 8672
rect 26132 8632 26141 8672
rect 26563 8632 26572 8672
rect 26612 8632 27052 8672
rect 27092 8632 27101 8672
rect 27907 8632 27916 8672
rect 27956 8632 29068 8672
rect 29108 8632 29117 8672
rect 31651 8632 31660 8672
rect 31700 8632 31709 8672
rect 31939 8632 31948 8672
rect 31988 8632 32716 8672
rect 32756 8632 32765 8672
rect 33667 8632 33676 8672
rect 33716 8632 33908 8672
rect 33955 8632 33964 8672
rect 34004 8632 35308 8672
rect 35348 8632 35357 8672
rect 31660 8588 31700 8632
rect 34435 8588 34493 8589
rect 24067 8548 24076 8588
rect 24116 8548 24748 8588
rect 24788 8548 25132 8588
rect 25172 8548 25181 8588
rect 25603 8548 25612 8588
rect 25652 8548 27244 8588
rect 27284 8548 27293 8588
rect 29827 8548 29836 8588
rect 29876 8548 30124 8588
rect 30164 8548 31508 8588
rect 31660 8548 33196 8588
rect 33236 8548 33245 8588
rect 34435 8548 34444 8588
rect 34484 8548 34828 8588
rect 34868 8548 34877 8588
rect 31468 8504 31508 8548
rect 32908 8504 32948 8548
rect 34435 8547 34493 8548
rect 8899 8464 8908 8504
rect 8948 8464 10540 8504
rect 10580 8464 10589 8504
rect 14659 8464 14668 8504
rect 14708 8464 16012 8504
rect 16052 8464 16061 8504
rect 22915 8464 22924 8504
rect 22964 8464 23596 8504
rect 23636 8464 23645 8504
rect 25027 8464 25036 8504
rect 25076 8464 25228 8504
rect 25268 8464 25277 8504
rect 25891 8464 25900 8504
rect 25940 8464 26188 8504
rect 26228 8464 26237 8504
rect 27139 8464 27148 8504
rect 27188 8464 31084 8504
rect 31124 8464 31133 8504
rect 31459 8464 31468 8504
rect 31508 8464 31517 8504
rect 31651 8464 31660 8504
rect 31700 8464 32140 8504
rect 32180 8464 32189 8504
rect 32899 8464 32908 8504
rect 32948 8464 32988 8504
rect 33091 8464 33100 8504
rect 33140 8464 33484 8504
rect 33524 8464 33533 8504
rect 14947 8420 15005 8421
rect 14275 8380 14284 8420
rect 14324 8380 14956 8420
rect 14996 8380 16684 8420
rect 16724 8380 19276 8420
rect 19316 8380 20180 8420
rect 23011 8380 23020 8420
rect 23060 8380 24844 8420
rect 24884 8380 25612 8420
rect 25652 8380 25661 8420
rect 26371 8380 26380 8420
rect 26420 8380 27532 8420
rect 27572 8380 31852 8420
rect 31892 8380 32812 8420
rect 32852 8380 32861 8420
rect 14947 8379 15005 8380
rect 15715 8336 15773 8337
rect 20140 8336 20180 8380
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 14755 8296 14764 8336
rect 14804 8296 15724 8336
rect 15764 8296 15773 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 20140 8296 20620 8336
rect 20660 8296 27916 8336
rect 27956 8296 27965 8336
rect 28387 8296 28396 8336
rect 28436 8296 29000 8336
rect 15715 8295 15773 8296
rect 7747 8212 7756 8252
rect 7796 8212 8332 8252
rect 8372 8212 9388 8252
rect 9428 8212 9437 8252
rect 25027 8212 25036 8252
rect 25076 8212 25612 8252
rect 25652 8212 25661 8252
rect 0 8168 80 8188
rect 28960 8168 29000 8296
rect 29068 8296 29740 8336
rect 29780 8296 29789 8336
rect 31852 8296 32620 8336
rect 32660 8296 32669 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 35011 8296 35020 8336
rect 35060 8296 36652 8336
rect 36692 8296 36701 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 29068 8252 29108 8296
rect 31852 8252 31892 8296
rect 35020 8252 35060 8296
rect 29059 8212 29068 8252
rect 29108 8212 29117 8252
rect 31843 8212 31852 8252
rect 31892 8212 31901 8252
rect 33283 8212 33292 8252
rect 33332 8212 35060 8252
rect 29068 8168 29108 8212
rect 34051 8168 34109 8169
rect 0 8128 556 8168
rect 596 8128 605 8168
rect 6691 8128 6700 8168
rect 6740 8128 8236 8168
rect 8276 8128 8285 8168
rect 13123 8128 13132 8168
rect 13172 8128 13181 8168
rect 23395 8128 23404 8168
rect 23444 8128 24172 8168
rect 24212 8128 24221 8168
rect 28960 8128 29108 8168
rect 30211 8128 30220 8168
rect 30260 8128 30700 8168
rect 30740 8128 30749 8168
rect 32428 8128 34060 8168
rect 34100 8128 34109 8168
rect 34243 8128 34252 8168
rect 34292 8128 35692 8168
rect 35732 8128 35741 8168
rect 0 8108 80 8128
rect 4867 8044 4876 8084
rect 4916 8044 5452 8084
rect 5492 8044 5501 8084
rect 4675 7960 4684 8000
rect 4724 7960 5164 8000
rect 5204 7960 5213 8000
rect 7555 7960 7564 8000
rect 7604 7960 9196 8000
rect 9236 7960 9245 8000
rect 13132 7916 13172 8128
rect 28867 8044 28876 8084
rect 28916 8044 30548 8084
rect 31171 8044 31180 8084
rect 31220 8044 31412 8084
rect 30508 8000 30548 8044
rect 15331 7960 15340 8000
rect 15380 7960 16492 8000
rect 16532 7960 16541 8000
rect 16963 7960 16972 8000
rect 17012 7960 18796 8000
rect 18836 7960 19180 8000
rect 19220 7960 19229 8000
rect 20515 7960 20524 8000
rect 20564 7960 21196 8000
rect 21236 7960 21245 8000
rect 22051 7960 22060 8000
rect 22100 7960 22540 8000
rect 22580 7960 22589 8000
rect 23107 7960 23116 8000
rect 23156 7960 23540 8000
rect 24163 7960 24172 8000
rect 24212 7960 25228 8000
rect 25268 7960 25277 8000
rect 25758 7960 25767 8000
rect 25807 7960 25996 8000
rect 26036 7960 26668 8000
rect 26708 7960 26717 8000
rect 28291 7960 28300 8000
rect 28340 7960 29260 8000
rect 29300 7960 29309 8000
rect 30499 7960 30508 8000
rect 30548 7960 30557 8000
rect 23500 7916 23540 7960
rect 25027 7916 25085 7917
rect 31372 7916 31412 8044
rect 32428 8000 32468 8128
rect 34051 8127 34109 8128
rect 33763 8044 33772 8084
rect 33812 8044 34060 8084
rect 34100 8044 37420 8084
rect 37460 8044 37469 8084
rect 31459 7960 31468 8000
rect 31508 7960 31948 8000
rect 31988 7960 32428 8000
rect 32468 7960 32477 8000
rect 33475 7960 33484 8000
rect 33524 7960 34348 8000
rect 34388 7960 34397 8000
rect 36739 7960 36748 8000
rect 36788 7960 37804 8000
rect 37844 7960 37853 8000
rect 6211 7876 6220 7916
rect 6260 7876 7660 7916
rect 7700 7876 7709 7916
rect 13027 7876 13036 7916
rect 13076 7876 13804 7916
rect 13844 7876 14188 7916
rect 14228 7876 14668 7916
rect 14708 7876 15532 7916
rect 15572 7876 15581 7916
rect 23011 7876 23020 7916
rect 23060 7876 23308 7916
rect 23348 7876 23357 7916
rect 23491 7876 23500 7916
rect 23540 7876 23692 7916
rect 23732 7876 25036 7916
rect 25076 7876 25085 7916
rect 25315 7876 25324 7916
rect 25364 7876 28492 7916
rect 28532 7876 28541 7916
rect 30883 7876 30892 7916
rect 30932 7876 31180 7916
rect 31220 7876 31229 7916
rect 31363 7876 31372 7916
rect 31412 7876 31421 7916
rect 32131 7876 32140 7916
rect 32180 7876 32620 7916
rect 32660 7876 32669 7916
rect 25027 7875 25085 7876
rect 4963 7792 4972 7832
rect 5012 7792 5356 7832
rect 5396 7792 5932 7832
rect 5972 7792 6316 7832
rect 6356 7792 6365 7832
rect 26659 7792 26668 7832
rect 26708 7792 28108 7832
rect 28148 7792 28157 7832
rect 28771 7792 28780 7832
rect 28820 7792 30028 7832
rect 30068 7792 30077 7832
rect 30272 7792 30281 7832
rect 30321 7792 31660 7832
rect 31700 7792 31709 7832
rect 33763 7792 33772 7832
rect 33812 7792 36364 7832
rect 36404 7792 36413 7832
rect 25219 7748 25277 7749
rect 31939 7748 31997 7749
rect 2371 7708 2380 7748
rect 2420 7708 3820 7748
rect 3860 7708 3869 7748
rect 7747 7708 7756 7748
rect 7796 7708 8908 7748
rect 8948 7708 8957 7748
rect 9187 7708 9196 7748
rect 9236 7708 10252 7748
rect 10292 7708 10444 7748
rect 10484 7708 10493 7748
rect 21475 7708 21484 7748
rect 21524 7708 23020 7748
rect 23060 7708 23069 7748
rect 25134 7708 25228 7748
rect 25268 7708 25277 7748
rect 29443 7708 29452 7748
rect 29492 7708 31564 7748
rect 31604 7708 31756 7748
rect 31796 7708 31805 7748
rect 31939 7708 31948 7748
rect 31988 7708 32082 7748
rect 33667 7708 33676 7748
rect 33716 7708 34060 7748
rect 34100 7708 34109 7748
rect 25219 7707 25277 7708
rect 31939 7707 31997 7708
rect 7651 7624 7660 7664
rect 7700 7624 9868 7664
rect 9908 7624 9917 7664
rect 10723 7624 10732 7664
rect 10772 7624 11212 7664
rect 11252 7624 11261 7664
rect 26755 7624 26764 7664
rect 26804 7624 30796 7664
rect 30836 7624 30988 7664
rect 31028 7624 31037 7664
rect 30595 7580 30653 7581
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 5827 7540 5836 7580
rect 5876 7540 6220 7580
rect 6260 7540 6796 7580
rect 6836 7540 7372 7580
rect 7412 7540 7421 7580
rect 9955 7540 9964 7580
rect 10004 7540 10348 7580
rect 10388 7540 10397 7580
rect 10627 7540 10636 7580
rect 10676 7540 12844 7580
rect 12884 7540 12893 7580
rect 13987 7540 13996 7580
rect 14036 7540 15244 7580
rect 15284 7540 15293 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 22243 7540 22252 7580
rect 22292 7540 22924 7580
rect 22964 7540 22973 7580
rect 23203 7540 23212 7580
rect 23252 7540 23884 7580
rect 23924 7540 23933 7580
rect 27235 7540 27244 7580
rect 27284 7540 28012 7580
rect 28052 7540 28061 7580
rect 28771 7540 28780 7580
rect 28820 7540 29356 7580
rect 29396 7540 29405 7580
rect 30510 7540 30604 7580
rect 30644 7540 30653 7580
rect 31747 7540 31756 7580
rect 31796 7540 32620 7580
rect 32660 7540 32812 7580
rect 32852 7540 32861 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 34339 7540 34348 7580
rect 34388 7540 35212 7580
rect 35252 7540 35261 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 30595 7539 30653 7540
rect 4771 7456 4780 7496
rect 4820 7456 5164 7496
rect 5204 7456 7468 7496
rect 7508 7456 8428 7496
rect 8468 7456 8477 7496
rect 26563 7456 26572 7496
rect 26612 7456 27052 7496
rect 27092 7456 27101 7496
rect 27144 7456 27153 7496
rect 27193 7456 28052 7496
rect 28675 7456 28684 7496
rect 28724 7456 28972 7496
rect 29012 7456 33812 7496
rect 28012 7412 28052 7456
rect 33772 7412 33812 7456
rect 5443 7372 5452 7412
rect 5492 7372 5836 7412
rect 5876 7372 5885 7412
rect 8131 7372 8140 7412
rect 8180 7372 9100 7412
rect 9140 7372 9149 7412
rect 22243 7372 22252 7412
rect 22292 7372 25516 7412
rect 25556 7372 25565 7412
rect 28012 7372 31276 7412
rect 31316 7372 32332 7412
rect 32372 7372 32524 7412
rect 32564 7372 33484 7412
rect 33524 7372 33533 7412
rect 33763 7372 33772 7412
rect 33812 7372 33964 7412
rect 34004 7372 34013 7412
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 22147 7288 22156 7328
rect 22196 7288 23465 7328
rect 23505 7288 24713 7328
rect 24753 7288 25420 7328
rect 25460 7288 25469 7328
rect 25987 7288 25996 7328
rect 26036 7288 26380 7328
rect 26420 7288 26429 7328
rect 29251 7288 29260 7328
rect 29300 7288 29836 7328
rect 29876 7288 29885 7328
rect 32035 7288 32044 7328
rect 32084 7288 35788 7328
rect 35828 7288 36940 7328
rect 36980 7288 36989 7328
rect 0 7268 80 7288
rect 24547 7244 24605 7245
rect 24462 7204 24556 7244
rect 24596 7204 24605 7244
rect 26380 7244 26420 7288
rect 26380 7204 28780 7244
rect 28820 7204 28829 7244
rect 31651 7204 31660 7244
rect 31700 7204 38092 7244
rect 38132 7204 38956 7244
rect 38996 7204 39005 7244
rect 24547 7203 24605 7204
rect 11491 7160 11549 7161
rect 18883 7160 18941 7161
rect 29251 7160 29309 7161
rect 3619 7120 3628 7160
rect 3668 7120 4972 7160
rect 5012 7120 6508 7160
rect 6548 7120 6557 7160
rect 7459 7120 7468 7160
rect 7508 7120 9004 7160
rect 9044 7120 10924 7160
rect 10964 7120 10973 7160
rect 11395 7120 11404 7160
rect 11444 7120 11500 7160
rect 11540 7120 11549 7160
rect 11875 7120 11884 7160
rect 11924 7120 12748 7160
rect 12788 7120 12797 7160
rect 13219 7120 13228 7160
rect 13268 7120 14284 7160
rect 14324 7120 14333 7160
rect 15043 7120 15052 7160
rect 15092 7120 17548 7160
rect 17588 7120 18028 7160
rect 18068 7120 18077 7160
rect 18883 7120 18892 7160
rect 18932 7120 18988 7160
rect 19028 7120 19037 7160
rect 22627 7120 22636 7160
rect 22676 7120 23788 7160
rect 23828 7120 23980 7160
rect 24020 7120 25036 7160
rect 25076 7120 25085 7160
rect 25411 7120 25420 7160
rect 25460 7120 26668 7160
rect 26708 7120 26717 7160
rect 27198 7120 27207 7160
rect 27247 7120 28108 7160
rect 28148 7120 28157 7160
rect 28675 7120 28684 7160
rect 28724 7120 28876 7160
rect 28916 7120 29000 7160
rect 29166 7120 29260 7160
rect 29300 7120 29309 7160
rect 29731 7120 29740 7160
rect 29780 7120 30124 7160
rect 30164 7120 30892 7160
rect 30932 7120 30941 7160
rect 32323 7120 32332 7160
rect 32372 7120 33868 7160
rect 33908 7120 34924 7160
rect 34964 7120 34973 7160
rect 11491 7119 11549 7120
rect 18883 7119 18941 7120
rect 28960 7076 29000 7120
rect 29251 7119 29309 7120
rect 23500 7036 23884 7076
rect 23924 7036 25228 7076
rect 25268 7036 26860 7076
rect 26900 7036 26909 7076
rect 28960 7036 29452 7076
rect 29492 7036 30220 7076
rect 30260 7036 37228 7076
rect 37268 7036 37900 7076
rect 37940 7036 37949 7076
rect 23500 6992 23540 7036
rect 8611 6952 8620 6992
rect 8660 6952 9100 6992
rect 9140 6952 9149 6992
rect 11587 6952 11596 6992
rect 11636 6952 12940 6992
rect 12980 6952 13612 6992
rect 13652 6952 13661 6992
rect 21379 6952 21388 6992
rect 21428 6952 21772 6992
rect 21812 6952 23308 6992
rect 23348 6952 23357 6992
rect 23491 6952 23500 6992
rect 23540 6952 23549 6992
rect 23779 6952 23788 6992
rect 23828 6952 24268 6992
rect 24308 6952 24317 6992
rect 28195 6952 28204 6992
rect 28244 6952 28492 6992
rect 28532 6952 28541 6992
rect 8419 6868 8428 6908
rect 8468 6868 9428 6908
rect 11299 6868 11308 6908
rect 11348 6868 11884 6908
rect 11924 6868 11933 6908
rect 25027 6868 25036 6908
rect 25076 6868 26516 6908
rect 26659 6868 26668 6908
rect 26708 6868 33100 6908
rect 33140 6868 33149 6908
rect 9388 6824 9428 6868
rect 26476 6824 26516 6868
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 6307 6784 6316 6824
rect 6356 6784 7756 6824
rect 7796 6784 8716 6824
rect 8756 6784 8765 6824
rect 9379 6784 9388 6824
rect 9428 6784 9437 6824
rect 10051 6784 10060 6824
rect 10100 6784 13804 6824
rect 13844 6784 13853 6824
rect 15427 6784 15436 6824
rect 15476 6784 16108 6824
rect 16148 6784 16157 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 23395 6784 23404 6824
rect 23444 6784 26188 6824
rect 26228 6784 26237 6824
rect 26467 6784 26476 6824
rect 26516 6784 27340 6824
rect 27380 6784 27389 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 23779 6740 23837 6741
rect 8323 6700 8332 6740
rect 8372 6700 9772 6740
rect 9812 6700 9821 6740
rect 9955 6700 9964 6740
rect 10004 6700 11788 6740
rect 11828 6700 11837 6740
rect 14563 6700 14572 6740
rect 14612 6700 15052 6740
rect 15092 6700 17740 6740
rect 17780 6700 17789 6740
rect 23107 6700 23116 6740
rect 23156 6700 23788 6740
rect 23828 6700 26572 6740
rect 26612 6700 26621 6740
rect 23779 6699 23837 6700
rect 8419 6616 8428 6656
rect 8468 6616 8812 6656
rect 8852 6616 8861 6656
rect 9475 6616 9484 6656
rect 9524 6616 9868 6656
rect 9908 6616 9917 6656
rect 10339 6616 10348 6656
rect 10388 6616 10397 6656
rect 13603 6616 13612 6656
rect 13652 6616 14476 6656
rect 14516 6616 14525 6656
rect 15331 6616 15340 6656
rect 15380 6616 15628 6656
rect 15668 6616 15677 6656
rect 23875 6616 23884 6656
rect 23924 6616 26764 6656
rect 26804 6616 26813 6656
rect 35299 6616 35308 6656
rect 35348 6616 36172 6656
rect 36212 6616 36221 6656
rect 10348 6572 10388 6616
rect 6211 6532 6220 6572
rect 6260 6532 9292 6572
rect 9332 6532 9772 6572
rect 9812 6532 10388 6572
rect 15715 6532 15724 6572
rect 15764 6532 16300 6572
rect 16340 6532 16349 6572
rect 22723 6532 22732 6572
rect 22772 6532 23692 6572
rect 23732 6532 23741 6572
rect 26563 6532 26572 6572
rect 26612 6532 27092 6572
rect 29059 6532 29068 6572
rect 29108 6532 29452 6572
rect 29492 6532 31852 6572
rect 31892 6532 31901 6572
rect 0 6488 80 6508
rect 6412 6488 6452 6532
rect 27052 6488 27092 6532
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 3715 6448 3724 6488
rect 3764 6448 4876 6488
rect 4916 6448 4925 6488
rect 6403 6448 6412 6488
rect 6452 6448 6492 6488
rect 7843 6448 7852 6488
rect 7892 6448 8524 6488
rect 8564 6448 9004 6488
rect 9044 6448 9053 6488
rect 9475 6448 9484 6488
rect 9524 6448 10540 6488
rect 10580 6448 10589 6488
rect 12067 6448 12076 6488
rect 12116 6448 12844 6488
rect 12884 6448 12893 6488
rect 14184 6448 14193 6488
rect 14233 6448 14380 6488
rect 14420 6448 14429 6488
rect 18115 6448 18124 6488
rect 18164 6448 19372 6488
rect 19412 6448 19564 6488
rect 19604 6448 19613 6488
rect 21571 6448 21580 6488
rect 21620 6448 22444 6488
rect 22484 6448 23212 6488
rect 23252 6448 23261 6488
rect 23587 6448 23596 6488
rect 23636 6448 24076 6488
rect 24116 6448 24268 6488
rect 24308 6448 24317 6488
rect 25219 6448 25228 6488
rect 25268 6448 26668 6488
rect 26708 6448 26717 6488
rect 27043 6448 27052 6488
rect 27092 6448 27101 6488
rect 28771 6448 28780 6488
rect 28820 6448 29164 6488
rect 29204 6448 29213 6488
rect 29731 6448 29740 6488
rect 29780 6448 29789 6488
rect 31555 6448 31564 6488
rect 31604 6448 32044 6488
rect 32084 6448 32093 6488
rect 33859 6448 33868 6488
rect 33908 6448 34636 6488
rect 34676 6448 34685 6488
rect 0 6428 80 6448
rect 25219 6404 25277 6405
rect 29740 6404 29780 6448
rect 5635 6364 5644 6404
rect 5684 6364 5836 6404
rect 5876 6364 7564 6404
rect 7604 6364 10004 6404
rect 9964 6320 10004 6364
rect 25219 6364 25228 6404
rect 25268 6364 25420 6404
rect 25460 6364 26284 6404
rect 26324 6364 26333 6404
rect 28291 6364 28300 6404
rect 28340 6364 28972 6404
rect 29012 6364 29780 6404
rect 25219 6363 25277 6364
rect 24931 6320 24989 6321
rect 6019 6280 6028 6320
rect 6068 6280 7084 6320
rect 7124 6280 7660 6320
rect 7700 6280 7709 6320
rect 7756 6280 8236 6320
rect 8276 6280 8908 6320
rect 8948 6280 9196 6320
rect 9236 6280 9868 6320
rect 9908 6280 9917 6320
rect 9964 6280 10348 6320
rect 10388 6280 10397 6320
rect 13795 6280 13804 6320
rect 13844 6280 14668 6320
rect 14708 6280 14717 6320
rect 16291 6280 16300 6320
rect 16340 6280 16876 6320
rect 16916 6280 16925 6320
rect 18403 6280 18412 6320
rect 18452 6280 18461 6320
rect 22243 6280 22252 6320
rect 22292 6280 22924 6320
rect 22964 6280 22973 6320
rect 24846 6280 24940 6320
rect 24980 6280 24989 6320
rect 7756 6236 7796 6280
rect 7363 6196 7372 6236
rect 7412 6196 7796 6236
rect 7939 6196 7948 6236
rect 7988 6196 10636 6236
rect 10676 6196 10685 6236
rect 18412 6152 18452 6280
rect 24931 6279 24989 6280
rect 25996 6280 26476 6320
rect 26516 6280 26525 6320
rect 26659 6280 26668 6320
rect 26708 6280 28204 6320
rect 28244 6280 28253 6320
rect 25996 6236 26036 6280
rect 25987 6196 25996 6236
rect 26036 6196 26045 6236
rect 29251 6196 29260 6236
rect 29300 6196 30028 6236
rect 30068 6196 30077 6236
rect 11683 6112 11692 6152
rect 11732 6112 14764 6152
rect 14804 6112 14813 6152
rect 18115 6112 18124 6152
rect 18164 6112 18452 6152
rect 24835 6112 24844 6152
rect 24884 6112 25612 6152
rect 25652 6112 26956 6152
rect 26996 6112 27005 6152
rect 25132 6068 25172 6112
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 11107 6028 11116 6068
rect 11156 6028 12364 6068
rect 12404 6028 13036 6068
rect 13076 6028 13085 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 25123 6028 25132 6068
rect 25172 6028 25181 6068
rect 29347 6028 29356 6068
rect 29396 6028 29436 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 29356 5984 29396 6028
rect 11203 5944 11212 5984
rect 11252 5944 13516 5984
rect 13556 5944 13565 5984
rect 27619 5944 27628 5984
rect 27668 5944 31124 5984
rect 11779 5900 11837 5901
rect 31084 5900 31124 5944
rect 6211 5860 6220 5900
rect 6260 5860 11596 5900
rect 11636 5860 11645 5900
rect 11779 5860 11788 5900
rect 11828 5860 12556 5900
rect 12596 5860 12605 5900
rect 25315 5860 25324 5900
rect 25364 5860 25612 5900
rect 25652 5860 25661 5900
rect 31075 5860 31084 5900
rect 31124 5860 31133 5900
rect 11779 5859 11837 5860
rect 4675 5776 4684 5816
rect 4724 5776 5548 5816
rect 5588 5776 5597 5816
rect 10723 5776 10732 5816
rect 10772 5776 14380 5816
rect 14420 5776 14429 5816
rect 15619 5776 15628 5816
rect 15668 5776 16396 5816
rect 16436 5776 16445 5816
rect 24931 5776 24940 5816
rect 24980 5776 25708 5816
rect 25748 5776 25757 5816
rect 15715 5732 15773 5733
rect 5827 5692 5836 5732
rect 5876 5692 7948 5732
rect 7988 5692 7997 5732
rect 10051 5692 10060 5732
rect 10100 5692 10828 5732
rect 10868 5692 10877 5732
rect 11395 5692 11404 5732
rect 11444 5692 11692 5732
rect 11732 5692 11741 5732
rect 11875 5692 11884 5732
rect 11924 5692 12268 5732
rect 12308 5692 12317 5732
rect 15630 5692 15724 5732
rect 15764 5692 15773 5732
rect 33955 5692 33964 5732
rect 34004 5692 34732 5732
rect 34772 5692 35020 5732
rect 35060 5692 35069 5732
rect 15715 5691 15773 5692
rect 0 5648 80 5668
rect 11491 5648 11549 5649
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 4579 5608 4588 5648
rect 4628 5608 6124 5648
rect 6164 5608 6173 5648
rect 8419 5608 8428 5648
rect 8468 5608 10444 5648
rect 10484 5608 10493 5648
rect 10723 5608 10732 5648
rect 10772 5608 11360 5648
rect 0 5588 80 5608
rect 11320 5564 11360 5608
rect 11491 5608 11500 5648
rect 11540 5608 12172 5648
rect 12212 5608 12221 5648
rect 13411 5608 13420 5648
rect 13460 5608 14860 5648
rect 14900 5608 14909 5648
rect 15043 5608 15052 5648
rect 15092 5608 17932 5648
rect 17972 5608 17981 5648
rect 18115 5608 18124 5648
rect 18164 5608 19180 5648
rect 19220 5608 20236 5648
rect 20276 5608 21868 5648
rect 21908 5608 22156 5648
rect 22196 5608 22205 5648
rect 23299 5608 23308 5648
rect 23348 5608 24268 5648
rect 24308 5608 25132 5648
rect 25172 5608 25420 5648
rect 25460 5608 25469 5648
rect 30883 5608 30892 5648
rect 30932 5608 31564 5648
rect 31604 5608 31613 5648
rect 33187 5608 33196 5648
rect 33236 5608 35308 5648
rect 35348 5608 35357 5648
rect 11491 5607 11549 5608
rect 34435 5564 34493 5565
rect 11320 5524 12748 5564
rect 12788 5524 12797 5564
rect 13603 5524 13612 5564
rect 13652 5524 14956 5564
rect 14996 5524 15005 5564
rect 25996 5524 34060 5564
rect 34100 5524 34444 5564
rect 34484 5524 34636 5564
rect 34676 5524 34685 5564
rect 4387 5440 4396 5480
rect 4436 5440 4445 5480
rect 4675 5440 4684 5480
rect 4724 5440 6412 5480
rect 6452 5440 7180 5480
rect 7220 5440 7468 5480
rect 7508 5440 7517 5480
rect 11299 5440 11308 5480
rect 11348 5440 12460 5480
rect 12500 5440 13132 5480
rect 13172 5440 13181 5480
rect 4396 5396 4436 5440
rect 13612 5396 13652 5524
rect 25027 5480 25085 5481
rect 14179 5440 14188 5480
rect 14228 5440 15532 5480
rect 15572 5440 16204 5480
rect 16244 5440 16253 5480
rect 25027 5440 25036 5480
rect 25076 5440 25324 5480
rect 25364 5440 25373 5480
rect 25027 5439 25085 5440
rect 15331 5396 15389 5397
rect 25996 5396 26036 5524
rect 34435 5523 34493 5524
rect 27811 5440 27820 5480
rect 27860 5440 28684 5480
rect 28724 5440 30220 5480
rect 30260 5440 30269 5480
rect 33475 5440 33484 5480
rect 33524 5440 34444 5480
rect 34484 5440 34924 5480
rect 34964 5440 34973 5480
rect 4195 5356 4204 5396
rect 4244 5356 5740 5396
rect 5780 5356 6124 5396
rect 6164 5356 6173 5396
rect 11107 5356 11116 5396
rect 11156 5356 11404 5396
rect 11444 5356 11453 5396
rect 11587 5356 11596 5396
rect 11636 5356 13652 5396
rect 13987 5356 13996 5396
rect 14036 5356 14764 5396
rect 14804 5356 14813 5396
rect 15246 5356 15340 5396
rect 15380 5356 15389 5396
rect 20323 5356 20332 5396
rect 20372 5356 21484 5396
rect 21524 5356 26036 5396
rect 27043 5356 27052 5396
rect 27092 5356 27340 5396
rect 27380 5356 27389 5396
rect 15331 5355 15389 5356
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 11491 5272 11500 5312
rect 11540 5272 11692 5312
rect 11732 5272 11741 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 9571 5104 9580 5144
rect 9620 5104 11788 5144
rect 11828 5104 11837 5144
rect 13795 5104 13804 5144
rect 13844 5104 14284 5144
rect 14324 5104 14333 5144
rect 25603 5104 25612 5144
rect 25652 5104 25900 5144
rect 25940 5104 25949 5144
rect 26371 5104 26380 5144
rect 26420 5104 27052 5144
rect 27092 5104 27340 5144
rect 27380 5104 27389 5144
rect 27907 5104 27916 5144
rect 27956 5104 27965 5144
rect 28579 5104 28588 5144
rect 28628 5104 28637 5144
rect 27916 5060 27956 5104
rect 28588 5060 28628 5104
rect 5923 5020 5932 5060
rect 5972 5020 6796 5060
rect 6836 5020 6845 5060
rect 7171 5020 7180 5060
rect 7220 5020 7756 5060
rect 7796 5020 9676 5060
rect 9716 5020 9725 5060
rect 10339 5020 10348 5060
rect 10388 5020 11116 5060
rect 11156 5020 11165 5060
rect 11491 5020 11500 5060
rect 11540 5020 11884 5060
rect 11924 5020 11933 5060
rect 14467 5020 14476 5060
rect 14516 5020 14956 5060
rect 14996 5020 15005 5060
rect 15523 5020 15532 5060
rect 15572 5020 16108 5060
rect 16148 5020 17740 5060
rect 17780 5020 17789 5060
rect 22339 5020 22348 5060
rect 22388 5020 22732 5060
rect 22772 5020 23212 5060
rect 23252 5020 23261 5060
rect 25699 5020 25708 5060
rect 25748 5020 26284 5060
rect 26324 5020 26333 5060
rect 27427 5020 27436 5060
rect 27476 5020 27820 5060
rect 27860 5020 27869 5060
rect 27916 5020 28628 5060
rect 26083 4976 26141 4977
rect 4387 4936 4396 4976
rect 4436 4936 6220 4976
rect 6260 4936 6269 4976
rect 9955 4936 9964 4976
rect 10004 4936 11020 4976
rect 11060 4936 11308 4976
rect 11348 4936 11357 4976
rect 12355 4936 12364 4976
rect 12404 4936 12940 4976
rect 12980 4936 12989 4976
rect 13123 4936 13132 4976
rect 13172 4936 13181 4976
rect 14083 4936 14092 4976
rect 14132 4936 16012 4976
rect 16052 4936 16396 4976
rect 16436 4936 16445 4976
rect 21955 4936 21964 4976
rect 22004 4936 23020 4976
rect 23060 4936 23692 4976
rect 23732 4936 23741 4976
rect 25998 4936 26092 4976
rect 26132 4936 26141 4976
rect 26659 4936 26668 4976
rect 26708 4936 26956 4976
rect 26996 4936 27340 4976
rect 27380 4936 27389 4976
rect 27523 4936 27532 4976
rect 27572 4936 29068 4976
rect 29108 4936 29117 4976
rect 0 4808 80 4828
rect 13132 4808 13172 4936
rect 26083 4935 26141 4936
rect 13987 4852 13996 4892
rect 14036 4852 14572 4892
rect 14612 4852 14621 4892
rect 22147 4852 22156 4892
rect 22196 4852 23596 4892
rect 23636 4852 23645 4892
rect 27235 4852 27244 4892
rect 27284 4852 28204 4892
rect 28244 4852 30220 4892
rect 30260 4852 30269 4892
rect 23779 4808 23837 4809
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 4483 4768 4492 4808
rect 4532 4768 5356 4808
rect 5396 4768 5405 4808
rect 11683 4768 11692 4808
rect 11732 4768 13172 4808
rect 14755 4768 14764 4808
rect 14804 4768 15148 4808
rect 15188 4768 15436 4808
rect 15476 4768 15820 4808
rect 15860 4768 15869 4808
rect 18403 4768 18412 4808
rect 18452 4768 19372 4808
rect 19412 4768 19421 4808
rect 21475 4768 21484 4808
rect 21524 4768 22060 4808
rect 22100 4768 23788 4808
rect 23828 4768 23837 4808
rect 27139 4768 27148 4808
rect 27188 4768 27628 4808
rect 27668 4768 28012 4808
rect 28052 4768 28061 4808
rect 0 4748 80 4768
rect 23779 4767 23837 4768
rect 15715 4724 15773 4725
rect 14179 4684 14188 4724
rect 14228 4684 15724 4724
rect 15764 4684 15773 4724
rect 18019 4684 18028 4724
rect 18068 4684 18892 4724
rect 18932 4684 20428 4724
rect 20468 4684 22156 4724
rect 22196 4684 22205 4724
rect 15715 4683 15773 4684
rect 15331 4640 15389 4641
rect 11971 4600 11980 4640
rect 12020 4600 13324 4640
rect 13364 4600 15340 4640
rect 15380 4600 15389 4640
rect 25315 4600 25324 4640
rect 25364 4600 29548 4640
rect 29588 4600 29740 4640
rect 29780 4600 29789 4640
rect 15331 4599 15389 4600
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 4579 4348 4588 4388
rect 4628 4348 7564 4388
rect 7604 4348 7613 4388
rect 11203 4348 11212 4388
rect 11252 4348 11884 4388
rect 11924 4348 13420 4388
rect 13460 4348 13469 4388
rect 7363 4264 7372 4304
rect 7412 4264 7852 4304
rect 7892 4264 7901 4304
rect 8515 4264 8524 4304
rect 8564 4264 9388 4304
rect 9428 4264 9437 4304
rect 10627 4264 10636 4304
rect 10676 4264 11404 4304
rect 11444 4264 12460 4304
rect 12500 4264 12509 4304
rect 14563 4264 14572 4304
rect 14612 4264 15244 4304
rect 15284 4264 15293 4304
rect 26179 4264 26188 4304
rect 26228 4264 26237 4304
rect 23779 4220 23837 4221
rect 26188 4220 26228 4264
rect 3331 4180 3340 4220
rect 3380 4180 4684 4220
rect 4724 4180 4733 4220
rect 5827 4180 5836 4220
rect 5876 4180 6124 4220
rect 6164 4180 6173 4220
rect 6307 4180 6316 4220
rect 6356 4180 6988 4220
rect 7028 4180 7037 4220
rect 23694 4180 23788 4220
rect 23828 4180 23837 4220
rect 23779 4179 23837 4180
rect 25612 4180 26228 4220
rect 4579 4096 4588 4136
rect 4628 4096 4972 4136
rect 5012 4096 6700 4136
rect 6740 4096 6749 4136
rect 7075 4096 7084 4136
rect 7124 4096 7276 4136
rect 7316 4096 8140 4136
rect 8180 4096 8189 4136
rect 9667 4096 9676 4136
rect 9716 4096 10252 4136
rect 10292 4096 10301 4136
rect 11011 4096 11020 4136
rect 11060 4096 11788 4136
rect 11828 4096 11837 4136
rect 14371 4096 14380 4136
rect 14420 4096 14764 4136
rect 14804 4096 14813 4136
rect 16099 4096 16108 4136
rect 16148 4096 16300 4136
rect 16340 4096 16349 4136
rect 19747 4096 19756 4136
rect 19796 4096 20044 4136
rect 20084 4096 20093 4136
rect 20707 4096 20716 4136
rect 20756 4096 21676 4136
rect 21716 4096 21725 4136
rect 22147 4096 22156 4136
rect 22196 4096 24844 4136
rect 24884 4096 24893 4136
rect 7276 4052 7316 4096
rect 25612 4052 25652 4180
rect 25699 4136 25757 4137
rect 25699 4096 25708 4136
rect 25748 4096 25842 4136
rect 26179 4096 26188 4136
rect 26228 4096 26668 4136
rect 26708 4096 26717 4136
rect 27331 4096 27340 4136
rect 27380 4096 28204 4136
rect 28244 4096 28253 4136
rect 28771 4096 28780 4136
rect 28820 4096 29260 4136
rect 29300 4096 29309 4136
rect 29731 4096 29740 4136
rect 29780 4096 30508 4136
rect 30548 4096 30557 4136
rect 31363 4096 31372 4136
rect 31412 4096 32332 4136
rect 32372 4096 32381 4136
rect 25699 4095 25757 4096
rect 6499 4012 6508 4052
rect 6548 4012 7316 4052
rect 9955 4012 9964 4052
rect 10004 4012 10540 4052
rect 10580 4012 10589 4052
rect 19843 4012 19852 4052
rect 19892 4012 20332 4052
rect 20372 4012 23924 4052
rect 25603 4012 25612 4052
rect 25652 4012 25661 4052
rect 26083 4012 26092 4052
rect 26132 4012 27284 4052
rect 0 3968 80 3988
rect 23884 3968 23924 4012
rect 27244 3968 27284 4012
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 9667 3928 9676 3968
rect 9716 3928 10636 3968
rect 10676 3928 10685 3968
rect 14275 3928 14284 3968
rect 14324 3928 15916 3968
rect 15956 3928 15965 3968
rect 19555 3928 19564 3968
rect 19604 3928 20180 3968
rect 23875 3928 23884 3968
rect 23924 3928 25996 3968
rect 26036 3928 26045 3968
rect 27235 3928 27244 3968
rect 27284 3928 27916 3968
rect 27956 3928 27965 3968
rect 0 3908 80 3928
rect 20140 3884 20180 3928
rect 25219 3884 25277 3885
rect 20140 3844 20716 3884
rect 20756 3844 20765 3884
rect 23587 3844 23596 3884
rect 23636 3844 25228 3884
rect 25268 3844 25277 3884
rect 26563 3844 26572 3884
rect 26612 3844 28396 3884
rect 28436 3844 28445 3884
rect 25219 3843 25277 3844
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 7651 3760 7660 3800
rect 7700 3760 7948 3800
rect 7988 3760 9196 3800
rect 9236 3760 9245 3800
rect 10819 3760 10828 3800
rect 10868 3760 11308 3800
rect 11348 3760 11884 3800
rect 11924 3760 13420 3800
rect 13460 3760 13469 3800
rect 14860 3760 15724 3800
rect 15764 3760 15773 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 20995 3760 21004 3800
rect 21044 3760 21292 3800
rect 21332 3760 22060 3800
rect 22100 3760 22109 3800
rect 25507 3760 25516 3800
rect 25556 3760 26476 3800
rect 26516 3760 26525 3800
rect 26851 3760 26860 3800
rect 26900 3760 27628 3800
rect 27668 3760 27677 3800
rect 28291 3760 28300 3800
rect 28340 3760 29164 3800
rect 29204 3760 29213 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 14860 3716 14900 3760
rect 9379 3676 9388 3716
rect 9428 3676 10444 3716
rect 10484 3676 14516 3716
rect 14851 3676 14860 3716
rect 14900 3676 14909 3716
rect 25123 3676 25132 3716
rect 25172 3676 25804 3716
rect 25844 3676 26764 3716
rect 26804 3676 26813 3716
rect 14476 3632 14516 3676
rect 9091 3592 9100 3632
rect 9140 3592 9580 3632
rect 9620 3592 11404 3632
rect 11444 3592 11453 3632
rect 14467 3592 14476 3632
rect 14516 3592 14525 3632
rect 14755 3508 14764 3548
rect 14804 3508 16588 3548
rect 16628 3508 16637 3548
rect 15331 3464 15389 3465
rect 9283 3424 9292 3464
rect 9332 3424 9484 3464
rect 9524 3424 9533 3464
rect 11299 3424 11308 3464
rect 11348 3424 12268 3464
rect 12308 3424 12317 3464
rect 15331 3424 15340 3464
rect 15380 3424 15436 3464
rect 15476 3424 15485 3464
rect 15811 3424 15820 3464
rect 15860 3424 16300 3464
rect 16340 3424 16349 3464
rect 26659 3424 26668 3464
rect 26708 3424 28492 3464
rect 28532 3424 28541 3464
rect 28675 3424 28684 3464
rect 28724 3424 30412 3464
rect 30452 3424 30461 3464
rect 15331 3423 15389 3424
rect 11779 3380 11837 3381
rect 7843 3340 7852 3380
rect 7892 3340 8716 3380
rect 8756 3340 8765 3380
rect 11779 3340 11788 3380
rect 11828 3340 12076 3380
rect 12116 3340 13132 3380
rect 13172 3340 13181 3380
rect 15235 3340 15244 3380
rect 15284 3340 16396 3380
rect 16436 3340 16445 3380
rect 25411 3340 25420 3380
rect 25460 3340 25708 3380
rect 25748 3340 26380 3380
rect 26420 3340 26429 3380
rect 11779 3339 11837 3340
rect 15619 3256 15628 3296
rect 15668 3256 16684 3296
rect 16724 3256 16733 3296
rect 11491 3172 11500 3212
rect 11540 3172 12460 3212
rect 12500 3172 15724 3212
rect 15764 3172 15773 3212
rect 20227 3172 20236 3212
rect 20276 3172 23980 3212
rect 24020 3172 27052 3212
rect 27092 3172 27101 3212
rect 0 3128 80 3148
rect 15715 3128 15773 3129
rect 0 3088 652 3128
rect 692 3088 701 3128
rect 15715 3088 15724 3128
rect 15764 3088 16492 3128
rect 16532 3088 16541 3128
rect 0 3068 80 3088
rect 15715 3087 15773 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 15427 3004 15436 3044
rect 15476 3004 16108 3044
rect 16148 3004 16157 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 29347 3004 29356 3044
rect 29396 3004 29836 3044
rect 29876 3004 29885 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 16387 2836 16396 2876
rect 16436 2836 16876 2876
rect 16916 2836 16925 2876
rect 22051 2836 22060 2876
rect 22100 2836 23980 2876
rect 24020 2836 25228 2876
rect 25268 2836 25277 2876
rect 25795 2836 25804 2876
rect 25844 2836 26572 2876
rect 26612 2836 26621 2876
rect 28291 2836 28300 2876
rect 28340 2836 29452 2876
rect 29492 2836 29836 2876
rect 29876 2836 29885 2876
rect 5827 2752 5836 2792
rect 5876 2752 6892 2792
rect 6932 2752 6941 2792
rect 8227 2752 8236 2792
rect 8276 2752 9100 2792
rect 9140 2752 9149 2792
rect 16003 2752 16012 2792
rect 16052 2752 16204 2792
rect 16244 2752 16253 2792
rect 23308 2752 24172 2792
rect 24212 2752 24221 2792
rect 23308 2708 23348 2752
rect 5443 2668 5452 2708
rect 5492 2668 6124 2708
rect 6164 2668 6173 2708
rect 16291 2668 16300 2708
rect 16340 2668 16972 2708
rect 17012 2668 17836 2708
rect 17876 2668 17885 2708
rect 18019 2668 18028 2708
rect 18068 2668 18077 2708
rect 21955 2668 21964 2708
rect 22004 2668 23308 2708
rect 23348 2668 23357 2708
rect 23587 2668 23596 2708
rect 23636 2668 24556 2708
rect 24596 2668 24605 2708
rect 18028 2624 18068 2668
rect 25219 2624 25277 2625
rect 8035 2584 8044 2624
rect 8084 2584 8428 2624
rect 8468 2584 8477 2624
rect 14083 2584 14092 2624
rect 14132 2584 16012 2624
rect 16052 2584 18068 2624
rect 18691 2584 18700 2624
rect 18740 2584 19180 2624
rect 19220 2584 19229 2624
rect 21859 2584 21868 2624
rect 21908 2584 23116 2624
rect 23156 2584 24460 2624
rect 24500 2584 24509 2624
rect 25219 2584 25228 2624
rect 25268 2584 25420 2624
rect 25460 2584 25469 2624
rect 26275 2584 26284 2624
rect 26324 2584 27244 2624
rect 27284 2584 28780 2624
rect 28820 2584 28829 2624
rect 30883 2584 30892 2624
rect 30932 2584 31852 2624
rect 31892 2584 31901 2624
rect 25219 2583 25277 2584
rect 8131 2416 8140 2456
rect 8180 2416 9292 2456
rect 9332 2416 9676 2456
rect 9716 2416 9725 2456
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 0 2228 80 2248
rect 20035 2080 20044 2120
rect 20084 2080 20812 2120
rect 20852 2080 20861 2120
rect 23920 1996 23980 2036
rect 24020 1996 26668 2036
rect 26708 1996 27724 2036
rect 27764 1996 27773 2036
rect 23920 1952 23960 1996
rect 9475 1912 9484 1952
rect 9524 1912 10732 1952
rect 10772 1912 10781 1952
rect 20995 1912 21004 1952
rect 21044 1912 22252 1952
rect 22292 1912 22301 1952
rect 22531 1912 22540 1952
rect 22580 1912 23960 1952
rect 27523 1912 27532 1952
rect 27572 1912 28684 1952
rect 28724 1912 28733 1952
rect 9955 1744 9964 1784
rect 10004 1744 10540 1784
rect 10580 1744 10589 1784
rect 835 1660 844 1700
rect 884 1660 17452 1700
rect 17492 1660 17501 1700
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 9763 1240 9772 1280
rect 9812 1240 10156 1280
rect 10196 1240 10205 1280
rect 25699 1112 25757 1113
rect 23971 1072 23980 1112
rect 24020 1072 25516 1112
rect 25556 1072 25708 1112
rect 25748 1072 25757 1112
rect 25699 1071 25757 1072
rect 25603 904 25612 944
rect 25652 904 25996 944
rect 26036 904 26476 944
rect 26516 904 26525 944
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 76 36688 116 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 28492 34000 28532 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 4780 32152 4820 32192
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 13132 31564 13172 31604
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 4780 30472 4820 30512
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 13132 29884 13172 29924
rect 5644 29800 5684 29840
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 14092 29128 14132 29168
rect 20236 29128 20276 29168
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 5644 28288 5684 28328
rect 20236 28288 20276 28328
rect 20620 28120 20660 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 31180 27868 31220 27908
rect 28492 27616 28532 27656
rect 20620 27532 20660 27572
rect 28588 27532 28628 27572
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 13036 26440 13076 26480
rect 14092 26440 14132 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 31180 26356 31220 26396
rect 47596 26356 47636 26396
rect 19180 26272 19220 26312
rect 39148 26188 39188 26228
rect 25996 26104 26036 26144
rect 29836 26104 29876 26144
rect 47596 26104 47636 26144
rect 30604 25852 30644 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 13036 25684 13076 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 25516 25516 25556 25556
rect 41260 25516 41300 25556
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 19180 24508 19220 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 24460 24172 24500 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 19180 24004 19220 24044
rect 25324 23752 25364 23792
rect 25708 23752 25748 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 24364 23500 24404 23540
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 28204 23332 28244 23372
rect 25132 23248 25172 23288
rect 25420 23248 25460 23288
rect 24460 23080 24500 23120
rect 25132 22996 25172 23036
rect 35500 22828 35540 22868
rect 24748 22744 24788 22784
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 25324 22576 25364 22616
rect 25516 22576 25556 22616
rect 24748 22408 24788 22448
rect 25708 21988 25748 22028
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 25420 21904 25460 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 24364 21652 24404 21692
rect 35212 21568 35252 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 16684 20056 16724 20096
rect 31948 20056 31988 20096
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4204 19300 4244 19340
rect 28588 19300 28628 19340
rect 26668 19216 26708 19256
rect 32428 19132 32468 19172
rect 18700 19048 18740 19088
rect 34252 19048 34292 19088
rect 25708 18964 25748 19004
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 23116 18880 23156 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 34252 18460 34292 18500
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 23788 18040 23828 18080
rect 24076 17956 24116 17996
rect 34444 17704 34484 17744
rect 23116 17620 23156 17660
rect 26188 17620 26228 17660
rect 4204 17536 4244 17576
rect 23788 17536 23828 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 36556 17284 36596 17324
rect 24076 17200 24116 17240
rect 37324 17200 37364 17240
rect 21580 16780 21620 16820
rect 32044 16696 32084 16736
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 18988 16444 19028 16484
rect 31564 16444 31604 16484
rect 36556 16444 36596 16484
rect 32428 16360 32468 16400
rect 20140 16192 20180 16232
rect 21196 16192 21236 16232
rect 24268 16192 24308 16232
rect 37324 16108 37364 16148
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 15436 15856 15476 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 24460 15856 24500 15896
rect 32428 16024 32468 16064
rect 37708 16024 37748 16064
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 20236 15772 20276 15812
rect 21676 15688 21716 15728
rect 31564 15604 31604 15644
rect 37132 15604 37172 15644
rect 27724 15520 27764 15560
rect 32044 15352 32084 15392
rect 37708 15436 37748 15476
rect 32524 15268 32564 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 20812 15100 20852 15140
rect 24268 15100 24308 15140
rect 25708 15100 25748 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 5932 15016 5972 15056
rect 17644 15016 17684 15056
rect 20140 15016 20180 15056
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 27724 15016 27764 15056
rect 18796 14932 18836 14972
rect 31948 14932 31988 14972
rect 37132 14932 37172 14972
rect 19948 14848 19988 14888
rect 20236 14764 20276 14804
rect 21676 14596 21716 14636
rect 32044 14512 32084 14552
rect 32620 14512 32660 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 18796 14176 18836 14216
rect 20044 14176 20084 14216
rect 29932 14176 29972 14216
rect 19180 14092 19220 14132
rect 26188 14092 26228 14132
rect 14956 14008 14996 14048
rect 31948 14008 31988 14048
rect 15244 13924 15284 13964
rect 19948 13924 19988 13964
rect 28204 13924 28244 13964
rect 20044 13840 20084 13880
rect 28972 13756 29012 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 18028 13504 18068 13544
rect 26764 13504 26804 13544
rect 15340 13336 15380 13376
rect 19180 13336 19220 13376
rect 21580 13420 21614 13460
rect 21614 13420 21620 13460
rect 28012 13336 28052 13376
rect 20044 13252 20084 13292
rect 17740 13168 17780 13208
rect 18028 13168 18068 13208
rect 28012 13168 28052 13208
rect 28204 13084 28244 13124
rect 19852 13000 19892 13040
rect 14956 12916 14996 12956
rect 15724 12916 15764 12956
rect 29740 12916 29780 12956
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 15628 12832 15668 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 28972 12832 29012 12872
rect 26668 12748 26708 12788
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 5932 12496 5972 12536
rect 20812 12496 20852 12536
rect 15724 12412 15764 12452
rect 18796 12412 18836 12452
rect 18988 12412 19028 12452
rect 19756 12412 19796 12452
rect 25996 12412 26036 12452
rect 15628 12328 15668 12368
rect 11788 12244 11828 12284
rect 14956 12244 14996 12284
rect 18892 12244 18932 12284
rect 19756 12244 19796 12284
rect 20044 12244 20084 12284
rect 34444 12160 34484 12200
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 19948 12076 19988 12116
rect 20140 12076 20180 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 26668 11992 26708 12032
rect 26764 11908 26804 11948
rect 17932 11824 17972 11864
rect 35020 11824 35060 11864
rect 21580 11740 21620 11780
rect 29740 11740 29780 11780
rect 26092 11656 26132 11696
rect 17932 11572 17972 11612
rect 15244 11488 15284 11528
rect 16108 11488 16148 11528
rect 15436 11404 15476 11444
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 15340 11320 15380 11360
rect 16396 11320 16436 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 29932 11320 29972 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 25996 11152 26036 11192
rect 35020 11152 35060 11192
rect 15724 11068 15764 11108
rect 32524 10984 32564 11024
rect 15916 10900 15956 10940
rect 18700 10900 18740 10940
rect 26668 10900 26708 10940
rect 17740 10816 17780 10856
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33100 10564 33140 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 16108 10312 16148 10352
rect 32524 10228 32564 10268
rect 18028 9892 18068 9932
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 15724 9808 15764 9848
rect 16204 9808 16244 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 14956 9640 14996 9680
rect 34828 9556 34868 9596
rect 31852 9472 31892 9512
rect 32620 9472 32660 9512
rect 33100 9472 33140 9512
rect 34828 9388 34868 9428
rect 15916 9304 15956 9344
rect 33868 9304 33908 9344
rect 16204 9136 16244 9176
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 34060 9052 34100 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 18796 8800 18836 8840
rect 25036 8800 25076 8840
rect 27724 8800 27764 8840
rect 31948 8800 31988 8840
rect 33868 8800 33908 8840
rect 34444 8548 34484 8588
rect 14956 8380 14996 8420
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 15724 8296 15764 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 34060 8128 34100 8168
rect 25036 7876 25076 7916
rect 25228 7708 25268 7748
rect 31948 7708 31988 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 30604 7540 30644 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 24556 7204 24596 7244
rect 11500 7120 11540 7160
rect 18892 7120 18932 7160
rect 29260 7120 29300 7160
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 23788 6700 23828 6740
rect 25228 6364 25268 6404
rect 24940 6280 24980 6320
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 11788 5860 11828 5900
rect 15724 5692 15764 5732
rect 11500 5608 11540 5648
rect 34444 5524 34484 5564
rect 25036 5440 25076 5480
rect 15340 5356 15380 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 26092 4936 26132 4976
rect 23788 4768 23828 4808
rect 15724 4684 15764 4724
rect 15340 4600 15380 4640
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 23788 4180 23828 4220
rect 25708 4096 25748 4136
rect 25228 3844 25268 3884
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 15340 3424 15380 3464
rect 11788 3340 11828 3380
rect 15724 3088 15764 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 25228 2584 25268 2624
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 25708 1072 25748 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 76 36728 116 36737
rect 76 19265 116 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 28492 34040 28532 34049
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 4780 32192 4820 32201
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4780 30512 4820 32152
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 4780 30463 4820 30472
rect 13132 31604 13172 31613
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 13132 29924 13172 31564
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 13132 29875 13172 29884
rect 5644 29840 5684 29849
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 5644 28328 5684 29800
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 5644 28279 5684 28288
rect 14092 29168 14132 29177
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 13036 26480 13076 26489
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 13036 25724 13076 26440
rect 14092 26480 14132 29128
rect 20236 29168 20276 29177
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 20236 28328 20276 29128
rect 20236 28279 20276 28288
rect 20620 28160 20660 28169
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 20620 27572 20660 28120
rect 28492 27656 28532 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 28492 27607 28532 27616
rect 31180 27908 31220 27917
rect 20620 27523 20660 27532
rect 28588 27572 28628 27581
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 14092 26431 14132 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 19180 26312 19220 26321
rect 13036 25675 13076 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19180 24548 19220 26272
rect 25995 26144 26037 26153
rect 25995 26104 25996 26144
rect 26036 26104 26037 26144
rect 25995 26095 26037 26104
rect 25996 26010 26036 26095
rect 25516 25556 25556 25565
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 19180 24044 19220 24508
rect 19180 23995 19220 24004
rect 24460 24212 24500 24221
rect 24364 23540 24404 23549
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 24364 21692 24404 23500
rect 24460 23120 24500 24172
rect 25324 23792 25364 23801
rect 24460 23071 24500 23080
rect 25132 23288 25172 23297
rect 25132 23036 25172 23248
rect 25132 22987 25172 22996
rect 24748 22784 24788 22793
rect 24748 22448 24788 22744
rect 25324 22616 25364 23752
rect 25324 22567 25364 22576
rect 25420 23288 25460 23297
rect 24748 22399 24788 22408
rect 25420 21944 25460 23248
rect 25516 22616 25556 25516
rect 25516 22567 25556 22576
rect 25708 23792 25748 23801
rect 25708 22028 25748 23752
rect 28203 23372 28245 23381
rect 28203 23332 28204 23372
rect 28244 23332 28245 23372
rect 28203 23323 28245 23332
rect 28491 23372 28533 23381
rect 28491 23332 28492 23372
rect 28532 23332 28533 23372
rect 28491 23323 28533 23332
rect 28204 23238 28244 23323
rect 25708 21979 25748 21988
rect 25420 21895 25460 21904
rect 24364 21643 24404 21652
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 28492 20180 28532 23323
rect 28588 22877 28628 27532
rect 31180 26396 31220 27868
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 31180 26347 31220 26356
rect 47596 26396 47636 26405
rect 39147 26228 39189 26237
rect 39147 26188 39148 26228
rect 39188 26188 39189 26228
rect 39147 26179 39189 26188
rect 29835 26144 29877 26153
rect 29835 26104 29836 26144
rect 29876 26104 29877 26144
rect 29835 26095 29877 26104
rect 29836 26010 29876 26095
rect 39148 26094 39188 26179
rect 47596 26144 47636 26356
rect 47596 26095 47636 26104
rect 41259 26060 41301 26069
rect 41259 26020 41260 26060
rect 41300 26020 41301 26060
rect 41259 26011 41301 26020
rect 30604 25892 30644 25901
rect 30604 23381 30644 25852
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 41260 25556 41300 26011
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 41260 25507 41300 25516
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 30603 23372 30645 23381
rect 30603 23332 30604 23372
rect 30644 23332 30645 23372
rect 30603 23323 30645 23332
rect 28587 22868 28629 22877
rect 28587 22828 28588 22868
rect 28628 22828 28629 22868
rect 28587 22819 28629 22828
rect 35499 22868 35541 22877
rect 35499 22828 35500 22868
rect 35540 22828 35541 22868
rect 35499 22819 35541 22828
rect 35500 22734 35540 22819
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 35212 21608 35252 21617
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 28492 20140 28628 20180
rect 16683 20096 16725 20105
rect 16683 20056 16684 20096
rect 16724 20056 16725 20096
rect 16683 20047 16725 20056
rect 16684 19962 16724 20047
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 4204 19340 4244 19349
rect 75 19256 117 19265
rect 75 19216 76 19256
rect 116 19216 117 19256
rect 75 19207 117 19216
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4204 17576 4244 19300
rect 28588 19340 28628 20140
rect 35212 20105 35252 21568
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 28588 19291 28628 19300
rect 31948 20096 31988 20105
rect 26667 19256 26709 19265
rect 26667 19216 26668 19256
rect 26708 19216 26709 19256
rect 26667 19207 26709 19216
rect 26668 19122 26708 19207
rect 18700 19088 18740 19097
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 4204 17527 4244 17536
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 15436 15896 15476 15905
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 5932 15056 5972 15065
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 5932 12536 5972 15016
rect 14955 14048 14997 14057
rect 14955 14008 14956 14048
rect 14996 14008 14997 14048
rect 14955 13999 14997 14008
rect 14956 13914 14996 13999
rect 15244 13964 15284 13973
rect 5932 12487 5972 12496
rect 14956 12956 14996 12965
rect 11788 12284 11828 12293
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 11788 11033 11828 12244
rect 14956 12284 14996 12916
rect 14956 12235 14996 12244
rect 15244 11528 15284 13924
rect 15244 11479 15284 11488
rect 15340 13376 15380 13385
rect 15340 11360 15380 13336
rect 15436 12545 15476 15856
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 17644 15056 17684 15065
rect 17644 14057 17684 15016
rect 16395 14048 16437 14057
rect 16395 14008 16396 14048
rect 16436 14008 16437 14048
rect 16395 13999 16437 14008
rect 17643 14048 17685 14057
rect 17643 14008 17644 14048
rect 17684 14008 17685 14048
rect 17643 13999 17685 14008
rect 15724 12956 15764 12965
rect 15628 12872 15668 12881
rect 15435 12536 15477 12545
rect 15435 12496 15436 12536
rect 15476 12496 15477 12536
rect 15435 12487 15477 12496
rect 15436 11444 15476 12487
rect 15628 12368 15668 12832
rect 15724 12452 15764 12916
rect 15724 12403 15764 12412
rect 15628 12319 15668 12328
rect 15436 11395 15476 11404
rect 16108 11528 16148 11537
rect 15340 11311 15380 11320
rect 15724 11108 15764 11117
rect 11787 11024 11829 11033
rect 11787 10984 11788 11024
rect 11828 10984 11829 11024
rect 11787 10975 11829 10984
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 15724 9848 15764 11068
rect 14956 9680 14996 9689
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 14956 8420 14996 9640
rect 14956 8371 14996 8380
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 15724 8336 15764 9808
rect 15916 10940 15956 10949
rect 15916 9344 15956 10900
rect 16108 10352 16148 11488
rect 16396 11360 16436 13999
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18028 13544 18068 13553
rect 16396 11311 16436 11320
rect 17740 13208 17780 13217
rect 17740 10856 17780 13168
rect 18028 13208 18068 13504
rect 17932 11864 17972 11873
rect 17932 11612 17972 11824
rect 17932 11563 17972 11572
rect 17740 10807 17780 10816
rect 16108 10303 16148 10312
rect 18028 9932 18068 13168
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 18700 10940 18740 19048
rect 25708 19004 25748 19013
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 23116 18920 23156 18929
rect 23116 17660 23156 18880
rect 23116 17611 23156 17620
rect 23788 18080 23828 18089
rect 23788 17576 23828 18040
rect 23788 17527 23828 17536
rect 24076 17996 24116 18005
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 24076 17240 24116 17956
rect 24076 17191 24116 17200
rect 21580 16820 21620 16829
rect 18988 16484 19028 16493
rect 18700 10891 18740 10900
rect 18796 14972 18836 14981
rect 18796 14216 18836 14932
rect 18796 12452 18836 14176
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 18028 9883 18068 9892
rect 15916 9295 15956 9304
rect 16204 9848 16244 9857
rect 16204 9176 16244 9808
rect 16204 9127 16244 9136
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 18796 8840 18836 12412
rect 18988 12452 19028 16444
rect 20140 16232 20180 16241
rect 21195 16232 21237 16241
rect 20180 16192 20276 16232
rect 20140 16183 20180 16192
rect 20236 16064 20276 16192
rect 21195 16192 21196 16232
rect 21236 16192 21237 16232
rect 21195 16183 21237 16192
rect 21196 16098 21236 16183
rect 20236 16024 20372 16064
rect 20332 15905 20372 16024
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 20331 15896 20373 15905
rect 20331 15856 20332 15896
rect 20372 15856 20373 15896
rect 20331 15847 20373 15856
rect 20236 15812 20276 15821
rect 20139 15224 20181 15233
rect 20139 15184 20140 15224
rect 20180 15184 20181 15224
rect 20139 15175 20181 15184
rect 20140 15056 20180 15175
rect 20140 15007 20180 15016
rect 19948 14888 19988 14897
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19948 14216 19988 14848
rect 20236 14804 20276 15772
rect 20332 15233 20372 15847
rect 20331 15224 20373 15233
rect 20331 15184 20332 15224
rect 20372 15184 20373 15224
rect 20331 15175 20373 15184
rect 20811 15140 20853 15149
rect 20811 15100 20812 15140
rect 20852 15100 20853 15140
rect 20811 15091 20853 15100
rect 20812 15006 20852 15091
rect 20236 14755 20276 14764
rect 19852 14176 19988 14216
rect 20044 14216 20084 14225
rect 19180 14132 19220 14141
rect 19180 13376 19220 14092
rect 19180 13327 19220 13336
rect 19852 13040 19892 14176
rect 19852 12991 19892 13000
rect 19948 13964 19988 13973
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 18988 12403 19028 12412
rect 19756 12452 19796 12461
rect 18796 8791 18836 8800
rect 18892 12284 18932 12293
rect 15724 8287 15764 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 11500 7160 11540 7169
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 11500 5648 11540 7120
rect 18892 7160 18932 12244
rect 19756 12284 19796 12412
rect 19756 12235 19796 12244
rect 19948 12116 19988 13924
rect 20044 13880 20084 14176
rect 20044 13831 20084 13840
rect 21580 13460 21620 16780
rect 24267 16232 24309 16241
rect 24267 16192 24268 16232
rect 24308 16192 24309 16232
rect 24267 16183 24309 16192
rect 24268 16098 24308 16183
rect 24459 15896 24501 15905
rect 24459 15856 24460 15896
rect 24500 15856 24501 15896
rect 24459 15847 24501 15856
rect 24460 15762 24500 15847
rect 21676 15728 21716 15737
rect 21676 14636 21716 15688
rect 24267 15140 24309 15149
rect 24267 15100 24268 15140
rect 24308 15100 24309 15140
rect 24267 15091 24309 15100
rect 25708 15140 25748 18964
rect 25708 15091 25748 15100
rect 26188 17660 26228 17669
rect 24268 15006 24308 15091
rect 21676 14587 21716 14596
rect 26188 14132 26228 17620
rect 31564 16484 31604 16493
rect 31564 15644 31604 16444
rect 31564 15595 31604 15604
rect 26188 14083 26228 14092
rect 27724 15560 27764 15569
rect 27724 15056 27764 15520
rect 20044 13292 20084 13301
rect 20044 12284 20084 13252
rect 20811 12536 20853 12545
rect 20811 12496 20812 12536
rect 20852 12496 20853 12536
rect 20811 12487 20853 12496
rect 20812 12402 20852 12487
rect 20044 12235 20084 12244
rect 20140 12116 20180 12125
rect 19988 12076 20140 12116
rect 19948 11981 19988 12076
rect 20140 12067 20180 12076
rect 21580 11780 21620 13420
rect 26764 13544 26804 13553
rect 26668 12788 26708 12797
rect 21580 11731 21620 11740
rect 25996 12452 26036 12461
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 25996 11192 26036 12412
rect 26668 12032 26708 12748
rect 26668 11983 26708 11992
rect 26764 11948 26804 13504
rect 26764 11899 26804 11908
rect 25996 11143 26036 11152
rect 26092 11696 26132 11705
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 25036 8840 25076 8849
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 25036 7916 25076 8800
rect 25227 8168 25269 8177
rect 25227 8128 25228 8168
rect 25268 8128 25269 8168
rect 25227 8119 25269 8128
rect 24556 7244 24596 7255
rect 24556 7169 24596 7204
rect 18892 7111 18932 7120
rect 24555 7160 24597 7169
rect 24555 7120 24556 7160
rect 24596 7120 24597 7160
rect 24555 7111 24597 7120
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 23788 6740 23828 6749
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 11500 5599 11540 5608
rect 11788 5900 11828 5909
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 11788 3380 11828 5860
rect 15724 5732 15764 5741
rect 15340 5396 15380 5405
rect 15340 4640 15380 5356
rect 15340 3464 15380 4600
rect 15340 3415 15380 3424
rect 15724 4724 15764 5692
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 11788 3331 11828 3340
rect 15724 3128 15764 4684
rect 23788 4808 23828 6700
rect 24939 6320 24981 6329
rect 24939 6280 24940 6320
rect 24980 6280 24981 6320
rect 24939 6271 24981 6280
rect 24940 6186 24980 6271
rect 25036 5480 25076 7876
rect 25228 7748 25268 8119
rect 25228 7699 25268 7708
rect 25036 5431 25076 5440
rect 25228 6404 25268 6413
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 23788 4220 23828 4768
rect 23788 4171 23828 4180
rect 25228 3884 25268 6364
rect 26092 4976 26132 11656
rect 26667 11024 26709 11033
rect 26667 10984 26668 11024
rect 26708 10984 26709 11024
rect 26667 10975 26709 10984
rect 26668 10940 26708 10975
rect 26668 10889 26708 10900
rect 27724 8840 27764 15016
rect 31948 14972 31988 20056
rect 35211 20096 35253 20105
rect 35211 20056 35212 20096
rect 35252 20056 35253 20096
rect 35211 20047 35253 20056
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 32428 19172 32468 19181
rect 29932 14216 29972 14225
rect 28204 13964 28244 13973
rect 28012 13376 28052 13385
rect 28012 13208 28052 13336
rect 28012 13159 28052 13168
rect 28204 13124 28244 13924
rect 28204 13075 28244 13084
rect 28972 13796 29012 13805
rect 28972 12872 29012 13756
rect 28972 12823 29012 12832
rect 29740 12956 29780 12965
rect 29740 11780 29780 12916
rect 29740 11731 29780 11740
rect 29932 11360 29972 14176
rect 31948 14048 31988 14932
rect 32044 16736 32084 16745
rect 32044 15392 32084 16696
rect 32428 16400 32468 19132
rect 34252 19088 34292 19097
rect 34252 18500 34292 19048
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 34252 18451 34292 18460
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 34444 17744 34484 17753
rect 34444 17669 34484 17704
rect 34443 17660 34485 17669
rect 34443 17620 34444 17660
rect 34484 17620 34485 17660
rect 34443 17611 34485 17620
rect 36555 17660 36597 17669
rect 36555 17620 36556 17660
rect 36596 17620 36597 17660
rect 36555 17611 36597 17620
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 32428 16064 32468 16360
rect 32428 16015 32468 16024
rect 32044 14552 32084 15352
rect 32044 14503 32084 14512
rect 32524 15308 32564 15317
rect 31948 13999 31988 14008
rect 29932 11311 29972 11320
rect 32524 11024 32564 15268
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 32524 10268 32564 10984
rect 32524 10219 32564 10228
rect 32620 14552 32660 14561
rect 27724 8791 27764 8800
rect 31852 9512 31892 9521
rect 31852 8177 31892 9472
rect 32620 9512 32660 14512
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 34444 12200 34484 17611
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 36556 17324 36596 17611
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 36556 16484 36596 17284
rect 36556 16435 36596 16444
rect 37324 17240 37364 17249
rect 37324 16148 37364 17200
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 37324 16099 37364 16108
rect 37708 16064 37748 16073
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 37132 15644 37172 15653
rect 37132 14972 37172 15604
rect 37708 15476 37748 16024
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 37708 15427 37748 15436
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 37132 14923 37172 14932
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 34444 12151 34484 12160
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 35020 11864 35060 11873
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 35020 11192 35060 11824
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 35020 11143 35060 11152
rect 32620 9463 32660 9472
rect 33100 10604 33140 10613
rect 33100 9512 33140 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 33100 9463 33140 9472
rect 34828 9596 34868 9605
rect 34828 9428 34868 9556
rect 34828 9379 34868 9388
rect 33868 9344 33908 9353
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 31948 8840 31988 8849
rect 31851 8168 31893 8177
rect 31851 8128 31852 8168
rect 31892 8128 31893 8168
rect 31851 8119 31893 8128
rect 31948 7748 31988 8800
rect 33868 8840 33908 9304
rect 33868 8791 33908 8800
rect 34060 9092 34100 9101
rect 34060 8168 34100 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 34060 8119 34100 8128
rect 34444 8588 34484 8597
rect 31948 7699 31988 7708
rect 30604 7580 30644 7589
rect 29259 7160 29301 7169
rect 29259 7120 29260 7160
rect 29300 7120 29301 7160
rect 29259 7111 29301 7120
rect 29260 7026 29300 7111
rect 30604 6329 30644 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 30603 6320 30645 6329
rect 30603 6280 30604 6320
rect 30644 6280 30645 6320
rect 30603 6271 30645 6280
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 34444 5564 34484 8548
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 34444 5515 34484 5524
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 26092 4927 26132 4936
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 15724 3079 15764 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 25228 2624 25268 3844
rect 25228 2575 25268 2584
rect 25708 4136 25748 4145
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 25708 1112 25748 4096
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 25708 1063 25748 1072
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 25996 26104 26036 26144
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 28204 23332 28244 23372
rect 28492 23332 28532 23372
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 39148 26188 39188 26228
rect 29836 26104 29876 26144
rect 41260 26020 41300 26060
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 30604 23332 30644 23372
rect 28588 22828 28628 22868
rect 35500 22828 35540 22868
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 16684 20056 16724 20096
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 76 19216 116 19256
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 26668 19216 26708 19256
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 14956 14008 14996 14048
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 16396 14008 16436 14048
rect 17644 14008 17684 14048
rect 15436 12496 15476 12536
rect 11788 10984 11828 11024
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 21196 16192 21236 16232
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 20332 15856 20372 15896
rect 20140 15184 20180 15224
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 20332 15184 20372 15224
rect 20812 15100 20852 15140
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 24268 16192 24308 16232
rect 24460 15856 24500 15896
rect 24268 15100 24308 15140
rect 20812 12496 20852 12536
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 25228 8128 25268 8168
rect 24556 7120 24596 7160
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 24940 6280 24980 6320
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 26668 10984 26708 11024
rect 35212 20056 35252 20096
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 34444 17620 34484 17660
rect 36556 17620 36596 17660
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 31852 8128 31892 8168
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 29260 7120 29300 7160
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 30604 6280 30644 6320
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 29492 26188 39148 26228
rect 39188 26188 39197 26228
rect 29492 26144 29532 26188
rect 25987 26104 25996 26144
rect 26036 26104 29532 26144
rect 29827 26104 29836 26144
rect 29876 26104 32780 26144
rect 32740 26060 32780 26104
rect 32740 26020 41260 26060
rect 41300 26020 41309 26060
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 28195 23332 28204 23372
rect 28244 23332 28492 23372
rect 28532 23332 30604 23372
rect 30644 23332 30653 23372
rect 28579 22828 28588 22868
rect 28628 22828 35500 22868
rect 35540 22828 35549 22868
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 16675 20056 16684 20096
rect 16724 20056 35212 20096
rect 35252 20056 35261 20096
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 67 19216 76 19256
rect 116 19216 26668 19256
rect 26708 19216 26717 19256
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 34435 17620 34444 17660
rect 34484 17620 36556 17660
rect 36596 17620 36605 17660
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 21187 16192 21196 16232
rect 21236 16192 24268 16232
rect 24308 16192 24317 16232
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 20323 15856 20332 15896
rect 20372 15856 24460 15896
rect 24500 15856 24509 15896
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 20131 15184 20140 15224
rect 20180 15184 20332 15224
rect 20372 15184 20381 15224
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 20803 15100 20812 15140
rect 20852 15100 24268 15140
rect 24308 15100 24317 15140
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 14947 14008 14956 14048
rect 14996 14008 16396 14048
rect 16436 14008 17644 14048
rect 17684 14008 17693 14048
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 15427 12496 15436 12536
rect 15476 12496 20812 12536
rect 20852 12496 20861 12536
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 11779 10984 11788 11024
rect 11828 10984 26668 11024
rect 26708 10984 26717 11024
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 25219 8128 25228 8168
rect 25268 8128 31852 8168
rect 31892 8128 31901 8168
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 24547 7120 24556 7160
rect 24596 7120 29260 7160
rect 29300 7120 29309 7160
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 24931 6280 24940 6320
rect 24980 6280 30604 6320
rect 30644 6280 30653 6320
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 37843 94236 38600
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 38599 95476 38682
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676451365
transform 1 0 26496 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_0_0_clk
timestamp 1676451365
transform -1 0 9888 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk
timestamp 1676451365
transform -1 0 9888 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk
timestamp 1676451365
transform 1 0 17376 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk
timestamp 1676451365
transform -1 0 18816 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk
timestamp 1676451365
transform -1 0 7200 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk
timestamp 1676451365
transform -1 0 7296 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk
timestamp 1676451365
transform 1 0 12672 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk
timestamp 1676451365
transform -1 0 14016 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk
timestamp 1676451365
transform -1 0 32736 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk
timestamp 1676451365
transform -1 0 31200 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk
timestamp 1676451365
transform -1 0 39840 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk
timestamp 1676451365
transform 1 0 40320 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk
timestamp 1676451365
transform -1 0 30720 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk
timestamp 1676451365
transform -1 0 30720 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk
timestamp 1676451365
transform 1 0 40320 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk
timestamp 1676451365
transform 1 0 40320 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_0__f_clk
timestamp 1676451365
transform -1 0 7680 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_1__f_clk
timestamp 1676451365
transform 1 0 10752 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_2__f_clk
timestamp 1676451365
transform -1 0 7008 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_3__f_clk
timestamp 1676451365
transform 1 0 11136 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_4__f_clk
timestamp 1676451365
transform -1 0 19776 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_5__f_clk
timestamp 1676451365
transform 1 0 19392 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_6__f_clk
timestamp 1676451365
transform -1 0 17472 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_7__f_clk
timestamp 1676451365
transform 1 0 19680 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_8__f_clk
timestamp 1676451365
transform -1 0 4320 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_9__f_clk
timestamp 1676451365
transform 1 0 7488 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_10__f_clk
timestamp 1676451365
transform -1 0 4896 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_11__f_clk
timestamp 1676451365
transform 1 0 5856 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_12__f_clk
timestamp 1676451365
transform -1 0 12480 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_13__f_clk
timestamp 1676451365
transform 1 0 14400 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_14__f_clk
timestamp 1676451365
transform -1 0 13440 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_15__f_clk
timestamp 1676451365
transform 1 0 14784 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_16__f_clk
timestamp 1676451365
transform -1 0 31584 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_17__f_clk
timestamp 1676451365
transform 1 0 33120 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_18__f_clk
timestamp 1676451365
transform -1 0 28128 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_19__f_clk
timestamp 1676451365
transform 1 0 30240 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_20__f_clk
timestamp 1676451365
transform -1 0 39264 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_21__f_clk
timestamp 1676451365
transform 1 0 39072 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_22__f_clk
timestamp 1676451365
transform -1 0 40512 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_23__f_clk
timestamp 1676451365
transform 1 0 43104 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_24__f_clk
timestamp 1676451365
transform -1 0 27168 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_25__f_clk
timestamp 1676451365
transform 1 0 32256 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_26__f_clk
timestamp 1676451365
transform -1 0 27072 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_27__f_clk
timestamp 1676451365
transform 1 0 31776 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_28__f_clk
timestamp 1676451365
transform 1 0 44448 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_29__f_clk
timestamp 1676451365
transform -1 0 44448 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_30__f_clk
timestamp 1676451365
transform -1 0 38304 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_31__f_clk
timestamp 1676451365
transform 1 0 43296 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_1  clkload0
timestamp 1676381911
transform 1 0 10656 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  clkload1
timestamp 1676381911
transform 1 0 11136 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  clkload2
timestamp 1676381911
transform 1 0 18720 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  clkload3
timestamp 1676381911
transform 1 0 19200 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  clkload4
timestamp 1676381911
transform 1 0 9600 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  clkload5
timestamp 1676381911
transform -1 0 10944 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  clkload6
timestamp 1676381911
transform -1 0 38112 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  clkload7
timestamp 1676381911
transform 1 0 37920 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  clkload8
timestamp 1676381911
transform 1 0 31872 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  clkload9
timestamp 1676381911
transform 1 0 24960 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_8  fanout307
timestamp 1676451365
transform -1 0 33408 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_1  fanout308
timestamp 1676381911
transform 1 0 33504 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_8  fanout309
timestamp 1676451365
transform -1 0 23232 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout310
timestamp 1676451365
transform -1 0 24480 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout311
timestamp 1676451365
transform -1 0 23232 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout312
timestamp 1676451365
transform 1 0 33600 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout313
timestamp 1676451365
transform 1 0 21216 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout314
timestamp 1676451365
transform -1 0 33504 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout315
timestamp 1676451365
transform -1 0 33504 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout316
timestamp 1676451365
transform -1 0 33600 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout317
timestamp 1676451365
transform 1 0 24864 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout318
timestamp 1676451365
transform -1 0 17184 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout319
timestamp 1676451365
transform -1 0 21984 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout320
timestamp 1676451365
transform -1 0 26784 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout321
timestamp 1676451365
transform 1 0 34464 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout322
timestamp 1676451365
transform 1 0 26784 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout323
timestamp 1676451365
transform 1 0 24192 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_1  fanout324
timestamp 1676381911
transform 1 0 24768 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_8  fanout325
timestamp 1676451365
transform -1 0 22848 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout326
timestamp 1676451365
transform 1 0 27744 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout327
timestamp 1676451365
transform -1 0 30240 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout328
timestamp 1676451365
transform -1 0 12960 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_1  fanout329
timestamp 1676381911
transform -1 0 13920 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_8  fanout330
timestamp 1676451365
transform 1 0 12192 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_2  fanout331
timestamp 1676381867
transform -1 0 33888 0 1 8316
box -48 -56 528 834
use sg13g2_buf_8  fanout332
timestamp 1676451365
transform 1 0 26592 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout333
timestamp 1676451365
transform -1 0 26592 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout334
timestamp 1676451365
transform -1 0 18144 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout335
timestamp 1676451365
transform 1 0 39168 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout336
timestamp 1676451365
transform 1 0 20832 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  fanout337
timestamp 1676451365
transform 1 0 7680 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_8  fanout338
timestamp 1676451365
transform 1 0 7200 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_2  fanout339
timestamp 1676381867
transform 1 0 8640 0 1 20412
box -48 -56 528 834
use sg13g2_buf_8  fanout340
timestamp 1676451365
transform -1 0 6336 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_1  fanout341
timestamp 1676381911
transform -1 0 5760 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_8  fanout342
timestamp 1676451365
transform 1 0 7200 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout343
timestamp 1676451365
transform -1 0 10368 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout344
timestamp 1676451365
transform -1 0 17184 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout345
timestamp 1676451365
transform 1 0 16416 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout346
timestamp 1676451365
transform 1 0 4032 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout347
timestamp 1676451365
transform 1 0 8448 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout348
timestamp 1676451365
transform -1 0 10176 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_1  fanout349
timestamp 1676381911
transform -1 0 9792 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_8  fanout350
timestamp 1676451365
transform 1 0 10944 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_2  fanout351
timestamp 1676381867
transform -1 0 10848 0 -1 34020
box -48 -56 528 834
use sg13g2_buf_2  fanout352
timestamp 1676381867
transform -1 0 10656 0 1 32508
box -48 -56 528 834
use sg13g2_buf_8  fanout353
timestamp 1676451365
transform 1 0 19008 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_1  fanout354
timestamp 1676381911
transform 1 0 19104 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_8  fanout355
timestamp 1676451365
transform 1 0 19872 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  fanout356
timestamp 1676451365
transform 1 0 19008 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout357
timestamp 1676451365
transform 1 0 13920 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout358
timestamp 1676451365
transform -1 0 37056 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_1  fanout359
timestamp 1676381911
transform 1 0 34560 0 1 23436
box -48 -56 432 834
use sg13g2_buf_8  fanout360
timestamp 1676451365
transform -1 0 47232 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_1  fanout361
timestamp 1676381911
transform -1 0 45984 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_8  fanout362
timestamp 1676451365
transform 1 0 40224 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout363
timestamp 1676451365
transform 1 0 35616 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout364
timestamp 1676451365
transform -1 0 33120 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_1  fanout365
timestamp 1676381911
transform -1 0 35904 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_8  fanout366
timestamp 1676451365
transform -1 0 31488 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_1  fanout367
timestamp 1676381911
transform -1 0 28608 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_8  fanout368
timestamp 1676451365
transform 1 0 32064 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout369
timestamp 1676451365
transform -1 0 33504 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout370
timestamp 1676451365
transform 1 0 46944 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout371
timestamp 1676451365
transform 1 0 45984 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout372
timestamp 1676451365
transform 1 0 38016 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout373
timestamp 1676451365
transform -1 0 43200 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_2  fanout374
timestamp 1676381867
transform 1 0 37824 0 -1 32508
box -48 -56 528 834
use sg13g2_buf_8  fanout375
timestamp 1676451365
transform -1 0 35136 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout376
timestamp 1676451365
transform 1 0 11328 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout377
timestamp 1676451365
transform 1 0 25920 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout378
timestamp 1676451365
transform -1 0 39072 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout379
timestamp 1676451365
transform -1 0 37248 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout380
timestamp 1676451365
transform -1 0 40704 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout381
timestamp 1676451365
transform -1 0 38016 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout382
timestamp 1676451365
transform 1 0 34464 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout383
timestamp 1676451365
transform 1 0 30240 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout384
timestamp 1676451365
transform -1 0 30624 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout385
timestamp 1676451365
transform 1 0 23232 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout386
timestamp 1676451365
transform -1 0 25920 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout387
timestamp 1676451365
transform -1 0 12768 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_1  fanout388
timestamp 1676381911
transform 1 0 11520 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_8  fanout389
timestamp 1676451365
transform -1 0 14112 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_2  fanout390
timestamp 1676381867
transform -1 0 12864 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_8  fanout391
timestamp 1676451365
transform -1 0 21312 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  fanout392
timestamp 1676451365
transform -1 0 21408 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_2  fanout393
timestamp 1676381867
transform -1 0 21888 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_8  fanout394
timestamp 1676451365
transform -1 0 25344 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_1  fanout395
timestamp 1676381911
transform 1 0 25056 0 1 9828
box -48 -56 432 834
use sg13g2_buf_8  fanout396
timestamp 1676451365
transform -1 0 23904 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_1  fanout397
timestamp 1676381911
transform 1 0 23232 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_8  fanout398
timestamp 1676451365
transform -1 0 22752 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_1  fanout399
timestamp 1676381911
transform 1 0 23232 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_8  fanout400
timestamp 1676451365
transform 1 0 30240 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_1  fanout401
timestamp 1676381911
transform -1 0 30240 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_8  fanout402
timestamp 1676451365
transform -1 0 25056 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout403
timestamp 1676451365
transform -1 0 23808 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout404
timestamp 1676451365
transform -1 0 16416 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_1  fanout405
timestamp 1676381911
transform -1 0 16416 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_8  fanout406
timestamp 1676451365
transform -1 0 25344 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout407
timestamp 1676451365
transform 1 0 27072 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout408
timestamp 1676451365
transform 1 0 28224 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout409
timestamp 1676451365
transform -1 0 32448 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout410
timestamp 1676451365
transform -1 0 9024 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout411
timestamp 1676451365
transform 1 0 8832 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout412
timestamp 1676451365
transform -1 0 23616 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout413
timestamp 1676451365
transform 1 0 22848 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout414
timestamp 1676451365
transform -1 0 25536 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout415
timestamp 1676451365
transform 1 0 34944 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout416
timestamp 1676451365
transform -1 0 28032 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout417
timestamp 1676451365
transform 1 0 40032 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout418
timestamp 1676451365
transform 1 0 41760 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_1  fanout419
timestamp 1676381911
transform -1 0 41568 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_2  fanout420
timestamp 1676381867
transform -1 0 40320 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_8  fanout421
timestamp 1676451365
transform 1 0 33696 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout422
timestamp 1676451365
transform -1 0 14400 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout423
timestamp 1676451365
transform -1 0 13824 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout424
timestamp 1676451365
transform -1 0 15840 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_1  fanout425
timestamp 1676381911
transform -1 0 15744 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_8  fanout426
timestamp 1676451365
transform 1 0 15168 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout427
timestamp 1676451365
transform 1 0 15744 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout428
timestamp 1676451365
transform -1 0 7296 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout429
timestamp 1676451365
transform -1 0 8736 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout430
timestamp 1676451365
transform -1 0 8064 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout431
timestamp 1676451365
transform -1 0 12192 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout432
timestamp 1676451365
transform -1 0 12864 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout433
timestamp 1676451365
transform -1 0 13248 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout434
timestamp 1676451365
transform -1 0 19872 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout435
timestamp 1676451365
transform 1 0 17280 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout436
timestamp 1676451365
transform -1 0 14304 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout437
timestamp 1676451365
transform -1 0 18336 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout438
timestamp 1676451365
transform -1 0 22752 0 -1 2268
box -48 -56 1296 834
use sg13g2_buf_8  fanout439
timestamp 1676451365
transform 1 0 24480 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout440
timestamp 1676451365
transform 1 0 31872 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout441
timestamp 1676451365
transform 1 0 31680 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout442
timestamp 1676451365
transform -1 0 33504 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout443
timestamp 1676451365
transform 1 0 31008 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout444
timestamp 1676451365
transform -1 0 27936 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout445
timestamp 1676451365
transform -1 0 34560 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  fanout446
timestamp 1676451365
transform -1 0 33312 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout447
timestamp 1676451365
transform 1 0 44448 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout448
timestamp 1676451365
transform -1 0 43680 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout449
timestamp 1676451365
transform -1 0 40032 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout450
timestamp 1676451365
transform -1 0 43200 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout451
timestamp 1676451365
transform 1 0 33312 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout452
timestamp 1676451365
transform 1 0 33120 0 1 20412
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_98
timestamp 1677579658
transform 1 0 9984 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_102
timestamp 1679581782
transform 1 0 10368 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_109
timestamp 1677579658
transform 1 0 11040 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_154
timestamp 1677579658
transform 1 0 15360 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_159
timestamp 1679581782
transform 1 0 15840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_166
timestamp 1679581782
transform 1 0 16512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_173
timestamp 1679581782
transform 1 0 17184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_180
timestamp 1679581782
transform 1 0 17856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_187
timestamp 1679581782
transform 1 0 18528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_194
timestamp 1679581782
transform 1 0 19200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_201
timestamp 1679581782
transform 1 0 19872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_208
timestamp 1679581782
transform 1 0 20544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_215
timestamp 1679581782
transform 1 0 21216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_222
timestamp 1679581782
transform 1 0 21888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_229
timestamp 1679581782
transform 1 0 22560 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_245
timestamp 1677580104
transform 1 0 24096 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_274
timestamp 1679581782
transform 1 0 26880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_281
timestamp 1679581782
transform 1 0 27552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_288
timestamp 1679581782
transform 1 0 28224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_295
timestamp 1679581782
transform 1 0 28896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_302
timestamp 1679581782
transform 1 0 29568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_309
timestamp 1679581782
transform 1 0 30240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_316
timestamp 1679581782
transform 1 0 30912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_323
timestamp 1679581782
transform 1 0 31584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_330
timestamp 1679581782
transform 1 0 32256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_337
timestamp 1679581782
transform 1 0 32928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_344
timestamp 1679581782
transform 1 0 33600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_351
timestamp 1679581782
transform 1 0 34272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_358
timestamp 1679581782
transform 1 0 34944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_365
timestamp 1679581782
transform 1 0 35616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_372
timestamp 1679581782
transform 1 0 36288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_379
timestamp 1679581782
transform 1 0 36960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_386
timestamp 1679581782
transform 1 0 37632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_393
timestamp 1679581782
transform 1 0 38304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_400
timestamp 1679581782
transform 1 0 38976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_407
timestamp 1679581782
transform 1 0 39648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_414
timestamp 1679581782
transform 1 0 40320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_421
timestamp 1679581782
transform 1 0 40992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_428
timestamp 1679581782
transform 1 0 41664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_435
timestamp 1679581782
transform 1 0 42336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_442
timestamp 1679581782
transform 1 0 43008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_449
timestamp 1679581782
transform 1 0 43680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_456
timestamp 1679581782
transform 1 0 44352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_463
timestamp 1679581782
transform 1 0 45024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_470
timestamp 1679581782
transform 1 0 45696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_477
timestamp 1679581782
transform 1 0 46368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_484
timestamp 1679581782
transform 1 0 47040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_491
timestamp 1679581782
transform 1 0 47712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_498
timestamp 1679581782
transform 1 0 48384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_505
timestamp 1679581782
transform 1 0 49056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_512
timestamp 1679581782
transform 1 0 49728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_519
timestamp 1679581782
transform 1 0 50400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_526
timestamp 1679581782
transform 1 0 51072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_533
timestamp 1679581782
transform 1 0 51744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_540
timestamp 1679581782
transform 1 0 52416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_547
timestamp 1679581782
transform 1 0 53088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_554
timestamp 1679581782
transform 1 0 53760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_561
timestamp 1679581782
transform 1 0 54432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_568
timestamp 1679581782
transform 1 0 55104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_575
timestamp 1679581782
transform 1 0 55776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_582
timestamp 1679581782
transform 1 0 56448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_589
timestamp 1679581782
transform 1 0 57120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_596
timestamp 1679581782
transform 1 0 57792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_603
timestamp 1679581782
transform 1 0 58464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_610
timestamp 1679581782
transform 1 0 59136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_617
timestamp 1679581782
transform 1 0 59808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_624
timestamp 1679581782
transform 1 0 60480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_631
timestamp 1679581782
transform 1 0 61152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_638
timestamp 1679581782
transform 1 0 61824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_645
timestamp 1679581782
transform 1 0 62496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_652
timestamp 1679581782
transform 1 0 63168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_659
timestamp 1679581782
transform 1 0 63840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_666
timestamp 1679581782
transform 1 0 64512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_673
timestamp 1679581782
transform 1 0 65184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_680
timestamp 1679581782
transform 1 0 65856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_687
timestamp 1679581782
transform 1 0 66528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_694
timestamp 1679581782
transform 1 0 67200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_701
timestamp 1679581782
transform 1 0 67872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_708
timestamp 1679581782
transform 1 0 68544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_715
timestamp 1679581782
transform 1 0 69216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_722
timestamp 1679581782
transform 1 0 69888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_729
timestamp 1679581782
transform 1 0 70560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_736
timestamp 1679581782
transform 1 0 71232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_743
timestamp 1679581782
transform 1 0 71904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_750
timestamp 1679581782
transform 1 0 72576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_757
timestamp 1679581782
transform 1 0 73248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_764
timestamp 1679581782
transform 1 0 73920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_771
timestamp 1679581782
transform 1 0 74592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_778
timestamp 1679581782
transform 1 0 75264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_785
timestamp 1679581782
transform 1 0 75936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_792
timestamp 1679581782
transform 1 0 76608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_799
timestamp 1679581782
transform 1 0 77280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_806
timestamp 1679581782
transform 1 0 77952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_813
timestamp 1679581782
transform 1 0 78624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_820
timestamp 1679581782
transform 1 0 79296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_827
timestamp 1679581782
transform 1 0 79968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_834
timestamp 1679581782
transform 1 0 80640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_841
timestamp 1679581782
transform 1 0 81312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_848
timestamp 1679581782
transform 1 0 81984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_855
timestamp 1679581782
transform 1 0 82656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_862
timestamp 1679581782
transform 1 0 83328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_869
timestamp 1679581782
transform 1 0 84000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_876
timestamp 1679581782
transform 1 0 84672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_883
timestamp 1679581782
transform 1 0 85344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_890
timestamp 1679581782
transform 1 0 86016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_897
timestamp 1679581782
transform 1 0 86688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_904
timestamp 1679581782
transform 1 0 87360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_911
timestamp 1679581782
transform 1 0 88032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_918
timestamp 1679581782
transform 1 0 88704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_925
timestamp 1679581782
transform 1 0 89376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_932
timestamp 1679581782
transform 1 0 90048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_939
timestamp 1679581782
transform 1 0 90720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_946
timestamp 1679581782
transform 1 0 91392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_953
timestamp 1679581782
transform 1 0 92064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_960
timestamp 1679581782
transform 1 0 92736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_967
timestamp 1679581782
transform 1 0 93408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_974
timestamp 1679581782
transform 1 0 94080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_981
timestamp 1679581782
transform 1 0 94752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_988
timestamp 1679581782
transform 1 0 95424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_995
timestamp 1679581782
transform 1 0 96096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1002
timestamp 1679581782
transform 1 0 96768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1009
timestamp 1679581782
transform 1 0 97440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1016
timestamp 1679581782
transform 1 0 98112 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_1023
timestamp 1679577901
transform 1 0 98784 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_1027
timestamp 1677580104
transform 1 0 99168 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_91
timestamp 1677580104
transform 1 0 9312 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_93
timestamp 1677579658
transform 1 0 9504 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_103
timestamp 1677580104
transform 1 0 10464 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_147
timestamp 1677580104
transform 1 0 14688 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_149
timestamp 1677579658
transform 1 0 14880 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_177
timestamp 1679581782
transform 1 0 17568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_184
timestamp 1679581782
transform 1 0 18240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_191
timestamp 1679581782
transform 1 0 18912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_198
timestamp 1679581782
transform 1 0 19584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_205
timestamp 1679577901
transform 1 0 20256 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_217
timestamp 1677579658
transform 1 0 21408 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_238
timestamp 1677579658
transform 1 0 23424 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_295
timestamp 1677580104
transform 1 0 28896 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_297
timestamp 1677579658
transform 1 0 29088 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_302
timestamp 1679581782
transform 1 0 29568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_309
timestamp 1679581782
transform 1 0 30240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_316
timestamp 1679581782
transform 1 0 30912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_323
timestamp 1679581782
transform 1 0 31584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_330
timestamp 1679581782
transform 1 0 32256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_337
timestamp 1679581782
transform 1 0 32928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_344
timestamp 1679581782
transform 1 0 33600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_351
timestamp 1679581782
transform 1 0 34272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_358
timestamp 1679581782
transform 1 0 34944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_365
timestamp 1679581782
transform 1 0 35616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_372
timestamp 1679581782
transform 1 0 36288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_379
timestamp 1679581782
transform 1 0 36960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_386
timestamp 1679581782
transform 1 0 37632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_393
timestamp 1679581782
transform 1 0 38304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_400
timestamp 1679581782
transform 1 0 38976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_407
timestamp 1679581782
transform 1 0 39648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_414
timestamp 1679581782
transform 1 0 40320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_421
timestamp 1679581782
transform 1 0 40992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_428
timestamp 1679581782
transform 1 0 41664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_435
timestamp 1679581782
transform 1 0 42336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_442
timestamp 1679581782
transform 1 0 43008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_449
timestamp 1679581782
transform 1 0 43680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_456
timestamp 1679581782
transform 1 0 44352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_463
timestamp 1679581782
transform 1 0 45024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_470
timestamp 1679581782
transform 1 0 45696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_477
timestamp 1679581782
transform 1 0 46368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_484
timestamp 1679581782
transform 1 0 47040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_491
timestamp 1679581782
transform 1 0 47712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_498
timestamp 1679581782
transform 1 0 48384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_505
timestamp 1679581782
transform 1 0 49056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_512
timestamp 1679581782
transform 1 0 49728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_519
timestamp 1679581782
transform 1 0 50400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_526
timestamp 1679581782
transform 1 0 51072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_533
timestamp 1679581782
transform 1 0 51744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_540
timestamp 1679581782
transform 1 0 52416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_547
timestamp 1679581782
transform 1 0 53088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_554
timestamp 1679581782
transform 1 0 53760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_561
timestamp 1679581782
transform 1 0 54432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_568
timestamp 1679581782
transform 1 0 55104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_575
timestamp 1679581782
transform 1 0 55776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_582
timestamp 1679581782
transform 1 0 56448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_589
timestamp 1679581782
transform 1 0 57120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_596
timestamp 1679581782
transform 1 0 57792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_603
timestamp 1679581782
transform 1 0 58464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_610
timestamp 1679581782
transform 1 0 59136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_617
timestamp 1679581782
transform 1 0 59808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_624
timestamp 1679581782
transform 1 0 60480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_631
timestamp 1679581782
transform 1 0 61152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_638
timestamp 1679581782
transform 1 0 61824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_645
timestamp 1679581782
transform 1 0 62496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_652
timestamp 1679581782
transform 1 0 63168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_659
timestamp 1679581782
transform 1 0 63840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_666
timestamp 1679581782
transform 1 0 64512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_673
timestamp 1679581782
transform 1 0 65184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_680
timestamp 1679581782
transform 1 0 65856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_687
timestamp 1679581782
transform 1 0 66528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_694
timestamp 1679581782
transform 1 0 67200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_701
timestamp 1679581782
transform 1 0 67872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_708
timestamp 1679581782
transform 1 0 68544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_715
timestamp 1679581782
transform 1 0 69216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_722
timestamp 1679581782
transform 1 0 69888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_729
timestamp 1679581782
transform 1 0 70560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_736
timestamp 1679581782
transform 1 0 71232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_743
timestamp 1679581782
transform 1 0 71904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_750
timestamp 1679581782
transform 1 0 72576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_757
timestamp 1679581782
transform 1 0 73248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_764
timestamp 1679581782
transform 1 0 73920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_771
timestamp 1679581782
transform 1 0 74592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_778
timestamp 1679581782
transform 1 0 75264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_785
timestamp 1679581782
transform 1 0 75936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_792
timestamp 1679581782
transform 1 0 76608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_799
timestamp 1679581782
transform 1 0 77280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_806
timestamp 1679581782
transform 1 0 77952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_813
timestamp 1679581782
transform 1 0 78624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_820
timestamp 1679581782
transform 1 0 79296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_827
timestamp 1679581782
transform 1 0 79968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_834
timestamp 1679581782
transform 1 0 80640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_841
timestamp 1679581782
transform 1 0 81312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_848
timestamp 1679581782
transform 1 0 81984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_855
timestamp 1679581782
transform 1 0 82656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_862
timestamp 1679581782
transform 1 0 83328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_869
timestamp 1679581782
transform 1 0 84000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_876
timestamp 1679581782
transform 1 0 84672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_883
timestamp 1679581782
transform 1 0 85344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_890
timestamp 1679581782
transform 1 0 86016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_897
timestamp 1679581782
transform 1 0 86688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_904
timestamp 1679581782
transform 1 0 87360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_911
timestamp 1679581782
transform 1 0 88032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_918
timestamp 1679581782
transform 1 0 88704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_925
timestamp 1679581782
transform 1 0 89376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_932
timestamp 1679581782
transform 1 0 90048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_939
timestamp 1679581782
transform 1 0 90720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_946
timestamp 1679581782
transform 1 0 91392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_953
timestamp 1679581782
transform 1 0 92064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_960
timestamp 1679581782
transform 1 0 92736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_967
timestamp 1679581782
transform 1 0 93408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_974
timestamp 1679581782
transform 1 0 94080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_981
timestamp 1679581782
transform 1 0 94752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_988
timestamp 1679581782
transform 1 0 95424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_995
timestamp 1679581782
transform 1 0 96096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1002
timestamp 1679581782
transform 1 0 96768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1009
timestamp 1679581782
transform 1 0 97440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1016
timestamp 1679581782
transform 1 0 98112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_1023
timestamp 1679577901
transform 1 0 98784 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_1027
timestamp 1677580104
transform 1 0 99168 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_53
timestamp 1677580104
transform 1 0 5664 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_55
timestamp 1677579658
transform 1 0 5856 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_69
timestamp 1679581782
transform 1 0 7200 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_76
timestamp 1677579658
transform 1 0 7872 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_85
timestamp 1677580104
transform 1 0 8736 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_87
timestamp 1677579658
transform 1 0 8928 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_121
timestamp 1679577901
transform 1 0 12192 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_125
timestamp 1677580104
transform 1 0 12576 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_154
timestamp 1677580104
transform 1 0 15360 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_156
timestamp 1677579658
transform 1 0 15552 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_172
timestamp 1677579658
transform 1 0 17088 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_177
timestamp 1679577901
transform 1 0 17568 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_190
timestamp 1679581782
transform 1 0 18816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_197
timestamp 1679577901
transform 1 0 19488 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_218
timestamp 1677580104
transform 1 0 21504 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_220
timestamp 1677579658
transform 1 0 21696 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_307
timestamp 1677579658
transform 1 0 30048 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_317
timestamp 1679581782
transform 1 0 31008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_324
timestamp 1679581782
transform 1 0 31680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_331
timestamp 1679581782
transform 1 0 32352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_338
timestamp 1679581782
transform 1 0 33024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_345
timestamp 1679581782
transform 1 0 33696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_352
timestamp 1679581782
transform 1 0 34368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_359
timestamp 1679581782
transform 1 0 35040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_366
timestamp 1679581782
transform 1 0 35712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_373
timestamp 1679581782
transform 1 0 36384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_380
timestamp 1679581782
transform 1 0 37056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_387
timestamp 1679581782
transform 1 0 37728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_394
timestamp 1679581782
transform 1 0 38400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_401
timestamp 1679581782
transform 1 0 39072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_408
timestamp 1679581782
transform 1 0 39744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_415
timestamp 1679581782
transform 1 0 40416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_422
timestamp 1679581782
transform 1 0 41088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_429
timestamp 1679581782
transform 1 0 41760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_436
timestamp 1679581782
transform 1 0 42432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_443
timestamp 1679581782
transform 1 0 43104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_450
timestamp 1679581782
transform 1 0 43776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_457
timestamp 1679581782
transform 1 0 44448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_464
timestamp 1679581782
transform 1 0 45120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_471
timestamp 1679581782
transform 1 0 45792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_478
timestamp 1679581782
transform 1 0 46464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_485
timestamp 1679581782
transform 1 0 47136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_492
timestamp 1679581782
transform 1 0 47808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_499
timestamp 1679581782
transform 1 0 48480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_506
timestamp 1679581782
transform 1 0 49152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_513
timestamp 1679581782
transform 1 0 49824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_520
timestamp 1679581782
transform 1 0 50496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_527
timestamp 1679581782
transform 1 0 51168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_534
timestamp 1679581782
transform 1 0 51840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_541
timestamp 1679581782
transform 1 0 52512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_548
timestamp 1679581782
transform 1 0 53184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_555
timestamp 1679581782
transform 1 0 53856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_562
timestamp 1679581782
transform 1 0 54528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_569
timestamp 1679581782
transform 1 0 55200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_576
timestamp 1679581782
transform 1 0 55872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_583
timestamp 1679581782
transform 1 0 56544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_590
timestamp 1679581782
transform 1 0 57216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_597
timestamp 1679581782
transform 1 0 57888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_604
timestamp 1679581782
transform 1 0 58560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_611
timestamp 1679581782
transform 1 0 59232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_618
timestamp 1679581782
transform 1 0 59904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_639
timestamp 1679581782
transform 1 0 61920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_646
timestamp 1679581782
transform 1 0 62592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_653
timestamp 1679581782
transform 1 0 63264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_660
timestamp 1679581782
transform 1 0 63936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_667
timestamp 1679581782
transform 1 0 64608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_674
timestamp 1679581782
transform 1 0 65280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_681
timestamp 1679581782
transform 1 0 65952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_688
timestamp 1679581782
transform 1 0 66624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_695
timestamp 1679581782
transform 1 0 67296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_702
timestamp 1679581782
transform 1 0 67968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_709
timestamp 1679581782
transform 1 0 68640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_730
timestamp 1679581782
transform 1 0 70656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_737
timestamp 1679581782
transform 1 0 71328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_744
timestamp 1679581782
transform 1 0 72000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_751
timestamp 1679581782
transform 1 0 72672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_758
timestamp 1679581782
transform 1 0 73344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_765
timestamp 1679581782
transform 1 0 74016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_772
timestamp 1679581782
transform 1 0 74688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_779
timestamp 1679581782
transform 1 0 75360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_786
timestamp 1679581782
transform 1 0 76032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_793
timestamp 1679581782
transform 1 0 76704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_800
timestamp 1679581782
transform 1 0 77376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_807
timestamp 1679581782
transform 1 0 78048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_814
timestamp 1679581782
transform 1 0 78720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_821
timestamp 1679581782
transform 1 0 79392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_828
timestamp 1679581782
transform 1 0 80064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_835
timestamp 1679581782
transform 1 0 80736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_842
timestamp 1679581782
transform 1 0 81408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_849
timestamp 1679581782
transform 1 0 82080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_856
timestamp 1679581782
transform 1 0 82752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_863
timestamp 1679581782
transform 1 0 83424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_870
timestamp 1679581782
transform 1 0 84096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_877
timestamp 1679581782
transform 1 0 84768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_884
timestamp 1679581782
transform 1 0 85440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_891
timestamp 1679581782
transform 1 0 86112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_898
timestamp 1679581782
transform 1 0 86784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_905
timestamp 1679581782
transform 1 0 87456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_912
timestamp 1679581782
transform 1 0 88128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_919
timestamp 1679581782
transform 1 0 88800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_926
timestamp 1679581782
transform 1 0 89472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_933
timestamp 1679581782
transform 1 0 90144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_940
timestamp 1679581782
transform 1 0 90816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_947
timestamp 1679581782
transform 1 0 91488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_954
timestamp 1679581782
transform 1 0 92160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_961
timestamp 1679581782
transform 1 0 92832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_968
timestamp 1679581782
transform 1 0 93504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_975
timestamp 1679581782
transform 1 0 94176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_982
timestamp 1679581782
transform 1 0 94848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_989
timestamp 1679581782
transform 1 0 95520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_996
timestamp 1679581782
transform 1 0 96192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1003
timestamp 1679581782
transform 1 0 96864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1010
timestamp 1679581782
transform 1 0 97536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1017
timestamp 1679581782
transform 1 0 98208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_1024
timestamp 1679577901
transform 1 0 98880 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_46
timestamp 1679577901
transform 1 0 4992 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_86
timestamp 1677580104
transform 1 0 8832 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_88
timestamp 1677579658
transform 1 0 9024 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_105
timestamp 1677580104
transform 1 0 10656 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_107
timestamp 1677579658
transform 1 0 10848 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_130
timestamp 1677580104
transform 1 0 13056 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_136
timestamp 1679581782
transform 1 0 13632 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_143
timestamp 1677579658
transform 1 0 14304 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_160
timestamp 1677580104
transform 1 0 15936 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_167
timestamp 1677579658
transform 1 0 16608 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_195
timestamp 1679577901
transform 1 0 19296 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_267
timestamp 1677580104
transform 1 0 26208 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_327
timestamp 1679581782
transform 1 0 31968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_334
timestamp 1679581782
transform 1 0 32640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_341
timestamp 1679581782
transform 1 0 33312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_348
timestamp 1679581782
transform 1 0 33984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_355
timestamp 1679581782
transform 1 0 34656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_362
timestamp 1679581782
transform 1 0 35328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_369
timestamp 1679581782
transform 1 0 36000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_376
timestamp 1679581782
transform 1 0 36672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_383
timestamp 1679581782
transform 1 0 37344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_390
timestamp 1679581782
transform 1 0 38016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_397
timestamp 1679581782
transform 1 0 38688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_404
timestamp 1679581782
transform 1 0 39360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_411
timestamp 1679581782
transform 1 0 40032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_418
timestamp 1679581782
transform 1 0 40704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_425
timestamp 1679581782
transform 1 0 41376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_432
timestamp 1679581782
transform 1 0 42048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_439
timestamp 1679581782
transform 1 0 42720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_446
timestamp 1679581782
transform 1 0 43392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_453
timestamp 1679581782
transform 1 0 44064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_460
timestamp 1679581782
transform 1 0 44736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_467
timestamp 1679581782
transform 1 0 45408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_474
timestamp 1679581782
transform 1 0 46080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_481
timestamp 1679581782
transform 1 0 46752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_488
timestamp 1679581782
transform 1 0 47424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_495
timestamp 1679581782
transform 1 0 48096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_502
timestamp 1679581782
transform 1 0 48768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_509
timestamp 1679581782
transform 1 0 49440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_516
timestamp 1679581782
transform 1 0 50112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_523
timestamp 1679581782
transform 1 0 50784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_530
timestamp 1679581782
transform 1 0 51456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_537
timestamp 1679581782
transform 1 0 52128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_544
timestamp 1679581782
transform 1 0 52800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_551
timestamp 1679581782
transform 1 0 53472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_558
timestamp 1679581782
transform 1 0 54144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_565
timestamp 1679581782
transform 1 0 54816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_572
timestamp 1679581782
transform 1 0 55488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_579
timestamp 1679581782
transform 1 0 56160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_586
timestamp 1679581782
transform 1 0 56832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_593
timestamp 1679581782
transform 1 0 57504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_600
timestamp 1679581782
transform 1 0 58176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_607
timestamp 1679581782
transform 1 0 58848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_614
timestamp 1679581782
transform 1 0 59520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_621
timestamp 1679581782
transform 1 0 60192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_628
timestamp 1679581782
transform 1 0 60864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_635
timestamp 1679581782
transform 1 0 61536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_642
timestamp 1679581782
transform 1 0 62208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_649
timestamp 1679581782
transform 1 0 62880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_656
timestamp 1679581782
transform 1 0 63552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_663
timestamp 1679581782
transform 1 0 64224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_670
timestamp 1679581782
transform 1 0 64896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_677
timestamp 1679581782
transform 1 0 65568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_684
timestamp 1679581782
transform 1 0 66240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_691
timestamp 1679581782
transform 1 0 66912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_698
timestamp 1679581782
transform 1 0 67584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_705
timestamp 1679581782
transform 1 0 68256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_712
timestamp 1679581782
transform 1 0 68928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_719
timestamp 1679581782
transform 1 0 69600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_726
timestamp 1679581782
transform 1 0 70272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_733
timestamp 1679581782
transform 1 0 70944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_740
timestamp 1679581782
transform 1 0 71616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_747
timestamp 1679581782
transform 1 0 72288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_754
timestamp 1679581782
transform 1 0 72960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_761
timestamp 1679581782
transform 1 0 73632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_768
timestamp 1679581782
transform 1 0 74304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_775
timestamp 1679581782
transform 1 0 74976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_782
timestamp 1679581782
transform 1 0 75648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_789
timestamp 1679581782
transform 1 0 76320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_796
timestamp 1679581782
transform 1 0 76992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_803
timestamp 1679581782
transform 1 0 77664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_810
timestamp 1679581782
transform 1 0 78336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_817
timestamp 1679581782
transform 1 0 79008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_824
timestamp 1679581782
transform 1 0 79680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_831
timestamp 1679581782
transform 1 0 80352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_838
timestamp 1679581782
transform 1 0 81024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_845
timestamp 1679581782
transform 1 0 81696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_852
timestamp 1679581782
transform 1 0 82368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_859
timestamp 1679581782
transform 1 0 83040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_866
timestamp 1679581782
transform 1 0 83712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_873
timestamp 1679581782
transform 1 0 84384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_880
timestamp 1679581782
transform 1 0 85056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_887
timestamp 1679581782
transform 1 0 85728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_894
timestamp 1679581782
transform 1 0 86400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_901
timestamp 1679581782
transform 1 0 87072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_908
timestamp 1679581782
transform 1 0 87744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_915
timestamp 1679581782
transform 1 0 88416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_922
timestamp 1679581782
transform 1 0 89088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_929
timestamp 1679581782
transform 1 0 89760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_936
timestamp 1679581782
transform 1 0 90432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_943
timestamp 1679581782
transform 1 0 91104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_950
timestamp 1679581782
transform 1 0 91776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_957
timestamp 1679581782
transform 1 0 92448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_964
timestamp 1679581782
transform 1 0 93120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_971
timestamp 1679581782
transform 1 0 93792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_978
timestamp 1679581782
transform 1 0 94464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_985
timestamp 1679581782
transform 1 0 95136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_992
timestamp 1679581782
transform 1 0 95808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_999
timestamp 1679581782
transform 1 0 96480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1006
timestamp 1679581782
transform 1 0 97152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1013
timestamp 1679581782
transform 1 0 97824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1020
timestamp 1679581782
transform 1 0 98496 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1027
timestamp 1677580104
transform 1 0 99168 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_25
timestamp 1677580104
transform 1 0 2976 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_27
timestamp 1677579658
transform 1 0 3168 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_56
timestamp 1677580104
transform 1 0 5952 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_96
timestamp 1679577901
transform 1 0 9792 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_100
timestamp 1677580104
transform 1 0 10176 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_244
timestamp 1679581782
transform 1 0 24000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_251
timestamp 1679577901
transform 1 0 24672 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_277
timestamp 1677580104
transform 1 0 27168 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_279
timestamp 1677579658
transform 1 0 27360 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_335
timestamp 1679581782
transform 1 0 32736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_342
timestamp 1679581782
transform 1 0 33408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_349
timestamp 1679581782
transform 1 0 34080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_356
timestamp 1679581782
transform 1 0 34752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_363
timestamp 1679581782
transform 1 0 35424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_370
timestamp 1679581782
transform 1 0 36096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_377
timestamp 1679581782
transform 1 0 36768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_384
timestamp 1679581782
transform 1 0 37440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_391
timestamp 1679581782
transform 1 0 38112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_398
timestamp 1679581782
transform 1 0 38784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_405
timestamp 1679581782
transform 1 0 39456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_412
timestamp 1679581782
transform 1 0 40128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_419
timestamp 1679581782
transform 1 0 40800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_426
timestamp 1679581782
transform 1 0 41472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_433
timestamp 1679581782
transform 1 0 42144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_440
timestamp 1679581782
transform 1 0 42816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_447
timestamp 1679581782
transform 1 0 43488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_454
timestamp 1679581782
transform 1 0 44160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_461
timestamp 1679581782
transform 1 0 44832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_468
timestamp 1679581782
transform 1 0 45504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_475
timestamp 1679581782
transform 1 0 46176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_482
timestamp 1679581782
transform 1 0 46848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_489
timestamp 1679581782
transform 1 0 47520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_496
timestamp 1679581782
transform 1 0 48192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_503
timestamp 1679581782
transform 1 0 48864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_510
timestamp 1679581782
transform 1 0 49536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_517
timestamp 1679581782
transform 1 0 50208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_524
timestamp 1679581782
transform 1 0 50880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_531
timestamp 1679581782
transform 1 0 51552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_538
timestamp 1679581782
transform 1 0 52224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_545
timestamp 1679581782
transform 1 0 52896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_552
timestamp 1679581782
transform 1 0 53568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_559
timestamp 1679581782
transform 1 0 54240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_566
timestamp 1679581782
transform 1 0 54912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_573
timestamp 1679581782
transform 1 0 55584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_580
timestamp 1679581782
transform 1 0 56256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_587
timestamp 1679581782
transform 1 0 56928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_594
timestamp 1679581782
transform 1 0 57600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_601
timestamp 1679581782
transform 1 0 58272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_608
timestamp 1679581782
transform 1 0 58944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_615
timestamp 1679581782
transform 1 0 59616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_622
timestamp 1679581782
transform 1 0 60288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_629
timestamp 1679581782
transform 1 0 60960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_636
timestamp 1679581782
transform 1 0 61632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_643
timestamp 1679581782
transform 1 0 62304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_650
timestamp 1679581782
transform 1 0 62976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_657
timestamp 1679581782
transform 1 0 63648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_664
timestamp 1679581782
transform 1 0 64320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_671
timestamp 1679581782
transform 1 0 64992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_678
timestamp 1679581782
transform 1 0 65664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_685
timestamp 1679581782
transform 1 0 66336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_692
timestamp 1679581782
transform 1 0 67008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_699
timestamp 1679581782
transform 1 0 67680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_706
timestamp 1679581782
transform 1 0 68352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_713
timestamp 1679581782
transform 1 0 69024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_720
timestamp 1679581782
transform 1 0 69696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_727
timestamp 1679581782
transform 1 0 70368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_734
timestamp 1679581782
transform 1 0 71040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_741
timestamp 1679581782
transform 1 0 71712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_748
timestamp 1679581782
transform 1 0 72384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_755
timestamp 1679581782
transform 1 0 73056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_762
timestamp 1679581782
transform 1 0 73728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_769
timestamp 1679581782
transform 1 0 74400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_776
timestamp 1679581782
transform 1 0 75072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_783
timestamp 1679581782
transform 1 0 75744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_790
timestamp 1679581782
transform 1 0 76416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_797
timestamp 1679581782
transform 1 0 77088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_804
timestamp 1679581782
transform 1 0 77760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_811
timestamp 1679581782
transform 1 0 78432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_818
timestamp 1679581782
transform 1 0 79104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_825
timestamp 1679581782
transform 1 0 79776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_832
timestamp 1679581782
transform 1 0 80448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_839
timestamp 1679581782
transform 1 0 81120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_846
timestamp 1679581782
transform 1 0 81792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_853
timestamp 1679581782
transform 1 0 82464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_860
timestamp 1679581782
transform 1 0 83136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_867
timestamp 1679581782
transform 1 0 83808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_874
timestamp 1679581782
transform 1 0 84480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_881
timestamp 1679581782
transform 1 0 85152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_888
timestamp 1679581782
transform 1 0 85824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_895
timestamp 1679581782
transform 1 0 86496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_902
timestamp 1679581782
transform 1 0 87168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_909
timestamp 1679581782
transform 1 0 87840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_916
timestamp 1679581782
transform 1 0 88512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_923
timestamp 1679581782
transform 1 0 89184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_930
timestamp 1679581782
transform 1 0 89856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_937
timestamp 1679581782
transform 1 0 90528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_944
timestamp 1679581782
transform 1 0 91200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_951
timestamp 1679581782
transform 1 0 91872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_958
timestamp 1679581782
transform 1 0 92544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_965
timestamp 1679581782
transform 1 0 93216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_972
timestamp 1679581782
transform 1 0 93888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_979
timestamp 1679581782
transform 1 0 94560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_986
timestamp 1679581782
transform 1 0 95232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_993
timestamp 1679581782
transform 1 0 95904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1000
timestamp 1679581782
transform 1 0 96576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1007
timestamp 1679581782
transform 1 0 97248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1014
timestamp 1679581782
transform 1 0 97920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1021
timestamp 1679581782
transform 1 0 98592 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_1028
timestamp 1677579658
transform 1 0 99264 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_32
timestamp 1677579658
transform 1 0 3648 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_51
timestamp 1677580104
transform 1 0 5472 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_112
timestamp 1677580104
transform 1 0 11328 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_114
timestamp 1677579658
transform 1 0 11520 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_135
timestamp 1677579658
transform 1 0 13536 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_150
timestamp 1677579658
transform 1 0 14976 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_177
timestamp 1677579658
transform 1 0 17568 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_200
timestamp 1677579658
transform 1 0 19776 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_263
timestamp 1677579658
transform 1 0 25824 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_283
timestamp 1677579658
transform 1 0 27744 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_325
timestamp 1679581782
transform 1 0 31776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_332
timestamp 1679581782
transform 1 0 32448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_339
timestamp 1679581782
transform 1 0 33120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_346
timestamp 1679581782
transform 1 0 33792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_353
timestamp 1679581782
transform 1 0 34464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_360
timestamp 1679581782
transform 1 0 35136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_367
timestamp 1679581782
transform 1 0 35808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_374
timestamp 1679581782
transform 1 0 36480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_381
timestamp 1679581782
transform 1 0 37152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_388
timestamp 1679581782
transform 1 0 37824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_395
timestamp 1679581782
transform 1 0 38496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_402
timestamp 1679581782
transform 1 0 39168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_409
timestamp 1679581782
transform 1 0 39840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_416
timestamp 1679581782
transform 1 0 40512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_423
timestamp 1679581782
transform 1 0 41184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_430
timestamp 1679581782
transform 1 0 41856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_437
timestamp 1679581782
transform 1 0 42528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_444
timestamp 1679581782
transform 1 0 43200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_451
timestamp 1679581782
transform 1 0 43872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_458
timestamp 1679581782
transform 1 0 44544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_465
timestamp 1679581782
transform 1 0 45216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_472
timestamp 1679581782
transform 1 0 45888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_479
timestamp 1679581782
transform 1 0 46560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_486
timestamp 1679581782
transform 1 0 47232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_493
timestamp 1679581782
transform 1 0 47904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_500
timestamp 1679581782
transform 1 0 48576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_507
timestamp 1679581782
transform 1 0 49248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_514
timestamp 1679581782
transform 1 0 49920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_521
timestamp 1679581782
transform 1 0 50592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_528
timestamp 1679581782
transform 1 0 51264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_535
timestamp 1679581782
transform 1 0 51936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_542
timestamp 1679581782
transform 1 0 52608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_549
timestamp 1679581782
transform 1 0 53280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_556
timestamp 1679581782
transform 1 0 53952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_563
timestamp 1679581782
transform 1 0 54624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_570
timestamp 1679581782
transform 1 0 55296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_577
timestamp 1679581782
transform 1 0 55968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_584
timestamp 1679581782
transform 1 0 56640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_591
timestamp 1679581782
transform 1 0 57312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_598
timestamp 1679581782
transform 1 0 57984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_605
timestamp 1679581782
transform 1 0 58656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_612
timestamp 1679581782
transform 1 0 59328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_619
timestamp 1679581782
transform 1 0 60000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_626
timestamp 1679581782
transform 1 0 60672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_633
timestamp 1679581782
transform 1 0 61344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_640
timestamp 1679581782
transform 1 0 62016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_647
timestamp 1679581782
transform 1 0 62688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_654
timestamp 1679581782
transform 1 0 63360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_661
timestamp 1679581782
transform 1 0 64032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_668
timestamp 1679581782
transform 1 0 64704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_675
timestamp 1679581782
transform 1 0 65376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_682
timestamp 1679581782
transform 1 0 66048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_689
timestamp 1679581782
transform 1 0 66720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_696
timestamp 1679581782
transform 1 0 67392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_703
timestamp 1679581782
transform 1 0 68064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_710
timestamp 1679581782
transform 1 0 68736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_717
timestamp 1679581782
transform 1 0 69408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_724
timestamp 1679581782
transform 1 0 70080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_731
timestamp 1679581782
transform 1 0 70752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_738
timestamp 1679581782
transform 1 0 71424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_745
timestamp 1679581782
transform 1 0 72096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_752
timestamp 1679581782
transform 1 0 72768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_759
timestamp 1679581782
transform 1 0 73440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_766
timestamp 1679581782
transform 1 0 74112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_773
timestamp 1679581782
transform 1 0 74784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_780
timestamp 1679581782
transform 1 0 75456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_787
timestamp 1679581782
transform 1 0 76128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_794
timestamp 1679581782
transform 1 0 76800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_801
timestamp 1679581782
transform 1 0 77472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679581782
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679581782
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_822
timestamp 1679581782
transform 1 0 79488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_829
timestamp 1679581782
transform 1 0 80160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_836
timestamp 1679581782
transform 1 0 80832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_843
timestamp 1679581782
transform 1 0 81504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_850
timestamp 1679581782
transform 1 0 82176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_857
timestamp 1679581782
transform 1 0 82848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_864
timestamp 1679581782
transform 1 0 83520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_871
timestamp 1679581782
transform 1 0 84192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_878
timestamp 1679581782
transform 1 0 84864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_885
timestamp 1679581782
transform 1 0 85536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_892
timestamp 1679581782
transform 1 0 86208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_899
timestamp 1679581782
transform 1 0 86880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_906
timestamp 1679581782
transform 1 0 87552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_913
timestamp 1679581782
transform 1 0 88224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_920
timestamp 1679581782
transform 1 0 88896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_927
timestamp 1679581782
transform 1 0 89568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_934
timestamp 1679581782
transform 1 0 90240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_941
timestamp 1679581782
transform 1 0 90912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_948
timestamp 1679581782
transform 1 0 91584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_955
timestamp 1679581782
transform 1 0 92256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_962
timestamp 1679581782
transform 1 0 92928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_969
timestamp 1679581782
transform 1 0 93600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_976
timestamp 1679581782
transform 1 0 94272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_983
timestamp 1679581782
transform 1 0 94944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_990
timestamp 1679581782
transform 1 0 95616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_997
timestamp 1679581782
transform 1 0 96288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1004
timestamp 1679581782
transform 1 0 96960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1011
timestamp 1679581782
transform 1 0 97632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1018
timestamp 1679581782
transform 1 0 98304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_1025
timestamp 1679577901
transform 1 0 98976 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_32
timestamp 1677580104
transform 1 0 3648 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_34
timestamp 1677579658
transform 1 0 3840 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_56
timestamp 1677579658
transform 1 0 5952 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_93
timestamp 1677579658
transform 1 0 9504 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_108
timestamp 1677579658
transform 1 0 10944 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_119
timestamp 1677579658
transform 1 0 12000 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_125
timestamp 1677579658
transform 1 0 12576 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_156
timestamp 1677579658
transform 1 0 15552 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16416 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_172
timestamp 1677580104
transform 1 0 17088 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_174
timestamp 1677579658
transform 1 0 17280 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_179
timestamp 1677579658
transform 1 0 17760 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_208
timestamp 1677580104
transform 1 0 20544 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_210
timestamp 1677579658
transform 1 0 20736 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_239
timestamp 1677579658
transform 1 0 23520 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_245
timestamp 1677579658
transform 1 0 24096 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_269
timestamp 1679577901
transform 1 0 26400 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_279
timestamp 1679577901
transform 1 0 27360 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 31872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 32544 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_340
timestamp 1677580104
transform 1 0 33216 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_363
timestamp 1679581782
transform 1 0 35424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_370
timestamp 1679581782
transform 1 0 36096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_377
timestamp 1679581782
transform 1 0 36768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_384
timestamp 1679581782
transform 1 0 37440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_391
timestamp 1679581782
transform 1 0 38112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_398
timestamp 1679581782
transform 1 0 38784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_405
timestamp 1679581782
transform 1 0 39456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_412
timestamp 1679581782
transform 1 0 40128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_419
timestamp 1679581782
transform 1 0 40800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_426
timestamp 1679581782
transform 1 0 41472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_433
timestamp 1679581782
transform 1 0 42144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_440
timestamp 1679581782
transform 1 0 42816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_447
timestamp 1679581782
transform 1 0 43488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_454
timestamp 1679581782
transform 1 0 44160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_461
timestamp 1679581782
transform 1 0 44832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_468
timestamp 1679581782
transform 1 0 45504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_475
timestamp 1679581782
transform 1 0 46176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_482
timestamp 1679581782
transform 1 0 46848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_489
timestamp 1679581782
transform 1 0 47520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_496
timestamp 1679581782
transform 1 0 48192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_503
timestamp 1679581782
transform 1 0 48864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_510
timestamp 1679581782
transform 1 0 49536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_517
timestamp 1679581782
transform 1 0 50208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_524
timestamp 1679581782
transform 1 0 50880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_531
timestamp 1679581782
transform 1 0 51552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_538
timestamp 1679581782
transform 1 0 52224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_545
timestamp 1679581782
transform 1 0 52896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_552
timestamp 1679581782
transform 1 0 53568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_559
timestamp 1679581782
transform 1 0 54240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_566
timestamp 1679581782
transform 1 0 54912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_573
timestamp 1679581782
transform 1 0 55584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_580
timestamp 1679581782
transform 1 0 56256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_587
timestamp 1679581782
transform 1 0 56928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_594
timestamp 1679581782
transform 1 0 57600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_601
timestamp 1679581782
transform 1 0 58272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_608
timestamp 1679581782
transform 1 0 58944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_615
timestamp 1679581782
transform 1 0 59616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_622
timestamp 1679581782
transform 1 0 60288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_629
timestamp 1679581782
transform 1 0 60960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_636
timestamp 1679581782
transform 1 0 61632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_643
timestamp 1679581782
transform 1 0 62304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_650
timestamp 1679581782
transform 1 0 62976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_657
timestamp 1679581782
transform 1 0 63648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_664
timestamp 1679581782
transform 1 0 64320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_671
timestamp 1679581782
transform 1 0 64992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_678
timestamp 1679581782
transform 1 0 65664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_685
timestamp 1679581782
transform 1 0 66336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_692
timestamp 1679581782
transform 1 0 67008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_699
timestamp 1679581782
transform 1 0 67680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_706
timestamp 1679581782
transform 1 0 68352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_713
timestamp 1679581782
transform 1 0 69024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_720
timestamp 1679581782
transform 1 0 69696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_727
timestamp 1679581782
transform 1 0 70368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_734
timestamp 1679581782
transform 1 0 71040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_741
timestamp 1679581782
transform 1 0 71712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_748
timestamp 1679581782
transform 1 0 72384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_755
timestamp 1679581782
transform 1 0 73056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_762
timestamp 1679581782
transform 1 0 73728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_769
timestamp 1679581782
transform 1 0 74400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_776
timestamp 1679581782
transform 1 0 75072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_783
timestamp 1679581782
transform 1 0 75744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_790
timestamp 1679581782
transform 1 0 76416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_797
timestamp 1679581782
transform 1 0 77088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_804
timestamp 1679581782
transform 1 0 77760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_811
timestamp 1679581782
transform 1 0 78432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_818
timestamp 1679581782
transform 1 0 79104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_825
timestamp 1679581782
transform 1 0 79776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_832
timestamp 1679581782
transform 1 0 80448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_839
timestamp 1679581782
transform 1 0 81120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_846
timestamp 1679581782
transform 1 0 81792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_853
timestamp 1679581782
transform 1 0 82464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_860
timestamp 1679581782
transform 1 0 83136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_867
timestamp 1679581782
transform 1 0 83808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_874
timestamp 1679581782
transform 1 0 84480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_881
timestamp 1679581782
transform 1 0 85152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_888
timestamp 1679581782
transform 1 0 85824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_895
timestamp 1679581782
transform 1 0 86496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_902
timestamp 1679581782
transform 1 0 87168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_909
timestamp 1679581782
transform 1 0 87840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_916
timestamp 1679581782
transform 1 0 88512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_923
timestamp 1679581782
transform 1 0 89184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_930
timestamp 1679581782
transform 1 0 89856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_937
timestamp 1679581782
transform 1 0 90528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_944
timestamp 1679581782
transform 1 0 91200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_951
timestamp 1679581782
transform 1 0 91872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_958
timestamp 1679581782
transform 1 0 92544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_965
timestamp 1679581782
transform 1 0 93216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_972
timestamp 1679581782
transform 1 0 93888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_979
timestamp 1679581782
transform 1 0 94560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_986
timestamp 1679581782
transform 1 0 95232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_993
timestamp 1679581782
transform 1 0 95904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1000
timestamp 1679581782
transform 1 0 96576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1007
timestamp 1679581782
transform 1 0 97248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1014
timestamp 1679581782
transform 1 0 97920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1021
timestamp 1679581782
transform 1 0 98592 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677579658
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_28
timestamp 1679577901
transform 1 0 3264 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_77
timestamp 1677580104
transform 1 0 7968 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_119
timestamp 1677580104
transform 1 0 12000 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_121
timestamp 1677579658
transform 1 0 12192 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_133
timestamp 1677580104
transform 1 0 13344 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_135
timestamp 1677579658
transform 1 0 13536 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_144
timestamp 1677579658
transform 1 0 14400 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_184
timestamp 1677579658
transform 1 0 18240 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_193
timestamp 1677580104
transform 1 0 19104 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_195
timestamp 1677579658
transform 1 0 19296 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_209
timestamp 1677580104
transform 1 0 20640 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_278
timestamp 1679581782
transform 1 0 27264 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_285
timestamp 1677580104
transform 1 0 27936 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_287
timestamp 1677579658
transform 1 0 28128 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_391
timestamp 1679581782
transform 1 0 38112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_398
timestamp 1679581782
transform 1 0 38784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_405
timestamp 1679581782
transform 1 0 39456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_412
timestamp 1679581782
transform 1 0 40128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_419
timestamp 1679581782
transform 1 0 40800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_426
timestamp 1679581782
transform 1 0 41472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_433
timestamp 1679581782
transform 1 0 42144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_440
timestamp 1679581782
transform 1 0 42816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_447
timestamp 1679581782
transform 1 0 43488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_454
timestamp 1679581782
transform 1 0 44160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_461
timestamp 1679581782
transform 1 0 44832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_468
timestamp 1679581782
transform 1 0 45504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_475
timestamp 1679581782
transform 1 0 46176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_482
timestamp 1679581782
transform 1 0 46848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_489
timestamp 1679581782
transform 1 0 47520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_496
timestamp 1679581782
transform 1 0 48192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_503
timestamp 1679581782
transform 1 0 48864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_510
timestamp 1679581782
transform 1 0 49536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_517
timestamp 1679581782
transform 1 0 50208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_524
timestamp 1679581782
transform 1 0 50880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_531
timestamp 1679581782
transform 1 0 51552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_538
timestamp 1679581782
transform 1 0 52224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_545
timestamp 1679581782
transform 1 0 52896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_552
timestamp 1679581782
transform 1 0 53568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_559
timestamp 1679581782
transform 1 0 54240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_566
timestamp 1679581782
transform 1 0 54912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_573
timestamp 1679581782
transform 1 0 55584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_580
timestamp 1679581782
transform 1 0 56256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_587
timestamp 1679581782
transform 1 0 56928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_594
timestamp 1679581782
transform 1 0 57600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_601
timestamp 1679581782
transform 1 0 58272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_608
timestamp 1679581782
transform 1 0 58944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_615
timestamp 1679581782
transform 1 0 59616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_622
timestamp 1679581782
transform 1 0 60288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_629
timestamp 1679581782
transform 1 0 60960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_636
timestamp 1679581782
transform 1 0 61632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_643
timestamp 1679581782
transform 1 0 62304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_650
timestamp 1679581782
transform 1 0 62976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_657
timestamp 1679581782
transform 1 0 63648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_664
timestamp 1679581782
transform 1 0 64320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_671
timestamp 1679581782
transform 1 0 64992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_678
timestamp 1679581782
transform 1 0 65664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_685
timestamp 1679581782
transform 1 0 66336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_692
timestamp 1679581782
transform 1 0 67008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_699
timestamp 1679581782
transform 1 0 67680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_706
timestamp 1679581782
transform 1 0 68352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_713
timestamp 1679581782
transform 1 0 69024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_720
timestamp 1679581782
transform 1 0 69696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_727
timestamp 1679581782
transform 1 0 70368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_734
timestamp 1679581782
transform 1 0 71040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_741
timestamp 1679581782
transform 1 0 71712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_748
timestamp 1679581782
transform 1 0 72384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_755
timestamp 1679581782
transform 1 0 73056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_762
timestamp 1679581782
transform 1 0 73728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_769
timestamp 1679581782
transform 1 0 74400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_776
timestamp 1679581782
transform 1 0 75072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_783
timestamp 1679581782
transform 1 0 75744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_790
timestamp 1679581782
transform 1 0 76416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_797
timestamp 1679581782
transform 1 0 77088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_804
timestamp 1679581782
transform 1 0 77760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_811
timestamp 1679581782
transform 1 0 78432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_818
timestamp 1679581782
transform 1 0 79104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_825
timestamp 1679581782
transform 1 0 79776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_832
timestamp 1679581782
transform 1 0 80448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_839
timestamp 1679581782
transform 1 0 81120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_846
timestamp 1679581782
transform 1 0 81792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_853
timestamp 1679581782
transform 1 0 82464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_860
timestamp 1679581782
transform 1 0 83136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_867
timestamp 1679581782
transform 1 0 83808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_874
timestamp 1679581782
transform 1 0 84480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_881
timestamp 1679581782
transform 1 0 85152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_888
timestamp 1679581782
transform 1 0 85824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_895
timestamp 1679581782
transform 1 0 86496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_902
timestamp 1679581782
transform 1 0 87168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_909
timestamp 1679581782
transform 1 0 87840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_916
timestamp 1679581782
transform 1 0 88512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_923
timestamp 1679581782
transform 1 0 89184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_930
timestamp 1679581782
transform 1 0 89856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_937
timestamp 1679581782
transform 1 0 90528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_944
timestamp 1679581782
transform 1 0 91200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_951
timestamp 1679581782
transform 1 0 91872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_958
timestamp 1679581782
transform 1 0 92544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_965
timestamp 1679581782
transform 1 0 93216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_972
timestamp 1679581782
transform 1 0 93888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_979
timestamp 1679581782
transform 1 0 94560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_986
timestamp 1679581782
transform 1 0 95232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_993
timestamp 1679581782
transform 1 0 95904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1000
timestamp 1679581782
transform 1 0 96576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1007
timestamp 1679581782
transform 1 0 97248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1014
timestamp 1679581782
transform 1 0 97920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1021
timestamp 1679581782
transform 1 0 98592 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677579658
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_46
timestamp 1677579658
transform 1 0 4992 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_74
timestamp 1677579658
transform 1 0 7680 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_109
timestamp 1677580104
transform 1 0 11040 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_139
timestamp 1677580104
transform 1 0 13920 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_181
timestamp 1679581782
transform 1 0 17952 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_188
timestamp 1677580104
transform 1 0 18624 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_190
timestamp 1677579658
transform 1 0 18816 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_231
timestamp 1677579658
transform 1 0 22752 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_253
timestamp 1677580104
transform 1 0 24864 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_255
timestamp 1677579658
transform 1 0 25056 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_279
timestamp 1679577901
transform 1 0 27360 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_283
timestamp 1677580104
transform 1 0 27744 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_310
timestamp 1679581782
transform 1 0 30336 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_317
timestamp 1677579658
transform 1 0 31008 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_321
timestamp 1677579658
transform 1 0 31392 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_334
timestamp 1679581782
transform 1 0 32640 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_341
timestamp 1677580104
transform 1 0 33312 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_343
timestamp 1677579658
transform 1 0 33504 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_372
timestamp 1677580104
transform 1 0 36288 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679581782
transform 1 0 38208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_399
timestamp 1679581782
transform 1 0 38880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679581782
transform 1 0 39552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679581782
transform 1 0 40224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679581782
transform 1 0 40896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679581782
transform 1 0 41568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679581782
transform 1 0 42240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 42912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 43584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 44256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 44928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 45600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 46272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 46944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679581782
transform 1 0 47616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679581782
transform 1 0 48288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679581782
transform 1 0 48960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679581782
transform 1 0 49632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_518
timestamp 1679581782
transform 1 0 50304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_525
timestamp 1679581782
transform 1 0 50976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_532
timestamp 1679581782
transform 1 0 51648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_539
timestamp 1679581782
transform 1 0 52320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_546
timestamp 1679581782
transform 1 0 52992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_553
timestamp 1679581782
transform 1 0 53664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_560
timestamp 1679581782
transform 1 0 54336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_567
timestamp 1679581782
transform 1 0 55008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_574
timestamp 1679581782
transform 1 0 55680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_581
timestamp 1679581782
transform 1 0 56352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_588
timestamp 1679581782
transform 1 0 57024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_595
timestamp 1679581782
transform 1 0 57696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_602
timestamp 1679581782
transform 1 0 58368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_609
timestamp 1679581782
transform 1 0 59040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_616
timestamp 1679581782
transform 1 0 59712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_623
timestamp 1679581782
transform 1 0 60384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_630
timestamp 1679581782
transform 1 0 61056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_637
timestamp 1679581782
transform 1 0 61728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_644
timestamp 1679581782
transform 1 0 62400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_651
timestamp 1679581782
transform 1 0 63072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_658
timestamp 1679581782
transform 1 0 63744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_665
timestamp 1679581782
transform 1 0 64416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_672
timestamp 1679581782
transform 1 0 65088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_679
timestamp 1679581782
transform 1 0 65760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_686
timestamp 1679581782
transform 1 0 66432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_693
timestamp 1679581782
transform 1 0 67104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_700
timestamp 1679581782
transform 1 0 67776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_707
timestamp 1679581782
transform 1 0 68448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_714
timestamp 1679581782
transform 1 0 69120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_721
timestamp 1679581782
transform 1 0 69792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 70464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_735
timestamp 1679581782
transform 1 0 71136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_742
timestamp 1679581782
transform 1 0 71808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_749
timestamp 1679581782
transform 1 0 72480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_756
timestamp 1679581782
transform 1 0 73152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_763
timestamp 1679581782
transform 1 0 73824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_770
timestamp 1679581782
transform 1 0 74496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_777
timestamp 1679581782
transform 1 0 75168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_784
timestamp 1679581782
transform 1 0 75840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_791
timestamp 1679581782
transform 1 0 76512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_798
timestamp 1679581782
transform 1 0 77184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_805
timestamp 1679581782
transform 1 0 77856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_812
timestamp 1679581782
transform 1 0 78528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_819
timestamp 1679581782
transform 1 0 79200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_826
timestamp 1679581782
transform 1 0 79872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_833
timestamp 1679581782
transform 1 0 80544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_840
timestamp 1679581782
transform 1 0 81216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_847
timestamp 1679581782
transform 1 0 81888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_854
timestamp 1679581782
transform 1 0 82560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_861
timestamp 1679581782
transform 1 0 83232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_868
timestamp 1679581782
transform 1 0 83904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_875
timestamp 1679581782
transform 1 0 84576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_882
timestamp 1679581782
transform 1 0 85248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_889
timestamp 1679581782
transform 1 0 85920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_896
timestamp 1679581782
transform 1 0 86592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_903
timestamp 1679581782
transform 1 0 87264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_910
timestamp 1679581782
transform 1 0 87936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_917
timestamp 1679581782
transform 1 0 88608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_924
timestamp 1679581782
transform 1 0 89280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_931
timestamp 1679581782
transform 1 0 89952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_938
timestamp 1679581782
transform 1 0 90624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_945
timestamp 1679581782
transform 1 0 91296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_952
timestamp 1679581782
transform 1 0 91968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_959
timestamp 1679581782
transform 1 0 92640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_966
timestamp 1679581782
transform 1 0 93312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_973
timestamp 1679581782
transform 1 0 93984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_980
timestamp 1679581782
transform 1 0 94656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_987
timestamp 1679581782
transform 1 0 95328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_994
timestamp 1679581782
transform 1 0 96000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1001
timestamp 1679581782
transform 1 0 96672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1008
timestamp 1679581782
transform 1 0 97344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1015
timestamp 1679581782
transform 1 0 98016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1022
timestamp 1679581782
transform 1 0 98688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_18
timestamp 1679577901
transform 1 0 2304 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_22
timestamp 1677579658
transform 1 0 2688 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_27
timestamp 1679577901
transform 1 0 3168 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_31
timestamp 1677580104
transform 1 0 3552 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_66
timestamp 1679577901
transform 1 0 6912 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_70
timestamp 1677579658
transform 1 0 7296 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_109
timestamp 1677580104
transform 1 0 11040 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_111
timestamp 1677579658
transform 1 0 11232 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_132
timestamp 1677580104
transform 1 0 13248 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_134
timestamp 1677579658
transform 1 0 13440 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_203
timestamp 1677579658
transform 1 0 20064 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_213
timestamp 1677579658
transform 1 0 21024 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_233
timestamp 1677580104
transform 1 0 22944 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_240
timestamp 1677579658
transform 1 0 23616 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_246
timestamp 1679577901
transform 1 0 24192 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_250
timestamp 1677579658
transform 1 0 24576 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_264
timestamp 1679577901
transform 1 0 25920 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_281
timestamp 1679577901
transform 1 0 27552 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_285
timestamp 1677579658
transform 1 0 27936 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_302
timestamp 1677579658
transform 1 0 29568 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_316
timestamp 1677579658
transform 1 0 30912 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_323
timestamp 1677579658
transform 1 0 31584 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_338
timestamp 1677579658
transform 1 0 33024 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_402
timestamp 1679581782
transform 1 0 39168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_409
timestamp 1679581782
transform 1 0 39840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_416
timestamp 1679581782
transform 1 0 40512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_423
timestamp 1679581782
transform 1 0 41184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_430
timestamp 1679581782
transform 1 0 41856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_437
timestamp 1679581782
transform 1 0 42528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_444
timestamp 1679581782
transform 1 0 43200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_451
timestamp 1679581782
transform 1 0 43872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_458
timestamp 1679581782
transform 1 0 44544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_465
timestamp 1679581782
transform 1 0 45216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_472
timestamp 1679581782
transform 1 0 45888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_479
timestamp 1679581782
transform 1 0 46560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_486
timestamp 1679581782
transform 1 0 47232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_493
timestamp 1679581782
transform 1 0 47904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_500
timestamp 1679581782
transform 1 0 48576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_507
timestamp 1679581782
transform 1 0 49248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_514
timestamp 1679581782
transform 1 0 49920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_521
timestamp 1679581782
transform 1 0 50592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_528
timestamp 1679581782
transform 1 0 51264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_535
timestamp 1679581782
transform 1 0 51936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_542
timestamp 1679581782
transform 1 0 52608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_549
timestamp 1679581782
transform 1 0 53280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_556
timestamp 1679581782
transform 1 0 53952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_563
timestamp 1679581782
transform 1 0 54624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_570
timestamp 1679581782
transform 1 0 55296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_577
timestamp 1679581782
transform 1 0 55968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_584
timestamp 1679581782
transform 1 0 56640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_591
timestamp 1679581782
transform 1 0 57312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_598
timestamp 1679581782
transform 1 0 57984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_605
timestamp 1679581782
transform 1 0 58656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_612
timestamp 1679581782
transform 1 0 59328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_619
timestamp 1679581782
transform 1 0 60000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_626
timestamp 1679581782
transform 1 0 60672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_633
timestamp 1679581782
transform 1 0 61344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_640
timestamp 1679581782
transform 1 0 62016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_647
timestamp 1679581782
transform 1 0 62688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_654
timestamp 1679581782
transform 1 0 63360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_661
timestamp 1679581782
transform 1 0 64032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_668
timestamp 1679581782
transform 1 0 64704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_675
timestamp 1679581782
transform 1 0 65376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_682
timestamp 1679581782
transform 1 0 66048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_689
timestamp 1679581782
transform 1 0 66720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_696
timestamp 1679581782
transform 1 0 67392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_703
timestamp 1679581782
transform 1 0 68064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_710
timestamp 1679581782
transform 1 0 68736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_717
timestamp 1679581782
transform 1 0 69408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_724
timestamp 1679581782
transform 1 0 70080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_731
timestamp 1679581782
transform 1 0 70752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_738
timestamp 1679581782
transform 1 0 71424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_745
timestamp 1679581782
transform 1 0 72096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_752
timestamp 1679581782
transform 1 0 72768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_759
timestamp 1679581782
transform 1 0 73440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_766
timestamp 1679581782
transform 1 0 74112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_773
timestamp 1679581782
transform 1 0 74784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_780
timestamp 1679581782
transform 1 0 75456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_787
timestamp 1679581782
transform 1 0 76128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_794
timestamp 1679581782
transform 1 0 76800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_801
timestamp 1679581782
transform 1 0 77472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_808
timestamp 1679581782
transform 1 0 78144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_815
timestamp 1679581782
transform 1 0 78816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_822
timestamp 1679581782
transform 1 0 79488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_829
timestamp 1679581782
transform 1 0 80160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_836
timestamp 1679581782
transform 1 0 80832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_843
timestamp 1679581782
transform 1 0 81504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_850
timestamp 1679581782
transform 1 0 82176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_857
timestamp 1679581782
transform 1 0 82848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_864
timestamp 1679581782
transform 1 0 83520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_871
timestamp 1679581782
transform 1 0 84192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_878
timestamp 1679581782
transform 1 0 84864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_885
timestamp 1679581782
transform 1 0 85536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_892
timestamp 1679581782
transform 1 0 86208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_899
timestamp 1679581782
transform 1 0 86880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_906
timestamp 1679581782
transform 1 0 87552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_913
timestamp 1679581782
transform 1 0 88224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_920
timestamp 1679581782
transform 1 0 88896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_927
timestamp 1679581782
transform 1 0 89568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_934
timestamp 1679581782
transform 1 0 90240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_941
timestamp 1679581782
transform 1 0 90912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_948
timestamp 1679581782
transform 1 0 91584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_955
timestamp 1679581782
transform 1 0 92256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_962
timestamp 1679581782
transform 1 0 92928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_969
timestamp 1679581782
transform 1 0 93600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_976
timestamp 1679581782
transform 1 0 94272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_983
timestamp 1679581782
transform 1 0 94944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_990
timestamp 1679581782
transform 1 0 95616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_997
timestamp 1679581782
transform 1 0 96288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1004
timestamp 1679581782
transform 1 0 96960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1011
timestamp 1679581782
transform 1 0 97632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1018
timestamp 1679581782
transform 1 0 98304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_1025
timestamp 1679577901
transform 1 0 98976 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_25
timestamp 1679577901
transform 1 0 2976 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_61
timestamp 1677580104
transform 1 0 6432 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_90
timestamp 1677580104
transform 1 0 9216 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_106
timestamp 1677580104
transform 1 0 10752 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_144
timestamp 1677580104
transform 1 0 14400 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_165
timestamp 1677580104
transform 1 0 16416 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_185
timestamp 1679581782
transform 1 0 18336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_192
timestamp 1679581782
transform 1 0 19008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_216
timestamp 1679581782
transform 1 0 21312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_228
timestamp 1679577901
transform 1 0 22464 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_247
timestamp 1677580104
transform 1 0 24288 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_249
timestamp 1677579658
transform 1 0 24480 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_259
timestamp 1677579658
transform 1 0 25440 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679581782
transform 1 0 27456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_287
timestamp 1679577901
transform 1 0 28128 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_291
timestamp 1677580104
transform 1 0 28512 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_309
timestamp 1679581782
transform 1 0 30240 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_316
timestamp 1677579658
transform 1 0 30912 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_341
timestamp 1677579658
transform 1 0 33312 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_359
timestamp 1677580104
transform 1 0 35040 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_403
timestamp 1679581782
transform 1 0 39264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_410
timestamp 1679581782
transform 1 0 39936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_417
timestamp 1679581782
transform 1 0 40608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679581782
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679581782
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679581782
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679581782
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_452
timestamp 1679581782
transform 1 0 43968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679581782
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_466
timestamp 1679581782
transform 1 0 45312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_473
timestamp 1679581782
transform 1 0 45984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_480
timestamp 1679581782
transform 1 0 46656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_487
timestamp 1679581782
transform 1 0 47328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_494
timestamp 1679581782
transform 1 0 48000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_501
timestamp 1679581782
transform 1 0 48672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_508
timestamp 1679581782
transform 1 0 49344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679581782
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_522
timestamp 1679581782
transform 1 0 50688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_529
timestamp 1679581782
transform 1 0 51360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_536
timestamp 1679581782
transform 1 0 52032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_543
timestamp 1679581782
transform 1 0 52704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_550
timestamp 1679581782
transform 1 0 53376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_557
timestamp 1679581782
transform 1 0 54048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_564
timestamp 1679581782
transform 1 0 54720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_571
timestamp 1679581782
transform 1 0 55392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_578
timestamp 1679581782
transform 1 0 56064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_585
timestamp 1679581782
transform 1 0 56736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_592
timestamp 1679581782
transform 1 0 57408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_599
timestamp 1679581782
transform 1 0 58080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_606
timestamp 1679581782
transform 1 0 58752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_613
timestamp 1679581782
transform 1 0 59424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_620
timestamp 1679581782
transform 1 0 60096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679581782
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679581782
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679581782
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679581782
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_655
timestamp 1679581782
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_662
timestamp 1679581782
transform 1 0 64128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_669
timestamp 1679581782
transform 1 0 64800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_676
timestamp 1679581782
transform 1 0 65472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_683
timestamp 1679581782
transform 1 0 66144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679581782
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679581782
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_704
timestamp 1679581782
transform 1 0 68160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_711
timestamp 1679581782
transform 1 0 68832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_718
timestamp 1679581782
transform 1 0 69504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_725
timestamp 1679581782
transform 1 0 70176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_732
timestamp 1679581782
transform 1 0 70848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_739
timestamp 1679581782
transform 1 0 71520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_746
timestamp 1679581782
transform 1 0 72192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_753
timestamp 1679581782
transform 1 0 72864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_760
timestamp 1679581782
transform 1 0 73536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_767
timestamp 1679581782
transform 1 0 74208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_774
timestamp 1679581782
transform 1 0 74880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_781
timestamp 1679581782
transform 1 0 75552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_788
timestamp 1679581782
transform 1 0 76224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_795
timestamp 1679581782
transform 1 0 76896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_802
timestamp 1679581782
transform 1 0 77568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_809
timestamp 1679581782
transform 1 0 78240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_816
timestamp 1679581782
transform 1 0 78912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_823
timestamp 1679581782
transform 1 0 79584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_830
timestamp 1679581782
transform 1 0 80256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_837
timestamp 1679581782
transform 1 0 80928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_844
timestamp 1679581782
transform 1 0 81600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_851
timestamp 1679581782
transform 1 0 82272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_858
timestamp 1679581782
transform 1 0 82944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_865
timestamp 1679581782
transform 1 0 83616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_872
timestamp 1679581782
transform 1 0 84288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_879
timestamp 1679581782
transform 1 0 84960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_886
timestamp 1679581782
transform 1 0 85632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_893
timestamp 1679581782
transform 1 0 86304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_900
timestamp 1679581782
transform 1 0 86976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_907
timestamp 1679581782
transform 1 0 87648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_914
timestamp 1679581782
transform 1 0 88320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_921
timestamp 1679581782
transform 1 0 88992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_928
timestamp 1679581782
transform 1 0 89664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_935
timestamp 1679581782
transform 1 0 90336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_942
timestamp 1679581782
transform 1 0 91008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_949
timestamp 1679581782
transform 1 0 91680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_956
timestamp 1679581782
transform 1 0 92352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_963
timestamp 1679581782
transform 1 0 93024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_970
timestamp 1679581782
transform 1 0 93696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_977
timestamp 1679581782
transform 1 0 94368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_984
timestamp 1679581782
transform 1 0 95040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_991
timestamp 1679581782
transform 1 0 95712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_998
timestamp 1679581782
transform 1 0 96384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1005
timestamp 1679581782
transform 1 0 97056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1012
timestamp 1679581782
transform 1 0 97728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1019
timestamp 1679581782
transform 1 0 98400 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_1026
timestamp 1677580104
transform 1 0 99072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677579658
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_32
timestamp 1677580104
transform 1 0 3648 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_38
timestamp 1679581782
transform 1 0 4224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_45
timestamp 1679577901
transform 1 0 4896 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_49
timestamp 1677580104
transform 1 0 5280 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_95
timestamp 1677579658
transform 1 0 9696 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_104
timestamp 1679577901
transform 1 0 10560 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_167
timestamp 1677580104
transform 1 0 16608 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_169
timestamp 1677579658
transform 1 0 16800 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_192
timestamp 1679581782
transform 1 0 19008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_199
timestamp 1679577901
transform 1 0 19680 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_203
timestamp 1677579658
transform 1 0 20064 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_222
timestamp 1679577901
transform 1 0 21888 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_226
timestamp 1677579658
transform 1 0 22272 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_243
timestamp 1677579658
transform 1 0 23904 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_254
timestamp 1677580104
transform 1 0 24960 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_260
timestamp 1679581782
transform 1 0 25536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_267
timestamp 1679581782
transform 1 0 26208 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_274
timestamp 1677580104
transform 1 0 26880 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_276
timestamp 1677579658
transform 1 0 27072 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_286
timestamp 1677579658
transform 1 0 28032 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679581782
transform 1 0 30816 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_322
timestamp 1677580104
transform 1 0 31488 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_324
timestamp 1677579658
transform 1 0 31680 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_330
timestamp 1677580104
transform 1 0 32256 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_332
timestamp 1677579658
transform 1 0 32448 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_341
timestamp 1679581782
transform 1 0 33312 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_348
timestamp 1677579658
transform 1 0 33984 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_369
timestamp 1677580104
transform 1 0 36000 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_380
timestamp 1677580104
transform 1 0 37056 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_400
timestamp 1679581782
transform 1 0 38976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_407
timestamp 1679581782
transform 1 0 39648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_414
timestamp 1679581782
transform 1 0 40320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_421
timestamp 1679581782
transform 1 0 40992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_428
timestamp 1679581782
transform 1 0 41664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_435
timestamp 1679581782
transform 1 0 42336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_442
timestamp 1679581782
transform 1 0 43008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_449
timestamp 1679581782
transform 1 0 43680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_456
timestamp 1679581782
transform 1 0 44352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_463
timestamp 1679581782
transform 1 0 45024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_470
timestamp 1679581782
transform 1 0 45696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_477
timestamp 1679581782
transform 1 0 46368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_484
timestamp 1679581782
transform 1 0 47040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_491
timestamp 1679581782
transform 1 0 47712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_498
timestamp 1679581782
transform 1 0 48384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_505
timestamp 1679581782
transform 1 0 49056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_512
timestamp 1679581782
transform 1 0 49728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_519
timestamp 1679581782
transform 1 0 50400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_526
timestamp 1679581782
transform 1 0 51072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_533
timestamp 1679581782
transform 1 0 51744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_540
timestamp 1679581782
transform 1 0 52416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_547
timestamp 1679581782
transform 1 0 53088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_554
timestamp 1679581782
transform 1 0 53760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_561
timestamp 1679581782
transform 1 0 54432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_568
timestamp 1679581782
transform 1 0 55104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_575
timestamp 1679581782
transform 1 0 55776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_582
timestamp 1679581782
transform 1 0 56448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_589
timestamp 1679581782
transform 1 0 57120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_596
timestamp 1679581782
transform 1 0 57792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_603
timestamp 1679581782
transform 1 0 58464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_610
timestamp 1679581782
transform 1 0 59136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_617
timestamp 1679581782
transform 1 0 59808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_624
timestamp 1679581782
transform 1 0 60480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_631
timestamp 1679581782
transform 1 0 61152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_638
timestamp 1679581782
transform 1 0 61824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_645
timestamp 1679581782
transform 1 0 62496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_652
timestamp 1679581782
transform 1 0 63168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_659
timestamp 1679581782
transform 1 0 63840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_666
timestamp 1679581782
transform 1 0 64512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_673
timestamp 1679581782
transform 1 0 65184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_680
timestamp 1679581782
transform 1 0 65856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_687
timestamp 1679581782
transform 1 0 66528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_694
timestamp 1679581782
transform 1 0 67200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_701
timestamp 1679581782
transform 1 0 67872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_708
timestamp 1679581782
transform 1 0 68544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_715
timestamp 1679581782
transform 1 0 69216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_722
timestamp 1679581782
transform 1 0 69888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_729
timestamp 1679581782
transform 1 0 70560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_736
timestamp 1679581782
transform 1 0 71232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_743
timestamp 1679581782
transform 1 0 71904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_750
timestamp 1679581782
transform 1 0 72576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_757
timestamp 1679581782
transform 1 0 73248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_764
timestamp 1679581782
transform 1 0 73920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_771
timestamp 1679581782
transform 1 0 74592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_778
timestamp 1679581782
transform 1 0 75264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_785
timestamp 1679581782
transform 1 0 75936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_792
timestamp 1679581782
transform 1 0 76608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_799
timestamp 1679581782
transform 1 0 77280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_806
timestamp 1679581782
transform 1 0 77952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_813
timestamp 1679581782
transform 1 0 78624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_820
timestamp 1679581782
transform 1 0 79296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_827
timestamp 1679581782
transform 1 0 79968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_834
timestamp 1679581782
transform 1 0 80640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_841
timestamp 1679581782
transform 1 0 81312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_848
timestamp 1679581782
transform 1 0 81984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_855
timestamp 1679581782
transform 1 0 82656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_862
timestamp 1679581782
transform 1 0 83328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_869
timestamp 1679581782
transform 1 0 84000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_876
timestamp 1679581782
transform 1 0 84672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_883
timestamp 1679581782
transform 1 0 85344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_890
timestamp 1679581782
transform 1 0 86016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_897
timestamp 1679581782
transform 1 0 86688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_904
timestamp 1679581782
transform 1 0 87360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_911
timestamp 1679581782
transform 1 0 88032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_918
timestamp 1679581782
transform 1 0 88704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_925
timestamp 1679581782
transform 1 0 89376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_932
timestamp 1679581782
transform 1 0 90048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_939
timestamp 1679581782
transform 1 0 90720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_946
timestamp 1679581782
transform 1 0 91392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_953
timestamp 1679581782
transform 1 0 92064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_960
timestamp 1679581782
transform 1 0 92736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_967
timestamp 1679581782
transform 1 0 93408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_974
timestamp 1679581782
transform 1 0 94080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_981
timestamp 1679581782
transform 1 0 94752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_988
timestamp 1679581782
transform 1 0 95424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_995
timestamp 1679581782
transform 1 0 96096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1002
timestamp 1679581782
transform 1 0 96768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1009
timestamp 1679581782
transform 1 0 97440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1016
timestamp 1679581782
transform 1 0 98112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_1023
timestamp 1679577901
transform 1 0 98784 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_1027
timestamp 1677580104
transform 1 0 99168 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679581782
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679581782
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679581782
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679581782
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_53
timestamp 1677580104
transform 1 0 5664 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_55
timestamp 1677579658
transform 1 0 5856 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_60
timestamp 1677580104
transform 1 0 6336 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_136
timestamp 1679581782
transform 1 0 13632 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_143
timestamp 1677580104
transform 1 0 14304 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_145
timestamp 1677579658
transform 1 0 14496 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_159
timestamp 1677580104
transform 1 0 15840 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_207
timestamp 1677580104
transform 1 0 20448 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_259
timestamp 1679581782
transform 1 0 25440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_279
timestamp 1679581782
transform 1 0 27360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_286
timestamp 1679581782
transform 1 0 28032 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_293
timestamp 1677579658
transform 1 0 28704 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_312
timestamp 1677580104
transform 1 0 30528 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_322
timestamp 1679577901
transform 1 0 31488 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_326
timestamp 1677580104
transform 1 0 31872 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679581782
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_347
timestamp 1679577901
transform 1 0 33888 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_411
timestamp 1679581782
transform 1 0 40032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_418
timestamp 1679581782
transform 1 0 40704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_425
timestamp 1679581782
transform 1 0 41376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_432
timestamp 1679581782
transform 1 0 42048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_439
timestamp 1679581782
transform 1 0 42720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_446
timestamp 1679581782
transform 1 0 43392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_453
timestamp 1679581782
transform 1 0 44064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_460
timestamp 1679581782
transform 1 0 44736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_467
timestamp 1679581782
transform 1 0 45408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_474
timestamp 1679581782
transform 1 0 46080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_481
timestamp 1679581782
transform 1 0 46752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_488
timestamp 1679581782
transform 1 0 47424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_495
timestamp 1679581782
transform 1 0 48096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_502
timestamp 1679581782
transform 1 0 48768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_509
timestamp 1679581782
transform 1 0 49440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_516
timestamp 1679581782
transform 1 0 50112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_523
timestamp 1679581782
transform 1 0 50784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_530
timestamp 1679581782
transform 1 0 51456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_537
timestamp 1679581782
transform 1 0 52128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_544
timestamp 1679581782
transform 1 0 52800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_551
timestamp 1679581782
transform 1 0 53472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_558
timestamp 1679581782
transform 1 0 54144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_565
timestamp 1679581782
transform 1 0 54816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_572
timestamp 1679581782
transform 1 0 55488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_579
timestamp 1679581782
transform 1 0 56160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_586
timestamp 1679581782
transform 1 0 56832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_593
timestamp 1679581782
transform 1 0 57504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_600
timestamp 1679581782
transform 1 0 58176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_607
timestamp 1679581782
transform 1 0 58848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_614
timestamp 1679581782
transform 1 0 59520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_621
timestamp 1679581782
transform 1 0 60192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_628
timestamp 1679581782
transform 1 0 60864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_635
timestamp 1679581782
transform 1 0 61536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_642
timestamp 1679581782
transform 1 0 62208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_649
timestamp 1679581782
transform 1 0 62880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_656
timestamp 1679581782
transform 1 0 63552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_663
timestamp 1679581782
transform 1 0 64224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_670
timestamp 1679581782
transform 1 0 64896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_677
timestamp 1679581782
transform 1 0 65568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_684
timestamp 1679581782
transform 1 0 66240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_691
timestamp 1679581782
transform 1 0 66912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_698
timestamp 1679581782
transform 1 0 67584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_705
timestamp 1679581782
transform 1 0 68256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_712
timestamp 1679581782
transform 1 0 68928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_719
timestamp 1679581782
transform 1 0 69600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_726
timestamp 1679581782
transform 1 0 70272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_733
timestamp 1679581782
transform 1 0 70944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_740
timestamp 1679581782
transform 1 0 71616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_747
timestamp 1679581782
transform 1 0 72288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_754
timestamp 1679581782
transform 1 0 72960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_761
timestamp 1679581782
transform 1 0 73632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_768
timestamp 1679581782
transform 1 0 74304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_775
timestamp 1679581782
transform 1 0 74976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_782
timestamp 1679581782
transform 1 0 75648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_789
timestamp 1679581782
transform 1 0 76320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_796
timestamp 1679581782
transform 1 0 76992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_803
timestamp 1679581782
transform 1 0 77664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_810
timestamp 1679581782
transform 1 0 78336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_817
timestamp 1679581782
transform 1 0 79008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_824
timestamp 1679581782
transform 1 0 79680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_831
timestamp 1679581782
transform 1 0 80352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_838
timestamp 1679581782
transform 1 0 81024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_845
timestamp 1679581782
transform 1 0 81696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_852
timestamp 1679581782
transform 1 0 82368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_859
timestamp 1679581782
transform 1 0 83040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_866
timestamp 1679581782
transform 1 0 83712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_873
timestamp 1679581782
transform 1 0 84384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_880
timestamp 1679581782
transform 1 0 85056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_887
timestamp 1679581782
transform 1 0 85728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_894
timestamp 1679581782
transform 1 0 86400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_901
timestamp 1679581782
transform 1 0 87072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_908
timestamp 1679581782
transform 1 0 87744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_915
timestamp 1679581782
transform 1 0 88416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_922
timestamp 1679581782
transform 1 0 89088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_929
timestamp 1679581782
transform 1 0 89760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_936
timestamp 1679581782
transform 1 0 90432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_943
timestamp 1679581782
transform 1 0 91104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_950
timestamp 1679581782
transform 1 0 91776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_957
timestamp 1679581782
transform 1 0 92448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_964
timestamp 1679581782
transform 1 0 93120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_971
timestamp 1679581782
transform 1 0 93792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_978
timestamp 1679581782
transform 1 0 94464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_985
timestamp 1679581782
transform 1 0 95136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_992
timestamp 1679581782
transform 1 0 95808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_999
timestamp 1679581782
transform 1 0 96480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1006
timestamp 1679581782
transform 1 0 97152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1013
timestamp 1679581782
transform 1 0 97824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1020
timestamp 1679581782
transform 1 0 98496 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_1027
timestamp 1677580104
transform 1 0 99168 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679581782
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679581782
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679581782
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679581782
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679581782
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679581782
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679581782
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_67
timestamp 1677580104
transform 1 0 7008 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_96
timestamp 1677580104
transform 1 0 9792 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_121
timestamp 1677580104
transform 1 0 12192 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_141
timestamp 1679577901
transform 1 0 14112 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_145
timestamp 1677579658
transform 1 0 14496 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_165
timestamp 1679577901
transform 1 0 16416 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_198
timestamp 1677579658
transform 1 0 19584 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_230
timestamp 1679577901
transform 1 0 22656 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_234
timestamp 1677580104
transform 1 0 23040 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_243
timestamp 1677580104
transform 1 0 23904 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_258
timestamp 1677580104
transform 1 0 25344 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_260
timestamp 1677579658
transform 1 0 25536 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_281
timestamp 1679581782
transform 1 0 27552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_288
timestamp 1679577901
transform 1 0 28224 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_315
timestamp 1677580104
transform 1 0 30816 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_317
timestamp 1677579658
transform 1 0 31008 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_326
timestamp 1679577901
transform 1 0 31872 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_330
timestamp 1677579658
transform 1 0 32256 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_340
timestamp 1679581782
transform 1 0 33216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_347
timestamp 1679577901
transform 1 0 33888 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_399
timestamp 1679581782
transform 1 0 38880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_406
timestamp 1679581782
transform 1 0 39552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_413
timestamp 1679581782
transform 1 0 40224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_420
timestamp 1679581782
transform 1 0 40896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_427
timestamp 1679581782
transform 1 0 41568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_434
timestamp 1679581782
transform 1 0 42240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_441
timestamp 1679581782
transform 1 0 42912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_448
timestamp 1679581782
transform 1 0 43584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_455
timestamp 1679581782
transform 1 0 44256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_462
timestamp 1679581782
transform 1 0 44928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_469
timestamp 1679581782
transform 1 0 45600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_476
timestamp 1679581782
transform 1 0 46272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_483
timestamp 1679581782
transform 1 0 46944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_490
timestamp 1679581782
transform 1 0 47616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_497
timestamp 1679581782
transform 1 0 48288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_504
timestamp 1679581782
transform 1 0 48960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_511
timestamp 1679581782
transform 1 0 49632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_518
timestamp 1679581782
transform 1 0 50304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_525
timestamp 1679581782
transform 1 0 50976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_532
timestamp 1679581782
transform 1 0 51648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_539
timestamp 1679581782
transform 1 0 52320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_546
timestamp 1679581782
transform 1 0 52992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_553
timestamp 1679581782
transform 1 0 53664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_560
timestamp 1679581782
transform 1 0 54336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_567
timestamp 1679581782
transform 1 0 55008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_574
timestamp 1679581782
transform 1 0 55680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_581
timestamp 1679581782
transform 1 0 56352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_588
timestamp 1679581782
transform 1 0 57024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_595
timestamp 1679581782
transform 1 0 57696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_602
timestamp 1679581782
transform 1 0 58368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_609
timestamp 1679581782
transform 1 0 59040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_616
timestamp 1679581782
transform 1 0 59712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_623
timestamp 1679581782
transform 1 0 60384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_630
timestamp 1679581782
transform 1 0 61056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_637
timestamp 1679581782
transform 1 0 61728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_644
timestamp 1679581782
transform 1 0 62400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_651
timestamp 1679581782
transform 1 0 63072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_658
timestamp 1679581782
transform 1 0 63744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_665
timestamp 1679581782
transform 1 0 64416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_672
timestamp 1679581782
transform 1 0 65088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_679
timestamp 1679581782
transform 1 0 65760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_686
timestamp 1679581782
transform 1 0 66432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_693
timestamp 1679581782
transform 1 0 67104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_700
timestamp 1679581782
transform 1 0 67776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_707
timestamp 1679581782
transform 1 0 68448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_714
timestamp 1679581782
transform 1 0 69120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_721
timestamp 1679581782
transform 1 0 69792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_728
timestamp 1679581782
transform 1 0 70464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_735
timestamp 1679581782
transform 1 0 71136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_742
timestamp 1679581782
transform 1 0 71808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_749
timestamp 1679581782
transform 1 0 72480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_756
timestamp 1679581782
transform 1 0 73152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_763
timestamp 1679581782
transform 1 0 73824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_770
timestamp 1679581782
transform 1 0 74496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_777
timestamp 1679581782
transform 1 0 75168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_784
timestamp 1679581782
transform 1 0 75840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_791
timestamp 1679581782
transform 1 0 76512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_798
timestamp 1679581782
transform 1 0 77184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_805
timestamp 1679581782
transform 1 0 77856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_812
timestamp 1679581782
transform 1 0 78528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_819
timestamp 1679581782
transform 1 0 79200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_826
timestamp 1679581782
transform 1 0 79872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_833
timestamp 1679581782
transform 1 0 80544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_840
timestamp 1679581782
transform 1 0 81216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_847
timestamp 1679581782
transform 1 0 81888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_854
timestamp 1679581782
transform 1 0 82560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_861
timestamp 1679581782
transform 1 0 83232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_868
timestamp 1679581782
transform 1 0 83904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_875
timestamp 1679581782
transform 1 0 84576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_882
timestamp 1679581782
transform 1 0 85248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_889
timestamp 1679581782
transform 1 0 85920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_896
timestamp 1679581782
transform 1 0 86592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_903
timestamp 1679581782
transform 1 0 87264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_910
timestamp 1679581782
transform 1 0 87936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_917
timestamp 1679581782
transform 1 0 88608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_924
timestamp 1679581782
transform 1 0 89280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_931
timestamp 1679581782
transform 1 0 89952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_938
timestamp 1679581782
transform 1 0 90624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_945
timestamp 1679581782
transform 1 0 91296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_952
timestamp 1679581782
transform 1 0 91968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_959
timestamp 1679581782
transform 1 0 92640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_966
timestamp 1679581782
transform 1 0 93312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_973
timestamp 1679581782
transform 1 0 93984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_980
timestamp 1679581782
transform 1 0 94656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_987
timestamp 1679581782
transform 1 0 95328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_994
timestamp 1679581782
transform 1 0 96000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1001
timestamp 1679581782
transform 1 0 96672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1008
timestamp 1679581782
transform 1 0 97344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1015
timestamp 1679581782
transform 1 0 98016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1022
timestamp 1679581782
transform 1 0 98688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679581782
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679581782
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679581782
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_53
timestamp 1677580104
transform 1 0 5664 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_55
timestamp 1677579658
transform 1 0 5856 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_83
timestamp 1677579658
transform 1 0 8544 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_97
timestamp 1677579658
transform 1 0 9888 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_125
timestamp 1677580104
transform 1 0 12576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_141
timestamp 1677580104
transform 1 0 14112 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_143
timestamp 1677579658
transform 1 0 14304 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_171
timestamp 1679581782
transform 1 0 16992 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_178
timestamp 1677579658
transform 1 0 17664 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_187
timestamp 1679581782
transform 1 0 18528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_206
timestamp 1679581782
transform 1 0 20352 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_213
timestamp 1677579658
transform 1 0 21024 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_218
timestamp 1677580104
transform 1 0 21504 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_256
timestamp 1679577901
transform 1 0 25152 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_260
timestamp 1677580104
transform 1 0 25536 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_280
timestamp 1679581782
transform 1 0 27456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_287
timestamp 1679581782
transform 1 0 28128 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_294
timestamp 1677579658
transform 1 0 28800 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_323
timestamp 1679577901
transform 1 0 31584 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_327
timestamp 1677579658
transform 1 0 31968 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_352
timestamp 1679577901
transform 1 0 34368 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_408
timestamp 1679581782
transform 1 0 39744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_415
timestamp 1679581782
transform 1 0 40416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_422
timestamp 1679581782
transform 1 0 41088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_429
timestamp 1679581782
transform 1 0 41760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_436
timestamp 1679581782
transform 1 0 42432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_443
timestamp 1679581782
transform 1 0 43104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_450
timestamp 1679581782
transform 1 0 43776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_457
timestamp 1679581782
transform 1 0 44448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_464
timestamp 1679581782
transform 1 0 45120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_471
timestamp 1679581782
transform 1 0 45792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_478
timestamp 1679581782
transform 1 0 46464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_485
timestamp 1679581782
transform 1 0 47136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_492
timestamp 1679581782
transform 1 0 47808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_499
timestamp 1679581782
transform 1 0 48480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_506
timestamp 1679581782
transform 1 0 49152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_513
timestamp 1679581782
transform 1 0 49824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_520
timestamp 1679581782
transform 1 0 50496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_527
timestamp 1679581782
transform 1 0 51168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_534
timestamp 1679581782
transform 1 0 51840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_541
timestamp 1679581782
transform 1 0 52512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_548
timestamp 1679581782
transform 1 0 53184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_555
timestamp 1679581782
transform 1 0 53856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_562
timestamp 1679581782
transform 1 0 54528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_569
timestamp 1679581782
transform 1 0 55200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_576
timestamp 1679581782
transform 1 0 55872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_583
timestamp 1679581782
transform 1 0 56544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_590
timestamp 1679581782
transform 1 0 57216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_597
timestamp 1679581782
transform 1 0 57888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_604
timestamp 1679581782
transform 1 0 58560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_611
timestamp 1679581782
transform 1 0 59232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_618
timestamp 1679581782
transform 1 0 59904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_625
timestamp 1679581782
transform 1 0 60576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_632
timestamp 1679581782
transform 1 0 61248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_639
timestamp 1679581782
transform 1 0 61920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_646
timestamp 1679581782
transform 1 0 62592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_653
timestamp 1679581782
transform 1 0 63264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_660
timestamp 1679581782
transform 1 0 63936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_667
timestamp 1679581782
transform 1 0 64608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_674
timestamp 1679581782
transform 1 0 65280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_681
timestamp 1679581782
transform 1 0 65952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_688
timestamp 1679581782
transform 1 0 66624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_695
timestamp 1679581782
transform 1 0 67296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_702
timestamp 1679581782
transform 1 0 67968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_709
timestamp 1679581782
transform 1 0 68640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_716
timestamp 1679581782
transform 1 0 69312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_723
timestamp 1679581782
transform 1 0 69984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_730
timestamp 1679581782
transform 1 0 70656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_737
timestamp 1679581782
transform 1 0 71328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_744
timestamp 1679581782
transform 1 0 72000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_751
timestamp 1679581782
transform 1 0 72672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_758
timestamp 1679581782
transform 1 0 73344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679581782
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679581782
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679581782
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679581782
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679581782
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679581782
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679581782
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679581782
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_821
timestamp 1679581782
transform 1 0 79392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_828
timestamp 1679581782
transform 1 0 80064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_835
timestamp 1679581782
transform 1 0 80736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_842
timestamp 1679581782
transform 1 0 81408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_849
timestamp 1679581782
transform 1 0 82080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_856
timestamp 1679581782
transform 1 0 82752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_863
timestamp 1679581782
transform 1 0 83424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_870
timestamp 1679581782
transform 1 0 84096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_877
timestamp 1679581782
transform 1 0 84768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_884
timestamp 1679581782
transform 1 0 85440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_891
timestamp 1679581782
transform 1 0 86112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_898
timestamp 1679581782
transform 1 0 86784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_905
timestamp 1679581782
transform 1 0 87456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_912
timestamp 1679581782
transform 1 0 88128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_919
timestamp 1679581782
transform 1 0 88800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_926
timestamp 1679581782
transform 1 0 89472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_933
timestamp 1679581782
transform 1 0 90144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_940
timestamp 1679581782
transform 1 0 90816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_947
timestamp 1679581782
transform 1 0 91488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_954
timestamp 1679581782
transform 1 0 92160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_961
timestamp 1679581782
transform 1 0 92832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_968
timestamp 1679581782
transform 1 0 93504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_975
timestamp 1679581782
transform 1 0 94176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_982
timestamp 1679581782
transform 1 0 94848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_989
timestamp 1679581782
transform 1 0 95520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_996
timestamp 1679581782
transform 1 0 96192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1003
timestamp 1679581782
transform 1 0 96864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1010
timestamp 1679581782
transform 1 0 97536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1017
timestamp 1679581782
transform 1 0 98208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_1024
timestamp 1679577901
transform 1 0 98880 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_1028
timestamp 1677579658
transform 1 0 99264 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679581782
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_36
timestamp 1677579658
transform 1 0 4032 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_46
timestamp 1677579658
transform 1 0 4992 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_52
timestamp 1677579658
transform 1 0 5568 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_82
timestamp 1677579658
transform 1 0 8448 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_110
timestamp 1679577901
transform 1 0 11136 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_15_127
timestamp 1679577901
transform 1 0 12768 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_169
timestamp 1679581782
transform 1 0 16800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_176
timestamp 1679581782
transform 1 0 17472 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_183
timestamp 1677579658
transform 1 0 18144 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_207
timestamp 1677579658
transform 1 0 20448 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_227
timestamp 1679577901
transform 1 0 22368 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_231
timestamp 1677579658
transform 1 0 22752 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_236
timestamp 1679581782
transform 1 0 23232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_243
timestamp 1679581782
transform 1 0 23904 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_250
timestamp 1677579658
transform 1 0 24576 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_286
timestamp 1677580104
transform 1 0 28032 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_288
timestamp 1677579658
transform 1 0 28224 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_311
timestamp 1679581782
transform 1 0 30432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_318
timestamp 1679581782
transform 1 0 31104 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_325
timestamp 1677579658
transform 1 0 31776 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_357
timestamp 1679577901
transform 1 0 34848 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_361
timestamp 1677579658
transform 1 0 35232 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_387
timestamp 1677580104
transform 1 0 37728 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_389
timestamp 1677579658
transform 1 0 37920 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_403
timestamp 1679581782
transform 1 0 39264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_410
timestamp 1679581782
transform 1 0 39936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_417
timestamp 1679581782
transform 1 0 40608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_424
timestamp 1679581782
transform 1 0 41280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_431
timestamp 1679581782
transform 1 0 41952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_438
timestamp 1679581782
transform 1 0 42624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_445
timestamp 1679581782
transform 1 0 43296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_452
timestamp 1679581782
transform 1 0 43968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_459
timestamp 1679581782
transform 1 0 44640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_466
timestamp 1679581782
transform 1 0 45312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_473
timestamp 1679581782
transform 1 0 45984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_480
timestamp 1679581782
transform 1 0 46656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_487
timestamp 1679581782
transform 1 0 47328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_494
timestamp 1679581782
transform 1 0 48000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_501
timestamp 1679581782
transform 1 0 48672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_508
timestamp 1679581782
transform 1 0 49344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_515
timestamp 1679581782
transform 1 0 50016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_522
timestamp 1679581782
transform 1 0 50688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_529
timestamp 1679581782
transform 1 0 51360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_536
timestamp 1679581782
transform 1 0 52032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_543
timestamp 1679581782
transform 1 0 52704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_550
timestamp 1679581782
transform 1 0 53376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_557
timestamp 1679581782
transform 1 0 54048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_564
timestamp 1679581782
transform 1 0 54720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_571
timestamp 1679581782
transform 1 0 55392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_578
timestamp 1679581782
transform 1 0 56064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_585
timestamp 1679581782
transform 1 0 56736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_592
timestamp 1679581782
transform 1 0 57408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_599
timestamp 1679581782
transform 1 0 58080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_606
timestamp 1679581782
transform 1 0 58752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_613
timestamp 1679581782
transform 1 0 59424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_620
timestamp 1679581782
transform 1 0 60096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_627
timestamp 1679581782
transform 1 0 60768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_634
timestamp 1679581782
transform 1 0 61440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_641
timestamp 1679581782
transform 1 0 62112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_648
timestamp 1679581782
transform 1 0 62784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_655
timestamp 1679581782
transform 1 0 63456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_662
timestamp 1679581782
transform 1 0 64128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_669
timestamp 1679581782
transform 1 0 64800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_676
timestamp 1679581782
transform 1 0 65472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_683
timestamp 1679581782
transform 1 0 66144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_690
timestamp 1679581782
transform 1 0 66816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_697
timestamp 1679581782
transform 1 0 67488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_704
timestamp 1679581782
transform 1 0 68160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_711
timestamp 1679581782
transform 1 0 68832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_718
timestamp 1679581782
transform 1 0 69504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_725
timestamp 1679581782
transform 1 0 70176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_732
timestamp 1679581782
transform 1 0 70848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_739
timestamp 1679581782
transform 1 0 71520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_746
timestamp 1679581782
transform 1 0 72192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_753
timestamp 1679581782
transform 1 0 72864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_760
timestamp 1679581782
transform 1 0 73536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_767
timestamp 1679581782
transform 1 0 74208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_774
timestamp 1679581782
transform 1 0 74880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_781
timestamp 1679581782
transform 1 0 75552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_788
timestamp 1679581782
transform 1 0 76224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_795
timestamp 1679581782
transform 1 0 76896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_802
timestamp 1679581782
transform 1 0 77568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_809
timestamp 1679581782
transform 1 0 78240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_816
timestamp 1679581782
transform 1 0 78912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_823
timestamp 1679581782
transform 1 0 79584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_830
timestamp 1679581782
transform 1 0 80256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_837
timestamp 1679581782
transform 1 0 80928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_844
timestamp 1679581782
transform 1 0 81600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_851
timestamp 1679581782
transform 1 0 82272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_858
timestamp 1679581782
transform 1 0 82944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_865
timestamp 1679581782
transform 1 0 83616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_872
timestamp 1679581782
transform 1 0 84288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_879
timestamp 1679581782
transform 1 0 84960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_886
timestamp 1679581782
transform 1 0 85632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_893
timestamp 1679581782
transform 1 0 86304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_900
timestamp 1679581782
transform 1 0 86976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_907
timestamp 1679581782
transform 1 0 87648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_914
timestamp 1679581782
transform 1 0 88320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_921
timestamp 1679581782
transform 1 0 88992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_928
timestamp 1679581782
transform 1 0 89664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_935
timestamp 1679581782
transform 1 0 90336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_942
timestamp 1679581782
transform 1 0 91008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_949
timestamp 1679581782
transform 1 0 91680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_956
timestamp 1679581782
transform 1 0 92352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_963
timestamp 1679581782
transform 1 0 93024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_970
timestamp 1679581782
transform 1 0 93696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_977
timestamp 1679581782
transform 1 0 94368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_984
timestamp 1679581782
transform 1 0 95040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_991
timestamp 1679581782
transform 1 0 95712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_998
timestamp 1679581782
transform 1 0 96384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1005
timestamp 1679581782
transform 1 0 97056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1012
timestamp 1679581782
transform 1 0 97728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1019
timestamp 1679581782
transform 1 0 98400 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_1026
timestamp 1677580104
transform 1 0 99072 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_1028
timestamp 1677579658
transform 1 0 99264 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679581782
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_18
timestamp 1679581782
transform 1 0 2304 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_25
timestamp 1677580104
transform 1 0 2976 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_67
timestamp 1677579658
transform 1 0 7008 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_96
timestamp 1677580104
transform 1 0 9792 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_102
timestamp 1679581782
transform 1 0 10368 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_109
timestamp 1677579658
transform 1 0 11040 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_127
timestamp 1677580104
transform 1 0 12768 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_158
timestamp 1677580104
transform 1 0 15744 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_165
timestamp 1679577901
transform 1 0 16416 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_169
timestamp 1677579658
transform 1 0 16800 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_175
timestamp 1677580104
transform 1 0 17376 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_185
timestamp 1679581782
transform 1 0 18336 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_202
timestamp 1677579658
transform 1 0 19968 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_208
timestamp 1679577901
transform 1 0 20544 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_212
timestamp 1677579658
transform 1 0 20928 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_226
timestamp 1677579658
transform 1 0 22272 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_255
timestamp 1677580104
transform 1 0 25056 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_257
timestamp 1677579658
transform 1 0 25248 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_267
timestamp 1677580104
transform 1 0 26208 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_280
timestamp 1677580104
transform 1 0 27456 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_316
timestamp 1679577901
transform 1 0 30912 0 1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_16_325
timestamp 1679577901
transform 1 0 31776 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_334
timestamp 1677579658
transform 1 0 32640 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_373
timestamp 1679577901
transform 1 0 36384 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_377
timestamp 1677579658
transform 1 0 36768 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_406
timestamp 1679581782
transform 1 0 39552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_413
timestamp 1679581782
transform 1 0 40224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_420
timestamp 1679581782
transform 1 0 40896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_427
timestamp 1679581782
transform 1 0 41568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_434
timestamp 1679581782
transform 1 0 42240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_441
timestamp 1679581782
transform 1 0 42912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_448
timestamp 1679581782
transform 1 0 43584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_455
timestamp 1679581782
transform 1 0 44256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_462
timestamp 1679581782
transform 1 0 44928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_469
timestamp 1679581782
transform 1 0 45600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_476
timestamp 1679581782
transform 1 0 46272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_483
timestamp 1679581782
transform 1 0 46944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_490
timestamp 1679581782
transform 1 0 47616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_497
timestamp 1679581782
transform 1 0 48288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_504
timestamp 1679581782
transform 1 0 48960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_511
timestamp 1679581782
transform 1 0 49632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_518
timestamp 1679581782
transform 1 0 50304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_525
timestamp 1679581782
transform 1 0 50976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_532
timestamp 1679581782
transform 1 0 51648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_539
timestamp 1679581782
transform 1 0 52320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_546
timestamp 1679581782
transform 1 0 52992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_553
timestamp 1679581782
transform 1 0 53664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_560
timestamp 1679581782
transform 1 0 54336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_567
timestamp 1679581782
transform 1 0 55008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_574
timestamp 1679581782
transform 1 0 55680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_581
timestamp 1679581782
transform 1 0 56352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_588
timestamp 1679581782
transform 1 0 57024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_595
timestamp 1679581782
transform 1 0 57696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_602
timestamp 1679581782
transform 1 0 58368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679581782
transform 1 0 59040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679581782
transform 1 0 59712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_623
timestamp 1679581782
transform 1 0 60384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_630
timestamp 1679581782
transform 1 0 61056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_637
timestamp 1679581782
transform 1 0 61728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_644
timestamp 1679581782
transform 1 0 62400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_651
timestamp 1679581782
transform 1 0 63072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_658
timestamp 1679581782
transform 1 0 63744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_665
timestamp 1679581782
transform 1 0 64416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_672
timestamp 1679581782
transform 1 0 65088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_679
timestamp 1679581782
transform 1 0 65760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_686
timestamp 1679581782
transform 1 0 66432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_693
timestamp 1679581782
transform 1 0 67104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_700
timestamp 1679581782
transform 1 0 67776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_707
timestamp 1679581782
transform 1 0 68448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_714
timestamp 1679581782
transform 1 0 69120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_721
timestamp 1679581782
transform 1 0 69792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_728
timestamp 1679581782
transform 1 0 70464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_735
timestamp 1679581782
transform 1 0 71136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_742
timestamp 1679581782
transform 1 0 71808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_749
timestamp 1679581782
transform 1 0 72480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_756
timestamp 1679581782
transform 1 0 73152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_763
timestamp 1679581782
transform 1 0 73824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_770
timestamp 1679581782
transform 1 0 74496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_777
timestamp 1679581782
transform 1 0 75168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_784
timestamp 1679581782
transform 1 0 75840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_791
timestamp 1679581782
transform 1 0 76512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_798
timestamp 1679581782
transform 1 0 77184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_805
timestamp 1679581782
transform 1 0 77856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_812
timestamp 1679581782
transform 1 0 78528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_819
timestamp 1679581782
transform 1 0 79200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_826
timestamp 1679581782
transform 1 0 79872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_833
timestamp 1679581782
transform 1 0 80544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_840
timestamp 1679581782
transform 1 0 81216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_847
timestamp 1679581782
transform 1 0 81888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_854
timestamp 1679581782
transform 1 0 82560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_861
timestamp 1679581782
transform 1 0 83232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_868
timestamp 1679581782
transform 1 0 83904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_875
timestamp 1679581782
transform 1 0 84576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_882
timestamp 1679581782
transform 1 0 85248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_889
timestamp 1679581782
transform 1 0 85920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_896
timestamp 1679581782
transform 1 0 86592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_903
timestamp 1679581782
transform 1 0 87264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_910
timestamp 1679581782
transform 1 0 87936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_917
timestamp 1679581782
transform 1 0 88608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_924
timestamp 1679581782
transform 1 0 89280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_931
timestamp 1679581782
transform 1 0 89952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_938
timestamp 1679581782
transform 1 0 90624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_945
timestamp 1679581782
transform 1 0 91296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_952
timestamp 1679581782
transform 1 0 91968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_959
timestamp 1679581782
transform 1 0 92640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_966
timestamp 1679581782
transform 1 0 93312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_973
timestamp 1679581782
transform 1 0 93984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_980
timestamp 1679581782
transform 1 0 94656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_987
timestamp 1679581782
transform 1 0 95328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_994
timestamp 1679581782
transform 1 0 96000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1001
timestamp 1679581782
transform 1 0 96672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1008
timestamp 1679581782
transform 1 0 97344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1015
timestamp 1679581782
transform 1 0 98016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1022
timestamp 1679581782
transform 1 0 98688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_0
timestamp 1679577901
transform 1 0 576 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_32
timestamp 1677580104
transform 1 0 3648 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_83
timestamp 1677579658
transform 1 0 8544 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_182
timestamp 1679581782
transform 1 0 18048 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_210
timestamp 1677580104
transform 1 0 20736 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_217
timestamp 1677579658
transform 1 0 21408 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_236
timestamp 1679581782
transform 1 0 23232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_243
timestamp 1679581782
transform 1 0 23904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_250
timestamp 1679581782
transform 1 0 24576 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_257
timestamp 1677579658
transform 1 0 25248 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_268
timestamp 1679577901
transform 1 0 26304 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_293
timestamp 1677579658
transform 1 0 28704 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_308
timestamp 1679581782
transform 1 0 30144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_315
timestamp 1679581782
transform 1 0 30816 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_322
timestamp 1677580104
transform 1 0 31488 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_337
timestamp 1677580104
transform 1 0 32928 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_339
timestamp 1677579658
transform 1 0 33120 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_366
timestamp 1679581782
transform 1 0 35712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_373
timestamp 1679577901
transform 1 0 36384 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_417
timestamp 1679581782
transform 1 0 40608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_424
timestamp 1679581782
transform 1 0 41280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_431
timestamp 1679581782
transform 1 0 41952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_438
timestamp 1679581782
transform 1 0 42624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_445
timestamp 1679581782
transform 1 0 43296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_452
timestamp 1679581782
transform 1 0 43968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_459
timestamp 1679581782
transform 1 0 44640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_466
timestamp 1679581782
transform 1 0 45312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_473
timestamp 1679581782
transform 1 0 45984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_480
timestamp 1679581782
transform 1 0 46656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_487
timestamp 1679581782
transform 1 0 47328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_494
timestamp 1679581782
transform 1 0 48000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_501
timestamp 1679581782
transform 1 0 48672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_508
timestamp 1679581782
transform 1 0 49344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_515
timestamp 1679581782
transform 1 0 50016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_522
timestamp 1679581782
transform 1 0 50688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_529
timestamp 1679581782
transform 1 0 51360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_536
timestamp 1679581782
transform 1 0 52032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_543
timestamp 1679581782
transform 1 0 52704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_550
timestamp 1679581782
transform 1 0 53376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_557
timestamp 1679581782
transform 1 0 54048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_564
timestamp 1679581782
transform 1 0 54720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_571
timestamp 1679581782
transform 1 0 55392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_578
timestamp 1679581782
transform 1 0 56064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_585
timestamp 1679581782
transform 1 0 56736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_592
timestamp 1679581782
transform 1 0 57408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_599
timestamp 1679581782
transform 1 0 58080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_606
timestamp 1679581782
transform 1 0 58752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_613
timestamp 1679581782
transform 1 0 59424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_620
timestamp 1679581782
transform 1 0 60096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_627
timestamp 1679581782
transform 1 0 60768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_634
timestamp 1679581782
transform 1 0 61440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_641
timestamp 1679581782
transform 1 0 62112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_648
timestamp 1679581782
transform 1 0 62784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_655
timestamp 1679581782
transform 1 0 63456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_662
timestamp 1679581782
transform 1 0 64128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_669
timestamp 1679581782
transform 1 0 64800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_676
timestamp 1679581782
transform 1 0 65472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_683
timestamp 1679581782
transform 1 0 66144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_690
timestamp 1679581782
transform 1 0 66816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_697
timestamp 1679581782
transform 1 0 67488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_704
timestamp 1679581782
transform 1 0 68160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_711
timestamp 1679581782
transform 1 0 68832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_718
timestamp 1679581782
transform 1 0 69504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_725
timestamp 1679581782
transform 1 0 70176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_732
timestamp 1679581782
transform 1 0 70848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_739
timestamp 1679581782
transform 1 0 71520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_746
timestamp 1679581782
transform 1 0 72192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_753
timestamp 1679581782
transform 1 0 72864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_760
timestamp 1679581782
transform 1 0 73536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_767
timestamp 1679581782
transform 1 0 74208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_774
timestamp 1679581782
transform 1 0 74880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_781
timestamp 1679581782
transform 1 0 75552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_788
timestamp 1679581782
transform 1 0 76224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_795
timestamp 1679581782
transform 1 0 76896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_802
timestamp 1679581782
transform 1 0 77568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_809
timestamp 1679581782
transform 1 0 78240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_816
timestamp 1679581782
transform 1 0 78912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_823
timestamp 1679581782
transform 1 0 79584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_830
timestamp 1679581782
transform 1 0 80256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_837
timestamp 1679581782
transform 1 0 80928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_844
timestamp 1679581782
transform 1 0 81600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_851
timestamp 1679581782
transform 1 0 82272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_858
timestamp 1679581782
transform 1 0 82944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_865
timestamp 1679581782
transform 1 0 83616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_872
timestamp 1679581782
transform 1 0 84288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_879
timestamp 1679581782
transform 1 0 84960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_886
timestamp 1679581782
transform 1 0 85632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_893
timestamp 1679581782
transform 1 0 86304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_900
timestamp 1679581782
transform 1 0 86976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_907
timestamp 1679581782
transform 1 0 87648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_914
timestamp 1679581782
transform 1 0 88320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_921
timestamp 1679581782
transform 1 0 88992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_928
timestamp 1679581782
transform 1 0 89664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_935
timestamp 1679581782
transform 1 0 90336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_942
timestamp 1679581782
transform 1 0 91008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_949
timestamp 1679581782
transform 1 0 91680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_956
timestamp 1679581782
transform 1 0 92352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_963
timestamp 1679581782
transform 1 0 93024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_970
timestamp 1679581782
transform 1 0 93696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_977
timestamp 1679581782
transform 1 0 94368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_984
timestamp 1679581782
transform 1 0 95040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_991
timestamp 1679581782
transform 1 0 95712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_998
timestamp 1679581782
transform 1 0 96384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1005
timestamp 1679581782
transform 1 0 97056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1012
timestamp 1679581782
transform 1 0 97728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1019
timestamp 1679581782
transform 1 0 98400 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_1026
timestamp 1677580104
transform 1 0 99072 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_1028
timestamp 1677579658
transform 1 0 99264 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_8
timestamp 1677579658
transform 1 0 1344 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_13
timestamp 1679581782
transform 1 0 1824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_20
timestamp 1679577901
transform 1 0 2496 0 1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_18_81
timestamp 1679577901
transform 1 0 8352 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_103
timestamp 1679581782
transform 1 0 10464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_123
timestamp 1679581782
transform 1 0 12384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_130
timestamp 1679577901
transform 1 0 13056 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_134
timestamp 1677580104
transform 1 0 13440 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_141
timestamp 1677580104
transform 1 0 14112 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_189
timestamp 1679581782
transform 1 0 18720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_196
timestamp 1679577901
transform 1 0 19392 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_275
timestamp 1679581782
transform 1 0 26976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_282
timestamp 1679577901
transform 1 0 27648 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_298
timestamp 1677579658
transform 1 0 29184 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_304
timestamp 1677580104
transform 1 0 29760 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_311
timestamp 1679581782
transform 1 0 30432 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_318
timestamp 1677580104
transform 1 0 31104 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_354
timestamp 1679581782
transform 1 0 34560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_361
timestamp 1679577901
transform 1 0 35232 0 1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_18_376
timestamp 1679577901
transform 1 0 36672 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_393
timestamp 1677580104
transform 1 0 38304 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_395
timestamp 1677579658
transform 1 0 38496 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_400
timestamp 1677579658
transform 1 0 38976 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_429
timestamp 1679581782
transform 1 0 41760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_436
timestamp 1679581782
transform 1 0 42432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_443
timestamp 1679581782
transform 1 0 43104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_450
timestamp 1679581782
transform 1 0 43776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_457
timestamp 1679581782
transform 1 0 44448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_464
timestamp 1679581782
transform 1 0 45120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_471
timestamp 1679581782
transform 1 0 45792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_478
timestamp 1679581782
transform 1 0 46464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_485
timestamp 1679581782
transform 1 0 47136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_492
timestamp 1679581782
transform 1 0 47808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_499
timestamp 1679581782
transform 1 0 48480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_506
timestamp 1679581782
transform 1 0 49152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_513
timestamp 1679581782
transform 1 0 49824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_520
timestamp 1679581782
transform 1 0 50496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_527
timestamp 1679581782
transform 1 0 51168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_534
timestamp 1679581782
transform 1 0 51840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_541
timestamp 1679581782
transform 1 0 52512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_548
timestamp 1679581782
transform 1 0 53184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_555
timestamp 1679581782
transform 1 0 53856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_562
timestamp 1679581782
transform 1 0 54528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_569
timestamp 1679581782
transform 1 0 55200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_576
timestamp 1679581782
transform 1 0 55872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_583
timestamp 1679581782
transform 1 0 56544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_590
timestamp 1679581782
transform 1 0 57216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_597
timestamp 1679581782
transform 1 0 57888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_604
timestamp 1679581782
transform 1 0 58560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_611
timestamp 1679581782
transform 1 0 59232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_618
timestamp 1679581782
transform 1 0 59904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_625
timestamp 1679581782
transform 1 0 60576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_632
timestamp 1679581782
transform 1 0 61248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_639
timestamp 1679581782
transform 1 0 61920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_646
timestamp 1679581782
transform 1 0 62592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_653
timestamp 1679581782
transform 1 0 63264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_660
timestamp 1679581782
transform 1 0 63936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_667
timestamp 1679581782
transform 1 0 64608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_674
timestamp 1679581782
transform 1 0 65280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_681
timestamp 1679581782
transform 1 0 65952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_688
timestamp 1679581782
transform 1 0 66624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_695
timestamp 1679581782
transform 1 0 67296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_702
timestamp 1679581782
transform 1 0 67968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_709
timestamp 1679581782
transform 1 0 68640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_716
timestamp 1679581782
transform 1 0 69312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_723
timestamp 1679581782
transform 1 0 69984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_730
timestamp 1679581782
transform 1 0 70656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_737
timestamp 1679581782
transform 1 0 71328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_744
timestamp 1679581782
transform 1 0 72000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_751
timestamp 1679581782
transform 1 0 72672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_758
timestamp 1679581782
transform 1 0 73344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_765
timestamp 1679581782
transform 1 0 74016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_772
timestamp 1679581782
transform 1 0 74688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_779
timestamp 1679581782
transform 1 0 75360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_786
timestamp 1679581782
transform 1 0 76032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_793
timestamp 1679581782
transform 1 0 76704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_800
timestamp 1679581782
transform 1 0 77376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_807
timestamp 1679581782
transform 1 0 78048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_821
timestamp 1679581782
transform 1 0 79392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_828
timestamp 1679581782
transform 1 0 80064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_835
timestamp 1679581782
transform 1 0 80736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_842
timestamp 1679581782
transform 1 0 81408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_849
timestamp 1679581782
transform 1 0 82080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_856
timestamp 1679581782
transform 1 0 82752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_863
timestamp 1679581782
transform 1 0 83424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_870
timestamp 1679581782
transform 1 0 84096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_877
timestamp 1679581782
transform 1 0 84768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_884
timestamp 1679581782
transform 1 0 85440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_891
timestamp 1679581782
transform 1 0 86112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_898
timestamp 1679581782
transform 1 0 86784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_905
timestamp 1679581782
transform 1 0 87456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_912
timestamp 1679581782
transform 1 0 88128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_919
timestamp 1679581782
transform 1 0 88800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_926
timestamp 1679581782
transform 1 0 89472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_933
timestamp 1679581782
transform 1 0 90144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_940
timestamp 1679581782
transform 1 0 90816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_947
timestamp 1679581782
transform 1 0 91488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_954
timestamp 1679581782
transform 1 0 92160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_961
timestamp 1679581782
transform 1 0 92832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_968
timestamp 1679581782
transform 1 0 93504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_975
timestamp 1679581782
transform 1 0 94176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_982
timestamp 1679581782
transform 1 0 94848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_989
timestamp 1679581782
transform 1 0 95520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_996
timestamp 1679581782
transform 1 0 96192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1003
timestamp 1679581782
transform 1 0 96864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1010
timestamp 1679581782
transform 1 0 97536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1017
timestamp 1679581782
transform 1 0 98208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_1024
timestamp 1679577901
transform 1 0 98880 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_1028
timestamp 1677579658
transform 1 0 99264 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_0
timestamp 1677580104
transform 1 0 576 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_2
timestamp 1677579658
transform 1 0 768 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_31
timestamp 1677580104
transform 1 0 3552 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_67
timestamp 1677579658
transform 1 0 7008 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_117
timestamp 1679581782
transform 1 0 11808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_124
timestamp 1679577901
transform 1 0 12480 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_173
timestamp 1679581782
transform 1 0 17184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_180
timestamp 1679581782
transform 1 0 17856 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_207
timestamp 1677580104
transform 1 0 20448 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_236
timestamp 1677580104
transform 1 0 23232 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_238
timestamp 1677579658
transform 1 0 23424 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_248
timestamp 1677580104
transform 1 0 24384 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_250
timestamp 1677579658
transform 1 0 24576 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_268
timestamp 1679581782
transform 1 0 26304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_275
timestamp 1679577901
transform 1 0 26976 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_308
timestamp 1677580104
transform 1 0 30144 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_310
timestamp 1677579658
transform 1 0 30336 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_314
timestamp 1679581782
transform 1 0 30720 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_321
timestamp 1677579658
transform 1 0 31392 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_338
timestamp 1677580104
transform 1 0 33024 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_340
timestamp 1677579658
transform 1 0 33216 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_360
timestamp 1677580104
transform 1 0 35136 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_382
timestamp 1677579658
transform 1 0 37248 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_418
timestamp 1679581782
transform 1 0 40704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_425
timestamp 1679581782
transform 1 0 41376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_432
timestamp 1679581782
transform 1 0 42048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_439
timestamp 1679581782
transform 1 0 42720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_446
timestamp 1679581782
transform 1 0 43392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_453
timestamp 1679581782
transform 1 0 44064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_460
timestamp 1679581782
transform 1 0 44736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_467
timestamp 1679581782
transform 1 0 45408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_474
timestamp 1679581782
transform 1 0 46080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_481
timestamp 1679581782
transform 1 0 46752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_488
timestamp 1679581782
transform 1 0 47424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_495
timestamp 1679581782
transform 1 0 48096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_502
timestamp 1679581782
transform 1 0 48768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_509
timestamp 1679581782
transform 1 0 49440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_516
timestamp 1679581782
transform 1 0 50112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_523
timestamp 1679581782
transform 1 0 50784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_530
timestamp 1679581782
transform 1 0 51456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_537
timestamp 1679581782
transform 1 0 52128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_544
timestamp 1679581782
transform 1 0 52800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_551
timestamp 1679581782
transform 1 0 53472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_558
timestamp 1679581782
transform 1 0 54144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_565
timestamp 1679581782
transform 1 0 54816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_572
timestamp 1679581782
transform 1 0 55488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_579
timestamp 1679581782
transform 1 0 56160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_586
timestamp 1679581782
transform 1 0 56832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_593
timestamp 1679581782
transform 1 0 57504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_600
timestamp 1679581782
transform 1 0 58176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_607
timestamp 1679581782
transform 1 0 58848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_614
timestamp 1679581782
transform 1 0 59520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_621
timestamp 1679581782
transform 1 0 60192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_628
timestamp 1679581782
transform 1 0 60864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_635
timestamp 1679581782
transform 1 0 61536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_642
timestamp 1679581782
transform 1 0 62208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_649
timestamp 1679581782
transform 1 0 62880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_656
timestamp 1679581782
transform 1 0 63552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_663
timestamp 1679581782
transform 1 0 64224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_670
timestamp 1679581782
transform 1 0 64896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_677
timestamp 1679581782
transform 1 0 65568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_684
timestamp 1679581782
transform 1 0 66240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_691
timestamp 1679581782
transform 1 0 66912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_698
timestamp 1679581782
transform 1 0 67584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_705
timestamp 1679581782
transform 1 0 68256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_712
timestamp 1679581782
transform 1 0 68928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_719
timestamp 1679581782
transform 1 0 69600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_726
timestamp 1679581782
transform 1 0 70272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_733
timestamp 1679581782
transform 1 0 70944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_740
timestamp 1679581782
transform 1 0 71616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_747
timestamp 1679581782
transform 1 0 72288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_754
timestamp 1679581782
transform 1 0 72960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_761
timestamp 1679581782
transform 1 0 73632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_768
timestamp 1679581782
transform 1 0 74304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_775
timestamp 1679581782
transform 1 0 74976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_782
timestamp 1679581782
transform 1 0 75648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_789
timestamp 1679581782
transform 1 0 76320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_796
timestamp 1679581782
transform 1 0 76992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_803
timestamp 1679581782
transform 1 0 77664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_810
timestamp 1679581782
transform 1 0 78336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_817
timestamp 1679581782
transform 1 0 79008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_824
timestamp 1679581782
transform 1 0 79680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_831
timestamp 1679581782
transform 1 0 80352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_838
timestamp 1679581782
transform 1 0 81024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_845
timestamp 1679581782
transform 1 0 81696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_852
timestamp 1679581782
transform 1 0 82368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_859
timestamp 1679581782
transform 1 0 83040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_866
timestamp 1679581782
transform 1 0 83712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_873
timestamp 1679581782
transform 1 0 84384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_880
timestamp 1679581782
transform 1 0 85056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_887
timestamp 1679581782
transform 1 0 85728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_894
timestamp 1679581782
transform 1 0 86400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_901
timestamp 1679581782
transform 1 0 87072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_908
timestamp 1679581782
transform 1 0 87744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_915
timestamp 1679581782
transform 1 0 88416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_922
timestamp 1679581782
transform 1 0 89088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_929
timestamp 1679581782
transform 1 0 89760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_936
timestamp 1679581782
transform 1 0 90432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_943
timestamp 1679581782
transform 1 0 91104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_950
timestamp 1679581782
transform 1 0 91776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_957
timestamp 1679581782
transform 1 0 92448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_964
timestamp 1679581782
transform 1 0 93120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_971
timestamp 1679581782
transform 1 0 93792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_978
timestamp 1679581782
transform 1 0 94464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_985
timestamp 1679581782
transform 1 0 95136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_992
timestamp 1679581782
transform 1 0 95808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_999
timestamp 1679581782
transform 1 0 96480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1006
timestamp 1679581782
transform 1 0 97152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1013
timestamp 1679581782
transform 1 0 97824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1020
timestamp 1679581782
transform 1 0 98496 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_1027
timestamp 1677580104
transform 1 0 99168 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_4
timestamp 1679577901
transform 1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_12
timestamp 1679581782
transform 1 0 1728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_19
timestamp 1679577901
transform 1 0 2400 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_23
timestamp 1677580104
transform 1 0 2784 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_34
timestamp 1677579658
transform 1 0 3840 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_44
timestamp 1677579658
transform 1 0 4800 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_49
timestamp 1677579658
transform 1 0 5280 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_65
timestamp 1677579658
transform 1 0 6816 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_74
timestamp 1677579658
transform 1 0 7680 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_84
timestamp 1679581782
transform 1 0 8640 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_118
timestamp 1677579658
transform 1 0 11904 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_124
timestamp 1677580104
transform 1 0 12480 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_126
timestamp 1677579658
transform 1 0 12672 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_151
timestamp 1677579658
transform 1 0 15072 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_169
timestamp 1679581782
transform 1 0 16800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_176
timestamp 1679581782
transform 1 0 17472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_183
timestamp 1679577901
transform 1 0 18144 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_220
timestamp 1677579658
transform 1 0 21696 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_254
timestamp 1679581782
transform 1 0 24960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_261
timestamp 1679577901
transform 1 0 25632 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_265
timestamp 1677579658
transform 1 0 26016 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_294
timestamp 1677579658
transform 1 0 28800 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_300
timestamp 1679577901
transform 1 0 29376 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_350
timestamp 1677580104
transform 1 0 34176 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_352
timestamp 1677579658
transform 1 0 34368 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_376
timestamp 1677580104
transform 1 0 36672 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_387
timestamp 1677580104
transform 1 0 37728 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_396
timestamp 1677580104
transform 1 0 38592 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_398
timestamp 1677579658
transform 1 0 38784 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_426
timestamp 1679581782
transform 1 0 41472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_433
timestamp 1679581782
transform 1 0 42144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_440
timestamp 1679581782
transform 1 0 42816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_447
timestamp 1679581782
transform 1 0 43488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_454
timestamp 1679581782
transform 1 0 44160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_461
timestamp 1679581782
transform 1 0 44832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_468
timestamp 1679581782
transform 1 0 45504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_475
timestamp 1679581782
transform 1 0 46176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_482
timestamp 1679581782
transform 1 0 46848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_489
timestamp 1679581782
transform 1 0 47520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_496
timestamp 1679581782
transform 1 0 48192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_503
timestamp 1679581782
transform 1 0 48864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_510
timestamp 1679581782
transform 1 0 49536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_517
timestamp 1679581782
transform 1 0 50208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_524
timestamp 1679581782
transform 1 0 50880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_531
timestamp 1679581782
transform 1 0 51552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_538
timestamp 1679581782
transform 1 0 52224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_545
timestamp 1679581782
transform 1 0 52896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_552
timestamp 1679581782
transform 1 0 53568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_559
timestamp 1679581782
transform 1 0 54240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_566
timestamp 1679581782
transform 1 0 54912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_573
timestamp 1679581782
transform 1 0 55584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_580
timestamp 1679581782
transform 1 0 56256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_587
timestamp 1679581782
transform 1 0 56928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_594
timestamp 1679581782
transform 1 0 57600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_601
timestamp 1679581782
transform 1 0 58272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_608
timestamp 1679581782
transform 1 0 58944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_615
timestamp 1679581782
transform 1 0 59616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_622
timestamp 1679581782
transform 1 0 60288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_629
timestamp 1679581782
transform 1 0 60960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_636
timestamp 1679581782
transform 1 0 61632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_643
timestamp 1679581782
transform 1 0 62304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_650
timestamp 1679581782
transform 1 0 62976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_657
timestamp 1679581782
transform 1 0 63648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_664
timestamp 1679581782
transform 1 0 64320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_671
timestamp 1679581782
transform 1 0 64992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_678
timestamp 1679581782
transform 1 0 65664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_685
timestamp 1679581782
transform 1 0 66336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_692
timestamp 1679581782
transform 1 0 67008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_699
timestamp 1679581782
transform 1 0 67680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_706
timestamp 1679581782
transform 1 0 68352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_713
timestamp 1679581782
transform 1 0 69024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_720
timestamp 1679581782
transform 1 0 69696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_727
timestamp 1679581782
transform 1 0 70368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_734
timestamp 1679581782
transform 1 0 71040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_741
timestamp 1679581782
transform 1 0 71712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_748
timestamp 1679581782
transform 1 0 72384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_755
timestamp 1679581782
transform 1 0 73056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_762
timestamp 1679581782
transform 1 0 73728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_769
timestamp 1679581782
transform 1 0 74400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_776
timestamp 1679581782
transform 1 0 75072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_783
timestamp 1679581782
transform 1 0 75744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_790
timestamp 1679581782
transform 1 0 76416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_797
timestamp 1679581782
transform 1 0 77088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_804
timestamp 1679581782
transform 1 0 77760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_811
timestamp 1679581782
transform 1 0 78432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_818
timestamp 1679581782
transform 1 0 79104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_825
timestamp 1679581782
transform 1 0 79776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_832
timestamp 1679581782
transform 1 0 80448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_839
timestamp 1679581782
transform 1 0 81120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_846
timestamp 1679581782
transform 1 0 81792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_853
timestamp 1679581782
transform 1 0 82464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_860
timestamp 1679581782
transform 1 0 83136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_867
timestamp 1679581782
transform 1 0 83808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_874
timestamp 1679581782
transform 1 0 84480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_881
timestamp 1679581782
transform 1 0 85152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_888
timestamp 1679581782
transform 1 0 85824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_895
timestamp 1679581782
transform 1 0 86496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_902
timestamp 1679581782
transform 1 0 87168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_909
timestamp 1679581782
transform 1 0 87840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_916
timestamp 1679581782
transform 1 0 88512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_923
timestamp 1679581782
transform 1 0 89184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_930
timestamp 1679581782
transform 1 0 89856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_937
timestamp 1679581782
transform 1 0 90528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_944
timestamp 1679581782
transform 1 0 91200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_951
timestamp 1679581782
transform 1 0 91872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_958
timestamp 1679581782
transform 1 0 92544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_965
timestamp 1679581782
transform 1 0 93216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_972
timestamp 1679581782
transform 1 0 93888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_979
timestamp 1679581782
transform 1 0 94560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_986
timestamp 1679581782
transform 1 0 95232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_993
timestamp 1679581782
transform 1 0 95904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1000
timestamp 1679581782
transform 1 0 96576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1007
timestamp 1679581782
transform 1 0 97248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1014
timestamp 1679581782
transform 1 0 97920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1021
timestamp 1679581782
transform 1 0 98592 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_1028
timestamp 1677579658
transform 1 0 99264 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679581782
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_25
timestamp 1677580104
transform 1 0 2976 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_49
timestamp 1677580104
transform 1 0 5280 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_51
timestamp 1677579658
transform 1 0 5472 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_84
timestamp 1679581782
transform 1 0 8640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_91
timestamp 1679577901
transform 1 0 9312 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_95
timestamp 1677579658
transform 1 0 9696 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_100
timestamp 1677580104
transform 1 0 10176 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_102
timestamp 1677579658
transform 1 0 10368 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_138
timestamp 1677580104
transform 1 0 13824 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_140
timestamp 1677579658
transform 1 0 14016 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_182
timestamp 1677580104
transform 1 0 18048 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_193
timestamp 1677580104
transform 1 0 19104 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_204
timestamp 1677579658
transform 1 0 20160 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_252
timestamp 1679577901
transform 1 0 24768 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_261
timestamp 1679581782
transform 1 0 25632 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_268
timestamp 1677579658
transform 1 0 26304 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_289
timestamp 1677580104
transform 1 0 28320 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_291
timestamp 1677579658
transform 1 0 28512 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_313
timestamp 1679577901
transform 1 0 30624 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_21_361
timestamp 1679577901
transform 1 0 35232 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_365
timestamp 1677580104
transform 1 0 35616 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_437
timestamp 1679581782
transform 1 0 42528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_444
timestamp 1679581782
transform 1 0 43200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_451
timestamp 1679581782
transform 1 0 43872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_458
timestamp 1679581782
transform 1 0 44544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_465
timestamp 1679581782
transform 1 0 45216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_472
timestamp 1679581782
transform 1 0 45888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_479
timestamp 1679581782
transform 1 0 46560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_486
timestamp 1679581782
transform 1 0 47232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_493
timestamp 1679581782
transform 1 0 47904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_500
timestamp 1679581782
transform 1 0 48576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_507
timestamp 1679581782
transform 1 0 49248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_514
timestamp 1679581782
transform 1 0 49920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_521
timestamp 1679581782
transform 1 0 50592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_528
timestamp 1679581782
transform 1 0 51264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_535
timestamp 1679581782
transform 1 0 51936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_542
timestamp 1679581782
transform 1 0 52608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_549
timestamp 1679581782
transform 1 0 53280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_556
timestamp 1679581782
transform 1 0 53952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_563
timestamp 1679581782
transform 1 0 54624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_570
timestamp 1679581782
transform 1 0 55296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_577
timestamp 1679581782
transform 1 0 55968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_584
timestamp 1679581782
transform 1 0 56640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_591
timestamp 1679581782
transform 1 0 57312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_598
timestamp 1679581782
transform 1 0 57984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_605
timestamp 1679581782
transform 1 0 58656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_612
timestamp 1679581782
transform 1 0 59328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_619
timestamp 1679581782
transform 1 0 60000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_626
timestamp 1679581782
transform 1 0 60672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_633
timestamp 1679581782
transform 1 0 61344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_640
timestamp 1679581782
transform 1 0 62016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_647
timestamp 1679581782
transform 1 0 62688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_654
timestamp 1679581782
transform 1 0 63360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_661
timestamp 1679581782
transform 1 0 64032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_668
timestamp 1679581782
transform 1 0 64704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_675
timestamp 1679581782
transform 1 0 65376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_682
timestamp 1679581782
transform 1 0 66048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_689
timestamp 1679581782
transform 1 0 66720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_696
timestamp 1679581782
transform 1 0 67392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_703
timestamp 1679581782
transform 1 0 68064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_710
timestamp 1679581782
transform 1 0 68736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_717
timestamp 1679581782
transform 1 0 69408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_724
timestamp 1679581782
transform 1 0 70080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_731
timestamp 1679581782
transform 1 0 70752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_738
timestamp 1679581782
transform 1 0 71424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_745
timestamp 1679581782
transform 1 0 72096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_752
timestamp 1679581782
transform 1 0 72768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_759
timestamp 1679581782
transform 1 0 73440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_766
timestamp 1679581782
transform 1 0 74112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_773
timestamp 1679581782
transform 1 0 74784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_780
timestamp 1679581782
transform 1 0 75456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_787
timestamp 1679581782
transform 1 0 76128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_794
timestamp 1679581782
transform 1 0 76800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_801
timestamp 1679581782
transform 1 0 77472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_808
timestamp 1679581782
transform 1 0 78144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_815
timestamp 1679581782
transform 1 0 78816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_822
timestamp 1679581782
transform 1 0 79488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_829
timestamp 1679581782
transform 1 0 80160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_836
timestamp 1679581782
transform 1 0 80832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_843
timestamp 1679581782
transform 1 0 81504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_850
timestamp 1679581782
transform 1 0 82176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_857
timestamp 1679581782
transform 1 0 82848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_864
timestamp 1679581782
transform 1 0 83520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_871
timestamp 1679581782
transform 1 0 84192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_878
timestamp 1679581782
transform 1 0 84864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_885
timestamp 1679581782
transform 1 0 85536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_892
timestamp 1679581782
transform 1 0 86208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_899
timestamp 1679581782
transform 1 0 86880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_906
timestamp 1679581782
transform 1 0 87552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_913
timestamp 1679581782
transform 1 0 88224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_920
timestamp 1679581782
transform 1 0 88896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_927
timestamp 1679581782
transform 1 0 89568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_934
timestamp 1679581782
transform 1 0 90240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_941
timestamp 1679581782
transform 1 0 90912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_948
timestamp 1679581782
transform 1 0 91584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_955
timestamp 1679581782
transform 1 0 92256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_962
timestamp 1679581782
transform 1 0 92928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_969
timestamp 1679581782
transform 1 0 93600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_976
timestamp 1679581782
transform 1 0 94272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_983
timestamp 1679581782
transform 1 0 94944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_990
timestamp 1679581782
transform 1 0 95616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_997
timestamp 1679581782
transform 1 0 96288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1004
timestamp 1679581782
transform 1 0 96960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1011
timestamp 1679581782
transform 1 0 97632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1018
timestamp 1679581782
transform 1 0 98304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1025
timestamp 1679577901
transform 1 0 98976 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_4
timestamp 1677579658
transform 1 0 960 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_36
timestamp 1677580104
transform 1 0 4032 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_38
timestamp 1677579658
transform 1 0 4224 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_80
timestamp 1677579658
transform 1 0 8256 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_113
timestamp 1677580104
transform 1 0 11424 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_152
timestamp 1679577901
transform 1 0 15168 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_156
timestamp 1677580104
transform 1 0 15552 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_171
timestamp 1679581782
transform 1 0 16992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_206
timestamp 1679577901
transform 1 0 20352 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_255
timestamp 1679581782
transform 1 0 25056 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_262
timestamp 1677580104
transform 1 0 25728 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_264
timestamp 1677579658
transform 1 0 25920 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_274
timestamp 1677579658
transform 1 0 26880 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_328
timestamp 1677580104
transform 1 0 32064 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_343
timestamp 1679577901
transform 1 0 33504 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_347
timestamp 1677580104
transform 1 0 33888 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_367
timestamp 1679581782
transform 1 0 35808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_425
timestamp 1679581782
transform 1 0 41376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_432
timestamp 1679581782
transform 1 0 42048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_439
timestamp 1679581782
transform 1 0 42720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_446
timestamp 1679581782
transform 1 0 43392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_453
timestamp 1679581782
transform 1 0 44064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_460
timestamp 1679581782
transform 1 0 44736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_467
timestamp 1679581782
transform 1 0 45408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_474
timestamp 1679581782
transform 1 0 46080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_481
timestamp 1679581782
transform 1 0 46752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_488
timestamp 1679581782
transform 1 0 47424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_495
timestamp 1679581782
transform 1 0 48096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_502
timestamp 1679581782
transform 1 0 48768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_509
timestamp 1679581782
transform 1 0 49440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_516
timestamp 1679581782
transform 1 0 50112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_523
timestamp 1679581782
transform 1 0 50784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_530
timestamp 1679581782
transform 1 0 51456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_537
timestamp 1679581782
transform 1 0 52128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_544
timestamp 1679581782
transform 1 0 52800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_551
timestamp 1679581782
transform 1 0 53472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_558
timestamp 1679581782
transform 1 0 54144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_565
timestamp 1679581782
transform 1 0 54816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_572
timestamp 1679581782
transform 1 0 55488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_579
timestamp 1679581782
transform 1 0 56160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_586
timestamp 1679581782
transform 1 0 56832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_593
timestamp 1679581782
transform 1 0 57504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_600
timestamp 1679581782
transform 1 0 58176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_607
timestamp 1679581782
transform 1 0 58848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_614
timestamp 1679581782
transform 1 0 59520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_621
timestamp 1679581782
transform 1 0 60192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_628
timestamp 1679581782
transform 1 0 60864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_635
timestamp 1679581782
transform 1 0 61536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_642
timestamp 1679581782
transform 1 0 62208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_649
timestamp 1679581782
transform 1 0 62880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_656
timestamp 1679581782
transform 1 0 63552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_663
timestamp 1679581782
transform 1 0 64224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_670
timestamp 1679581782
transform 1 0 64896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_677
timestamp 1679581782
transform 1 0 65568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_684
timestamp 1679581782
transform 1 0 66240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_691
timestamp 1679581782
transform 1 0 66912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_698
timestamp 1679581782
transform 1 0 67584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_705
timestamp 1679581782
transform 1 0 68256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_712
timestamp 1679581782
transform 1 0 68928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_719
timestamp 1679581782
transform 1 0 69600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_726
timestamp 1679581782
transform 1 0 70272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_733
timestamp 1679581782
transform 1 0 70944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_740
timestamp 1679581782
transform 1 0 71616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_747
timestamp 1679581782
transform 1 0 72288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_754
timestamp 1679581782
transform 1 0 72960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_761
timestamp 1679581782
transform 1 0 73632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_768
timestamp 1679581782
transform 1 0 74304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_775
timestamp 1679581782
transform 1 0 74976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_782
timestamp 1679581782
transform 1 0 75648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_789
timestamp 1679581782
transform 1 0 76320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_796
timestamp 1679581782
transform 1 0 76992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_803
timestamp 1679581782
transform 1 0 77664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_810
timestamp 1679581782
transform 1 0 78336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_817
timestamp 1679581782
transform 1 0 79008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_824
timestamp 1679581782
transform 1 0 79680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_831
timestamp 1679581782
transform 1 0 80352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_838
timestamp 1679581782
transform 1 0 81024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_845
timestamp 1679581782
transform 1 0 81696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_852
timestamp 1679581782
transform 1 0 82368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_859
timestamp 1679581782
transform 1 0 83040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_866
timestamp 1679581782
transform 1 0 83712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_873
timestamp 1679581782
transform 1 0 84384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_880
timestamp 1679581782
transform 1 0 85056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_887
timestamp 1679581782
transform 1 0 85728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_894
timestamp 1679581782
transform 1 0 86400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_901
timestamp 1679581782
transform 1 0 87072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_908
timestamp 1679581782
transform 1 0 87744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_915
timestamp 1679581782
transform 1 0 88416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_922
timestamp 1679581782
transform 1 0 89088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_929
timestamp 1679581782
transform 1 0 89760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_936
timestamp 1679581782
transform 1 0 90432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_943
timestamp 1679581782
transform 1 0 91104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_950
timestamp 1679581782
transform 1 0 91776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_957
timestamp 1679581782
transform 1 0 92448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_964
timestamp 1679581782
transform 1 0 93120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_971
timestamp 1679581782
transform 1 0 93792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_978
timestamp 1679581782
transform 1 0 94464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_985
timestamp 1679581782
transform 1 0 95136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_992
timestamp 1679581782
transform 1 0 95808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_999
timestamp 1679581782
transform 1 0 96480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1006
timestamp 1679581782
transform 1 0 97152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1013
timestamp 1679581782
transform 1 0 97824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1020
timestamp 1679581782
transform 1 0 98496 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_1027
timestamp 1677580104
transform 1 0 99168 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_4
timestamp 1677580104
transform 1 0 960 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_6
timestamp 1677579658
transform 1 0 1152 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_48
timestamp 1677580104
transform 1 0 5184 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_50
timestamp 1677579658
transform 1 0 5376 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_78
timestamp 1679581782
transform 1 0 8064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_85
timestamp 1679577901
transform 1 0 8736 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_89
timestamp 1677580104
transform 1 0 9120 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_95
timestamp 1679577901
transform 1 0 9696 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_99
timestamp 1677579658
transform 1 0 10080 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_105
timestamp 1677579658
transform 1 0 10656 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_145
timestamp 1679577901
transform 1 0 14496 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_166
timestamp 1679581782
transform 1 0 16512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_173
timestamp 1679581782
transform 1 0 17184 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_180
timestamp 1677580104
transform 1 0 17856 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_182
timestamp 1677579658
transform 1 0 18048 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_187
timestamp 1679581782
transform 1 0 18528 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_194
timestamp 1677580104
transform 1 0 19200 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_196
timestamp 1677579658
transform 1 0 19392 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_206
timestamp 1677579658
transform 1 0 20352 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_231
timestamp 1677580104
transform 1 0 22752 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_233
timestamp 1677579658
transform 1 0 22944 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_266
timestamp 1677580104
transform 1 0 26112 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_274
timestamp 1677580104
transform 1 0 26880 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_328
timestamp 1677579658
transform 1 0 32064 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_342
timestamp 1677579658
transform 1 0 33408 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_386
timestamp 1677580104
transform 1 0 37632 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_427
timestamp 1679581782
transform 1 0 41568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_434
timestamp 1679581782
transform 1 0 42240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_441
timestamp 1679581782
transform 1 0 42912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_448
timestamp 1679581782
transform 1 0 43584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_455
timestamp 1679581782
transform 1 0 44256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_462
timestamp 1679581782
transform 1 0 44928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_469
timestamp 1679581782
transform 1 0 45600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_476
timestamp 1679581782
transform 1 0 46272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_483
timestamp 1679581782
transform 1 0 46944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_490
timestamp 1679581782
transform 1 0 47616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_497
timestamp 1679581782
transform 1 0 48288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_504
timestamp 1679581782
transform 1 0 48960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_511
timestamp 1679581782
transform 1 0 49632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_518
timestamp 1679581782
transform 1 0 50304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_525
timestamp 1679581782
transform 1 0 50976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_532
timestamp 1679581782
transform 1 0 51648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_539
timestamp 1679581782
transform 1 0 52320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_546
timestamp 1679581782
transform 1 0 52992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_553
timestamp 1679581782
transform 1 0 53664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_560
timestamp 1679581782
transform 1 0 54336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_567
timestamp 1679581782
transform 1 0 55008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_574
timestamp 1679581782
transform 1 0 55680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_581
timestamp 1679581782
transform 1 0 56352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_588
timestamp 1679581782
transform 1 0 57024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_595
timestamp 1679581782
transform 1 0 57696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_602
timestamp 1679581782
transform 1 0 58368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_609
timestamp 1679581782
transform 1 0 59040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_616
timestamp 1679581782
transform 1 0 59712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_623
timestamp 1679581782
transform 1 0 60384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_630
timestamp 1679581782
transform 1 0 61056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_637
timestamp 1679581782
transform 1 0 61728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_644
timestamp 1679581782
transform 1 0 62400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_651
timestamp 1679581782
transform 1 0 63072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_658
timestamp 1679581782
transform 1 0 63744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_665
timestamp 1679581782
transform 1 0 64416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_672
timestamp 1679581782
transform 1 0 65088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_679
timestamp 1679581782
transform 1 0 65760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_686
timestamp 1679581782
transform 1 0 66432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_693
timestamp 1679581782
transform 1 0 67104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_700
timestamp 1679581782
transform 1 0 67776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_707
timestamp 1679581782
transform 1 0 68448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_714
timestamp 1679581782
transform 1 0 69120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_721
timestamp 1679581782
transform 1 0 69792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_728
timestamp 1679581782
transform 1 0 70464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_735
timestamp 1679581782
transform 1 0 71136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_742
timestamp 1679581782
transform 1 0 71808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_749
timestamp 1679581782
transform 1 0 72480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_756
timestamp 1679581782
transform 1 0 73152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_763
timestamp 1679581782
transform 1 0 73824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_770
timestamp 1679581782
transform 1 0 74496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_777
timestamp 1679581782
transform 1 0 75168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_784
timestamp 1679581782
transform 1 0 75840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_791
timestamp 1679581782
transform 1 0 76512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_798
timestamp 1679581782
transform 1 0 77184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_805
timestamp 1679581782
transform 1 0 77856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_812
timestamp 1679581782
transform 1 0 78528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_819
timestamp 1679581782
transform 1 0 79200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_826
timestamp 1679581782
transform 1 0 79872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_833
timestamp 1679581782
transform 1 0 80544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_840
timestamp 1679581782
transform 1 0 81216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_847
timestamp 1679581782
transform 1 0 81888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_854
timestamp 1679581782
transform 1 0 82560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_861
timestamp 1679581782
transform 1 0 83232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_868
timestamp 1679581782
transform 1 0 83904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_875
timestamp 1679581782
transform 1 0 84576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_882
timestamp 1679581782
transform 1 0 85248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_889
timestamp 1679581782
transform 1 0 85920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_896
timestamp 1679581782
transform 1 0 86592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_903
timestamp 1679581782
transform 1 0 87264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_910
timestamp 1679581782
transform 1 0 87936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_917
timestamp 1679581782
transform 1 0 88608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_924
timestamp 1679581782
transform 1 0 89280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_931
timestamp 1679581782
transform 1 0 89952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_938
timestamp 1679581782
transform 1 0 90624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_945
timestamp 1679581782
transform 1 0 91296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_952
timestamp 1679581782
transform 1 0 91968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_959
timestamp 1679581782
transform 1 0 92640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_966
timestamp 1679581782
transform 1 0 93312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_973
timestamp 1679581782
transform 1 0 93984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_980
timestamp 1679581782
transform 1 0 94656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_987
timestamp 1679581782
transform 1 0 95328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_994
timestamp 1679581782
transform 1 0 96000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1001
timestamp 1679581782
transform 1 0 96672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1008
timestamp 1679581782
transform 1 0 97344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1015
timestamp 1679581782
transform 1 0 98016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1022
timestamp 1679581782
transform 1 0 98688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_11
timestamp 1677580104
transform 1 0 1632 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_13
timestamp 1677579658
transform 1 0 1824 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_25
timestamp 1679577901
transform 1 0 2976 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_29
timestamp 1677579658
transform 1 0 3360 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_39
timestamp 1677579658
transform 1 0 4320 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_95
timestamp 1679577901
transform 1 0 9696 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_99
timestamp 1677580104
transform 1 0 10080 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_113
timestamp 1677580104
transform 1 0 11424 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_221
timestamp 1677580104
transform 1 0 21792 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_223
timestamp 1677579658
transform 1 0 21984 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_252
timestamp 1679581782
transform 1 0 24768 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_268
timestamp 1677580104
transform 1 0 26304 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_291
timestamp 1677579658
transform 1 0 28512 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_329
timestamp 1677579658
transform 1 0 32160 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_343
timestamp 1677580104
transform 1 0 33504 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_367
timestamp 1677580104
transform 1 0 35808 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_419
timestamp 1679581782
transform 1 0 40800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_426
timestamp 1679581782
transform 1 0 41472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_433
timestamp 1679581782
transform 1 0 42144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_440
timestamp 1679581782
transform 1 0 42816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_447
timestamp 1679581782
transform 1 0 43488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_454
timestamp 1679581782
transform 1 0 44160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_461
timestamp 1679581782
transform 1 0 44832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_468
timestamp 1679581782
transform 1 0 45504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_475
timestamp 1679581782
transform 1 0 46176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_482
timestamp 1679581782
transform 1 0 46848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_489
timestamp 1679581782
transform 1 0 47520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_496
timestamp 1679581782
transform 1 0 48192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_503
timestamp 1679581782
transform 1 0 48864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_510
timestamp 1679581782
transform 1 0 49536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_517
timestamp 1679581782
transform 1 0 50208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_524
timestamp 1679581782
transform 1 0 50880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_531
timestamp 1679581782
transform 1 0 51552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_538
timestamp 1679581782
transform 1 0 52224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_545
timestamp 1679581782
transform 1 0 52896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_552
timestamp 1679581782
transform 1 0 53568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_559
timestamp 1679581782
transform 1 0 54240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_566
timestamp 1679581782
transform 1 0 54912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_573
timestamp 1679581782
transform 1 0 55584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_580
timestamp 1679581782
transform 1 0 56256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_587
timestamp 1679581782
transform 1 0 56928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_594
timestamp 1679581782
transform 1 0 57600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_601
timestamp 1679581782
transform 1 0 58272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_608
timestamp 1679581782
transform 1 0 58944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_615
timestamp 1679581782
transform 1 0 59616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_622
timestamp 1679581782
transform 1 0 60288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_629
timestamp 1679581782
transform 1 0 60960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_636
timestamp 1679581782
transform 1 0 61632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_643
timestamp 1679581782
transform 1 0 62304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_650
timestamp 1679581782
transform 1 0 62976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_657
timestamp 1679581782
transform 1 0 63648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_664
timestamp 1679581782
transform 1 0 64320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_671
timestamp 1679581782
transform 1 0 64992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_678
timestamp 1679581782
transform 1 0 65664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_685
timestamp 1679581782
transform 1 0 66336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_692
timestamp 1679581782
transform 1 0 67008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_699
timestamp 1679581782
transform 1 0 67680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_706
timestamp 1679581782
transform 1 0 68352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_713
timestamp 1679581782
transform 1 0 69024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_720
timestamp 1679581782
transform 1 0 69696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_727
timestamp 1679581782
transform 1 0 70368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_734
timestamp 1679581782
transform 1 0 71040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_741
timestamp 1679581782
transform 1 0 71712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_748
timestamp 1679581782
transform 1 0 72384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_755
timestamp 1679581782
transform 1 0 73056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_762
timestamp 1679581782
transform 1 0 73728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_769
timestamp 1679581782
transform 1 0 74400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_776
timestamp 1679581782
transform 1 0 75072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_783
timestamp 1679581782
transform 1 0 75744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_790
timestamp 1679581782
transform 1 0 76416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_797
timestamp 1679581782
transform 1 0 77088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_804
timestamp 1679581782
transform 1 0 77760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_811
timestamp 1679581782
transform 1 0 78432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_818
timestamp 1679581782
transform 1 0 79104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_825
timestamp 1679581782
transform 1 0 79776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_832
timestamp 1679581782
transform 1 0 80448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_839
timestamp 1679581782
transform 1 0 81120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_846
timestamp 1679581782
transform 1 0 81792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_853
timestamp 1679581782
transform 1 0 82464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_860
timestamp 1679581782
transform 1 0 83136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_867
timestamp 1679581782
transform 1 0 83808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_874
timestamp 1679581782
transform 1 0 84480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_881
timestamp 1679581782
transform 1 0 85152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_888
timestamp 1679581782
transform 1 0 85824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_895
timestamp 1679581782
transform 1 0 86496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_902
timestamp 1679581782
transform 1 0 87168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_909
timestamp 1679581782
transform 1 0 87840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_916
timestamp 1679581782
transform 1 0 88512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_923
timestamp 1679581782
transform 1 0 89184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_930
timestamp 1679581782
transform 1 0 89856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_937
timestamp 1679581782
transform 1 0 90528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_944
timestamp 1679581782
transform 1 0 91200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_951
timestamp 1679581782
transform 1 0 91872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_958
timestamp 1679581782
transform 1 0 92544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_965
timestamp 1679581782
transform 1 0 93216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_972
timestamp 1679581782
transform 1 0 93888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_979
timestamp 1679581782
transform 1 0 94560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_986
timestamp 1679581782
transform 1 0 95232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_993
timestamp 1679581782
transform 1 0 95904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1000
timestamp 1679581782
transform 1 0 96576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1007
timestamp 1679581782
transform 1 0 97248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1014
timestamp 1679581782
transform 1 0 97920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1021
timestamp 1679581782
transform 1 0 98592 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677579658
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_32
timestamp 1679577901
transform 1 0 3648 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_63
timestamp 1677579658
transform 1 0 6624 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_69
timestamp 1677580104
transform 1 0 7200 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_71
timestamp 1677579658
transform 1 0 7392 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_85
timestamp 1679577901
transform 1 0 8736 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_130
timestamp 1677579658
transform 1 0 13056 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_135
timestamp 1679581782
transform 1 0 13536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_142
timestamp 1679577901
transform 1 0 14208 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_146
timestamp 1677579658
transform 1 0 14592 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_178
timestamp 1679581782
transform 1 0 17664 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_185
timestamp 1677579658
transform 1 0 18336 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_215
timestamp 1677580104
transform 1 0 21216 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_227
timestamp 1677580104
transform 1 0 22368 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_242
timestamp 1677580104
transform 1 0 23808 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_248
timestamp 1677580104
transform 1 0 24384 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_250
timestamp 1677579658
transform 1 0 24576 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_318
timestamp 1677580104
transform 1 0 31104 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_320
timestamp 1677579658
transform 1 0 31296 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_329
timestamp 1677579658
transform 1 0 32160 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_347
timestamp 1679577901
transform 1 0 33888 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_379
timestamp 1679581782
transform 1 0 36960 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_386
timestamp 1677580104
transform 1 0 37632 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_392
timestamp 1679581782
transform 1 0 38208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_399
timestamp 1679577901
transform 1 0 38880 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_417
timestamp 1679581782
transform 1 0 40608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_424
timestamp 1679581782
transform 1 0 41280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_431
timestamp 1679581782
transform 1 0 41952 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_438
timestamp 1677579658
transform 1 0 42624 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_443
timestamp 1679581782
transform 1 0 43104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_450
timestamp 1679581782
transform 1 0 43776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_457
timestamp 1679581782
transform 1 0 44448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_464
timestamp 1679581782
transform 1 0 45120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_471
timestamp 1679581782
transform 1 0 45792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_478
timestamp 1679581782
transform 1 0 46464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_485
timestamp 1679581782
transform 1 0 47136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_492
timestamp 1679581782
transform 1 0 47808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_499
timestamp 1679581782
transform 1 0 48480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_506
timestamp 1679581782
transform 1 0 49152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_513
timestamp 1679581782
transform 1 0 49824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_520
timestamp 1679581782
transform 1 0 50496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_527
timestamp 1679581782
transform 1 0 51168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_534
timestamp 1679581782
transform 1 0 51840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_541
timestamp 1679581782
transform 1 0 52512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_548
timestamp 1679581782
transform 1 0 53184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_555
timestamp 1679581782
transform 1 0 53856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_562
timestamp 1679581782
transform 1 0 54528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_569
timestamp 1679581782
transform 1 0 55200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_576
timestamp 1679581782
transform 1 0 55872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_583
timestamp 1679581782
transform 1 0 56544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_590
timestamp 1679581782
transform 1 0 57216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_597
timestamp 1679581782
transform 1 0 57888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_604
timestamp 1679581782
transform 1 0 58560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_611
timestamp 1679581782
transform 1 0 59232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_618
timestamp 1679581782
transform 1 0 59904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_625
timestamp 1679581782
transform 1 0 60576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_632
timestamp 1679581782
transform 1 0 61248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_639
timestamp 1679581782
transform 1 0 61920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_646
timestamp 1679581782
transform 1 0 62592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_653
timestamp 1679581782
transform 1 0 63264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_660
timestamp 1679581782
transform 1 0 63936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_667
timestamp 1679581782
transform 1 0 64608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_674
timestamp 1679581782
transform 1 0 65280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_681
timestamp 1679581782
transform 1 0 65952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_688
timestamp 1679581782
transform 1 0 66624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_695
timestamp 1679581782
transform 1 0 67296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_702
timestamp 1679581782
transform 1 0 67968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_709
timestamp 1679581782
transform 1 0 68640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_716
timestamp 1679581782
transform 1 0 69312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_723
timestamp 1679581782
transform 1 0 69984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_730
timestamp 1679581782
transform 1 0 70656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_737
timestamp 1679581782
transform 1 0 71328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_744
timestamp 1679581782
transform 1 0 72000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_751
timestamp 1679581782
transform 1 0 72672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_758
timestamp 1679581782
transform 1 0 73344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_765
timestamp 1679581782
transform 1 0 74016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_772
timestamp 1679581782
transform 1 0 74688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_779
timestamp 1679581782
transform 1 0 75360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_786
timestamp 1679581782
transform 1 0 76032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_793
timestamp 1679581782
transform 1 0 76704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_800
timestamp 1679581782
transform 1 0 77376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_807
timestamp 1679581782
transform 1 0 78048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_814
timestamp 1679581782
transform 1 0 78720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_821
timestamp 1679581782
transform 1 0 79392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_828
timestamp 1679581782
transform 1 0 80064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_835
timestamp 1679581782
transform 1 0 80736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_842
timestamp 1679581782
transform 1 0 81408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_849
timestamp 1679581782
transform 1 0 82080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_856
timestamp 1679581782
transform 1 0 82752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_863
timestamp 1679581782
transform 1 0 83424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_870
timestamp 1679581782
transform 1 0 84096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_877
timestamp 1679581782
transform 1 0 84768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_884
timestamp 1679581782
transform 1 0 85440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_891
timestamp 1679581782
transform 1 0 86112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_898
timestamp 1679581782
transform 1 0 86784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_905
timestamp 1679581782
transform 1 0 87456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_912
timestamp 1679581782
transform 1 0 88128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_919
timestamp 1679581782
transform 1 0 88800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_926
timestamp 1679581782
transform 1 0 89472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_933
timestamp 1679581782
transform 1 0 90144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_940
timestamp 1679581782
transform 1 0 90816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_947
timestamp 1679581782
transform 1 0 91488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_954
timestamp 1679581782
transform 1 0 92160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_961
timestamp 1679581782
transform 1 0 92832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_968
timestamp 1679581782
transform 1 0 93504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_975
timestamp 1679581782
transform 1 0 94176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_982
timestamp 1679581782
transform 1 0 94848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_989
timestamp 1679581782
transform 1 0 95520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_996
timestamp 1679581782
transform 1 0 96192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1003
timestamp 1679581782
transform 1 0 96864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1010
timestamp 1679581782
transform 1 0 97536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1017
timestamp 1679581782
transform 1 0 98208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_1024
timestamp 1679577901
transform 1 0 98880 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_1028
timestamp 1677579658
transform 1 0 99264 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_38
timestamp 1677579658
transform 1 0 4224 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_57
timestamp 1677579658
transform 1 0 6048 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_67
timestamp 1677580104
transform 1 0 7008 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_82
timestamp 1677580104
transform 1 0 8448 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_92
timestamp 1677579658
transform 1 0 9408 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_98
timestamp 1677580104
transform 1 0 9984 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_100
timestamp 1677579658
transform 1 0 10176 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_125
timestamp 1679577901
transform 1 0 12576 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_129
timestamp 1677579658
transform 1 0 12960 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_143
timestamp 1679581782
transform 1 0 14304 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_150
timestamp 1677579658
transform 1 0 14976 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_165
timestamp 1677580104
transform 1 0 16416 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_185
timestamp 1679577901
transform 1 0 18336 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_189
timestamp 1677579658
transform 1 0 18720 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_231
timestamp 1679581782
transform 1 0 22752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_238
timestamp 1679581782
transform 1 0 23424 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_245
timestamp 1677579658
transform 1 0 24096 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_259
timestamp 1677579658
transform 1 0 25440 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_286
timestamp 1679581782
transform 1 0 28032 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_293
timestamp 1677580104
transform 1 0 28704 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_295
timestamp 1677579658
transform 1 0 28896 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_300
timestamp 1679581782
transform 1 0 29376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_307
timestamp 1679581782
transform 1 0 30048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_314
timestamp 1679581782
transform 1 0 30720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_321
timestamp 1679581782
transform 1 0 31392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_328
timestamp 1679581782
transform 1 0 32064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_335
timestamp 1679577901
transform 1 0 32736 0 1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_26_352
timestamp 1679577901
transform 1 0 34368 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_360
timestamp 1677579658
transform 1 0 35136 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_366
timestamp 1679581782
transform 1 0 35712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_373
timestamp 1679581782
transform 1 0 36384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_383
timestamp 1679577901
transform 1 0 37344 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_390
timestamp 1679581782
transform 1 0 38016 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_397
timestamp 1677580104
transform 1 0 38688 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_429
timestamp 1679577901
transform 1 0 41760 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_461
timestamp 1679581782
transform 1 0 44832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_468
timestamp 1679581782
transform 1 0 45504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_475
timestamp 1679581782
transform 1 0 46176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_482
timestamp 1679581782
transform 1 0 46848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_489
timestamp 1679581782
transform 1 0 47520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_496
timestamp 1679581782
transform 1 0 48192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_503
timestamp 1679581782
transform 1 0 48864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_510
timestamp 1679581782
transform 1 0 49536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_517
timestamp 1679581782
transform 1 0 50208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_524
timestamp 1679581782
transform 1 0 50880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_531
timestamp 1679581782
transform 1 0 51552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_538
timestamp 1679581782
transform 1 0 52224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_545
timestamp 1679581782
transform 1 0 52896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_552
timestamp 1679581782
transform 1 0 53568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_559
timestamp 1679581782
transform 1 0 54240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_566
timestamp 1679581782
transform 1 0 54912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_573
timestamp 1679581782
transform 1 0 55584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_580
timestamp 1679581782
transform 1 0 56256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_587
timestamp 1679581782
transform 1 0 56928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_594
timestamp 1679581782
transform 1 0 57600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_601
timestamp 1679581782
transform 1 0 58272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_608
timestamp 1679581782
transform 1 0 58944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_615
timestamp 1679581782
transform 1 0 59616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_622
timestamp 1679581782
transform 1 0 60288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_629
timestamp 1679581782
transform 1 0 60960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_636
timestamp 1679581782
transform 1 0 61632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_643
timestamp 1679581782
transform 1 0 62304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_650
timestamp 1679581782
transform 1 0 62976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_657
timestamp 1679581782
transform 1 0 63648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_664
timestamp 1679581782
transform 1 0 64320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_671
timestamp 1679581782
transform 1 0 64992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_678
timestamp 1679581782
transform 1 0 65664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_685
timestamp 1679581782
transform 1 0 66336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_692
timestamp 1679581782
transform 1 0 67008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_699
timestamp 1679581782
transform 1 0 67680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_706
timestamp 1679581782
transform 1 0 68352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_713
timestamp 1679581782
transform 1 0 69024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_720
timestamp 1679581782
transform 1 0 69696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_727
timestamp 1679581782
transform 1 0 70368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_734
timestamp 1679581782
transform 1 0 71040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_741
timestamp 1679581782
transform 1 0 71712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_748
timestamp 1679581782
transform 1 0 72384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_755
timestamp 1679581782
transform 1 0 73056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_762
timestamp 1679581782
transform 1 0 73728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_769
timestamp 1679581782
transform 1 0 74400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_776
timestamp 1679581782
transform 1 0 75072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_783
timestamp 1679581782
transform 1 0 75744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_790
timestamp 1679581782
transform 1 0 76416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_797
timestamp 1679581782
transform 1 0 77088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_804
timestamp 1679581782
transform 1 0 77760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_811
timestamp 1679581782
transform 1 0 78432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_818
timestamp 1679581782
transform 1 0 79104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_825
timestamp 1679581782
transform 1 0 79776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_832
timestamp 1679581782
transform 1 0 80448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_839
timestamp 1679581782
transform 1 0 81120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_846
timestamp 1679581782
transform 1 0 81792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_853
timestamp 1679581782
transform 1 0 82464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_860
timestamp 1679581782
transform 1 0 83136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_867
timestamp 1679581782
transform 1 0 83808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_874
timestamp 1679581782
transform 1 0 84480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_881
timestamp 1679581782
transform 1 0 85152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_888
timestamp 1679581782
transform 1 0 85824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_895
timestamp 1679581782
transform 1 0 86496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_902
timestamp 1679581782
transform 1 0 87168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_909
timestamp 1679581782
transform 1 0 87840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_916
timestamp 1679581782
transform 1 0 88512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_923
timestamp 1679581782
transform 1 0 89184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_930
timestamp 1679581782
transform 1 0 89856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_937
timestamp 1679581782
transform 1 0 90528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_944
timestamp 1679581782
transform 1 0 91200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_951
timestamp 1679581782
transform 1 0 91872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_958
timestamp 1679581782
transform 1 0 92544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_965
timestamp 1679581782
transform 1 0 93216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_972
timestamp 1679581782
transform 1 0 93888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_979
timestamp 1679581782
transform 1 0 94560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_986
timestamp 1679581782
transform 1 0 95232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_993
timestamp 1679581782
transform 1 0 95904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1000
timestamp 1679581782
transform 1 0 96576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1007
timestamp 1679581782
transform 1 0 97248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1014
timestamp 1679581782
transform 1 0 97920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1021
timestamp 1679581782
transform 1 0 98592 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677579658
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_7
timestamp 1679577901
transform 1 0 1248 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_15
timestamp 1677579658
transform 1 0 2016 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_20
timestamp 1677579658
transform 1 0 2496 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_39
timestamp 1677579658
transform 1 0 4320 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_120
timestamp 1679581782
transform 1 0 12096 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_127
timestamp 1677580104
transform 1 0 12768 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_159
timestamp 1677579658
transform 1 0 15840 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_200
timestamp 1679581782
transform 1 0 19776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_207
timestamp 1679581782
transform 1 0 20448 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_242
timestamp 1677580104
transform 1 0 23808 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_277
timestamp 1677579658
transform 1 0 27168 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_314
timestamp 1679581782
transform 1 0 30720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_321
timestamp 1679581782
transform 1 0 31392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_328
timestamp 1679581782
transform 1 0 32064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_335
timestamp 1679581782
transform 1 0 32736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_342
timestamp 1679581782
transform 1 0 33408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_349
timestamp 1679581782
transform 1 0 34080 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_356
timestamp 1677579658
transform 1 0 34752 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_361
timestamp 1679577901
transform 1 0 35232 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_405
timestamp 1677579658
transform 1 0 39456 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_441
timestamp 1677580104
transform 1 0 42912 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 45600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 46272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679581782
transform 1 0 75168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679581782
transform 1 0 75840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679581782
transform 1 0 76512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679581782
transform 1 0 77184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679581782
transform 1 0 77856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679581782
transform 1 0 78528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679581782
transform 1 0 79200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679581782
transform 1 0 79872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679581782
transform 1 0 80544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_840
timestamp 1679581782
transform 1 0 81216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_847
timestamp 1679581782
transform 1 0 81888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_854
timestamp 1679581782
transform 1 0 82560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_861
timestamp 1679581782
transform 1 0 83232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_868
timestamp 1679581782
transform 1 0 83904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_875
timestamp 1679581782
transform 1 0 84576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679581782
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679581782
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679581782
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679581782
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679581782
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679581782
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_924
timestamp 1679581782
transform 1 0 89280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_931
timestamp 1679581782
transform 1 0 89952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_938
timestamp 1679581782
transform 1 0 90624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679581782
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679581782
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_959
timestamp 1679581782
transform 1 0 92640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_966
timestamp 1679581782
transform 1 0 93312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_973
timestamp 1679581782
transform 1 0 93984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_980
timestamp 1679581782
transform 1 0 94656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_987
timestamp 1679581782
transform 1 0 95328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_994
timestamp 1679581782
transform 1 0 96000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1001
timestamp 1679581782
transform 1 0 96672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1008
timestamp 1679581782
transform 1 0 97344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1015
timestamp 1679581782
transform 1 0 98016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1022
timestamp 1679581782
transform 1 0 98688 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_4
timestamp 1677580104
transform 1 0 960 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_82
timestamp 1677580104
transform 1 0 8448 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_102
timestamp 1677579658
transform 1 0 10368 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_113
timestamp 1679577901
transform 1 0 11424 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_117
timestamp 1677580104
transform 1 0 11808 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_132
timestamp 1677580104
transform 1 0 13248 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_143
timestamp 1677579658
transform 1 0 14304 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_170
timestamp 1677580104
transform 1 0 16896 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_28_196
timestamp 1679577901
transform 1 0 19392 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_200
timestamp 1677579658
transform 1 0 19776 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_204
timestamp 1679581782
transform 1 0 20160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_211
timestamp 1679581782
transform 1 0 20832 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_218
timestamp 1677579658
transform 1 0 21504 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_223
timestamp 1679581782
transform 1 0 21984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_230
timestamp 1679577901
transform 1 0 22656 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_267
timestamp 1677580104
transform 1 0 26208 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_269
timestamp 1677579658
transform 1 0 26400 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_288
timestamp 1677580104
transform 1 0 28224 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_290
timestamp 1677579658
transform 1 0 28416 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_349
timestamp 1677580104
transform 1 0 34080 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_351
timestamp 1677579658
transform 1 0 34272 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_379
timestamp 1677579658
transform 1 0 36960 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_393
timestamp 1677579658
transform 1 0 38304 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_462
timestamp 1677579658
transform 1 0 44928 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_476
timestamp 1679577901
transform 1 0 46272 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_508
timestamp 1679581782
transform 1 0 49344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_515
timestamp 1679581782
transform 1 0 50016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_522
timestamp 1679581782
transform 1 0 50688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_529
timestamp 1679581782
transform 1 0 51360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_536
timestamp 1679581782
transform 1 0 52032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_543
timestamp 1679581782
transform 1 0 52704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_550
timestamp 1679581782
transform 1 0 53376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_557
timestamp 1679581782
transform 1 0 54048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_564
timestamp 1679581782
transform 1 0 54720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_571
timestamp 1679581782
transform 1 0 55392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_578
timestamp 1679581782
transform 1 0 56064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_585
timestamp 1679581782
transform 1 0 56736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_592
timestamp 1679581782
transform 1 0 57408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_599
timestamp 1679581782
transform 1 0 58080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_606
timestamp 1679581782
transform 1 0 58752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_613
timestamp 1679581782
transform 1 0 59424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_620
timestamp 1679581782
transform 1 0 60096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_627
timestamp 1679581782
transform 1 0 60768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_634
timestamp 1679581782
transform 1 0 61440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_641
timestamp 1679581782
transform 1 0 62112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_648
timestamp 1679581782
transform 1 0 62784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_655
timestamp 1679581782
transform 1 0 63456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_662
timestamp 1679581782
transform 1 0 64128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_669
timestamp 1679581782
transform 1 0 64800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_676
timestamp 1679581782
transform 1 0 65472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_683
timestamp 1679581782
transform 1 0 66144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_690
timestamp 1679581782
transform 1 0 66816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_697
timestamp 1679581782
transform 1 0 67488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_704
timestamp 1679581782
transform 1 0 68160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_711
timestamp 1679581782
transform 1 0 68832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_718
timestamp 1679581782
transform 1 0 69504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_725
timestamp 1679581782
transform 1 0 70176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_732
timestamp 1679581782
transform 1 0 70848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_739
timestamp 1679581782
transform 1 0 71520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_746
timestamp 1679581782
transform 1 0 72192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_753
timestamp 1679581782
transform 1 0 72864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_760
timestamp 1679581782
transform 1 0 73536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_767
timestamp 1679581782
transform 1 0 74208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_774
timestamp 1679581782
transform 1 0 74880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_781
timestamp 1679581782
transform 1 0 75552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_788
timestamp 1679581782
transform 1 0 76224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_795
timestamp 1679581782
transform 1 0 76896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_802
timestamp 1679581782
transform 1 0 77568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_809
timestamp 1679581782
transform 1 0 78240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_816
timestamp 1679581782
transform 1 0 78912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_823
timestamp 1679581782
transform 1 0 79584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_830
timestamp 1679581782
transform 1 0 80256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_837
timestamp 1679581782
transform 1 0 80928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_844
timestamp 1679581782
transform 1 0 81600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_851
timestamp 1679581782
transform 1 0 82272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_858
timestamp 1679581782
transform 1 0 82944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_865
timestamp 1679581782
transform 1 0 83616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_872
timestamp 1679581782
transform 1 0 84288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_879
timestamp 1679581782
transform 1 0 84960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_886
timestamp 1679581782
transform 1 0 85632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_893
timestamp 1679581782
transform 1 0 86304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_900
timestamp 1679581782
transform 1 0 86976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_907
timestamp 1679581782
transform 1 0 87648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_914
timestamp 1679581782
transform 1 0 88320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_921
timestamp 1679581782
transform 1 0 88992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_928
timestamp 1679581782
transform 1 0 89664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_935
timestamp 1679581782
transform 1 0 90336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_942
timestamp 1679581782
transform 1 0 91008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_949
timestamp 1679581782
transform 1 0 91680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_956
timestamp 1679581782
transform 1 0 92352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_963
timestamp 1679581782
transform 1 0 93024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_970
timestamp 1679581782
transform 1 0 93696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_977
timestamp 1679581782
transform 1 0 94368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_984
timestamp 1679581782
transform 1 0 95040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_991
timestamp 1679581782
transform 1 0 95712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_998
timestamp 1679581782
transform 1 0 96384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1005
timestamp 1679581782
transform 1 0 97056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1012
timestamp 1679581782
transform 1 0 97728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1019
timestamp 1679581782
transform 1 0 98400 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_1026
timestamp 1677580104
transform 1 0 99072 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_1028
timestamp 1677579658
transform 1 0 99264 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_4
timestamp 1677580104
transform 1 0 960 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_33
timestamp 1677579658
transform 1 0 3744 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_49
timestamp 1677579658
transform 1 0 5280 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_59
timestamp 1679577901
transform 1 0 6240 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_29_85
timestamp 1679577901
transform 1 0 8736 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_29_103
timestamp 1679577901
transform 1 0 10464 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_107
timestamp 1677580104
transform 1 0 10848 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_162
timestamp 1677579658
transform 1 0 16128 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_172
timestamp 1677580104
transform 1 0 17088 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_210
timestamp 1679581782
transform 1 0 20736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_217
timestamp 1679581782
transform 1 0 21408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_224
timestamp 1679581782
transform 1 0 22080 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_231
timestamp 1677580104
transform 1 0 22752 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_233
timestamp 1677579658
transform 1 0 22944 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_239
timestamp 1677579658
transform 1 0 23520 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_253
timestamp 1677579658
transform 1 0 24864 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_299
timestamp 1677579658
transform 1 0 29280 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_304
timestamp 1677579658
transform 1 0 29760 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_331
timestamp 1679577901
transform 1 0 32352 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_335
timestamp 1677579658
transform 1 0 32736 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_378
timestamp 1677580104
transform 1 0 36864 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_402
timestamp 1677579658
transform 1 0 39168 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_451
timestamp 1677580104
transform 1 0 43872 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_493
timestamp 1679581782
transform 1 0 47904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_528
timestamp 1679581782
transform 1 0 51264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_535
timestamp 1679581782
transform 1 0 51936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_542
timestamp 1679581782
transform 1 0 52608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_549
timestamp 1679581782
transform 1 0 53280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_556
timestamp 1679581782
transform 1 0 53952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_563
timestamp 1679581782
transform 1 0 54624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_570
timestamp 1679581782
transform 1 0 55296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_577
timestamp 1679581782
transform 1 0 55968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_584
timestamp 1679581782
transform 1 0 56640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_591
timestamp 1679581782
transform 1 0 57312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_598
timestamp 1679581782
transform 1 0 57984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_605
timestamp 1679581782
transform 1 0 58656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_612
timestamp 1679581782
transform 1 0 59328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_619
timestamp 1679581782
transform 1 0 60000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_626
timestamp 1679581782
transform 1 0 60672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_633
timestamp 1679581782
transform 1 0 61344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_640
timestamp 1679581782
transform 1 0 62016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_647
timestamp 1679581782
transform 1 0 62688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_654
timestamp 1679581782
transform 1 0 63360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_661
timestamp 1679581782
transform 1 0 64032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_668
timestamp 1679581782
transform 1 0 64704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_675
timestamp 1679581782
transform 1 0 65376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_682
timestamp 1679581782
transform 1 0 66048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_689
timestamp 1679581782
transform 1 0 66720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_696
timestamp 1679581782
transform 1 0 67392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_703
timestamp 1679581782
transform 1 0 68064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_710
timestamp 1679581782
transform 1 0 68736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_717
timestamp 1679581782
transform 1 0 69408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_724
timestamp 1679581782
transform 1 0 70080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_731
timestamp 1679581782
transform 1 0 70752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_738
timestamp 1679581782
transform 1 0 71424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_745
timestamp 1679581782
transform 1 0 72096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_752
timestamp 1679581782
transform 1 0 72768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_759
timestamp 1679581782
transform 1 0 73440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_766
timestamp 1679581782
transform 1 0 74112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_773
timestamp 1679581782
transform 1 0 74784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_780
timestamp 1679581782
transform 1 0 75456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_787
timestamp 1679581782
transform 1 0 76128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_794
timestamp 1679581782
transform 1 0 76800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_801
timestamp 1679581782
transform 1 0 77472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_808
timestamp 1679581782
transform 1 0 78144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_815
timestamp 1679581782
transform 1 0 78816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_822
timestamp 1679581782
transform 1 0 79488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_829
timestamp 1679581782
transform 1 0 80160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_836
timestamp 1679581782
transform 1 0 80832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_843
timestamp 1679581782
transform 1 0 81504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_850
timestamp 1679581782
transform 1 0 82176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_857
timestamp 1679581782
transform 1 0 82848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_864
timestamp 1679581782
transform 1 0 83520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_871
timestamp 1679581782
transform 1 0 84192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_878
timestamp 1679581782
transform 1 0 84864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_885
timestamp 1679581782
transform 1 0 85536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_892
timestamp 1679581782
transform 1 0 86208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_899
timestamp 1679581782
transform 1 0 86880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_906
timestamp 1679581782
transform 1 0 87552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_913
timestamp 1679581782
transform 1 0 88224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_920
timestamp 1679581782
transform 1 0 88896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_927
timestamp 1679581782
transform 1 0 89568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_934
timestamp 1679581782
transform 1 0 90240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_941
timestamp 1679581782
transform 1 0 90912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_948
timestamp 1679581782
transform 1 0 91584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_955
timestamp 1679581782
transform 1 0 92256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_962
timestamp 1679581782
transform 1 0 92928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_969
timestamp 1679581782
transform 1 0 93600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_976
timestamp 1679581782
transform 1 0 94272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_983
timestamp 1679581782
transform 1 0 94944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_990
timestamp 1679581782
transform 1 0 95616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_997
timestamp 1679581782
transform 1 0 96288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1004
timestamp 1679581782
transform 1 0 96960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1011
timestamp 1679581782
transform 1 0 97632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1018
timestamp 1679581782
transform 1 0 98304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_1025
timestamp 1679577901
transform 1 0 98976 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679581782
transform 1 0 576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_7
timestamp 1679577901
transform 1 0 1248 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_15
timestamp 1677580104
transform 1 0 2016 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_97
timestamp 1677579658
transform 1 0 9888 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_155
timestamp 1677579658
transform 1 0 15456 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_184
timestamp 1679581782
transform 1 0 18240 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_191
timestamp 1677579658
transform 1 0 18912 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_244
timestamp 1679577901
transform 1 0 24000 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_248
timestamp 1677580104
transform 1 0 24384 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_273
timestamp 1677580104
transform 1 0 26784 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_275
timestamp 1677579658
transform 1 0 26976 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_305
timestamp 1679581782
transform 1 0 29856 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_312
timestamp 1677580104
transform 1 0 30528 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_322
timestamp 1679577901
transform 1 0 31488 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_326
timestamp 1677580104
transform 1 0 31872 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_420
timestamp 1677579658
transform 1 0 40896 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_486
timestamp 1677580104
transform 1 0 47232 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_488
timestamp 1677579658
transform 1 0 47424 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_511
timestamp 1677580104
transform 1 0 49632 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_517
timestamp 1679581782
transform 1 0 50208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_524
timestamp 1679581782
transform 1 0 50880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_531
timestamp 1679581782
transform 1 0 51552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_538
timestamp 1679581782
transform 1 0 52224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_545
timestamp 1679581782
transform 1 0 52896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_552
timestamp 1679581782
transform 1 0 53568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_559
timestamp 1679581782
transform 1 0 54240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_566
timestamp 1679581782
transform 1 0 54912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_573
timestamp 1679581782
transform 1 0 55584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_580
timestamp 1679581782
transform 1 0 56256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_587
timestamp 1679581782
transform 1 0 56928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_594
timestamp 1679581782
transform 1 0 57600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_601
timestamp 1679581782
transform 1 0 58272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_608
timestamp 1679581782
transform 1 0 58944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_615
timestamp 1679581782
transform 1 0 59616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_622
timestamp 1679581782
transform 1 0 60288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_629
timestamp 1679581782
transform 1 0 60960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_636
timestamp 1679581782
transform 1 0 61632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_643
timestamp 1679581782
transform 1 0 62304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_650
timestamp 1679581782
transform 1 0 62976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_657
timestamp 1679581782
transform 1 0 63648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_664
timestamp 1679581782
transform 1 0 64320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_671
timestamp 1679581782
transform 1 0 64992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_678
timestamp 1679581782
transform 1 0 65664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_685
timestamp 1679581782
transform 1 0 66336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_692
timestamp 1679581782
transform 1 0 67008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_699
timestamp 1679581782
transform 1 0 67680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_706
timestamp 1679581782
transform 1 0 68352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_713
timestamp 1679581782
transform 1 0 69024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_720
timestamp 1679581782
transform 1 0 69696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_727
timestamp 1679581782
transform 1 0 70368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_734
timestamp 1679581782
transform 1 0 71040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_741
timestamp 1679581782
transform 1 0 71712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_748
timestamp 1679581782
transform 1 0 72384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_755
timestamp 1679581782
transform 1 0 73056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_762
timestamp 1679581782
transform 1 0 73728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_769
timestamp 1679581782
transform 1 0 74400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_776
timestamp 1679581782
transform 1 0 75072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_783
timestamp 1679581782
transform 1 0 75744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_790
timestamp 1679581782
transform 1 0 76416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_797
timestamp 1679581782
transform 1 0 77088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_804
timestamp 1679581782
transform 1 0 77760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_811
timestamp 1679581782
transform 1 0 78432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_818
timestamp 1679581782
transform 1 0 79104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_825
timestamp 1679581782
transform 1 0 79776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_832
timestamp 1679581782
transform 1 0 80448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_839
timestamp 1679581782
transform 1 0 81120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_846
timestamp 1679581782
transform 1 0 81792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_853
timestamp 1679581782
transform 1 0 82464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_860
timestamp 1679581782
transform 1 0 83136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_867
timestamp 1679581782
transform 1 0 83808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_874
timestamp 1679581782
transform 1 0 84480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_881
timestamp 1679581782
transform 1 0 85152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_888
timestamp 1679581782
transform 1 0 85824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_895
timestamp 1679581782
transform 1 0 86496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_902
timestamp 1679581782
transform 1 0 87168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_909
timestamp 1679581782
transform 1 0 87840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_916
timestamp 1679581782
transform 1 0 88512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_923
timestamp 1679581782
transform 1 0 89184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_930
timestamp 1679581782
transform 1 0 89856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_937
timestamp 1679581782
transform 1 0 90528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_944
timestamp 1679581782
transform 1 0 91200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_951
timestamp 1679581782
transform 1 0 91872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_958
timestamp 1679581782
transform 1 0 92544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_965
timestamp 1679581782
transform 1 0 93216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_972
timestamp 1679581782
transform 1 0 93888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_979
timestamp 1679581782
transform 1 0 94560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_986
timestamp 1679581782
transform 1 0 95232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_993
timestamp 1679581782
transform 1 0 95904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1000
timestamp 1679581782
transform 1 0 96576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1007
timestamp 1679581782
transform 1 0 97248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1014
timestamp 1679581782
transform 1 0 97920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1021
timestamp 1679581782
transform 1 0 98592 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_1028
timestamp 1677579658
transform 1 0 99264 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_0
timestamp 1679577901
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_4
timestamp 1677579658
transform 1 0 960 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_32
timestamp 1679577901
transform 1 0 3648 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_31_92
timestamp 1679577901
transform 1 0 9408 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_118
timestamp 1677580104
transform 1 0 11904 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_145
timestamp 1677580104
transform 1 0 14496 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_182
timestamp 1679577901
transform 1 0 18048 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_186
timestamp 1677579658
transform 1 0 18432 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_240
timestamp 1679581782
transform 1 0 23616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_247
timestamp 1679581782
transform 1 0 24288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_254
timestamp 1679581782
transform 1 0 24960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_265
timestamp 1679581782
transform 1 0 26016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_272
timestamp 1679581782
transform 1 0 26688 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_279
timestamp 1677580104
transform 1 0 27360 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_293
timestamp 1679577901
transform 1 0 28704 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_297
timestamp 1677580104
transform 1 0 29088 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_326
timestamp 1679581782
transform 1 0 31872 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_333
timestamp 1677580104
transform 1 0 32544 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_362
timestamp 1677580104
transform 1 0 35328 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_372
timestamp 1677580104
transform 1 0 36288 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_374
timestamp 1677579658
transform 1 0 36480 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_396
timestamp 1677580104
transform 1 0 38592 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_402
timestamp 1679577901
transform 1 0 39168 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_406
timestamp 1677580104
transform 1 0 39552 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_429
timestamp 1677580104
transform 1 0 41760 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_431
timestamp 1677579658
transform 1 0 41952 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_449
timestamp 1677579658
transform 1 0 43680 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_492
timestamp 1677579658
transform 1 0 47808 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_506
timestamp 1677580104
transform 1 0 49152 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_536
timestamp 1679581782
transform 1 0 52032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_543
timestamp 1679581782
transform 1 0 52704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_550
timestamp 1679581782
transform 1 0 53376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_557
timestamp 1679581782
transform 1 0 54048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_564
timestamp 1679581782
transform 1 0 54720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_571
timestamp 1679581782
transform 1 0 55392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_578
timestamp 1679581782
transform 1 0 56064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_585
timestamp 1679581782
transform 1 0 56736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_592
timestamp 1679581782
transform 1 0 57408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_599
timestamp 1679581782
transform 1 0 58080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_606
timestamp 1679581782
transform 1 0 58752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_613
timestamp 1679581782
transform 1 0 59424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_620
timestamp 1679581782
transform 1 0 60096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_627
timestamp 1679581782
transform 1 0 60768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_634
timestamp 1679581782
transform 1 0 61440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_641
timestamp 1679581782
transform 1 0 62112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_648
timestamp 1679581782
transform 1 0 62784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_655
timestamp 1679581782
transform 1 0 63456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_662
timestamp 1679581782
transform 1 0 64128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_669
timestamp 1679581782
transform 1 0 64800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_676
timestamp 1679581782
transform 1 0 65472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_683
timestamp 1679581782
transform 1 0 66144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_690
timestamp 1679581782
transform 1 0 66816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_697
timestamp 1679581782
transform 1 0 67488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_704
timestamp 1679581782
transform 1 0 68160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_711
timestamp 1679581782
transform 1 0 68832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_718
timestamp 1679581782
transform 1 0 69504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_725
timestamp 1679581782
transform 1 0 70176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_732
timestamp 1679581782
transform 1 0 70848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_739
timestamp 1679581782
transform 1 0 71520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_746
timestamp 1679581782
transform 1 0 72192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_753
timestamp 1679581782
transform 1 0 72864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_760
timestamp 1679581782
transform 1 0 73536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_767
timestamp 1679581782
transform 1 0 74208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_774
timestamp 1679581782
transform 1 0 74880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_781
timestamp 1679581782
transform 1 0 75552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_788
timestamp 1679581782
transform 1 0 76224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_795
timestamp 1679581782
transform 1 0 76896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_802
timestamp 1679581782
transform 1 0 77568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_809
timestamp 1679581782
transform 1 0 78240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_816
timestamp 1679581782
transform 1 0 78912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_823
timestamp 1679581782
transform 1 0 79584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_830
timestamp 1679581782
transform 1 0 80256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_837
timestamp 1679581782
transform 1 0 80928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_844
timestamp 1679581782
transform 1 0 81600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_851
timestamp 1679581782
transform 1 0 82272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_858
timestamp 1679581782
transform 1 0 82944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_865
timestamp 1679581782
transform 1 0 83616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_872
timestamp 1679581782
transform 1 0 84288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_879
timestamp 1679581782
transform 1 0 84960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_886
timestamp 1679581782
transform 1 0 85632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_893
timestamp 1679581782
transform 1 0 86304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_900
timestamp 1679581782
transform 1 0 86976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_907
timestamp 1679581782
transform 1 0 87648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_914
timestamp 1679581782
transform 1 0 88320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_921
timestamp 1679581782
transform 1 0 88992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_928
timestamp 1679581782
transform 1 0 89664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_935
timestamp 1679581782
transform 1 0 90336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_942
timestamp 1679581782
transform 1 0 91008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_949
timestamp 1679581782
transform 1 0 91680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_956
timestamp 1679581782
transform 1 0 92352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_963
timestamp 1679581782
transform 1 0 93024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_970
timestamp 1679581782
transform 1 0 93696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_977
timestamp 1679581782
transform 1 0 94368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_984
timestamp 1679581782
transform 1 0 95040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_991
timestamp 1679581782
transform 1 0 95712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_998
timestamp 1679581782
transform 1 0 96384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1005
timestamp 1679581782
transform 1 0 97056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1012
timestamp 1679581782
transform 1 0 97728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1019
timestamp 1679581782
transform 1 0 98400 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_1026
timestamp 1677580104
transform 1 0 99072 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_1028
timestamp 1677579658
transform 1 0 99264 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679581782
transform 1 0 576 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_7
timestamp 1677580104
transform 1 0 1248 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_9
timestamp 1677579658
transform 1 0 1440 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1679581782
transform 1 0 1920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_21
timestamp 1679581782
transform 1 0 2592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_69
timestamp 1679577901
transform 1 0 7200 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_73
timestamp 1677580104
transform 1 0 7584 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_124
timestamp 1677580104
transform 1 0 12480 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_144
timestamp 1677579658
transform 1 0 14400 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_182
timestamp 1679581782
transform 1 0 18048 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_189
timestamp 1677580104
transform 1 0 18720 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_191
timestamp 1677579658
transform 1 0 18912 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_222
timestamp 1679581782
transform 1 0 21888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_296
timestamp 1679581782
transform 1 0 28992 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_303
timestamp 1677579658
transform 1 0 29664 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_308
timestamp 1679581782
transform 1 0 30144 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_315
timestamp 1677580104
transform 1 0 30816 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_353
timestamp 1677580104
transform 1 0 34464 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_396
timestamp 1677580104
transform 1 0 38592 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_398
timestamp 1677579658
transform 1 0 38784 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_420
timestamp 1677580104
transform 1 0 40896 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_422
timestamp 1677579658
transform 1 0 41088 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_433
timestamp 1677579658
transform 1 0 42144 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_447
timestamp 1677580104
transform 1 0 43488 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_454
timestamp 1677579658
transform 1 0 44160 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_528
timestamp 1679581782
transform 1 0 51264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_535
timestamp 1679581782
transform 1 0 51936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_542
timestamp 1679581782
transform 1 0 52608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_549
timestamp 1679581782
transform 1 0 53280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_556
timestamp 1679581782
transform 1 0 53952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_563
timestamp 1679581782
transform 1 0 54624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_570
timestamp 1679581782
transform 1 0 55296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_577
timestamp 1679581782
transform 1 0 55968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_584
timestamp 1679581782
transform 1 0 56640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_591
timestamp 1679581782
transform 1 0 57312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_598
timestamp 1679581782
transform 1 0 57984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_605
timestamp 1679581782
transform 1 0 58656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_612
timestamp 1679581782
transform 1 0 59328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_619
timestamp 1679581782
transform 1 0 60000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_626
timestamp 1679581782
transform 1 0 60672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_633
timestamp 1679581782
transform 1 0 61344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_640
timestamp 1679581782
transform 1 0 62016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_647
timestamp 1679581782
transform 1 0 62688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_654
timestamp 1679581782
transform 1 0 63360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_661
timestamp 1679581782
transform 1 0 64032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_668
timestamp 1679581782
transform 1 0 64704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_675
timestamp 1679581782
transform 1 0 65376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_682
timestamp 1679581782
transform 1 0 66048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_689
timestamp 1679581782
transform 1 0 66720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_696
timestamp 1679581782
transform 1 0 67392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_703
timestamp 1679581782
transform 1 0 68064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_710
timestamp 1679581782
transform 1 0 68736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_717
timestamp 1679581782
transform 1 0 69408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_724
timestamp 1679581782
transform 1 0 70080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_731
timestamp 1679581782
transform 1 0 70752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_738
timestamp 1679581782
transform 1 0 71424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_745
timestamp 1679581782
transform 1 0 72096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_752
timestamp 1679581782
transform 1 0 72768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_759
timestamp 1679581782
transform 1 0 73440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_766
timestamp 1679581782
transform 1 0 74112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_773
timestamp 1679581782
transform 1 0 74784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_780
timestamp 1679581782
transform 1 0 75456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_787
timestamp 1679581782
transform 1 0 76128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_794
timestamp 1679581782
transform 1 0 76800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_801
timestamp 1679581782
transform 1 0 77472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_808
timestamp 1679581782
transform 1 0 78144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_815
timestamp 1679581782
transform 1 0 78816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_822
timestamp 1679581782
transform 1 0 79488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_829
timestamp 1679581782
transform 1 0 80160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_836
timestamp 1679581782
transform 1 0 80832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_843
timestamp 1679581782
transform 1 0 81504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_850
timestamp 1679581782
transform 1 0 82176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_857
timestamp 1679581782
transform 1 0 82848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_864
timestamp 1679581782
transform 1 0 83520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_871
timestamp 1679581782
transform 1 0 84192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_878
timestamp 1679581782
transform 1 0 84864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_885
timestamp 1679581782
transform 1 0 85536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_892
timestamp 1679581782
transform 1 0 86208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_899
timestamp 1679581782
transform 1 0 86880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_906
timestamp 1679581782
transform 1 0 87552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_913
timestamp 1679581782
transform 1 0 88224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_920
timestamp 1679581782
transform 1 0 88896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_927
timestamp 1679581782
transform 1 0 89568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_934
timestamp 1679581782
transform 1 0 90240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_941
timestamp 1679581782
transform 1 0 90912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_948
timestamp 1679581782
transform 1 0 91584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_955
timestamp 1679581782
transform 1 0 92256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_962
timestamp 1679581782
transform 1 0 92928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_969
timestamp 1679581782
transform 1 0 93600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_976
timestamp 1679581782
transform 1 0 94272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_983
timestamp 1679581782
transform 1 0 94944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_990
timestamp 1679581782
transform 1 0 95616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_997
timestamp 1679581782
transform 1 0 96288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1004
timestamp 1679581782
transform 1 0 96960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1011
timestamp 1679581782
transform 1 0 97632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1018
timestamp 1679581782
transform 1 0 98304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_1025
timestamp 1679577901
transform 1 0 98976 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_0
timestamp 1677580104
transform 1 0 576 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_43
timestamp 1677580104
transform 1 0 4704 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_50
timestamp 1677580104
transform 1 0 5376 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_56
timestamp 1677579658
transform 1 0 5952 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_80
timestamp 1679577901
transform 1 0 8256 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_93
timestamp 1677579658
transform 1 0 9504 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_140
timestamp 1677580104
transform 1 0 14016 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_158
timestamp 1677579658
transform 1 0 15744 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_179
timestamp 1677580104
transform 1 0 17760 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_181
timestamp 1677579658
transform 1 0 17952 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_187
timestamp 1677579658
transform 1 0 18528 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_238
timestamp 1677580104
transform 1 0 23424 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_266
timestamp 1677579658
transform 1 0 26112 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_284
timestamp 1679577901
transform 1 0 27840 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_306
timestamp 1679577901
transform 1 0 29952 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_310
timestamp 1677579658
transform 1 0 30336 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_332
timestamp 1679581782
transform 1 0 32448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_339
timestamp 1679577901
transform 1 0 33120 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_351
timestamp 1679581782
transform 1 0 34272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_358
timestamp 1679581782
transform 1 0 34944 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_365
timestamp 1677580104
transform 1 0 35616 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_367
timestamp 1677579658
transform 1 0 35808 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_381
timestamp 1679581782
transform 1 0 37152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_388
timestamp 1679581782
transform 1 0 37824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_395
timestamp 1679577901
transform 1 0 38496 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_399
timestamp 1677580104
transform 1 0 38880 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_422
timestamp 1679581782
transform 1 0 41088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_429
timestamp 1679577901
transform 1 0 41760 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_438
timestamp 1677579658
transform 1 0 42624 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_452
timestamp 1677580104
transform 1 0 43968 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_463
timestamp 1677580104
transform 1 0 45024 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_497
timestamp 1677580104
transform 1 0 48288 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_533
timestamp 1679581782
transform 1 0 51744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_540
timestamp 1679581782
transform 1 0 52416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_547
timestamp 1679581782
transform 1 0 53088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_554
timestamp 1679581782
transform 1 0 53760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_561
timestamp 1679581782
transform 1 0 54432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_568
timestamp 1679581782
transform 1 0 55104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_575
timestamp 1679581782
transform 1 0 55776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_582
timestamp 1679581782
transform 1 0 56448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_589
timestamp 1679581782
transform 1 0 57120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_596
timestamp 1679581782
transform 1 0 57792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_603
timestamp 1679581782
transform 1 0 58464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_610
timestamp 1679581782
transform 1 0 59136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_617
timestamp 1679581782
transform 1 0 59808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_624
timestamp 1679581782
transform 1 0 60480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_631
timestamp 1679581782
transform 1 0 61152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_638
timestamp 1679581782
transform 1 0 61824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_645
timestamp 1679581782
transform 1 0 62496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_652
timestamp 1679581782
transform 1 0 63168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_659
timestamp 1679581782
transform 1 0 63840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_666
timestamp 1679581782
transform 1 0 64512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_673
timestamp 1679581782
transform 1 0 65184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_680
timestamp 1679581782
transform 1 0 65856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_687
timestamp 1679581782
transform 1 0 66528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_694
timestamp 1679581782
transform 1 0 67200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_701
timestamp 1679581782
transform 1 0 67872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_708
timestamp 1679581782
transform 1 0 68544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_715
timestamp 1679581782
transform 1 0 69216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_722
timestamp 1679581782
transform 1 0 69888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_729
timestamp 1679581782
transform 1 0 70560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_736
timestamp 1679581782
transform 1 0 71232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_743
timestamp 1679581782
transform 1 0 71904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_750
timestamp 1679581782
transform 1 0 72576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_757
timestamp 1679581782
transform 1 0 73248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_764
timestamp 1679581782
transform 1 0 73920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_771
timestamp 1679581782
transform 1 0 74592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_778
timestamp 1679581782
transform 1 0 75264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_785
timestamp 1679581782
transform 1 0 75936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_792
timestamp 1679581782
transform 1 0 76608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_799
timestamp 1679581782
transform 1 0 77280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_806
timestamp 1679581782
transform 1 0 77952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_813
timestamp 1679581782
transform 1 0 78624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_820
timestamp 1679581782
transform 1 0 79296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_827
timestamp 1679581782
transform 1 0 79968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_834
timestamp 1679581782
transform 1 0 80640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_841
timestamp 1679581782
transform 1 0 81312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_848
timestamp 1679581782
transform 1 0 81984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_855
timestamp 1679581782
transform 1 0 82656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_862
timestamp 1679581782
transform 1 0 83328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_869
timestamp 1679581782
transform 1 0 84000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_876
timestamp 1679581782
transform 1 0 84672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_883
timestamp 1679581782
transform 1 0 85344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_890
timestamp 1679581782
transform 1 0 86016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_897
timestamp 1679581782
transform 1 0 86688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_904
timestamp 1679581782
transform 1 0 87360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_911
timestamp 1679581782
transform 1 0 88032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_918
timestamp 1679581782
transform 1 0 88704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_925
timestamp 1679581782
transform 1 0 89376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_932
timestamp 1679581782
transform 1 0 90048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_939
timestamp 1679581782
transform 1 0 90720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_946
timestamp 1679581782
transform 1 0 91392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_953
timestamp 1679581782
transform 1 0 92064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_960
timestamp 1679581782
transform 1 0 92736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_967
timestamp 1679581782
transform 1 0 93408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_974
timestamp 1679581782
transform 1 0 94080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_981
timestamp 1679581782
transform 1 0 94752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_988
timestamp 1679581782
transform 1 0 95424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_995
timestamp 1679581782
transform 1 0 96096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1002
timestamp 1679581782
transform 1 0 96768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1009
timestamp 1679581782
transform 1 0 97440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1016
timestamp 1679581782
transform 1 0 98112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_1023
timestamp 1679577901
transform 1 0 98784 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_1027
timestamp 1677580104
transform 1 0 99168 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_0
timestamp 1679577901
transform 1 0 576 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_4
timestamp 1677580104
transform 1 0 960 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_69
timestamp 1677580104
transform 1 0 7200 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_71
timestamp 1677579658
transform 1 0 7392 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_85
timestamp 1679577901
transform 1 0 8736 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_125
timestamp 1677580104
transform 1 0 12576 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_155
timestamp 1679581782
transform 1 0 15456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_162
timestamp 1679577901
transform 1 0 16128 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_166
timestamp 1677580104
transform 1 0 16512 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_190
timestamp 1679577901
transform 1 0 18816 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_204
timestamp 1677580104
transform 1 0 20160 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_228
timestamp 1679581782
transform 1 0 22464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_235
timestamp 1679581782
transform 1 0 23136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_242
timestamp 1679577901
transform 1 0 23808 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_256
timestamp 1679581782
transform 1 0 25152 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_263
timestamp 1677580104
transform 1 0 25824 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_265
timestamp 1677579658
transform 1 0 26016 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_270
timestamp 1679577901
transform 1 0 26496 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_274
timestamp 1677580104
transform 1 0 26880 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_289
timestamp 1679577901
transform 1 0 28320 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_298
timestamp 1677580104
transform 1 0 29184 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_304
timestamp 1677579658
transform 1 0 29760 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_313
timestamp 1677580104
transform 1 0 30624 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_408
timestamp 1677580104
transform 1 0 39744 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_410
timestamp 1677579658
transform 1 0 39936 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_424
timestamp 1679577901
transform 1 0 41280 0 1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_34_464
timestamp 1679577901
transform 1 0 45120 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_509
timestamp 1677579658
transform 1 0 49440 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_537
timestamp 1679581782
transform 1 0 52128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_544
timestamp 1679581782
transform 1 0 52800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_551
timestamp 1679581782
transform 1 0 53472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_558
timestamp 1679581782
transform 1 0 54144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_565
timestamp 1679581782
transform 1 0 54816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_572
timestamp 1679581782
transform 1 0 55488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_579
timestamp 1679581782
transform 1 0 56160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_586
timestamp 1679581782
transform 1 0 56832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_593
timestamp 1679581782
transform 1 0 57504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_600
timestamp 1679581782
transform 1 0 58176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_607
timestamp 1679581782
transform 1 0 58848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_614
timestamp 1679581782
transform 1 0 59520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_621
timestamp 1679581782
transform 1 0 60192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_628
timestamp 1679581782
transform 1 0 60864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_635
timestamp 1679581782
transform 1 0 61536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_642
timestamp 1679581782
transform 1 0 62208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_649
timestamp 1679581782
transform 1 0 62880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_656
timestamp 1679581782
transform 1 0 63552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_663
timestamp 1679581782
transform 1 0 64224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_670
timestamp 1679581782
transform 1 0 64896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_677
timestamp 1679581782
transform 1 0 65568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_684
timestamp 1679581782
transform 1 0 66240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_691
timestamp 1679581782
transform 1 0 66912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_698
timestamp 1679581782
transform 1 0 67584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_705
timestamp 1679581782
transform 1 0 68256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_712
timestamp 1679581782
transform 1 0 68928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_719
timestamp 1679581782
transform 1 0 69600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_726
timestamp 1679581782
transform 1 0 70272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_733
timestamp 1679581782
transform 1 0 70944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_740
timestamp 1679581782
transform 1 0 71616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_747
timestamp 1679581782
transform 1 0 72288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_754
timestamp 1679581782
transform 1 0 72960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_761
timestamp 1679581782
transform 1 0 73632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_768
timestamp 1679581782
transform 1 0 74304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_775
timestamp 1679581782
transform 1 0 74976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_782
timestamp 1679581782
transform 1 0 75648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_789
timestamp 1679581782
transform 1 0 76320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_796
timestamp 1679581782
transform 1 0 76992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_803
timestamp 1679581782
transform 1 0 77664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_810
timestamp 1679581782
transform 1 0 78336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_817
timestamp 1679581782
transform 1 0 79008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_824
timestamp 1679581782
transform 1 0 79680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_831
timestamp 1679581782
transform 1 0 80352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_838
timestamp 1679581782
transform 1 0 81024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_845
timestamp 1679581782
transform 1 0 81696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_852
timestamp 1679581782
transform 1 0 82368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_859
timestamp 1679581782
transform 1 0 83040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_866
timestamp 1679581782
transform 1 0 83712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_873
timestamp 1679581782
transform 1 0 84384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_880
timestamp 1679581782
transform 1 0 85056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_887
timestamp 1679581782
transform 1 0 85728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_894
timestamp 1679581782
transform 1 0 86400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_901
timestamp 1679581782
transform 1 0 87072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_908
timestamp 1679581782
transform 1 0 87744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_915
timestamp 1679581782
transform 1 0 88416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_922
timestamp 1679581782
transform 1 0 89088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_929
timestamp 1679581782
transform 1 0 89760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_936
timestamp 1679581782
transform 1 0 90432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_943
timestamp 1679581782
transform 1 0 91104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_950
timestamp 1679581782
transform 1 0 91776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_957
timestamp 1679581782
transform 1 0 92448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_964
timestamp 1679581782
transform 1 0 93120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_971
timestamp 1679581782
transform 1 0 93792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_978
timestamp 1679581782
transform 1 0 94464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_985
timestamp 1679581782
transform 1 0 95136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_992
timestamp 1679581782
transform 1 0 95808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_999
timestamp 1679581782
transform 1 0 96480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1006
timestamp 1679581782
transform 1 0 97152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1013
timestamp 1679581782
transform 1 0 97824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1020
timestamp 1679581782
transform 1 0 98496 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_1027
timestamp 1677580104
transform 1 0 99168 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_7
timestamp 1679577901
transform 1 0 1248 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_15
timestamp 1679577901
transform 1 0 2016 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_19
timestamp 1677580104
transform 1 0 2400 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_35
timestamp 1677579658
transform 1 0 3936 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_49
timestamp 1677579658
transform 1 0 5280 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_114
timestamp 1677579658
transform 1 0 11520 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_128
timestamp 1677580104
transform 1 0 12864 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_143
timestamp 1679577901
transform 1 0 14304 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_155
timestamp 1679577901
transform 1 0 15456 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_159
timestamp 1677579658
transform 1 0 15840 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_165
timestamp 1679581782
transform 1 0 16416 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_172
timestamp 1677580104
transform 1 0 17088 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_187
timestamp 1679577901
transform 1 0 18528 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_191
timestamp 1677580104
transform 1 0 18912 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_220
timestamp 1677579658
transform 1 0 21696 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_248
timestamp 1677580104
transform 1 0 24384 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_305
timestamp 1679577901
transform 1 0 29856 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_309
timestamp 1677580104
transform 1 0 30240 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_330
timestamp 1679577901
transform 1 0 32256 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_334
timestamp 1677580104
transform 1 0 32640 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_354
timestamp 1679577901
transform 1 0 34560 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_375
timestamp 1677580104
transform 1 0 36576 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_377
timestamp 1677579658
transform 1 0 36768 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_382
timestamp 1679577901
transform 1 0 37248 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_389
timestamp 1677580104
transform 1 0 37920 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_396
timestamp 1677580104
transform 1 0 38592 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_398
timestamp 1677579658
transform 1 0 38784 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_408
timestamp 1677579658
transform 1 0 39744 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_414
timestamp 1679581782
transform 1 0 40320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_421
timestamp 1679581782
transform 1 0 40992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_428
timestamp 1679577901
transform 1 0 41664 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_432
timestamp 1677579658
transform 1 0 42048 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_437
timestamp 1677580104
transform 1 0 42528 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_439
timestamp 1677579658
transform 1 0 42720 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_453
timestamp 1677580104
transform 1 0 44064 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_459
timestamp 1679577901
transform 1 0 44640 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_35_468
timestamp 1679577901
transform 1 0 45504 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_481
timestamp 1677579658
transform 1 0 46752 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_493
timestamp 1677580104
transform 1 0 47904 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_505
timestamp 1677579658
transform 1 0 49056 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_533
timestamp 1679581782
transform 1 0 51744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_540
timestamp 1679581782
transform 1 0 52416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_547
timestamp 1679581782
transform 1 0 53088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_554
timestamp 1679581782
transform 1 0 53760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_561
timestamp 1679581782
transform 1 0 54432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_568
timestamp 1679581782
transform 1 0 55104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_575
timestamp 1679581782
transform 1 0 55776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_582
timestamp 1679581782
transform 1 0 56448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_589
timestamp 1679581782
transform 1 0 57120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_596
timestamp 1679581782
transform 1 0 57792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_603
timestamp 1679581782
transform 1 0 58464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_610
timestamp 1679581782
transform 1 0 59136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_617
timestamp 1679581782
transform 1 0 59808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_624
timestamp 1679581782
transform 1 0 60480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_631
timestamp 1679581782
transform 1 0 61152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_638
timestamp 1679581782
transform 1 0 61824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_645
timestamp 1679581782
transform 1 0 62496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_652
timestamp 1679581782
transform 1 0 63168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_659
timestamp 1679581782
transform 1 0 63840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_666
timestamp 1679581782
transform 1 0 64512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_673
timestamp 1679581782
transform 1 0 65184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_680
timestamp 1679581782
transform 1 0 65856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_687
timestamp 1679581782
transform 1 0 66528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_694
timestamp 1679581782
transform 1 0 67200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_701
timestamp 1679581782
transform 1 0 67872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_708
timestamp 1679581782
transform 1 0 68544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_715
timestamp 1679581782
transform 1 0 69216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_722
timestamp 1679581782
transform 1 0 69888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_729
timestamp 1679581782
transform 1 0 70560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_736
timestamp 1679581782
transform 1 0 71232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_743
timestamp 1679581782
transform 1 0 71904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_750
timestamp 1679581782
transform 1 0 72576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_757
timestamp 1679581782
transform 1 0 73248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_764
timestamp 1679581782
transform 1 0 73920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_771
timestamp 1679581782
transform 1 0 74592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_778
timestamp 1679581782
transform 1 0 75264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_785
timestamp 1679581782
transform 1 0 75936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_792
timestamp 1679581782
transform 1 0 76608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_799
timestamp 1679581782
transform 1 0 77280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_806
timestamp 1679581782
transform 1 0 77952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_813
timestamp 1679581782
transform 1 0 78624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_820
timestamp 1679581782
transform 1 0 79296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_827
timestamp 1679581782
transform 1 0 79968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_834
timestamp 1679581782
transform 1 0 80640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_841
timestamp 1679581782
transform 1 0 81312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_848
timestamp 1679581782
transform 1 0 81984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_855
timestamp 1679581782
transform 1 0 82656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_862
timestamp 1679581782
transform 1 0 83328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_869
timestamp 1679581782
transform 1 0 84000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_876
timestamp 1679581782
transform 1 0 84672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_883
timestamp 1679581782
transform 1 0 85344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_890
timestamp 1679581782
transform 1 0 86016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_897
timestamp 1679581782
transform 1 0 86688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_904
timestamp 1679581782
transform 1 0 87360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_911
timestamp 1679581782
transform 1 0 88032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_918
timestamp 1679581782
transform 1 0 88704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_925
timestamp 1679581782
transform 1 0 89376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_932
timestamp 1679581782
transform 1 0 90048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_939
timestamp 1679581782
transform 1 0 90720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_946
timestamp 1679581782
transform 1 0 91392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_953
timestamp 1679581782
transform 1 0 92064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_960
timestamp 1679581782
transform 1 0 92736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_967
timestamp 1679581782
transform 1 0 93408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_974
timestamp 1679581782
transform 1 0 94080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_981
timestamp 1679581782
transform 1 0 94752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_988
timestamp 1679581782
transform 1 0 95424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_995
timestamp 1679581782
transform 1 0 96096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1002
timestamp 1679581782
transform 1 0 96768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1009
timestamp 1679581782
transform 1 0 97440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1016
timestamp 1679581782
transform 1 0 98112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_1023
timestamp 1679577901
transform 1 0 98784 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_1027
timestamp 1677580104
transform 1 0 99168 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_34
timestamp 1677579658
transform 1 0 3840 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_81
timestamp 1677579658
transform 1 0 8352 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_95
timestamp 1677580104
transform 1 0 9696 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_97
timestamp 1677579658
transform 1 0 9888 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_101
timestamp 1679581782
transform 1 0 10272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_108
timestamp 1679577901
transform 1 0 10944 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_116
timestamp 1677579658
transform 1 0 11712 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_152
timestamp 1679581782
transform 1 0 15168 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_159
timestamp 1677580104
transform 1 0 15840 0 1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_165
timestamp 1679577901
transform 1 0 16416 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_169
timestamp 1677579658
transform 1 0 16800 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_183
timestamp 1679577901
transform 1 0 18144 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_187
timestamp 1677579658
transform 1 0 18528 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_193
timestamp 1677579658
transform 1 0 19104 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_215
timestamp 1679581782
transform 1 0 21216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_222
timestamp 1679577901
transform 1 0 21888 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_239
timestamp 1679581782
transform 1 0 23520 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_246
timestamp 1677579658
transform 1 0 24192 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_260
timestamp 1679577901
transform 1 0 25536 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_286
timestamp 1677580104
transform 1 0 28032 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_298
timestamp 1679581782
transform 1 0 29184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_305
timestamp 1679581782
transform 1 0 29856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_344
timestamp 1679577901
transform 1 0 33600 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_348
timestamp 1677580104
transform 1 0 33984 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_353
timestamp 1679581782
transform 1 0 34464 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_360
timestamp 1677579658
transform 1 0 35136 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_371
timestamp 1677580104
transform 1 0 36192 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_377
timestamp 1677580104
transform 1 0 36768 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_379
timestamp 1677579658
transform 1 0 36960 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_385
timestamp 1679577901
transform 1 0 37536 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_389
timestamp 1677580104
transform 1 0 37920 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_406
timestamp 1677580104
transform 1 0 39552 0 1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_471
timestamp 1679577901
transform 1 0 45792 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_475
timestamp 1677580104
transform 1 0 46176 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_531
timestamp 1679581782
transform 1 0 51552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_538
timestamp 1679581782
transform 1 0 52224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_545
timestamp 1679581782
transform 1 0 52896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_552
timestamp 1679581782
transform 1 0 53568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_559
timestamp 1679581782
transform 1 0 54240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_566
timestamp 1679581782
transform 1 0 54912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_573
timestamp 1679581782
transform 1 0 55584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_580
timestamp 1679581782
transform 1 0 56256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_587
timestamp 1679581782
transform 1 0 56928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_594
timestamp 1679581782
transform 1 0 57600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_601
timestamp 1679581782
transform 1 0 58272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_608
timestamp 1679581782
transform 1 0 58944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_615
timestamp 1679581782
transform 1 0 59616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_622
timestamp 1679581782
transform 1 0 60288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_629
timestamp 1679581782
transform 1 0 60960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_636
timestamp 1679581782
transform 1 0 61632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_643
timestamp 1679581782
transform 1 0 62304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_650
timestamp 1679581782
transform 1 0 62976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_657
timestamp 1679581782
transform 1 0 63648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_664
timestamp 1679581782
transform 1 0 64320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_671
timestamp 1679581782
transform 1 0 64992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_678
timestamp 1679581782
transform 1 0 65664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_685
timestamp 1679581782
transform 1 0 66336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_692
timestamp 1679581782
transform 1 0 67008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_699
timestamp 1679581782
transform 1 0 67680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_706
timestamp 1679581782
transform 1 0 68352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_713
timestamp 1679581782
transform 1 0 69024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_720
timestamp 1679581782
transform 1 0 69696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_727
timestamp 1679581782
transform 1 0 70368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_734
timestamp 1679581782
transform 1 0 71040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_741
timestamp 1679581782
transform 1 0 71712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_748
timestamp 1679581782
transform 1 0 72384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_755
timestamp 1679581782
transform 1 0 73056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_762
timestamp 1679581782
transform 1 0 73728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_769
timestamp 1679581782
transform 1 0 74400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_776
timestamp 1679581782
transform 1 0 75072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_783
timestamp 1679581782
transform 1 0 75744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_790
timestamp 1679581782
transform 1 0 76416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_797
timestamp 1679581782
transform 1 0 77088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_804
timestamp 1679581782
transform 1 0 77760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_811
timestamp 1679581782
transform 1 0 78432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_818
timestamp 1679581782
transform 1 0 79104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_825
timestamp 1679581782
transform 1 0 79776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_832
timestamp 1679581782
transform 1 0 80448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_839
timestamp 1679581782
transform 1 0 81120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_846
timestamp 1679581782
transform 1 0 81792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_853
timestamp 1679581782
transform 1 0 82464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_860
timestamp 1679581782
transform 1 0 83136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_867
timestamp 1679581782
transform 1 0 83808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_874
timestamp 1679581782
transform 1 0 84480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_881
timestamp 1679581782
transform 1 0 85152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_888
timestamp 1679581782
transform 1 0 85824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_895
timestamp 1679581782
transform 1 0 86496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_902
timestamp 1679581782
transform 1 0 87168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_909
timestamp 1679581782
transform 1 0 87840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_916
timestamp 1679581782
transform 1 0 88512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_923
timestamp 1679581782
transform 1 0 89184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_930
timestamp 1679581782
transform 1 0 89856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_937
timestamp 1679581782
transform 1 0 90528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_944
timestamp 1679581782
transform 1 0 91200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_951
timestamp 1679581782
transform 1 0 91872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_958
timestamp 1679581782
transform 1 0 92544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_965
timestamp 1679581782
transform 1 0 93216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_972
timestamp 1679581782
transform 1 0 93888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_979
timestamp 1679581782
transform 1 0 94560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_986
timestamp 1679581782
transform 1 0 95232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_993
timestamp 1679581782
transform 1 0 95904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1000
timestamp 1679581782
transform 1 0 96576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1007
timestamp 1679581782
transform 1 0 97248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1014
timestamp 1679581782
transform 1 0 97920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1021
timestamp 1679581782
transform 1 0 98592 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_1028
timestamp 1677579658
transform 1 0 99264 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_7
timestamp 1679577901
transform 1 0 1248 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_11
timestamp 1677579658
transform 1 0 1632 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_16
timestamp 1679577901
transform 1 0 2112 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_20
timestamp 1677580104
transform 1 0 2496 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_45
timestamp 1677579658
transform 1 0 4896 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_99
timestamp 1679581782
transform 1 0 10080 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_106
timestamp 1677579658
transform 1 0 10752 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_134
timestamp 1679577901
transform 1 0 13440 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_148
timestamp 1677580104
transform 1 0 14784 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_163
timestamp 1677580104
transform 1 0 16224 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_234
timestamp 1679581782
transform 1 0 23040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_241
timestamp 1679581782
transform 1 0 23712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_248
timestamp 1679581782
transform 1 0 24384 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_255
timestamp 1677579658
transform 1 0 25056 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_260
timestamp 1679581782
transform 1 0 25536 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_282
timestamp 1677580104
transform 1 0 27648 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_292
timestamp 1679577901
transform 1 0 28608 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_301
timestamp 1677580104
transform 1 0 29472 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_303
timestamp 1677579658
transform 1 0 29664 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_395
timestamp 1677580104
transform 1 0 38496 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_397
timestamp 1677579658
transform 1 0 38688 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_411
timestamp 1679581782
transform 1 0 40032 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_418
timestamp 1677579658
transform 1 0 40704 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_473
timestamp 1679581782
transform 1 0 45984 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_480
timestamp 1677580104
transform 1 0 46656 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_482
timestamp 1677579658
transform 1 0 46848 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_496
timestamp 1677579658
transform 1 0 48192 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_533
timestamp 1679581782
transform 1 0 51744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_540
timestamp 1679581782
transform 1 0 52416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_547
timestamp 1679581782
transform 1 0 53088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_554
timestamp 1679581782
transform 1 0 53760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_561
timestamp 1679581782
transform 1 0 54432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_568
timestamp 1679581782
transform 1 0 55104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_575
timestamp 1679581782
transform 1 0 55776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_582
timestamp 1679581782
transform 1 0 56448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_589
timestamp 1679581782
transform 1 0 57120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_596
timestamp 1679581782
transform 1 0 57792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_603
timestamp 1679581782
transform 1 0 58464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_610
timestamp 1679581782
transform 1 0 59136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_617
timestamp 1679581782
transform 1 0 59808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_624
timestamp 1679581782
transform 1 0 60480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_631
timestamp 1679581782
transform 1 0 61152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_638
timestamp 1679581782
transform 1 0 61824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_645
timestamp 1679581782
transform 1 0 62496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_652
timestamp 1679581782
transform 1 0 63168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_659
timestamp 1679581782
transform 1 0 63840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_666
timestamp 1679581782
transform 1 0 64512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_673
timestamp 1679581782
transform 1 0 65184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_680
timestamp 1679581782
transform 1 0 65856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_687
timestamp 1679581782
transform 1 0 66528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_694
timestamp 1679581782
transform 1 0 67200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_701
timestamp 1679581782
transform 1 0 67872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_708
timestamp 1679581782
transform 1 0 68544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_715
timestamp 1679581782
transform 1 0 69216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_722
timestamp 1679581782
transform 1 0 69888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_729
timestamp 1679581782
transform 1 0 70560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_736
timestamp 1679581782
transform 1 0 71232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_743
timestamp 1679581782
transform 1 0 71904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_750
timestamp 1679581782
transform 1 0 72576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_757
timestamp 1679581782
transform 1 0 73248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_764
timestamp 1679581782
transform 1 0 73920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_771
timestamp 1679581782
transform 1 0 74592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_778
timestamp 1679581782
transform 1 0 75264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_785
timestamp 1679581782
transform 1 0 75936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_792
timestamp 1679581782
transform 1 0 76608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_799
timestamp 1679581782
transform 1 0 77280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_806
timestamp 1679581782
transform 1 0 77952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_813
timestamp 1679581782
transform 1 0 78624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_820
timestamp 1679581782
transform 1 0 79296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_827
timestamp 1679581782
transform 1 0 79968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_834
timestamp 1679581782
transform 1 0 80640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_841
timestamp 1679581782
transform 1 0 81312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_848
timestamp 1679581782
transform 1 0 81984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_855
timestamp 1679581782
transform 1 0 82656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_862
timestamp 1679581782
transform 1 0 83328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_869
timestamp 1679581782
transform 1 0 84000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_876
timestamp 1679581782
transform 1 0 84672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_883
timestamp 1679581782
transform 1 0 85344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_890
timestamp 1679581782
transform 1 0 86016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_897
timestamp 1679581782
transform 1 0 86688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_904
timestamp 1679581782
transform 1 0 87360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_911
timestamp 1679581782
transform 1 0 88032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_918
timestamp 1679581782
transform 1 0 88704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_925
timestamp 1679581782
transform 1 0 89376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_932
timestamp 1679581782
transform 1 0 90048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_939
timestamp 1679581782
transform 1 0 90720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_946
timestamp 1679581782
transform 1 0 91392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_953
timestamp 1679581782
transform 1 0 92064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_960
timestamp 1679581782
transform 1 0 92736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_967
timestamp 1679581782
transform 1 0 93408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_974
timestamp 1679581782
transform 1 0 94080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_981
timestamp 1679581782
transform 1 0 94752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_988
timestamp 1679581782
transform 1 0 95424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_995
timestamp 1679581782
transform 1 0 96096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1002
timestamp 1679581782
transform 1 0 96768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1009
timestamp 1679581782
transform 1 0 97440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1016
timestamp 1679581782
transform 1 0 98112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_1023
timestamp 1679577901
transform 1 0 98784 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_1027
timestamp 1677580104
transform 1 0 99168 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_0
timestamp 1677580104
transform 1 0 576 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_33
timestamp 1677580104
transform 1 0 3744 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_70
timestamp 1677580104
transform 1 0 7296 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_113
timestamp 1677579658
transform 1 0 11424 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_143
timestamp 1677579658
transform 1 0 14304 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_176
timestamp 1679581782
transform 1 0 17472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_183
timestamp 1679577901
transform 1 0 18144 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_205
timestamp 1677579658
transform 1 0 20256 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_228
timestamp 1679577901
transform 1 0 22464 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_272
timestamp 1677580104
transform 1 0 26688 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_293
timestamp 1677579658
transform 1 0 28704 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_366
timestamp 1677580104
transform 1 0 35712 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_382
timestamp 1677579658
transform 1 0 37248 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_388
timestamp 1679577901
transform 1 0 37824 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_493
timestamp 1677580104
transform 1 0 47904 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_522
timestamp 1679581782
transform 1 0 50688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_529
timestamp 1679581782
transform 1 0 51360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_536
timestamp 1679581782
transform 1 0 52032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_543
timestamp 1679581782
transform 1 0 52704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_550
timestamp 1679581782
transform 1 0 53376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_557
timestamp 1679581782
transform 1 0 54048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_564
timestamp 1679581782
transform 1 0 54720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_571
timestamp 1679581782
transform 1 0 55392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_578
timestamp 1679581782
transform 1 0 56064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_585
timestamp 1679581782
transform 1 0 56736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_592
timestamp 1679581782
transform 1 0 57408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_599
timestamp 1679581782
transform 1 0 58080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_606
timestamp 1679581782
transform 1 0 58752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_613
timestamp 1679581782
transform 1 0 59424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_620
timestamp 1679581782
transform 1 0 60096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_627
timestamp 1679581782
transform 1 0 60768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_634
timestamp 1679581782
transform 1 0 61440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_641
timestamp 1679581782
transform 1 0 62112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_648
timestamp 1679581782
transform 1 0 62784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_655
timestamp 1679581782
transform 1 0 63456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_662
timestamp 1679581782
transform 1 0 64128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_669
timestamp 1679581782
transform 1 0 64800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_676
timestamp 1679581782
transform 1 0 65472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_683
timestamp 1679581782
transform 1 0 66144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_690
timestamp 1679581782
transform 1 0 66816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_697
timestamp 1679581782
transform 1 0 67488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_704
timestamp 1679581782
transform 1 0 68160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_711
timestamp 1679581782
transform 1 0 68832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_718
timestamp 1679581782
transform 1 0 69504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_725
timestamp 1679581782
transform 1 0 70176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_732
timestamp 1679581782
transform 1 0 70848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_739
timestamp 1679581782
transform 1 0 71520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_746
timestamp 1679581782
transform 1 0 72192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_753
timestamp 1679581782
transform 1 0 72864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_760
timestamp 1679581782
transform 1 0 73536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_767
timestamp 1679581782
transform 1 0 74208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_774
timestamp 1679581782
transform 1 0 74880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_781
timestamp 1679581782
transform 1 0 75552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_788
timestamp 1679581782
transform 1 0 76224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_795
timestamp 1679581782
transform 1 0 76896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_802
timestamp 1679581782
transform 1 0 77568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_809
timestamp 1679581782
transform 1 0 78240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_816
timestamp 1679581782
transform 1 0 78912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_823
timestamp 1679581782
transform 1 0 79584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_830
timestamp 1679581782
transform 1 0 80256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_837
timestamp 1679581782
transform 1 0 80928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_844
timestamp 1679581782
transform 1 0 81600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_851
timestamp 1679581782
transform 1 0 82272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_858
timestamp 1679581782
transform 1 0 82944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_865
timestamp 1679581782
transform 1 0 83616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_872
timestamp 1679581782
transform 1 0 84288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_879
timestamp 1679581782
transform 1 0 84960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_886
timestamp 1679581782
transform 1 0 85632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_893
timestamp 1679581782
transform 1 0 86304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_900
timestamp 1679581782
transform 1 0 86976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_907
timestamp 1679581782
transform 1 0 87648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_914
timestamp 1679581782
transform 1 0 88320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_921
timestamp 1679581782
transform 1 0 88992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_928
timestamp 1679581782
transform 1 0 89664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_935
timestamp 1679581782
transform 1 0 90336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_942
timestamp 1679581782
transform 1 0 91008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_949
timestamp 1679581782
transform 1 0 91680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_956
timestamp 1679581782
transform 1 0 92352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_963
timestamp 1679581782
transform 1 0 93024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_970
timestamp 1679581782
transform 1 0 93696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_977
timestamp 1679581782
transform 1 0 94368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_984
timestamp 1679581782
transform 1 0 95040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_991
timestamp 1679581782
transform 1 0 95712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_998
timestamp 1679581782
transform 1 0 96384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1005
timestamp 1679581782
transform 1 0 97056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1012
timestamp 1679581782
transform 1 0 97728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1019
timestamp 1679581782
transform 1 0 98400 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_1026
timestamp 1677580104
transform 1 0 99072 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_1028
timestamp 1677579658
transform 1 0 99264 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_34
timestamp 1677579658
transform 1 0 3840 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_53
timestamp 1677580104
transform 1 0 5664 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_85
timestamp 1677580104
transform 1 0 8736 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_100
timestamp 1679581782
transform 1 0 10176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_165
timestamp 1679581782
transform 1 0 16416 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_172
timestamp 1677580104
transform 1 0 17088 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_174
timestamp 1677579658
transform 1 0 17280 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_179
timestamp 1679581782
transform 1 0 17760 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_186
timestamp 1677580104
transform 1 0 18432 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_256
timestamp 1677580104
transform 1 0 25152 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_258
timestamp 1677579658
transform 1 0 25344 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_287
timestamp 1677580104
transform 1 0 28128 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_294
timestamp 1677580104
transform 1 0 28800 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_325
timestamp 1677579658
transform 1 0 31776 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_366
timestamp 1677580104
transform 1 0 35712 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_377
timestamp 1677580104
transform 1 0 36768 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_383
timestamp 1679581782
transform 1 0 37344 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_432
timestamp 1677579658
transform 1 0 42048 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_476
timestamp 1677579658
transform 1 0 46272 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_488
timestamp 1677580104
transform 1 0 47424 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_495
timestamp 1677579658
transform 1 0 48096 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_501
timestamp 1677580104
transform 1 0 48672 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_520
timestamp 1679581782
transform 1 0 50496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_527
timestamp 1679581782
transform 1 0 51168 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_534
timestamp 1679581782
transform 1 0 51840 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_541
timestamp 1679581782
transform 1 0 52512 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_548
timestamp 1679581782
transform 1 0 53184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_555
timestamp 1679581782
transform 1 0 53856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_562
timestamp 1679581782
transform 1 0 54528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_569
timestamp 1679581782
transform 1 0 55200 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_576
timestamp 1679581782
transform 1 0 55872 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_583
timestamp 1679581782
transform 1 0 56544 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_590
timestamp 1679581782
transform 1 0 57216 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_597
timestamp 1679581782
transform 1 0 57888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_604
timestamp 1679581782
transform 1 0 58560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_611
timestamp 1679581782
transform 1 0 59232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_618
timestamp 1679581782
transform 1 0 59904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_625
timestamp 1679581782
transform 1 0 60576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_632
timestamp 1679581782
transform 1 0 61248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_639
timestamp 1679581782
transform 1 0 61920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_646
timestamp 1679581782
transform 1 0 62592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_653
timestamp 1679581782
transform 1 0 63264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_660
timestamp 1679581782
transform 1 0 63936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_667
timestamp 1679581782
transform 1 0 64608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_674
timestamp 1679581782
transform 1 0 65280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_681
timestamp 1679581782
transform 1 0 65952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_688
timestamp 1679581782
transform 1 0 66624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_695
timestamp 1679581782
transform 1 0 67296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_702
timestamp 1679581782
transform 1 0 67968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_709
timestamp 1679581782
transform 1 0 68640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_716
timestamp 1679581782
transform 1 0 69312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_723
timestamp 1679581782
transform 1 0 69984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_730
timestamp 1679581782
transform 1 0 70656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_737
timestamp 1679581782
transform 1 0 71328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_744
timestamp 1679581782
transform 1 0 72000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_751
timestamp 1679581782
transform 1 0 72672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_758
timestamp 1679581782
transform 1 0 73344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_765
timestamp 1679581782
transform 1 0 74016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_772
timestamp 1679581782
transform 1 0 74688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_779
timestamp 1679581782
transform 1 0 75360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_786
timestamp 1679581782
transform 1 0 76032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_793
timestamp 1679581782
transform 1 0 76704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_800
timestamp 1679581782
transform 1 0 77376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_807
timestamp 1679581782
transform 1 0 78048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_814
timestamp 1679581782
transform 1 0 78720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_821
timestamp 1679581782
transform 1 0 79392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_828
timestamp 1679581782
transform 1 0 80064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_835
timestamp 1679581782
transform 1 0 80736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_842
timestamp 1679581782
transform 1 0 81408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_849
timestamp 1679581782
transform 1 0 82080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_856
timestamp 1679581782
transform 1 0 82752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_863
timestamp 1679581782
transform 1 0 83424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_870
timestamp 1679581782
transform 1 0 84096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_877
timestamp 1679581782
transform 1 0 84768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_884
timestamp 1679581782
transform 1 0 85440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_891
timestamp 1679581782
transform 1 0 86112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_898
timestamp 1679581782
transform 1 0 86784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_905
timestamp 1679581782
transform 1 0 87456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_912
timestamp 1679581782
transform 1 0 88128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_919
timestamp 1679581782
transform 1 0 88800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_926
timestamp 1679581782
transform 1 0 89472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_933
timestamp 1679581782
transform 1 0 90144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_940
timestamp 1679581782
transform 1 0 90816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_947
timestamp 1679581782
transform 1 0 91488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_954
timestamp 1679581782
transform 1 0 92160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_961
timestamp 1679581782
transform 1 0 92832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_968
timestamp 1679581782
transform 1 0 93504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_975
timestamp 1679581782
transform 1 0 94176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_982
timestamp 1679581782
transform 1 0 94848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_989
timestamp 1679581782
transform 1 0 95520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_996
timestamp 1679581782
transform 1 0 96192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1003
timestamp 1679581782
transform 1 0 96864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1010
timestamp 1679581782
transform 1 0 97536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1017
timestamp 1679581782
transform 1 0 98208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_1024
timestamp 1679577901
transform 1 0 98880 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_1028
timestamp 1677579658
transform 1 0 99264 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_7
timestamp 1679577901
transform 1 0 1248 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_11
timestamp 1677580104
transform 1 0 1632 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_17
timestamp 1679581782
transform 1 0 2208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_24
timestamp 1679577901
transform 1 0 2880 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_28
timestamp 1677579658
transform 1 0 3264 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_53
timestamp 1677580104
transform 1 0 5664 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_96
timestamp 1677579658
transform 1 0 9792 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_150
timestamp 1677580104
transform 1 0 14976 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_164
timestamp 1677579658
transform 1 0 16320 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_218
timestamp 1679581782
transform 1 0 21504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_225
timestamp 1679577901
transform 1 0 22176 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_229
timestamp 1677580104
transform 1 0 22560 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_235
timestamp 1679581782
transform 1 0 23136 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_242
timestamp 1677580104
transform 1 0 23808 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_260
timestamp 1677580104
transform 1 0 25536 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_262
timestamp 1677579658
transform 1 0 25728 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_277
timestamp 1677579658
transform 1 0 27168 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_334
timestamp 1677580104
transform 1 0 32640 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_355
timestamp 1677580104
transform 1 0 34656 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_357
timestamp 1677579658
transform 1 0 34848 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_385
timestamp 1679577901
transform 1 0 37536 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_389
timestamp 1677579658
transform 1 0 37920 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_513
timestamp 1679581782
transform 1 0 49824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_520
timestamp 1679581782
transform 1 0 50496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_527
timestamp 1679581782
transform 1 0 51168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_534
timestamp 1679581782
transform 1 0 51840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_541
timestamp 1679581782
transform 1 0 52512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_548
timestamp 1679581782
transform 1 0 53184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_555
timestamp 1679581782
transform 1 0 53856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_562
timestamp 1679581782
transform 1 0 54528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_569
timestamp 1679581782
transform 1 0 55200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_576
timestamp 1679581782
transform 1 0 55872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_583
timestamp 1679581782
transform 1 0 56544 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_590
timestamp 1679581782
transform 1 0 57216 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_597
timestamp 1679581782
transform 1 0 57888 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_604
timestamp 1679581782
transform 1 0 58560 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_611
timestamp 1679581782
transform 1 0 59232 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_618
timestamp 1679581782
transform 1 0 59904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_625
timestamp 1679581782
transform 1 0 60576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_632
timestamp 1679581782
transform 1 0 61248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_639
timestamp 1679581782
transform 1 0 61920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_646
timestamp 1679581782
transform 1 0 62592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_653
timestamp 1679581782
transform 1 0 63264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_660
timestamp 1679581782
transform 1 0 63936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_667
timestamp 1679581782
transform 1 0 64608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_674
timestamp 1679581782
transform 1 0 65280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_681
timestamp 1679581782
transform 1 0 65952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_688
timestamp 1679581782
transform 1 0 66624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_695
timestamp 1679581782
transform 1 0 67296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_702
timestamp 1679581782
transform 1 0 67968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_709
timestamp 1679581782
transform 1 0 68640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_716
timestamp 1679581782
transform 1 0 69312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_723
timestamp 1679581782
transform 1 0 69984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_730
timestamp 1679581782
transform 1 0 70656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_737
timestamp 1679581782
transform 1 0 71328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_744
timestamp 1679581782
transform 1 0 72000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_751
timestamp 1679581782
transform 1 0 72672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_758
timestamp 1679581782
transform 1 0 73344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_765
timestamp 1679581782
transform 1 0 74016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_772
timestamp 1679581782
transform 1 0 74688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_779
timestamp 1679581782
transform 1 0 75360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_786
timestamp 1679581782
transform 1 0 76032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_793
timestamp 1679581782
transform 1 0 76704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_800
timestamp 1679581782
transform 1 0 77376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_807
timestamp 1679581782
transform 1 0 78048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_814
timestamp 1679581782
transform 1 0 78720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_821
timestamp 1679581782
transform 1 0 79392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_828
timestamp 1679581782
transform 1 0 80064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_835
timestamp 1679581782
transform 1 0 80736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_842
timestamp 1679581782
transform 1 0 81408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_849
timestamp 1679581782
transform 1 0 82080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_856
timestamp 1679581782
transform 1 0 82752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_863
timestamp 1679581782
transform 1 0 83424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_870
timestamp 1679581782
transform 1 0 84096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_877
timestamp 1679581782
transform 1 0 84768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_884
timestamp 1679581782
transform 1 0 85440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_891
timestamp 1679581782
transform 1 0 86112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_898
timestamp 1679581782
transform 1 0 86784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_905
timestamp 1679581782
transform 1 0 87456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_912
timestamp 1679581782
transform 1 0 88128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_919
timestamp 1679581782
transform 1 0 88800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_926
timestamp 1679581782
transform 1 0 89472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_933
timestamp 1679581782
transform 1 0 90144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_940
timestamp 1679581782
transform 1 0 90816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_947
timestamp 1679581782
transform 1 0 91488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_954
timestamp 1679581782
transform 1 0 92160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_961
timestamp 1679581782
transform 1 0 92832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_968
timestamp 1679581782
transform 1 0 93504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_975
timestamp 1679581782
transform 1 0 94176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_982
timestamp 1679581782
transform 1 0 94848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_989
timestamp 1679581782
transform 1 0 95520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_996
timestamp 1679581782
transform 1 0 96192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1003
timestamp 1679581782
transform 1 0 96864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1010
timestamp 1679581782
transform 1 0 97536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1017
timestamp 1679581782
transform 1 0 98208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_1024
timestamp 1679577901
transform 1 0 98880 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_1028
timestamp 1677579658
transform 1 0 99264 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_34
timestamp 1677580104
transform 1 0 3840 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_75
timestamp 1677579658
transform 1 0 7776 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_179
timestamp 1677579658
transform 1 0 17760 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_230
timestamp 1679581782
transform 1 0 22656 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_237
timestamp 1677579658
transform 1 0 23328 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_243
timestamp 1679581782
transform 1 0 23904 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_250
timestamp 1677580104
transform 1 0 24576 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_324
timestamp 1677579658
transform 1 0 31680 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_371
timestamp 1677580104
transform 1 0 36192 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_373
timestamp 1677579658
transform 1 0 36384 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_377
timestamp 1679581782
transform 1 0 36768 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_384
timestamp 1677579658
transform 1 0 37440 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_397
timestamp 1677579658
transform 1 0 38688 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_427
timestamp 1677580104
transform 1 0 41568 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_429
timestamp 1677579658
transform 1 0 41760 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_458
timestamp 1677579658
transform 1 0 44544 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_486
timestamp 1677579658
transform 1 0 47232 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_501
timestamp 1679577901
transform 1 0 48672 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_514
timestamp 1679581782
transform 1 0 49920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_521
timestamp 1679581782
transform 1 0 50592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_528
timestamp 1679581782
transform 1 0 51264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_535
timestamp 1679581782
transform 1 0 51936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_542
timestamp 1679581782
transform 1 0 52608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_549
timestamp 1679581782
transform 1 0 53280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_556
timestamp 1679581782
transform 1 0 53952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_563
timestamp 1679581782
transform 1 0 54624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_570
timestamp 1679581782
transform 1 0 55296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_577
timestamp 1679581782
transform 1 0 55968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_584
timestamp 1679581782
transform 1 0 56640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_591
timestamp 1679581782
transform 1 0 57312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_598
timestamp 1679581782
transform 1 0 57984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_605
timestamp 1679581782
transform 1 0 58656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_612
timestamp 1679581782
transform 1 0 59328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_619
timestamp 1679581782
transform 1 0 60000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_626
timestamp 1679581782
transform 1 0 60672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_633
timestamp 1679581782
transform 1 0 61344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_640
timestamp 1679581782
transform 1 0 62016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_647
timestamp 1679581782
transform 1 0 62688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_654
timestamp 1679581782
transform 1 0 63360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_661
timestamp 1679581782
transform 1 0 64032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_668
timestamp 1679581782
transform 1 0 64704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_675
timestamp 1679581782
transform 1 0 65376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_682
timestamp 1679581782
transform 1 0 66048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_689
timestamp 1679581782
transform 1 0 66720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_696
timestamp 1679581782
transform 1 0 67392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_703
timestamp 1679581782
transform 1 0 68064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_710
timestamp 1679581782
transform 1 0 68736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_717
timestamp 1679581782
transform 1 0 69408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_724
timestamp 1679581782
transform 1 0 70080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_731
timestamp 1679581782
transform 1 0 70752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_738
timestamp 1679581782
transform 1 0 71424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_745
timestamp 1679581782
transform 1 0 72096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_752
timestamp 1679581782
transform 1 0 72768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_759
timestamp 1679581782
transform 1 0 73440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_766
timestamp 1679581782
transform 1 0 74112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_773
timestamp 1679581782
transform 1 0 74784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_780
timestamp 1679581782
transform 1 0 75456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_787
timestamp 1679581782
transform 1 0 76128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_794
timestamp 1679581782
transform 1 0 76800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_801
timestamp 1679581782
transform 1 0 77472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_808
timestamp 1679581782
transform 1 0 78144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_815
timestamp 1679581782
transform 1 0 78816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_822
timestamp 1679581782
transform 1 0 79488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_829
timestamp 1679581782
transform 1 0 80160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_836
timestamp 1679581782
transform 1 0 80832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_843
timestamp 1679581782
transform 1 0 81504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_850
timestamp 1679581782
transform 1 0 82176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_857
timestamp 1679581782
transform 1 0 82848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_864
timestamp 1679581782
transform 1 0 83520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_871
timestamp 1679581782
transform 1 0 84192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_878
timestamp 1679581782
transform 1 0 84864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_885
timestamp 1679581782
transform 1 0 85536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_892
timestamp 1679581782
transform 1 0 86208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_899
timestamp 1679581782
transform 1 0 86880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_906
timestamp 1679581782
transform 1 0 87552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_913
timestamp 1679581782
transform 1 0 88224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_920
timestamp 1679581782
transform 1 0 88896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_927
timestamp 1679581782
transform 1 0 89568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_934
timestamp 1679581782
transform 1 0 90240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_941
timestamp 1679581782
transform 1 0 90912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_948
timestamp 1679581782
transform 1 0 91584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_955
timestamp 1679581782
transform 1 0 92256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_962
timestamp 1679581782
transform 1 0 92928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_969
timestamp 1679581782
transform 1 0 93600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_976
timestamp 1679581782
transform 1 0 94272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_983
timestamp 1679581782
transform 1 0 94944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_990
timestamp 1679581782
transform 1 0 95616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_997
timestamp 1679581782
transform 1 0 96288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1004
timestamp 1679581782
transform 1 0 96960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1011
timestamp 1679581782
transform 1 0 97632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1018
timestamp 1679581782
transform 1 0 98304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_1025
timestamp 1679577901
transform 1 0 98976 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_7
timestamp 1679577901
transform 1 0 1248 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_34
timestamp 1677579658
transform 1 0 3840 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_58
timestamp 1677579658
transform 1 0 6144 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_105
timestamp 1677580104
transform 1 0 10656 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_107
timestamp 1677579658
transform 1 0 10848 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_218
timestamp 1679581782
transform 1 0 21504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_225
timestamp 1679581782
transform 1 0 22176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_232
timestamp 1679577901
transform 1 0 22848 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_294
timestamp 1677580104
transform 1 0 28800 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_344
timestamp 1677579658
transform 1 0 33600 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_358
timestamp 1679581782
transform 1 0 34944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_365
timestamp 1679577901
transform 1 0 35616 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_455
timestamp 1677580104
transform 1 0 44256 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_457
timestamp 1677579658
transform 1 0 44448 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_471
timestamp 1679581782
transform 1 0 45792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_478
timestamp 1679577901
transform 1 0 46464 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_482
timestamp 1677579658
transform 1 0 46848 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_496
timestamp 1679581782
transform 1 0 48192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_503
timestamp 1679581782
transform 1 0 48864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_510
timestamp 1679581782
transform 1 0 49536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_517
timestamp 1679581782
transform 1 0 50208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_524
timestamp 1679581782
transform 1 0 50880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_531
timestamp 1679581782
transform 1 0 51552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_538
timestamp 1679581782
transform 1 0 52224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_545
timestamp 1679581782
transform 1 0 52896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_552
timestamp 1679581782
transform 1 0 53568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_559
timestamp 1679581782
transform 1 0 54240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_566
timestamp 1679581782
transform 1 0 54912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_573
timestamp 1679581782
transform 1 0 55584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_580
timestamp 1679581782
transform 1 0 56256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_587
timestamp 1679581782
transform 1 0 56928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_594
timestamp 1679581782
transform 1 0 57600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_601
timestamp 1679581782
transform 1 0 58272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_608
timestamp 1679581782
transform 1 0 58944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_615
timestamp 1679581782
transform 1 0 59616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_622
timestamp 1679581782
transform 1 0 60288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_629
timestamp 1679581782
transform 1 0 60960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_636
timestamp 1679581782
transform 1 0 61632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_643
timestamp 1679581782
transform 1 0 62304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_650
timestamp 1679581782
transform 1 0 62976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_657
timestamp 1679581782
transform 1 0 63648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_664
timestamp 1679581782
transform 1 0 64320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_671
timestamp 1679581782
transform 1 0 64992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_678
timestamp 1679581782
transform 1 0 65664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_685
timestamp 1679581782
transform 1 0 66336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_692
timestamp 1679581782
transform 1 0 67008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_699
timestamp 1679581782
transform 1 0 67680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_706
timestamp 1679581782
transform 1 0 68352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_713
timestamp 1679581782
transform 1 0 69024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_720
timestamp 1679581782
transform 1 0 69696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_727
timestamp 1679581782
transform 1 0 70368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_734
timestamp 1679581782
transform 1 0 71040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_741
timestamp 1679581782
transform 1 0 71712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_748
timestamp 1679581782
transform 1 0 72384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_755
timestamp 1679581782
transform 1 0 73056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_762
timestamp 1679581782
transform 1 0 73728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_769
timestamp 1679581782
transform 1 0 74400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_776
timestamp 1679581782
transform 1 0 75072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_783
timestamp 1679581782
transform 1 0 75744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_790
timestamp 1679581782
transform 1 0 76416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_797
timestamp 1679581782
transform 1 0 77088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_804
timestamp 1679581782
transform 1 0 77760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_811
timestamp 1679581782
transform 1 0 78432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_818
timestamp 1679581782
transform 1 0 79104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_825
timestamp 1679581782
transform 1 0 79776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_832
timestamp 1679581782
transform 1 0 80448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_839
timestamp 1679581782
transform 1 0 81120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_846
timestamp 1679581782
transform 1 0 81792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_853
timestamp 1679581782
transform 1 0 82464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_860
timestamp 1679581782
transform 1 0 83136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_867
timestamp 1679581782
transform 1 0 83808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_874
timestamp 1679581782
transform 1 0 84480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_881
timestamp 1679581782
transform 1 0 85152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_888
timestamp 1679581782
transform 1 0 85824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_895
timestamp 1679581782
transform 1 0 86496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_902
timestamp 1679581782
transform 1 0 87168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_909
timestamp 1679581782
transform 1 0 87840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_916
timestamp 1679581782
transform 1 0 88512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_923
timestamp 1679581782
transform 1 0 89184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_930
timestamp 1679581782
transform 1 0 89856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_937
timestamp 1679581782
transform 1 0 90528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_944
timestamp 1679581782
transform 1 0 91200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_951
timestamp 1679581782
transform 1 0 91872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_958
timestamp 1679581782
transform 1 0 92544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_965
timestamp 1679581782
transform 1 0 93216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_972
timestamp 1679581782
transform 1 0 93888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_979
timestamp 1679581782
transform 1 0 94560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_986
timestamp 1679581782
transform 1 0 95232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_993
timestamp 1679581782
transform 1 0 95904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1000
timestamp 1679581782
transform 1 0 96576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1007
timestamp 1679581782
transform 1 0 97248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1014
timestamp 1679581782
transform 1 0 97920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1021
timestamp 1679581782
transform 1 0 98592 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_1028
timestamp 1677579658
transform 1 0 99264 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_58
timestamp 1677579658
transform 1 0 6144 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_64
timestamp 1677579658
transform 1 0 6720 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_43_78
timestamp 1679577901
transform 1 0 8064 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_4  FILLER_43_96
timestamp 1679577901
transform 1 0 9792 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_100
timestamp 1677580104
transform 1 0 10176 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_168
timestamp 1679577901
transform 1 0 16704 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_172
timestamp 1677580104
transform 1 0 17088 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_184
timestamp 1677580104
transform 1 0 18240 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_186
timestamp 1677579658
transform 1 0 18432 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_208
timestamp 1677580104
transform 1 0 20544 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_223
timestamp 1679581782
transform 1 0 21984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_230
timestamp 1679581782
transform 1 0 22656 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_237
timestamp 1677579658
transform 1 0 23328 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_251
timestamp 1677580104
transform 1 0 24672 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_253
timestamp 1677579658
transform 1 0 24864 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_258
timestamp 1677579658
transform 1 0 25344 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_269
timestamp 1677580104
transform 1 0 26400 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_271
timestamp 1677579658
transform 1 0 26592 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_343
timestamp 1677579658
transform 1 0 33504 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_358
timestamp 1679581782
transform 1 0 34944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_365
timestamp 1679581782
transform 1 0 35616 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_386
timestamp 1677580104
transform 1 0 37632 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_388
timestamp 1677579658
transform 1 0 37824 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_420
timestamp 1677580104
transform 1 0 40896 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_474
timestamp 1679581782
transform 1 0 46080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_481
timestamp 1679581782
transform 1 0 46752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_488
timestamp 1679581782
transform 1 0 47424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_495
timestamp 1679581782
transform 1 0 48096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_502
timestamp 1679581782
transform 1 0 48768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_509
timestamp 1679581782
transform 1 0 49440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_516
timestamp 1679581782
transform 1 0 50112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_523
timestamp 1679581782
transform 1 0 50784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_530
timestamp 1679581782
transform 1 0 51456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_537
timestamp 1679581782
transform 1 0 52128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_544
timestamp 1679581782
transform 1 0 52800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_551
timestamp 1679581782
transform 1 0 53472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_558
timestamp 1679581782
transform 1 0 54144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_565
timestamp 1679581782
transform 1 0 54816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_572
timestamp 1679581782
transform 1 0 55488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_579
timestamp 1679581782
transform 1 0 56160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_586
timestamp 1679581782
transform 1 0 56832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_593
timestamp 1679581782
transform 1 0 57504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_600
timestamp 1679581782
transform 1 0 58176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_607
timestamp 1679581782
transform 1 0 58848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_614
timestamp 1679581782
transform 1 0 59520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_621
timestamp 1679581782
transform 1 0 60192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_628
timestamp 1679581782
transform 1 0 60864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_635
timestamp 1679581782
transform 1 0 61536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_642
timestamp 1679581782
transform 1 0 62208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_649
timestamp 1679581782
transform 1 0 62880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_656
timestamp 1679581782
transform 1 0 63552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_663
timestamp 1679581782
transform 1 0 64224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_670
timestamp 1679581782
transform 1 0 64896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_677
timestamp 1679581782
transform 1 0 65568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_684
timestamp 1679581782
transform 1 0 66240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_691
timestamp 1679581782
transform 1 0 66912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_698
timestamp 1679581782
transform 1 0 67584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_705
timestamp 1679581782
transform 1 0 68256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_712
timestamp 1679581782
transform 1 0 68928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_719
timestamp 1679581782
transform 1 0 69600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_726
timestamp 1679581782
transform 1 0 70272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_733
timestamp 1679581782
transform 1 0 70944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_740
timestamp 1679581782
transform 1 0 71616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_747
timestamp 1679581782
transform 1 0 72288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_754
timestamp 1679581782
transform 1 0 72960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_761
timestamp 1679581782
transform 1 0 73632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_768
timestamp 1679581782
transform 1 0 74304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_775
timestamp 1679581782
transform 1 0 74976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_782
timestamp 1679581782
transform 1 0 75648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_789
timestamp 1679581782
transform 1 0 76320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_796
timestamp 1679581782
transform 1 0 76992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_803
timestamp 1679581782
transform 1 0 77664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_810
timestamp 1679581782
transform 1 0 78336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_817
timestamp 1679581782
transform 1 0 79008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_824
timestamp 1679581782
transform 1 0 79680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_831
timestamp 1679581782
transform 1 0 80352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_838
timestamp 1679581782
transform 1 0 81024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_845
timestamp 1679581782
transform 1 0 81696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_852
timestamp 1679581782
transform 1 0 82368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_859
timestamp 1679581782
transform 1 0 83040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_866
timestamp 1679581782
transform 1 0 83712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_873
timestamp 1679581782
transform 1 0 84384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_880
timestamp 1679581782
transform 1 0 85056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_887
timestamp 1679581782
transform 1 0 85728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_894
timestamp 1679581782
transform 1 0 86400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_901
timestamp 1679581782
transform 1 0 87072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_908
timestamp 1679581782
transform 1 0 87744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_915
timestamp 1679581782
transform 1 0 88416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_922
timestamp 1679581782
transform 1 0 89088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_929
timestamp 1679581782
transform 1 0 89760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_936
timestamp 1679581782
transform 1 0 90432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_943
timestamp 1679581782
transform 1 0 91104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_950
timestamp 1679581782
transform 1 0 91776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_957
timestamp 1679581782
transform 1 0 92448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_964
timestamp 1679581782
transform 1 0 93120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_971
timestamp 1679581782
transform 1 0 93792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_978
timestamp 1679581782
transform 1 0 94464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_985
timestamp 1679581782
transform 1 0 95136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_992
timestamp 1679581782
transform 1 0 95808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_999
timestamp 1679581782
transform 1 0 96480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1006
timestamp 1679581782
transform 1 0 97152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1013
timestamp 1679581782
transform 1 0 97824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1020
timestamp 1679581782
transform 1 0 98496 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_1027
timestamp 1677580104
transform 1 0 99168 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_14
timestamp 1679577901
transform 1 0 1920 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_18
timestamp 1677580104
transform 1 0 2304 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_24
timestamp 1679581782
transform 1 0 2880 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_127
timestamp 1677579658
transform 1 0 12768 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_156
timestamp 1677579658
transform 1 0 15552 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_198
timestamp 1679581782
transform 1 0 19584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_205
timestamp 1679581782
transform 1 0 20256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_212
timestamp 1679577901
transform 1 0 20928 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_243
timestamp 1677579658
transform 1 0 23904 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_256
timestamp 1677580104
transform 1 0 25152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_276
timestamp 1677580104
transform 1 0 27072 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_302
timestamp 1677580104
transform 1 0 29568 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_322
timestamp 1677579658
transform 1 0 31488 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_395
timestamp 1677580104
transform 1 0 38496 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_397
timestamp 1677579658
transform 1 0 38688 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_444
timestamp 1677580104
transform 1 0 43200 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_459
timestamp 1679581782
transform 1 0 44640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_466
timestamp 1679581782
transform 1 0 45312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_473
timestamp 1679581782
transform 1 0 45984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_480
timestamp 1679581782
transform 1 0 46656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_487
timestamp 1679581782
transform 1 0 47328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_494
timestamp 1679581782
transform 1 0 48000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_501
timestamp 1679581782
transform 1 0 48672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_508
timestamp 1679581782
transform 1 0 49344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_515
timestamp 1679581782
transform 1 0 50016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_522
timestamp 1679581782
transform 1 0 50688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_529
timestamp 1679581782
transform 1 0 51360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_536
timestamp 1679581782
transform 1 0 52032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_543
timestamp 1679581782
transform 1 0 52704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_550
timestamp 1679581782
transform 1 0 53376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_557
timestamp 1679581782
transform 1 0 54048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_564
timestamp 1679581782
transform 1 0 54720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_571
timestamp 1679581782
transform 1 0 55392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_578
timestamp 1679581782
transform 1 0 56064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_585
timestamp 1679581782
transform 1 0 56736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_592
timestamp 1679581782
transform 1 0 57408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_599
timestamp 1679581782
transform 1 0 58080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_606
timestamp 1679581782
transform 1 0 58752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_613
timestamp 1679581782
transform 1 0 59424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_620
timestamp 1679581782
transform 1 0 60096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_627
timestamp 1679581782
transform 1 0 60768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_634
timestamp 1679581782
transform 1 0 61440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_641
timestamp 1679581782
transform 1 0 62112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_648
timestamp 1679581782
transform 1 0 62784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_655
timestamp 1679581782
transform 1 0 63456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_662
timestamp 1679581782
transform 1 0 64128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_669
timestamp 1679581782
transform 1 0 64800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_676
timestamp 1679581782
transform 1 0 65472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_683
timestamp 1679581782
transform 1 0 66144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_690
timestamp 1679581782
transform 1 0 66816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_697
timestamp 1679581782
transform 1 0 67488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_704
timestamp 1679581782
transform 1 0 68160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_711
timestamp 1679581782
transform 1 0 68832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_718
timestamp 1679581782
transform 1 0 69504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_725
timestamp 1679581782
transform 1 0 70176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_732
timestamp 1679581782
transform 1 0 70848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_739
timestamp 1679581782
transform 1 0 71520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_746
timestamp 1679581782
transform 1 0 72192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_753
timestamp 1679581782
transform 1 0 72864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_760
timestamp 1679581782
transform 1 0 73536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_767
timestamp 1679581782
transform 1 0 74208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_774
timestamp 1679581782
transform 1 0 74880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_781
timestamp 1679581782
transform 1 0 75552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_788
timestamp 1679581782
transform 1 0 76224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_795
timestamp 1679581782
transform 1 0 76896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_802
timestamp 1679581782
transform 1 0 77568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_809
timestamp 1679581782
transform 1 0 78240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_816
timestamp 1679581782
transform 1 0 78912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_823
timestamp 1679581782
transform 1 0 79584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_830
timestamp 1679581782
transform 1 0 80256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_837
timestamp 1679581782
transform 1 0 80928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_844
timestamp 1679581782
transform 1 0 81600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_851
timestamp 1679581782
transform 1 0 82272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_858
timestamp 1679581782
transform 1 0 82944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_865
timestamp 1679581782
transform 1 0 83616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_872
timestamp 1679581782
transform 1 0 84288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_879
timestamp 1679581782
transform 1 0 84960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_886
timestamp 1679581782
transform 1 0 85632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_893
timestamp 1679581782
transform 1 0 86304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_900
timestamp 1679581782
transform 1 0 86976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_907
timestamp 1679581782
transform 1 0 87648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_914
timestamp 1679581782
transform 1 0 88320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_921
timestamp 1679581782
transform 1 0 88992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_928
timestamp 1679581782
transform 1 0 89664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_935
timestamp 1679581782
transform 1 0 90336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_942
timestamp 1679581782
transform 1 0 91008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_949
timestamp 1679581782
transform 1 0 91680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_956
timestamp 1679581782
transform 1 0 92352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_963
timestamp 1679581782
transform 1 0 93024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_970
timestamp 1679581782
transform 1 0 93696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_977
timestamp 1679581782
transform 1 0 94368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_984
timestamp 1679581782
transform 1 0 95040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_991
timestamp 1679581782
transform 1 0 95712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_998
timestamp 1679581782
transform 1 0 96384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1005
timestamp 1679581782
transform 1 0 97056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1012
timestamp 1679581782
transform 1 0 97728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1019
timestamp 1679581782
transform 1 0 98400 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_1026
timestamp 1677580104
transform 1 0 99072 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_1028
timestamp 1677579658
transform 1 0 99264 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_35
timestamp 1679577901
transform 1 0 3936 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_39
timestamp 1677579658
transform 1 0 4320 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_44
timestamp 1679577901
transform 1 0 4800 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_48
timestamp 1677579658
transform 1 0 5184 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_72
timestamp 1677579658
transform 1 0 7488 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_82
timestamp 1677580104
transform 1 0 8448 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_84
timestamp 1677579658
transform 1 0 8640 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_179
timestamp 1679577901
transform 1 0 17760 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_183
timestamp 1677579658
transform 1 0 18144 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_187
timestamp 1677580104
transform 1 0 18528 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_216
timestamp 1677580104
transform 1 0 21312 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_231
timestamp 1679577901
transform 1 0 22752 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_235
timestamp 1677580104
transform 1 0 23136 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_286
timestamp 1677580104
transform 1 0 28032 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_300
timestamp 1677579658
transform 1 0 29376 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_398
timestamp 1677580104
transform 1 0 38784 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_408
timestamp 1677580104
transform 1 0 39744 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_410
timestamp 1677579658
transform 1 0 39936 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_447
timestamp 1677580104
transform 1 0 43488 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_458
timestamp 1679581782
transform 1 0 44544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_465
timestamp 1679581782
transform 1 0 45216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_472
timestamp 1679581782
transform 1 0 45888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_479
timestamp 1679581782
transform 1 0 46560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_486
timestamp 1679581782
transform 1 0 47232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_493
timestamp 1679581782
transform 1 0 47904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_500
timestamp 1679581782
transform 1 0 48576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_507
timestamp 1679581782
transform 1 0 49248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_514
timestamp 1679581782
transform 1 0 49920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_521
timestamp 1679581782
transform 1 0 50592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_528
timestamp 1679581782
transform 1 0 51264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_535
timestamp 1679581782
transform 1 0 51936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_542
timestamp 1679581782
transform 1 0 52608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_549
timestamp 1679581782
transform 1 0 53280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_556
timestamp 1679581782
transform 1 0 53952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_563
timestamp 1679581782
transform 1 0 54624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_570
timestamp 1679581782
transform 1 0 55296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_577
timestamp 1679581782
transform 1 0 55968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_584
timestamp 1679581782
transform 1 0 56640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_591
timestamp 1679581782
transform 1 0 57312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_598
timestamp 1679581782
transform 1 0 57984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_605
timestamp 1679581782
transform 1 0 58656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_612
timestamp 1679581782
transform 1 0 59328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_619
timestamp 1679581782
transform 1 0 60000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_626
timestamp 1679581782
transform 1 0 60672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_633
timestamp 1679581782
transform 1 0 61344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_640
timestamp 1679581782
transform 1 0 62016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_647
timestamp 1679581782
transform 1 0 62688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_654
timestamp 1679581782
transform 1 0 63360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_661
timestamp 1679581782
transform 1 0 64032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_668
timestamp 1679581782
transform 1 0 64704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_675
timestamp 1679581782
transform 1 0 65376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_682
timestamp 1679581782
transform 1 0 66048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_689
timestamp 1679581782
transform 1 0 66720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_696
timestamp 1679581782
transform 1 0 67392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_703
timestamp 1679581782
transform 1 0 68064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_710
timestamp 1679581782
transform 1 0 68736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_717
timestamp 1679581782
transform 1 0 69408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_724
timestamp 1679581782
transform 1 0 70080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_731
timestamp 1679581782
transform 1 0 70752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_738
timestamp 1679581782
transform 1 0 71424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_745
timestamp 1679581782
transform 1 0 72096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_752
timestamp 1679581782
transform 1 0 72768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_759
timestamp 1679581782
transform 1 0 73440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_766
timestamp 1679581782
transform 1 0 74112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_773
timestamp 1679581782
transform 1 0 74784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_780
timestamp 1679581782
transform 1 0 75456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_787
timestamp 1679581782
transform 1 0 76128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_794
timestamp 1679581782
transform 1 0 76800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_801
timestamp 1679581782
transform 1 0 77472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_808
timestamp 1679581782
transform 1 0 78144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_815
timestamp 1679581782
transform 1 0 78816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_822
timestamp 1679581782
transform 1 0 79488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_829
timestamp 1679581782
transform 1 0 80160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_836
timestamp 1679581782
transform 1 0 80832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_843
timestamp 1679581782
transform 1 0 81504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_850
timestamp 1679581782
transform 1 0 82176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_857
timestamp 1679581782
transform 1 0 82848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_864
timestamp 1679581782
transform 1 0 83520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_871
timestamp 1679581782
transform 1 0 84192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_878
timestamp 1679581782
transform 1 0 84864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_885
timestamp 1679581782
transform 1 0 85536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_892
timestamp 1679581782
transform 1 0 86208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_899
timestamp 1679581782
transform 1 0 86880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_906
timestamp 1679581782
transform 1 0 87552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_913
timestamp 1679581782
transform 1 0 88224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_920
timestamp 1679581782
transform 1 0 88896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_927
timestamp 1679581782
transform 1 0 89568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_934
timestamp 1679581782
transform 1 0 90240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_941
timestamp 1679581782
transform 1 0 90912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_948
timestamp 1679581782
transform 1 0 91584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_955
timestamp 1679581782
transform 1 0 92256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_962
timestamp 1679581782
transform 1 0 92928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_969
timestamp 1679581782
transform 1 0 93600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_976
timestamp 1679581782
transform 1 0 94272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_983
timestamp 1679581782
transform 1 0 94944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_990
timestamp 1679581782
transform 1 0 95616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_997
timestamp 1679581782
transform 1 0 96288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1004
timestamp 1679581782
transform 1 0 96960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1011
timestamp 1679581782
transform 1 0 97632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1018
timestamp 1679581782
transform 1 0 98304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_1025
timestamp 1679577901
transform 1 0 98976 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_91
timestamp 1677579658
transform 1 0 9312 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_119
timestamp 1679577901
transform 1 0 12000 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_180
timestamp 1679581782
transform 1 0 17856 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_187
timestamp 1677580104
transform 1 0 18528 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_189
timestamp 1677579658
transform 1 0 18720 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_210
timestamp 1677580104
transform 1 0 20736 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_212
timestamp 1677579658
transform 1 0 20928 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_222
timestamp 1679581782
transform 1 0 21888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_229
timestamp 1679581782
transform 1 0 22560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_236
timestamp 1679577901
transform 1 0 23232 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_240
timestamp 1677580104
transform 1 0 23616 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_246
timestamp 1677580104
transform 1 0 24192 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_362
timestamp 1677579658
transform 1 0 35328 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679581782
transform 1 0 74496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679581782
transform 1 0 76512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679581782
transform 1 0 77184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679581782
transform 1 0 77856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679581782
transform 1 0 78528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679581782
transform 1 0 79200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679581782
transform 1 0 79872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679581782
transform 1 0 80544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_840
timestamp 1679581782
transform 1 0 81216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_847
timestamp 1679581782
transform 1 0 81888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_854
timestamp 1679581782
transform 1 0 82560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_861
timestamp 1679581782
transform 1 0 83232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_868
timestamp 1679581782
transform 1 0 83904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_875
timestamp 1679581782
transform 1 0 84576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_882
timestamp 1679581782
transform 1 0 85248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_889
timestamp 1679581782
transform 1 0 85920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_896
timestamp 1679581782
transform 1 0 86592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_903
timestamp 1679581782
transform 1 0 87264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_910
timestamp 1679581782
transform 1 0 87936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_917
timestamp 1679581782
transform 1 0 88608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_924
timestamp 1679581782
transform 1 0 89280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_931
timestamp 1679581782
transform 1 0 89952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_938
timestamp 1679581782
transform 1 0 90624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_945
timestamp 1679581782
transform 1 0 91296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_952
timestamp 1679581782
transform 1 0 91968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_959
timestamp 1679581782
transform 1 0 92640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_966
timestamp 1679581782
transform 1 0 93312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_973
timestamp 1679581782
transform 1 0 93984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_980
timestamp 1679581782
transform 1 0 94656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_987
timestamp 1679581782
transform 1 0 95328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_994
timestamp 1679581782
transform 1 0 96000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1001
timestamp 1679581782
transform 1 0 96672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1008
timestamp 1679581782
transform 1 0 97344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1015
timestamp 1679581782
transform 1 0 98016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1022
timestamp 1679581782
transform 1 0 98688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_91
timestamp 1679577901
transform 1 0 9312 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_95
timestamp 1677580104
transform 1 0 9696 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_101
timestamp 1679581782
transform 1 0 10272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_108
timestamp 1679581782
transform 1 0 10944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_115
timestamp 1679581782
transform 1 0 11616 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_122
timestamp 1677580104
transform 1 0 12288 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_142
timestamp 1679581782
transform 1 0 14208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_149
timestamp 1679577901
transform 1 0 14880 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_153
timestamp 1677579658
transform 1 0 15264 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_167
timestamp 1679581782
transform 1 0 16608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_174
timestamp 1679581782
transform 1 0 17280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_181
timestamp 1679581782
transform 1 0 17952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_188
timestamp 1679581782
transform 1 0 18624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_195
timestamp 1679581782
transform 1 0 19296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_202
timestamp 1679581782
transform 1 0 19968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_209
timestamp 1679581782
transform 1 0 20640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_216
timestamp 1679581782
transform 1 0 21312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_223
timestamp 1679581782
transform 1 0 21984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_230
timestamp 1679581782
transform 1 0 22656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_237
timestamp 1679581782
transform 1 0 23328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_244
timestamp 1679581782
transform 1 0 24000 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_251
timestamp 1677580104
transform 1 0 24672 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_257
timestamp 1677580104
transform 1 0 25248 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_259
timestamp 1677579658
transform 1 0 25440 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_270
timestamp 1679577901
transform 1 0 26496 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_274
timestamp 1677579658
transform 1 0 26880 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_284
timestamp 1677579658
transform 1 0 27840 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_294
timestamp 1677579658
transform 1 0 28800 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_298
timestamp 1677580104
transform 1 0 29184 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_313
timestamp 1677579658
transform 1 0 30624 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_332
timestamp 1677579658
transform 1 0 32448 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_346
timestamp 1679581782
transform 1 0 33792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_353
timestamp 1679581782
transform 1 0 34464 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_360
timestamp 1677580104
transform 1 0 35136 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_375
timestamp 1679581782
transform 1 0 36576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_382
timestamp 1679581782
transform 1 0 37248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_389
timestamp 1679581782
transform 1 0 37920 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_396
timestamp 1677580104
transform 1 0 38592 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_398
timestamp 1677579658
transform 1 0 38784 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_412
timestamp 1677580104
transform 1 0 40128 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_423
timestamp 1679581782
transform 1 0 41184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_430
timestamp 1679581782
transform 1 0 41856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_437
timestamp 1679581782
transform 1 0 42528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_444
timestamp 1679581782
transform 1 0 43200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_451
timestamp 1679581782
transform 1 0 43872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_458
timestamp 1679581782
transform 1 0 44544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_465
timestamp 1679581782
transform 1 0 45216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_472
timestamp 1679581782
transform 1 0 45888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_479
timestamp 1679581782
transform 1 0 46560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_486
timestamp 1679581782
transform 1 0 47232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_493
timestamp 1679581782
transform 1 0 47904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_500
timestamp 1679581782
transform 1 0 48576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_507
timestamp 1679581782
transform 1 0 49248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_514
timestamp 1679581782
transform 1 0 49920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_521
timestamp 1679581782
transform 1 0 50592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_528
timestamp 1679581782
transform 1 0 51264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_535
timestamp 1679581782
transform 1 0 51936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_542
timestamp 1679581782
transform 1 0 52608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_549
timestamp 1679581782
transform 1 0 53280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_556
timestamp 1679581782
transform 1 0 53952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_563
timestamp 1679581782
transform 1 0 54624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_570
timestamp 1679581782
transform 1 0 55296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_577
timestamp 1679581782
transform 1 0 55968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_584
timestamp 1679581782
transform 1 0 56640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_591
timestamp 1679581782
transform 1 0 57312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_598
timestamp 1679581782
transform 1 0 57984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_605
timestamp 1679581782
transform 1 0 58656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_612
timestamp 1679581782
transform 1 0 59328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_619
timestamp 1679581782
transform 1 0 60000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_626
timestamp 1679581782
transform 1 0 60672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_633
timestamp 1679581782
transform 1 0 61344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_640
timestamp 1679581782
transform 1 0 62016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_647
timestamp 1679581782
transform 1 0 62688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_654
timestamp 1679581782
transform 1 0 63360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_661
timestamp 1679581782
transform 1 0 64032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_668
timestamp 1679581782
transform 1 0 64704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_675
timestamp 1679581782
transform 1 0 65376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_682
timestamp 1679581782
transform 1 0 66048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_689
timestamp 1679581782
transform 1 0 66720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_696
timestamp 1679581782
transform 1 0 67392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_703
timestamp 1679581782
transform 1 0 68064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_710
timestamp 1679581782
transform 1 0 68736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_717
timestamp 1679581782
transform 1 0 69408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_724
timestamp 1679581782
transform 1 0 70080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_731
timestamp 1679581782
transform 1 0 70752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_738
timestamp 1679581782
transform 1 0 71424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_745
timestamp 1679581782
transform 1 0 72096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_752
timestamp 1679581782
transform 1 0 72768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_759
timestamp 1679581782
transform 1 0 73440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_766
timestamp 1679581782
transform 1 0 74112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_773
timestamp 1679581782
transform 1 0 74784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_780
timestamp 1679581782
transform 1 0 75456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_787
timestamp 1679581782
transform 1 0 76128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_794
timestamp 1679581782
transform 1 0 76800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_801
timestamp 1679581782
transform 1 0 77472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_808
timestamp 1679581782
transform 1 0 78144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_815
timestamp 1679581782
transform 1 0 78816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_822
timestamp 1679581782
transform 1 0 79488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_829
timestamp 1679581782
transform 1 0 80160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_836
timestamp 1679581782
transform 1 0 80832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_843
timestamp 1679581782
transform 1 0 81504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_850
timestamp 1679581782
transform 1 0 82176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_857
timestamp 1679581782
transform 1 0 82848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_864
timestamp 1679581782
transform 1 0 83520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_871
timestamp 1679581782
transform 1 0 84192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_878
timestamp 1679581782
transform 1 0 84864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_885
timestamp 1679581782
transform 1 0 85536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_892
timestamp 1679581782
transform 1 0 86208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_899
timestamp 1679581782
transform 1 0 86880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_906
timestamp 1679581782
transform 1 0 87552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_913
timestamp 1679581782
transform 1 0 88224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_920
timestamp 1679581782
transform 1 0 88896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_927
timestamp 1679581782
transform 1 0 89568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_934
timestamp 1679581782
transform 1 0 90240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_941
timestamp 1679581782
transform 1 0 90912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_948
timestamp 1679581782
transform 1 0 91584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_955
timestamp 1679581782
transform 1 0 92256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_962
timestamp 1679581782
transform 1 0 92928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_969
timestamp 1679581782
transform 1 0 93600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_976
timestamp 1679581782
transform 1 0 94272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_983
timestamp 1679581782
transform 1 0 94944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_990
timestamp 1679581782
transform 1 0 95616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_997
timestamp 1679581782
transform 1 0 96288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1004
timestamp 1679581782
transform 1 0 96960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1011
timestamp 1679581782
transform 1 0 97632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1018
timestamp 1679581782
transform 1 0 98304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_1025
timestamp 1679577901
transform 1 0 98976 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_318
timestamp 1679577901
transform 1 0 31104 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_322
timestamp 1677580104
transform 1 0 31488 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_333
timestamp 1679581782
transform 1 0 32544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_340
timestamp 1679581782
transform 1 0 33216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_347
timestamp 1679581782
transform 1 0 33888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_354
timestamp 1679581782
transform 1 0 34560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_361
timestamp 1679581782
transform 1 0 35232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_368
timestamp 1679581782
transform 1 0 35904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_375
timestamp 1679581782
transform 1 0 36576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_382
timestamp 1679581782
transform 1 0 37248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_389
timestamp 1679581782
transform 1 0 37920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_396
timestamp 1679581782
transform 1 0 38592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_403
timestamp 1679581782
transform 1 0 39264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_410
timestamp 1679581782
transform 1 0 39936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_417
timestamp 1679581782
transform 1 0 40608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_424
timestamp 1679581782
transform 1 0 41280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_431
timestamp 1679581782
transform 1 0 41952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_438
timestamp 1679581782
transform 1 0 42624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_445
timestamp 1679581782
transform 1 0 43296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_452
timestamp 1679581782
transform 1 0 43968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_459
timestamp 1679581782
transform 1 0 44640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_466
timestamp 1679581782
transform 1 0 45312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_473
timestamp 1679581782
transform 1 0 45984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_480
timestamp 1679581782
transform 1 0 46656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_487
timestamp 1679581782
transform 1 0 47328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_494
timestamp 1679581782
transform 1 0 48000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_501
timestamp 1679581782
transform 1 0 48672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_508
timestamp 1679581782
transform 1 0 49344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_515
timestamp 1679581782
transform 1 0 50016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_522
timestamp 1679581782
transform 1 0 50688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_529
timestamp 1679581782
transform 1 0 51360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_536
timestamp 1679581782
transform 1 0 52032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_543
timestamp 1679581782
transform 1 0 52704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_550
timestamp 1679581782
transform 1 0 53376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_557
timestamp 1679581782
transform 1 0 54048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_564
timestamp 1679581782
transform 1 0 54720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_571
timestamp 1679581782
transform 1 0 55392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_578
timestamp 1679581782
transform 1 0 56064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_585
timestamp 1679581782
transform 1 0 56736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_592
timestamp 1679581782
transform 1 0 57408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_599
timestamp 1679581782
transform 1 0 58080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_606
timestamp 1679581782
transform 1 0 58752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_613
timestamp 1679581782
transform 1 0 59424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_620
timestamp 1679581782
transform 1 0 60096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_627
timestamp 1679581782
transform 1 0 60768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_634
timestamp 1679581782
transform 1 0 61440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_641
timestamp 1679581782
transform 1 0 62112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_648
timestamp 1679581782
transform 1 0 62784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_655
timestamp 1679581782
transform 1 0 63456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_662
timestamp 1679581782
transform 1 0 64128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_669
timestamp 1679581782
transform 1 0 64800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_676
timestamp 1679581782
transform 1 0 65472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_683
timestamp 1679581782
transform 1 0 66144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_690
timestamp 1679581782
transform 1 0 66816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_697
timestamp 1679581782
transform 1 0 67488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_704
timestamp 1679581782
transform 1 0 68160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_711
timestamp 1679581782
transform 1 0 68832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_718
timestamp 1679581782
transform 1 0 69504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_725
timestamp 1679581782
transform 1 0 70176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_732
timestamp 1679581782
transform 1 0 70848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_739
timestamp 1679581782
transform 1 0 71520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_746
timestamp 1679581782
transform 1 0 72192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_753
timestamp 1679581782
transform 1 0 72864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_760
timestamp 1679581782
transform 1 0 73536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_767
timestamp 1679581782
transform 1 0 74208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_774
timestamp 1679581782
transform 1 0 74880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_781
timestamp 1679581782
transform 1 0 75552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_788
timestamp 1679581782
transform 1 0 76224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_795
timestamp 1679581782
transform 1 0 76896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_802
timestamp 1679581782
transform 1 0 77568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_809
timestamp 1679581782
transform 1 0 78240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_816
timestamp 1679581782
transform 1 0 78912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_823
timestamp 1679581782
transform 1 0 79584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_830
timestamp 1679581782
transform 1 0 80256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_837
timestamp 1679581782
transform 1 0 80928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_844
timestamp 1679581782
transform 1 0 81600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_851
timestamp 1679581782
transform 1 0 82272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_858
timestamp 1679581782
transform 1 0 82944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_865
timestamp 1679581782
transform 1 0 83616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_872
timestamp 1679581782
transform 1 0 84288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_879
timestamp 1679581782
transform 1 0 84960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_886
timestamp 1679581782
transform 1 0 85632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_893
timestamp 1679581782
transform 1 0 86304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_900
timestamp 1679581782
transform 1 0 86976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_907
timestamp 1679581782
transform 1 0 87648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_914
timestamp 1679581782
transform 1 0 88320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_921
timestamp 1679581782
transform 1 0 88992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_928
timestamp 1679581782
transform 1 0 89664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_935
timestamp 1679581782
transform 1 0 90336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_942
timestamp 1679581782
transform 1 0 91008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_949
timestamp 1679581782
transform 1 0 91680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_956
timestamp 1679581782
transform 1 0 92352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_963
timestamp 1679581782
transform 1 0 93024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_970
timestamp 1679581782
transform 1 0 93696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_977
timestamp 1679581782
transform 1 0 94368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_984
timestamp 1679581782
transform 1 0 95040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_991
timestamp 1679581782
transform 1 0 95712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_998
timestamp 1679581782
transform 1 0 96384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1005
timestamp 1679581782
transform 1 0 97056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1012
timestamp 1679581782
transform 1 0 97728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1019
timestamp 1679581782
transform 1 0 98400 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_1026
timestamp 1677580104
transform 1 0 99072 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_1028
timestamp 1677579658
transform 1 0 99264 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 36192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 36864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 37536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 38208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 38880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 39552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 40224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 40896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 41568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 42240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 42912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 43584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 44256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 44928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 45600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 46272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 46944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 47616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 48288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 48960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 49632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 50304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 50976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 51648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 52320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 52992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 53664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 54336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 55008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 55680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 56352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 57696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 58368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 59040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 59712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 60384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 61056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 61728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 62400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 63072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 63744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 64416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 65088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 65760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 66432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 67104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 67776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 68448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 69120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 69792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 70464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 73824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 74496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 75168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 75840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 76512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 77184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 77856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 78528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 79200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 79872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 80544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_840
timestamp 1679581782
transform 1 0 81216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_847
timestamp 1679581782
transform 1 0 81888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_854
timestamp 1679581782
transform 1 0 82560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_861
timestamp 1679581782
transform 1 0 83232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_868
timestamp 1679581782
transform 1 0 83904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_875
timestamp 1679581782
transform 1 0 84576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_882
timestamp 1679581782
transform 1 0 85248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_889
timestamp 1679581782
transform 1 0 85920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_896
timestamp 1679581782
transform 1 0 86592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_903
timestamp 1679581782
transform 1 0 87264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_910
timestamp 1679581782
transform 1 0 87936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_917
timestamp 1679581782
transform 1 0 88608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_924
timestamp 1679581782
transform 1 0 89280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_931
timestamp 1679581782
transform 1 0 89952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_938
timestamp 1679581782
transform 1 0 90624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_945
timestamp 1679581782
transform 1 0 91296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_952
timestamp 1679581782
transform 1 0 91968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_959
timestamp 1679581782
transform 1 0 92640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_966
timestamp 1679581782
transform 1 0 93312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_973
timestamp 1679581782
transform 1 0 93984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_980
timestamp 1679581782
transform 1 0 94656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_987
timestamp 1679581782
transform 1 0 95328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_994
timestamp 1679581782
transform 1 0 96000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1001
timestamp 1679581782
transform 1 0 96672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1008
timestamp 1679581782
transform 1 0 97344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1015
timestamp 1679581782
transform 1 0 98016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1022
timestamp 1679581782
transform 1 0 98688 0 -1 38556
box -48 -56 720 834
use sg13g2_tielo  heichips25_ppwm_3
timestamp 1680000637
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_4
timestamp 1680000637
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_5
timestamp 1680000637
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_6
timestamp 1680000637
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_7
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_8
timestamp 1680000637
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_9
timestamp 1680000637
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_10
timestamp 1680000637
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_11
timestamp 1680000637
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_12
timestamp 1680000637
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_13
timestamp 1680000637
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_14
timestamp 1680000637
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_15
timestamp 1680000637
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_16
timestamp 1680000637
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_17
timestamp 1680000637
transform -1 0 1344 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_18
timestamp 1680000637
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_19
timestamp 1680000637
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_20
timestamp 1680000637
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_21
timestamp 1680000637
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_22
timestamp 1680000637
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_23
timestamp 1680000637
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_24
timestamp 1680000637
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_25
timestamp 1680000637
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677672058
transform -1 0 38976 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677672058
transform 1 0 36480 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677672058
transform -1 0 9408 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677672058
transform -1 0 8448 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677672058
transform -1 0 28416 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677672058
transform -1 0 28320 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677672058
transform -1 0 38880 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677672058
transform -1 0 37728 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677672058
transform -1 0 12384 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677672058
transform -1 0 13248 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677672058
transform -1 0 5664 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677672058
transform -1 0 6144 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677672058
transform 1 0 12864 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677672058
transform -1 0 14592 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677672058
transform 1 0 4224 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677672058
transform -1 0 5952 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677672058
transform -1 0 19104 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677672058
transform -1 0 19680 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677672058
transform 1 0 26304 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677672058
transform 1 0 28704 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677672058
transform 1 0 7776 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677672058
transform -1 0 10752 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677672058
transform -1 0 14400 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677672058
transform -1 0 12768 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677672058
transform -1 0 17664 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677672058
transform 1 0 15552 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677672058
transform -1 0 13920 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677672058
transform -1 0 5280 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677672058
transform 1 0 6432 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677672058
transform 1 0 23232 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677672058
transform -1 0 25152 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677672058
transform 1 0 19200 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677672058
transform -1 0 20736 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677672058
transform -1 0 22080 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677672058
transform -1 0 19968 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677672058
transform 1 0 5184 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677672058
transform -1 0 5184 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677672058
transform 1 0 33216 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677672058
transform -1 0 33984 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677672058
transform -1 0 40896 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677672058
transform -1 0 40128 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677672058
transform -1 0 8832 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677672058
transform -1 0 9792 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677672058
transform -1 0 48960 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677672058
transform 1 0 47808 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1677672058
transform 1 0 7200 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1677672058
transform -1 0 7104 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1677672058
transform 1 0 16224 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1677672058
transform 1 0 16992 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1677672058
transform -1 0 27840 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1677672058
transform -1 0 28032 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1677672058
transform 1 0 12480 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1677672058
transform 1 0 10464 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1677672058
transform 1 0 23232 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1677672058
transform 1 0 19680 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1677672058
transform -1 0 8448 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1677672058
transform 1 0 35136 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1677672058
transform 1 0 35904 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1677672058
transform 1 0 27936 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1677672058
transform -1 0 30624 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1677672058
transform -1 0 19872 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1677672058
transform 1 0 19584 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1677672058
transform -1 0 41184 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1677672058
transform -1 0 38976 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1677672058
transform -1 0 9408 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1677672058
transform 1 0 6432 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1677672058
transform -1 0 18528 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1677672058
transform 1 0 16704 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1677672058
transform 1 0 11616 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1677672058
transform -1 0 11904 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1677672058
transform 1 0 22368 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1677672058
transform 1 0 19872 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1677672058
transform -1 0 13056 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1677672058
transform -1 0 13824 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1677672058
transform -1 0 25536 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1677672058
transform -1 0 24288 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold77
timestamp 1677672058
transform -1 0 23520 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold78
timestamp 1677672058
transform 1 0 20352 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold79
timestamp 1677672058
transform -1 0 16896 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold80
timestamp 1677672058
transform 1 0 13920 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold81
timestamp 1677672058
transform -1 0 14784 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold82
timestamp 1677672058
transform -1 0 16032 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold83
timestamp 1677672058
transform 1 0 27936 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold84
timestamp 1677672058
transform -1 0 29472 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold85
timestamp 1677672058
transform -1 0 21888 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold86
timestamp 1677672058
transform -1 0 22368 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold87
timestamp 1677672058
transform -1 0 22080 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold88
timestamp 1677672058
transform 1 0 20352 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold89
timestamp 1677672058
transform -1 0 4320 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold90
timestamp 1677672058
transform -1 0 4896 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold91
timestamp 1677672058
transform -1 0 3840 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold92
timestamp 1677672058
transform -1 0 32736 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold93
timestamp 1677672058
transform -1 0 29856 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold94
timestamp 1677672058
transform 1 0 25632 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold95
timestamp 1677672058
transform -1 0 25344 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold96
timestamp 1677672058
transform -1 0 6720 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold97
timestamp 1677672058
transform 1 0 8064 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold98
timestamp 1677672058
transform -1 0 20736 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold99
timestamp 1677672058
transform 1 0 19872 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold100
timestamp 1677672058
transform 1 0 39168 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold101
timestamp 1677672058
transform 1 0 41088 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold102
timestamp 1677672058
transform -1 0 43104 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold103
timestamp 1677672058
transform -1 0 43008 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold104
timestamp 1677672058
transform 1 0 43008 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold105
timestamp 1677672058
transform -1 0 45792 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold106
timestamp 1677672058
transform 1 0 9504 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold107
timestamp 1677672058
transform 1 0 17088 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold108
timestamp 1677672058
transform -1 0 15936 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold109
timestamp 1677672058
transform 1 0 36768 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold110
timestamp 1677672058
transform -1 0 16032 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold111
timestamp 1677672058
transform -1 0 12192 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold112
timestamp 1677672058
transform 1 0 30720 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold113
timestamp 1677672058
transform 1 0 32544 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold114
timestamp 1677672058
transform -1 0 36192 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold115
timestamp 1677672058
transform -1 0 22368 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold116
timestamp 1677672058
transform -1 0 36768 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold117
timestamp 1677672058
transform -1 0 34368 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold118
timestamp 1677672058
transform -1 0 31008 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold119
timestamp 1677672058
transform -1 0 29280 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold120
timestamp 1677672058
transform 1 0 28320 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold121
timestamp 1677672058
transform 1 0 45600 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold122
timestamp 1677672058
transform 1 0 49056 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold123
timestamp 1677672058
transform 1 0 31488 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold124
timestamp 1677672058
transform -1 0 15552 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold125
timestamp 1677672058
transform -1 0 16224 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold126
timestamp 1677672058
transform -1 0 41856 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold127
timestamp 1677672058
transform 1 0 42144 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold128
timestamp 1677672058
transform -1 0 11616 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold129
timestamp 1677672058
transform 1 0 5664 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold130
timestamp 1677672058
transform 1 0 16032 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold131
timestamp 1677672058
transform 1 0 17088 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold132
timestamp 1677672058
transform -1 0 44736 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold133
timestamp 1677672058
transform 1 0 43584 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold134
timestamp 1677672058
transform -1 0 11424 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold135
timestamp 1677672058
transform 1 0 11616 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold136
timestamp 1677672058
transform -1 0 44928 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold137
timestamp 1677672058
transform -1 0 40224 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold138
timestamp 1677672058
transform -1 0 48384 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold139
timestamp 1677672058
transform 1 0 45024 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold140
timestamp 1677672058
transform -1 0 47808 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold141
timestamp 1677672058
transform -1 0 48192 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold142
timestamp 1677672058
transform -1 0 13920 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold143
timestamp 1677672058
transform -1 0 9984 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold144
timestamp 1677672058
transform -1 0 16416 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold145
timestamp 1677672058
transform -1 0 15168 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold146
timestamp 1677672058
transform 1 0 11328 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold147
timestamp 1677672058
transform 1 0 12672 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold148
timestamp 1677672058
transform -1 0 41280 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold149
timestamp 1677672058
transform -1 0 39168 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold150
timestamp 1677672058
transform -1 0 6144 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold151
timestamp 1677672058
transform -1 0 35232 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold152
timestamp 1677672058
transform 1 0 31008 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold153
timestamp 1677672058
transform -1 0 9216 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold154
timestamp 1677672058
transform -1 0 7776 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold155
timestamp 1677672058
transform -1 0 18816 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold156
timestamp 1677672058
transform -1 0 10848 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold157
timestamp 1677672058
transform -1 0 47328 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold158
timestamp 1677672058
transform -1 0 49152 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold159
timestamp 1677672058
transform 1 0 48864 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold160
timestamp 1677672058
transform 1 0 38880 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold161
timestamp 1677672058
transform 1 0 39168 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold162
timestamp 1677672058
transform -1 0 47904 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold163
timestamp 1677672058
transform -1 0 47328 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold164
timestamp 1677672058
transform -1 0 40416 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold165
timestamp 1677672058
transform 1 0 12192 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold166
timestamp 1677672058
transform -1 0 17760 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold167
timestamp 1677672058
transform 1 0 10944 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold168
timestamp 1677672058
transform -1 0 45120 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold169
timestamp 1677672058
transform -1 0 43488 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold170
timestamp 1677672058
transform -1 0 11328 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold171
timestamp 1677672058
transform -1 0 10080 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold172
timestamp 1677672058
transform -1 0 32544 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold173
timestamp 1677672058
transform -1 0 4608 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold174
timestamp 1677672058
transform 1 0 30528 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold175
timestamp 1677672058
transform -1 0 34560 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold176
timestamp 1677672058
transform -1 0 44544 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold177
timestamp 1677672058
transform 1 0 40704 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold178
timestamp 1677672058
transform 1 0 15360 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold179
timestamp 1677672058
transform -1 0 15552 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold180
timestamp 1677672058
transform -1 0 50784 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold181
timestamp 1677672058
transform -1 0 4800 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold182
timestamp 1677672058
transform -1 0 16224 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold183
timestamp 1677672058
transform -1 0 8352 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold184
timestamp 1677672058
transform 1 0 44736 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold185
timestamp 1677672058
transform -1 0 32640 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold186
timestamp 1677672058
transform 1 0 30144 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold187
timestamp 1677672058
transform 1 0 36000 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold188
timestamp 1677672058
transform -1 0 37248 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold189
timestamp 1677672058
transform -1 0 37920 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold190
timestamp 1677672058
transform 1 0 42048 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold191
timestamp 1677672058
transform -1 0 14112 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold192
timestamp 1677672058
transform 1 0 5088 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold193
timestamp 1677672058
transform -1 0 4608 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold194
timestamp 1677672058
transform 1 0 37440 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold195
timestamp 1677672058
transform 1 0 18336 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold196
timestamp 1677672058
transform -1 0 37056 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold197
timestamp 1677672058
transform -1 0 32256 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold198
timestamp 1677672058
transform -1 0 33600 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold199
timestamp 1677672058
transform -1 0 28704 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold200
timestamp 1677672058
transform 1 0 4224 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold201
timestamp 1677672058
transform 1 0 5280 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold202
timestamp 1677672058
transform 1 0 26304 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold203
timestamp 1677672058
transform -1 0 31008 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold204
timestamp 1677672058
transform 1 0 28416 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold205
timestamp 1677672058
transform -1 0 44640 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold206
timestamp 1677672058
transform -1 0 7872 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold207
timestamp 1677672058
transform -1 0 6528 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold208
timestamp 1677672058
transform -1 0 6432 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold209
timestamp 1677672058
transform -1 0 38208 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold210
timestamp 1677672058
transform -1 0 36480 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold211
timestamp 1677672058
transform 1 0 36192 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold212
timestamp 1677672058
transform 1 0 33888 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold213
timestamp 1677672058
transform -1 0 34560 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold214
timestamp 1677672058
transform 1 0 34560 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold215
timestamp 1677672058
transform -1 0 9504 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold216
timestamp 1677672058
transform -1 0 25152 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold217
timestamp 1677672058
transform -1 0 50880 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold218
timestamp 1677672058
transform 1 0 48384 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold219
timestamp 1677672058
transform 1 0 9408 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold220
timestamp 1677672058
transform -1 0 9024 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold221
timestamp 1677672058
transform -1 0 38880 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold222
timestamp 1677672058
transform 1 0 36192 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold223
timestamp 1677672058
transform -1 0 7008 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold224
timestamp 1677672058
transform -1 0 7584 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold225
timestamp 1677672058
transform -1 0 18816 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold226
timestamp 1677672058
transform 1 0 16032 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold227
timestamp 1677672058
transform 1 0 38880 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold228
timestamp 1677672058
transform 1 0 39456 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold229
timestamp 1677672058
transform -1 0 22272 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold230
timestamp 1677672058
transform -1 0 20544 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold231
timestamp 1677672058
transform -1 0 8928 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold232
timestamp 1677672058
transform -1 0 38976 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold233
timestamp 1677672058
transform -1 0 32448 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold234
timestamp 1677672058
transform -1 0 38112 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold235
timestamp 1677672058
transform 1 0 35712 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold236
timestamp 1677672058
transform -1 0 8256 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold237
timestamp 1677672058
transform -1 0 12000 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold238
timestamp 1677672058
transform -1 0 10656 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold239
timestamp 1677672058
transform -1 0 7776 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold240
timestamp 1677672058
transform 1 0 4800 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold241
timestamp 1677672058
transform -1 0 6720 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold242
timestamp 1677672058
transform -1 0 48288 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold243
timestamp 1677672058
transform -1 0 31872 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold244
timestamp 1677672058
transform -1 0 30144 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold245
timestamp 1677672058
transform 1 0 29184 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold246
timestamp 1677672058
transform -1 0 51744 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold247
timestamp 1677672058
transform 1 0 48864 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold248
timestamp 1677672058
transform -1 0 49920 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold249
timestamp 1677672058
transform -1 0 16416 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold250
timestamp 1677672058
transform 1 0 9504 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold251
timestamp 1677672058
transform 1 0 15072 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold252
timestamp 1677672058
transform -1 0 13536 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold253
timestamp 1677672058
transform 1 0 14304 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold254
timestamp 1677672058
transform -1 0 5568 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold255
timestamp 1677672058
transform -1 0 5664 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold256
timestamp 1677672058
transform -1 0 4704 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold257
timestamp 1677672058
transform -1 0 43872 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold258
timestamp 1677672058
transform -1 0 35808 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold259
timestamp 1677672058
transform 1 0 4704 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold260
timestamp 1677672058
transform 1 0 6048 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold261
timestamp 1677672058
transform 1 0 15168 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold262
timestamp 1677672058
transform -1 0 13056 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold263
timestamp 1677672058
transform -1 0 30720 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold264
timestamp 1677672058
transform 1 0 20928 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold265
timestamp 1677672058
transform -1 0 20352 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold266
timestamp 1677672058
transform 1 0 24192 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold267
timestamp 1677672058
transform 1 0 25536 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold268
timestamp 1677672058
transform 1 0 6336 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold269
timestamp 1677672058
transform -1 0 6912 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold270
timestamp 1677672058
transform -1 0 5664 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold271
timestamp 1677672058
transform -1 0 36192 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold272
timestamp 1677672058
transform -1 0 37344 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold273
timestamp 1677672058
transform 1 0 34752 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold274
timestamp 1677672058
transform -1 0 11712 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold275
timestamp 1677672058
transform 1 0 4416 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold276
timestamp 1677672058
transform 1 0 3840 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold277
timestamp 1677672058
transform -1 0 9792 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold278
timestamp 1677672058
transform 1 0 6144 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold279
timestamp 1677672058
transform -1 0 7008 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold280
timestamp 1677672058
transform -1 0 5472 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold281
timestamp 1677672058
transform -1 0 4800 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold282
timestamp 1677672058
transform -1 0 9504 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold283
timestamp 1677672058
transform -1 0 12192 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold284
timestamp 1677672058
transform -1 0 31488 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold285
timestamp 1677672058
transform 1 0 28320 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold286
timestamp 1677672058
transform 1 0 28224 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold287
timestamp 1677672058
transform 1 0 6048 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold288
timestamp 1677672058
transform 1 0 25344 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold289
timestamp 1677672058
transform -1 0 27360 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold290
timestamp 1677672058
transform 1 0 27360 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold291
timestamp 1677672058
transform 1 0 21312 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold292
timestamp 1677672058
transform -1 0 23424 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold293
timestamp 1677672058
transform -1 0 34464 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold294
timestamp 1677672058
transform 1 0 33216 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold295
timestamp 1677672058
transform -1 0 27072 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold296
timestamp 1677672058
transform -1 0 41088 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold297
timestamp 1677672058
transform 1 0 37824 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold298
timestamp 1677672058
transform 1 0 24000 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold299
timestamp 1677672058
transform -1 0 21600 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold300
timestamp 1677672058
transform -1 0 10464 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold301
timestamp 1677672058
transform 1 0 7776 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold302
timestamp 1677672058
transform -1 0 9504 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold303
timestamp 1677672058
transform -1 0 37152 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold304
timestamp 1677672058
transform 1 0 34176 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold305
timestamp 1677672058
transform -1 0 40800 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold306
timestamp 1677672058
transform 1 0 18240 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold307
timestamp 1677672058
transform -1 0 20160 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold308
timestamp 1677672058
transform -1 0 16416 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold309
timestamp 1677672058
transform -1 0 15360 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold310
timestamp 1677672058
transform -1 0 40224 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold311
timestamp 1677672058
transform 1 0 22272 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold312
timestamp 1677672058
transform -1 0 20832 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold313
timestamp 1677672058
transform 1 0 20640 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold314
timestamp 1677672058
transform -1 0 27360 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold315
timestamp 1677672058
transform 1 0 29760 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold316
timestamp 1677672058
transform 1 0 29088 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold317
timestamp 1677672058
transform -1 0 8832 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold318
timestamp 1677672058
transform -1 0 21600 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold319
timestamp 1677672058
transform 1 0 23232 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold320
timestamp 1677672058
transform -1 0 40608 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold321
timestamp 1677672058
transform 1 0 24288 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold322
timestamp 1677672058
transform 1 0 21504 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold323
timestamp 1677672058
transform -1 0 21792 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold324
timestamp 1677672058
transform 1 0 16992 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold325
timestamp 1677672058
transform 1 0 12768 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold326
timestamp 1677672058
transform -1 0 12768 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold327
timestamp 1677672058
transform 1 0 21600 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold328
timestamp 1677672058
transform 1 0 22464 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold329
timestamp 1677672058
transform 1 0 32832 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold330
timestamp 1677672058
transform -1 0 12960 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold331
timestamp 1677672058
transform -1 0 13824 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold332
timestamp 1677672058
transform 1 0 20160 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold333
timestamp 1677672058
transform -1 0 26208 0 1 12852
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_ex__415_
timestamp 1676382947
transform -1 0 32448 0 1 11340
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__416_
timestamp 1676382929
transform 1 0 32352 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__417_
timestamp 1676382929
transform 1 0 32544 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__418_
timestamp 1676382929
transform -1 0 30240 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__419_
timestamp 1676382929
transform -1 0 25440 0 1 8316
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__420_
timestamp 1676382947
transform 1 0 25152 0 -1 9828
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__421_
timestamp 1676382929
transform -1 0 29184 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__422_
timestamp 1676382929
transform 1 0 28320 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__423_
timestamp 1676382947
transform -1 0 28032 0 -1 9828
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__424_
timestamp 1676382929
transform 1 0 22368 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__425_
timestamp 1676382929
transform 1 0 23616 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__426_
timestamp 1676382929
transform 1 0 30720 0 1 23436
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__427_
timestamp 1676382947
transform 1 0 28608 0 1 18900
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__428_
timestamp 1676382929
transform -1 0 30720 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__429_
timestamp 1676382929
transform -1 0 20736 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__430_
timestamp 1676382929
transform -1 0 33216 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__431_
timestamp 1676382929
transform -1 0 31776 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__432_
timestamp 1676382929
transform 1 0 28704 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__433_
timestamp 1676382929
transform -1 0 28512 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__434_
timestamp 1676382929
transform 1 0 25728 0 1 11340
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__435_
timestamp 1676382947
transform 1 0 25920 0 -1 5292
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__436_
timestamp 1676382929
transform -1 0 25920 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__437_
timestamp 1676382947
transform -1 0 29568 0 -1 2268
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__438_
timestamp 1676382929
transform -1 0 31392 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__439_
timestamp 1676382929
transform 1 0 31008 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__440_
timestamp 1676382929
transform -1 0 22368 0 -1 6804
box -48 -56 336 834
use sg13g2_nand2_1  u_ppwm_u_ex__441_
timestamp 1676557249
transform 1 0 26400 0 1 23436
box -48 -56 432 834
use sg13g2_nand3_1  u_ppwm_u_ex__442_
timestamp 1683988354
transform 1 0 22560 0 1 23436
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__443_
timestamp 1685201930
transform -1 0 23616 0 1 23436
box -48 -56 624 834
use sg13g2_inv_1  u_ppwm_u_ex__444_
timestamp 1676382929
transform 1 0 20640 0 1 18900
box -48 -56 336 834
use sg13g2_nor2b_1  u_ppwm_u_ex__445_
timestamp 1685181386
transform -1 0 26976 0 1 14364
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__446_
timestamp 1676567195
transform -1 0 26304 0 -1 14364
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__447_
timestamp 1684236171
transform 1 0 24672 0 -1 20412
box -48 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__448_
timestamp 1676643125
transform -1 0 26880 0 -1 18900
box -48 -56 624 834
use sg13g2_nand2b_1  u_ppwm_u_ex__449_
timestamp 1676567195
transform -1 0 22368 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__450_
timestamp 1685175443
transform -1 0 19680 0 -1 20412
box -48 -56 538 834
use sg13g2_a21o_1  u_ppwm_u_ex__451_
timestamp 1677175127
transform 1 0 20544 0 -1 20412
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_ex__452_
timestamp 1685175443
transform -1 0 21216 0 -1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__453_
timestamp 1685175443
transform 1 0 22272 0 1 20412
box -48 -56 538 834
use sg13g2_and2_1  u_ppwm_u_ex__454_
timestamp 1676901763
transform -1 0 21888 0 -1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__455_
timestamp 1685173987
transform 1 0 20736 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2b_1  u_ppwm_u_ex__456_
timestamp 1685181386
transform 1 0 17568 0 1 18900
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__457_
timestamp 1676567195
transform -1 0 27744 0 -1 21924
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__458_
timestamp 1683988354
transform -1 0 27456 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__459_
timestamp 1685175443
transform 1 0 28512 0 1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__460_
timestamp 1685175443
transform 1 0 31008 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__461_
timestamp 1683973020
transform 1 0 31488 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__462_
timestamp 1676557249
transform 1 0 25152 0 -1 21924
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__463_
timestamp 1676557249
transform 1 0 27552 0 1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__464_
timestamp 1685175443
transform -1 0 29376 0 1 23436
box -48 -56 538 834
use sg13g2_xnor2_1  u_ppwm_u_ex__465_
timestamp 1677516600
transform 1 0 27456 0 -1 23436
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__466_
timestamp 1676557249
transform -1 0 29760 0 -1 23436
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__467_
timestamp 1676901763
transform 1 0 27936 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__468_
timestamp 1676627187
transform 1 0 28896 0 -1 23436
box -48 -56 432 834
use sg13g2_or3_1  u_ppwm_u_ex__469_
timestamp 1677141922
transform 1 0 28224 0 -1 23436
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_ex__470_
timestamp 1685175443
transform 1 0 28416 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__471_
timestamp 1683973020
transform 1 0 29376 0 1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__472_
timestamp 1676567195
transform -1 0 25920 0 1 23436
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__473_
timestamp 1676567195
transform 1 0 24864 0 1 21924
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__474_
timestamp 1683988354
transform 1 0 25920 0 1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__475_
timestamp 1683973020
transform -1 0 27552 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__476_
timestamp 1676557249
transform 1 0 23040 0 1 21924
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__477_
timestamp 1677516600
transform 1 0 24096 0 -1 23436
box -48 -56 816 834
use sg13g2_or2_1  u_ppwm_u_ex__478_
timestamp 1684236171
transform -1 0 24864 0 1 21924
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__479_
timestamp 1683973020
transform -1 0 26496 0 -1 23436
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__480_
timestamp 1685173987
transform 1 0 24960 0 -1 23436
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__481_
timestamp 1685175443
transform 1 0 25536 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__482_
timestamp 1676627187
transform 1 0 25632 0 -1 24948
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__483_
timestamp 1677516600
transform -1 0 24768 0 -1 21924
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__484_
timestamp 1683973020
transform -1 0 23904 0 1 21924
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__485_
timestamp 1683988354
transform -1 0 25440 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__486_
timestamp 1676627187
transform -1 0 24960 0 1 23436
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_ex__487_
timestamp 1685181386
transform 1 0 23040 0 -1 23436
box -54 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__488_
timestamp 1676557249
transform -1 0 24000 0 1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__489_
timestamp 1685175443
transform 1 0 23616 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__490_
timestamp 1683973020
transform 1 0 23904 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__491_
timestamp 1685175443
transform -1 0 26976 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__492_
timestamp 1676627187
transform 1 0 25536 0 -1 21924
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__493_
timestamp 1685173987
transform 1 0 32640 0 -1 11340
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__494_
timestamp 1676557249
transform 1 0 31680 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_ex__495_
timestamp 1685181386
transform 1 0 24672 0 -1 8316
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__496_
timestamp 1676567195
transform 1 0 24096 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__497_
timestamp 1676567195
transform -1 0 30336 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__498_
timestamp 1685175443
transform 1 0 28512 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__499_
timestamp 1676567195
transform -1 0 25536 0 1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__500_
timestamp 1683973020
transform -1 0 25056 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__501_
timestamp 1685181386
transform 1 0 28896 0 1 6804
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__502_
timestamp 1685181386
transform 1 0 29376 0 1 6804
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__503_
timestamp 1685197497
transform 1 0 29664 0 -1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__504_
timestamp 1685175443
transform 1 0 30432 0 -1 8316
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__505_
timestamp 1685173987
transform -1 0 32832 0 1 8316
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__506_
timestamp 1676557249
transform 1 0 32544 0 1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__507_
timestamp 1685175443
transform 1 0 32832 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__508_
timestamp 1685175443
transform -1 0 32544 0 1 9828
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__509_
timestamp 1685181386
transform 1 0 32736 0 1 12852
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__510_
timestamp 1676567195
transform -1 0 39360 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__511_
timestamp 1676567195
transform 1 0 34368 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__512_
timestamp 1685181386
transform 1 0 32832 0 1 11340
box -54 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__513_
timestamp 1676627187
transform 1 0 32448 0 1 11340
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_ex__514_
timestamp 1685181386
transform -1 0 34368 0 1 11340
box -54 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__515_
timestamp 1676643125
transform -1 0 33888 0 1 11340
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_ex__516_
timestamp 1683973020
transform 1 0 33216 0 1 12852
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__517_
timestamp 1683988354
transform -1 0 31776 0 1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__518_
timestamp 1683973020
transform 1 0 32160 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__519_
timestamp 1676557249
transform 1 0 30432 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_ex__520_
timestamp 1676627187
transform -1 0 28992 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_ex__521_
timestamp 1685181386
transform 1 0 23136 0 -1 8316
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__522_
timestamp 1676567195
transform 1 0 23328 0 1 8316
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__523_
timestamp 1676567195
transform -1 0 24576 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__524_
timestamp 1685175443
transform 1 0 24000 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__525_
timestamp 1676567195
transform -1 0 23328 0 1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__526_
timestamp 1683973020
transform -1 0 24288 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__527_
timestamp 1685173987
transform -1 0 25152 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__528_
timestamp 1685175443
transform 1 0 24480 0 -1 9828
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__529_
timestamp 1676639442
transform -1 0 25056 0 1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__530_
timestamp 1676567195
transform -1 0 29952 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__531_
timestamp 1685175443
transform -1 0 29088 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__532_
timestamp 1676567195
transform 1 0 28992 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__533_
timestamp 1685175443
transform -1 0 28608 0 -1 9828
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__534_
timestamp 1676639442
transform 1 0 28800 0 1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__535_
timestamp 1685181386
transform 1 0 30048 0 1 9828
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__536_
timestamp 1685197497
transform -1 0 29856 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__537_
timestamp 1685175443
transform 1 0 28992 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__538_
timestamp 1676627187
transform -1 0 30912 0 1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__539_
timestamp 1677516600
transform -1 0 29568 0 -1 14364
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__540_
timestamp 1676567195
transform 1 0 26688 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__541_
timestamp 1676627187
transform -1 0 30528 0 1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__542_
timestamp 1677516600
transform 1 0 27936 0 -1 14364
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_ex__543_
timestamp 1685201930
transform 1 0 29568 0 -1 14364
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_ex__544_
timestamp 1676639442
transform 1 0 29664 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__545_
timestamp 1683973020
transform -1 0 29088 0 1 12852
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__546_
timestamp 1676901763
transform 1 0 29952 0 1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__547_
timestamp 1683973020
transform 1 0 29280 0 1 14364
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_ex__548_
timestamp 1676985977
transform -1 0 28512 0 1 18900
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__549_
timestamp 1676567195
transform 1 0 22464 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__550_
timestamp 1685181386
transform 1 0 21120 0 -1 8316
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__551_
timestamp 1685181386
transform 1 0 21984 0 1 8316
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__552_
timestamp 1685197497
transform 1 0 22848 0 1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__553_
timestamp 1676567195
transform -1 0 26112 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__554_
timestamp 1685175443
transform 1 0 25536 0 1 8316
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__555_
timestamp 1685181386
transform 1 0 26016 0 1 8316
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__556_
timestamp 1685181386
transform 1 0 26304 0 -1 8316
box -54 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__557_
timestamp 1677577977
transform -1 0 27552 0 -1 8316
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_ex__558_
timestamp 1676639442
transform 1 0 26496 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__559_
timestamp 1685175443
transform 1 0 26112 0 1 6804
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__560_
timestamp 1676639442
transform -1 0 27456 0 1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__561_
timestamp 1683973020
transform 1 0 27168 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__562_
timestamp 1676627187
transform -1 0 27552 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__563_
timestamp 1676557249
transform -1 0 27168 0 -1 11340
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__564_
timestamp 1685175443
transform 1 0 26112 0 1 9828
box -48 -56 538 834
use sg13g2_a221oi_1  u_ppwm_u_ex__565_
timestamp 1685197497
transform 1 0 26592 0 1 9828
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__566_
timestamp 1676627187
transform -1 0 26784 0 -1 11340
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__567_
timestamp 1685175443
transform -1 0 26400 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__568_
timestamp 1685175443
transform 1 0 26016 0 1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__569_
timestamp 1685173987
transform 1 0 26400 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__570_
timestamp 1685175443
transform 1 0 26976 0 1 11340
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__571_
timestamp 1676627187
transform -1 0 28416 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__572_
timestamp 1683973020
transform 1 0 28128 0 1 12852
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__573_
timestamp 1683988354
transform -1 0 28128 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__574_
timestamp 1685173987
transform 1 0 29856 0 -1 9828
box -48 -56 624 834
use sg13g2_nand2b_1  u_ppwm_u_ex__575_
timestamp 1676567195
transform 1 0 26784 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__576_
timestamp 1685181386
transform 1 0 23616 0 -1 6804
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__577_
timestamp 1685181386
transform 1 0 25152 0 1 6804
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__578_
timestamp 1685197497
transform 1 0 26592 0 1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__579_
timestamp 1676567195
transform -1 0 28896 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__580_
timestamp 1685175443
transform 1 0 27936 0 1 6804
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__581_
timestamp 1685173987
transform 1 0 28992 0 -1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__582_
timestamp 1685175443
transform 1 0 28032 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__583_
timestamp 1676627187
transform 1 0 30432 0 -1 9828
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__584_
timestamp 1685197497
transform 1 0 29280 0 1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__585_
timestamp 1676567195
transform -1 0 30432 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__586_
timestamp 1685175443
transform -1 0 29952 0 -1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__587_
timestamp 1685173987
transform -1 0 29664 0 -1 12852
box -48 -56 624 834
use sg13g2_nand2b_1  u_ppwm_u_ex__588_
timestamp 1676567195
transform -1 0 29088 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__589_
timestamp 1676567195
transform -1 0 30336 0 1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__590_
timestamp 1676567195
transform 1 0 29664 0 1 12852
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_ex__591_
timestamp 1676985977
transform -1 0 30432 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__592_
timestamp 1685175443
transform -1 0 29376 0 1 11340
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__593_
timestamp 1676567195
transform -1 0 29856 0 1 11340
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__594_
timestamp 1685201930
transform -1 0 29664 0 1 12852
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__595_
timestamp 1676627187
transform 1 0 30720 0 1 9828
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_ex__596_
timestamp 1676567195
transform 1 0 23616 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__597_
timestamp 1685181386
transform -1 0 24096 0 1 5292
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__598_
timestamp 1685181386
transform 1 0 23712 0 -1 8316
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__599_
timestamp 1685197497
transform 1 0 24096 0 1 6804
box -48 -56 816 834
use sg13g2_a221oi_1  u_ppwm_u_ex__600_
timestamp 1685197497
transform 1 0 25152 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__601_
timestamp 1676567195
transform 1 0 32832 0 1 8316
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__602_
timestamp 1676567195
transform -1 0 32544 0 -1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__603_
timestamp 1685173987
transform -1 0 31584 0 -1 8316
box -48 -56 624 834
use sg13g2_nand3_1  u_ppwm_u_ex__604_
timestamp 1683988354
transform 1 0 31296 0 1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__605_
timestamp 1685181386
transform -1 0 33024 0 -1 8316
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__606_
timestamp 1683973020
transform -1 0 32256 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__607_
timestamp 1685175443
transform 1 0 31776 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__608_
timestamp 1676557249
transform 1 0 31104 0 1 9828
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__609_
timestamp 1685197497
transform 1 0 31104 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__610_
timestamp 1676567195
transform -1 0 27648 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__611_
timestamp 1685175443
transform 1 0 26496 0 1 11340
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__612_
timestamp 1676557249
transform 1 0 27648 0 -1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__613_
timestamp 1685173987
transform 1 0 25920 0 -1 12852
box -48 -56 624 834
use sg13g2_nand3b_1  u_ppwm_u_ex__614_
timestamp 1676573470
transform 1 0 26496 0 -1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  u_ppwm_u_ex__615_
timestamp 1683973020
transform -1 0 25824 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__616_
timestamp 1685175443
transform -1 0 27456 0 1 12852
box -48 -56 538 834
use sg13g2_and4_1  u_ppwm_u_ex__617_
timestamp 1676985977
transform -1 0 27936 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__618_
timestamp 1685175443
transform -1 0 28320 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__619_
timestamp 1683973020
transform -1 0 28896 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__620_
timestamp 1676557249
transform 1 0 26496 0 -1 20412
box -48 -56 432 834
use sg13g2_nor2_2  u_ppwm_u_ex__621_
timestamp 1683979924
transform 1 0 25920 0 -1 20412
box -48 -56 624 834
use sg13g2_nor3_2  u_ppwm_u_ex__622_
timestamp 1685180723
transform 1 0 25440 0 1 18900
box -48 -56 912 834
use sg13g2_nand2b_2  u_ppwm_u_ex__623_
timestamp 1685211885
transform -1 0 26496 0 1 14364
box -48 -56 816 834
use sg13g2_nand2b_2  u_ppwm_u_ex__624_
timestamp 1685211885
transform -1 0 25920 0 -1 20412
box -48 -56 816 834
use sg13g2_nor2_2  u_ppwm_u_ex__625_
timestamp 1683979924
transform 1 0 31488 0 -1 18900
box -48 -56 624 834
use sg13g2_nand2b_2  u_ppwm_u_ex__626_
timestamp 1685211885
transform 1 0 31392 0 -1 20412
box -48 -56 816 834
use sg13g2_and2_1  u_ppwm_u_ex__627_
timestamp 1676901763
transform -1 0 19968 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__628_
timestamp 1685175443
transform 1 0 19968 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__629_
timestamp 1685175443
transform 1 0 20640 0 1 15876
box -48 -56 538 834
use sg13g2_nor3_2  u_ppwm_u_ex__630_
timestamp 1685180723
transform 1 0 31200 0 1 17388
box -48 -56 912 834
use sg13g2_a22oi_1  u_ppwm_u_ex__631_
timestamp 1685173987
transform -1 0 21696 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__632_
timestamp 1685175443
transform 1 0 20640 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__633_
timestamp 1683973020
transform 1 0 20256 0 -1 17388
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__634_
timestamp 1676901763
transform -1 0 19488 0 -1 15876
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__635_
timestamp 1677577977
transform 1 0 18528 0 1 15876
box -48 -56 816 834
use sg13g2_xor2_1  u_ppwm_u_ex__636_
timestamp 1677577977
transform 1 0 19296 0 1 15876
box -48 -56 816 834
use sg13g2_nor3_2  u_ppwm_u_ex__637_
timestamp 1685180723
transform 1 0 31008 0 -1 17388
box -48 -56 912 834
use sg13g2_a22oi_1  u_ppwm_u_ex__638_
timestamp 1685173987
transform 1 0 20064 0 1 15876
box -48 -56 624 834
use sg13g2_a221oi_1  u_ppwm_u_ex__639_
timestamp 1685197497
transform 1 0 19584 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__640_
timestamp 1685175443
transform -1 0 20448 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__641_
timestamp 1683973020
transform 1 0 18720 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__642_
timestamp 1683973020
transform -1 0 19008 0 -1 15876
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__643_
timestamp 1677516600
transform 1 0 19200 0 -1 14364
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__644_
timestamp 1676627187
transform -1 0 22176 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__645_
timestamp 1683973020
transform -1 0 20256 0 1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__646_
timestamp 1685181386
transform 1 0 20256 0 1 14364
box -54 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__647_
timestamp 1676557249
transform -1 0 24384 0 -1 15876
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__648_
timestamp 1685173987
transform -1 0 23232 0 -1 15876
box -48 -56 624 834
use sg13g2_nand3_1  u_ppwm_u_ex__649_
timestamp 1683988354
transform -1 0 22656 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__650_
timestamp 1685175443
transform 1 0 21504 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__651_
timestamp 1683973020
transform 1 0 21792 0 -1 11340
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__652_
timestamp 1677577977
transform 1 0 19968 0 -1 14364
box -48 -56 816 834
use sg13g2_a21o_1  u_ppwm_u_ex__653_
timestamp 1677175127
transform 1 0 21120 0 -1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  u_ppwm_u_ex__654_
timestamp 1683973020
transform -1 0 21408 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__655_
timestamp 1685175443
transform 1 0 21024 0 1 12852
box -48 -56 538 834
use sg13g2_a221oi_1  u_ppwm_u_ex__656_
timestamp 1685197497
transform -1 0 22272 0 1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__657_
timestamp 1685175443
transform 1 0 20544 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__658_
timestamp 1683973020
transform 1 0 21024 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__659_
timestamp 1676567195
transform -1 0 20544 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__660_
timestamp 1685175443
transform 1 0 18720 0 -1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__661_
timestamp 1685175443
transform -1 0 19968 0 1 12852
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__662_
timestamp 1676557249
transform 1 0 15648 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__663_
timestamp 1677516600
transform 1 0 14880 0 1 11340
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__664_
timestamp 1676567195
transform 1 0 16512 0 1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__665_
timestamp 1676567195
transform -1 0 16512 0 1 11340
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__666_
timestamp 1683988354
transform 1 0 16032 0 1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__667_
timestamp 1685197497
transform 1 0 18816 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__668_
timestamp 1685175443
transform 1 0 15648 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__669_
timestamp 1683973020
transform 1 0 16512 0 1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__670_
timestamp 1677516600
transform 1 0 14592 0 -1 11340
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_ex__671_
timestamp 1683988354
transform 1 0 15936 0 1 8316
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_ex__672_
timestamp 1677175127
transform 1 0 15744 0 -1 11340
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__673_
timestamp 1683988354
transform 1 0 16128 0 -1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__674_
timestamp 1685197497
transform -1 0 17568 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__675_
timestamp 1685175443
transform 1 0 16608 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__676_
timestamp 1683973020
transform 1 0 16896 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__677_
timestamp 1676557249
transform -1 0 14688 0 1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__678_
timestamp 1677516600
transform 1 0 13440 0 1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__679_
timestamp 1685175443
transform 1 0 14400 0 1 11340
box -48 -56 538 834
use sg13g2_inv_1  u_ppwm_u_ex__680_
timestamp 1676382929
transform 1 0 16512 0 -1 12852
box -48 -56 336 834
use sg13g2_nor2_1  u_ppwm_u_ex__681_
timestamp 1676627187
transform -1 0 16512 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__682_
timestamp 1683973020
transform 1 0 15648 0 -1 12852
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__683_
timestamp 1684236171
transform -1 0 14592 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__684_
timestamp 1683973020
transform -1 0 15360 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__685_
timestamp 1676557249
transform -1 0 15456 0 -1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__686_
timestamp 1685197497
transform 1 0 17760 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__687_
timestamp 1685175443
transform 1 0 13152 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__688_
timestamp 1683973020
transform 1 0 13632 0 1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__689_
timestamp 1677516600
transform -1 0 14592 0 -1 14364
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_ex__690_
timestamp 1683988354
transform 1 0 12960 0 1 12852
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_ex__691_
timestamp 1677175127
transform -1 0 14880 0 1 12852
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__692_
timestamp 1683988354
transform 1 0 14592 0 -1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__693_
timestamp 1685197497
transform 1 0 17568 0 1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__694_
timestamp 1685175443
transform -1 0 14112 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__695_
timestamp 1683973020
transform 1 0 13632 0 -1 12852
box -48 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__696_
timestamp 1676643125
transform -1 0 15648 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__697_
timestamp 1685175443
transform 1 0 14592 0 -1 12852
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__698_
timestamp 1676557249
transform 1 0 15360 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__699_
timestamp 1683973020
transform -1 0 16416 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__700_
timestamp 1676557249
transform 1 0 17664 0 -1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__701_
timestamp 1677516600
transform 1 0 14688 0 1 14364
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__702_
timestamp 1683973020
transform -1 0 17376 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__703_
timestamp 1685175443
transform 1 0 17184 0 -1 14364
box -48 -56 538 834
use sg13g2_a221oi_1  u_ppwm_u_ex__704_
timestamp 1685197497
transform -1 0 19968 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__705_
timestamp 1685175443
transform 1 0 18240 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__706_
timestamp 1683973020
transform 1 0 19008 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__707_
timestamp 1685175443
transform 1 0 18240 0 1 14364
box -48 -56 538 834
use sg13g2_xnor2_1  u_ppwm_u_ex__708_
timestamp 1677516600
transform 1 0 15456 0 1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__709_
timestamp 1677516600
transform 1 0 16416 0 -1 15876
box -48 -56 816 834
use sg13g2_a221oi_1  u_ppwm_u_ex__710_
timestamp 1685197497
transform 1 0 17472 0 1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__711_
timestamp 1685175443
transform 1 0 15456 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__712_
timestamp 1676627187
transform -1 0 16800 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__713_
timestamp 1676901763
transform 1 0 26400 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_2  u_ppwm_u_ex__714_
timestamp 1685180049
transform -1 0 26304 0 -1 15876
box -48 -56 624 834
use sg13g2_and2_1  u_ppwm_u_ex__715_
timestamp 1676901763
transform -1 0 24000 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__716_
timestamp 1676557249
transform 1 0 24000 0 -1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__717_
timestamp 1685175443
transform -1 0 23808 0 -1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__718_
timestamp 1685175443
transform -1 0 23520 0 -1 18900
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__719_
timestamp 1685173987
transform 1 0 22176 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__720_
timestamp 1685175443
transform -1 0 24000 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__721_
timestamp 1683973020
transform -1 0 23328 0 1 17388
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__722_
timestamp 1676901763
transform -1 0 24960 0 1 15876
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__723_
timestamp 1684236171
transform 1 0 21792 0 1 15876
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__724_
timestamp 1676567195
transform 1 0 22752 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__725_
timestamp 1685175443
transform 1 0 24288 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__726_
timestamp 1683973020
transform -1 0 23808 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__727_
timestamp 1683973020
transform -1 0 25632 0 -1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__728_
timestamp 1685197497
transform 1 0 24288 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__729_
timestamp 1685175443
transform 1 0 23808 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__730_
timestamp 1683973020
transform 1 0 23808 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__731_
timestamp 1683973020
transform -1 0 22752 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__732_
timestamp 1676557249
transform 1 0 27360 0 1 17388
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__733_
timestamp 1677516600
transform 1 0 26880 0 -1 17388
box -48 -56 816 834
use sg13g2_or2_1  u_ppwm_u_ex__734_
timestamp 1684236171
transform -1 0 27840 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__735_
timestamp 1683973020
transform 1 0 26592 0 1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__736_
timestamp 1685173987
transform 1 0 24672 0 -1 15876
box -48 -56 624 834
use sg13g2_nand3_1  u_ppwm_u_ex__737_
timestamp 1683988354
transform 1 0 25248 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__738_
timestamp 1683973020
transform 1 0 26400 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__739_
timestamp 1685175443
transform -1 0 26592 0 1 15876
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__740_
timestamp 1676627187
transform -1 0 26400 0 1 17388
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__741_
timestamp 1677516600
transform 1 0 27072 0 1 15876
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_ex__742_
timestamp 1683988354
transform 1 0 27840 0 1 15876
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_ex__743_
timestamp 1677175127
transform -1 0 28320 0 -1 17388
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__744_
timestamp 1683988354
transform 1 0 28320 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__745_
timestamp 1685197497
transform -1 0 29376 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__746_
timestamp 1685175443
transform -1 0 29472 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__747_
timestamp 1683973020
transform -1 0 29376 0 1 15876
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__748_
timestamp 1684236171
transform 1 0 27744 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__749_
timestamp 1685175443
transform -1 0 30240 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__750_
timestamp 1685175443
transform 1 0 29184 0 -1 15876
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__751_
timestamp 1676557249
transform -1 0 35136 0 -1 15876
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__752_
timestamp 1677516600
transform 1 0 33984 0 -1 15876
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__753_
timestamp 1676567195
transform -1 0 34560 0 1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__754_
timestamp 1676567195
transform -1 0 33216 0 1 14364
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__755_
timestamp 1683988354
transform -1 0 32736 0 1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__756_
timestamp 1685197497
transform 1 0 31488 0 -1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__757_
timestamp 1685175443
transform -1 0 31776 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__758_
timestamp 1683973020
transform -1 0 32256 0 1 14364
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__759_
timestamp 1677516600
transform -1 0 36672 0 1 14364
box -48 -56 816 834
use sg13g2_a21o_1  u_ppwm_u_ex__760_
timestamp 1677175127
transform 1 0 33312 0 -1 15876
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__761_
timestamp 1683988354
transform -1 0 34176 0 1 15876
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__762_
timestamp 1683988354
transform -1 0 33696 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__763_
timestamp 1685197497
transform -1 0 33024 0 -1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__764_
timestamp 1685175443
transform 1 0 31872 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__765_
timestamp 1683973020
transform -1 0 33216 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__766_
timestamp 1676557249
transform 1 0 38592 0 1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__767_
timestamp 1677516600
transform -1 0 38304 0 1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__768_
timestamp 1685175443
transform -1 0 36192 0 -1 15876
box -48 -56 538 834
use sg13g2_inv_1  u_ppwm_u_ex__769_
timestamp 1676382929
transform -1 0 35904 0 1 14364
box -48 -56 336 834
use sg13g2_nor2_1  u_ppwm_u_ex__770_
timestamp 1676627187
transform 1 0 35328 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__771_
timestamp 1683973020
transform -1 0 36672 0 -1 15876
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__772_
timestamp 1684236171
transform 1 0 37344 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__773_
timestamp 1683973020
transform 1 0 37056 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__774_
timestamp 1676557249
transform 1 0 36864 0 1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__775_
timestamp 1685197497
transform -1 0 37728 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__776_
timestamp 1685175443
transform 1 0 37248 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__777_
timestamp 1683973020
transform 1 0 38112 0 -1 17388
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__778_
timestamp 1677516600
transform 1 0 37824 0 -1 15876
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_ex__779_
timestamp 1683988354
transform -1 0 39360 0 1 15876
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_ex__780_
timestamp 1677175127
transform -1 0 38592 0 1 15876
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__781_
timestamp 1683988354
transform -1 0 39072 0 -1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__782_
timestamp 1685197497
transform -1 0 36960 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__783_
timestamp 1685175443
transform -1 0 37344 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__784_
timestamp 1683973020
transform -1 0 37824 0 1 17388
box -48 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__785_
timestamp 1676643125
transform 1 0 36672 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__786_
timestamp 1685175443
transform -1 0 36672 0 1 15876
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__787_
timestamp 1676557249
transform -1 0 36192 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__788_
timestamp 1683973020
transform 1 0 35712 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__789_
timestamp 1676557249
transform 1 0 34848 0 -1 17388
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__790_
timestamp 1677516600
transform -1 0 35808 0 1 18900
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__791_
timestamp 1683973020
transform 1 0 34080 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__792_
timestamp 1685175443
transform -1 0 34176 0 1 18900
box -48 -56 538 834
use sg13g2_a221oi_1  u_ppwm_u_ex__793_
timestamp 1685197497
transform 1 0 34560 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__794_
timestamp 1685175443
transform -1 0 35808 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__795_
timestamp 1683973020
transform -1 0 33984 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__796_
timestamp 1685175443
transform -1 0 35712 0 1 20412
box -48 -56 538 834
use sg13g2_xnor2_1  u_ppwm_u_ex__797_
timestamp 1677516600
transform 1 0 33984 0 -1 18900
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__798_
timestamp 1677516600
transform 1 0 34752 0 -1 18900
box -48 -56 816 834
use sg13g2_a221oi_1  u_ppwm_u_ex__799_
timestamp 1685197497
transform -1 0 36288 0 -1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__800_
timestamp 1685175443
transform -1 0 37632 0 -1 18900
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__801_
timestamp 1676627187
transform 1 0 36480 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__802_
timestamp 1746535128
transform 1 0 31488 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__802__51
timestamp 1680000651
transform -1 0 32352 0 -1 23436
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__803__44
timestamp 1680000651
transform -1 0 30144 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__803_
timestamp 1746535128
transform 1 0 29280 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__804_
timestamp 1746535184
transform 1 0 25056 0 1 24948
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__804__42
timestamp 1680000651
transform -1 0 26496 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__805__40
timestamp 1680000651
transform 1 0 27744 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__805_
timestamp 1746535128
transform 1 0 28128 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__806__38
timestamp 1680000651
transform -1 0 29376 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__806_
timestamp 1746535128
transform 1 0 28512 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__807__36
timestamp 1680000651
transform 1 0 14112 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__807_
timestamp 1746535184
transform -1 0 18048 0 -1 17388
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__808_
timestamp 1746535128
transform 1 0 18912 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__808__34
timestamp 1680000651
transform -1 0 20064 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__809__32
timestamp 1680000651
transform -1 0 21504 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__809_
timestamp 1746535128
transform 1 0 20640 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__810_
timestamp 1746535128
transform 1 0 21696 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__810__30
timestamp 1680000651
transform -1 0 22656 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__811_
timestamp 1746535128
transform 1 0 17856 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__811__28
timestamp 1680000651
transform -1 0 19008 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__812__26
timestamp 1680000651
transform -1 0 18336 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__812_
timestamp 1746535128
transform 1 0 17472 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__813_
timestamp 1746535128
transform 1 0 9984 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__813__49
timestamp 1680000651
transform -1 0 11136 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__814__47
timestamp 1680000651
transform -1 0 10368 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__814_
timestamp 1746535128
transform 1 0 9504 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__815_
timestamp 1746535184
transform 1 0 22368 0 1 12852
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__815__45
timestamp 1680000651
transform -1 0 23232 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__816_
timestamp 1746535184
transform 1 0 12864 0 -1 15876
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__816__41
timestamp 1680000651
transform 1 0 12768 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__817_
timestamp 1746535184
transform 1 0 22080 0 1 18900
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__817__37
timestamp 1680000651
transform -1 0 23808 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__818_
timestamp 1746535184
transform 1 0 17664 0 1 17388
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__818__33
timestamp 1680000651
transform -1 0 18528 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__819__29
timestamp 1680000651
transform 1 0 26976 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__819_
timestamp 1746535184
transform 1 0 27072 0 -1 18900
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__820_
timestamp 1746535184
transform 1 0 29472 0 1 18900
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__820__50
timestamp 1680000651
transform 1 0 28128 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__821__46
timestamp 1680000651
transform 1 0 33216 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__821_
timestamp 1746535184
transform 1 0 33696 0 1 12852
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__822__39
timestamp 1680000651
transform 1 0 39360 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__822_
timestamp 1746535184
transform 1 0 39072 0 1 14364
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__823__31
timestamp 1680000651
transform -1 0 41472 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__823_
timestamp 1746535184
transform 1 0 39840 0 -1 17388
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__824_
timestamp 1746535184
transform 1 0 38688 0 1 17388
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__824__48
timestamp 1680000651
transform -1 0 39456 0 -1 15876
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__825__35
timestamp 1680000651
transform -1 0 35136 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__825_
timestamp 1746535184
transform 1 0 34272 0 -1 20412
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__826__52
timestamp 1680000651
transform -1 0 38208 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__826_
timestamp 1746535184
transform 1 0 37248 0 1 18900
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__827_
timestamp 1746535128
transform 1 0 18816 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__827__53
timestamp 1680000651
transform 1 0 18816 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__828_
timestamp 1746535128
transform 1 0 18048 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__828__27
timestamp 1680000651
transform -1 0 18816 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__829__43
timestamp 1680000651
transform -1 0 21984 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__829_
timestamp 1746535184
transform 1 0 21120 0 -1 21924
box -48 -56 2736 834
use sg13g2_inv_1  u_ppwm_u_global_counter__053_
timestamp 1676382929
transform 1 0 27744 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__054_
timestamp 1676382929
transform 1 0 25056 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__055_
timestamp 1676382929
transform -1 0 33408 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__056_
timestamp 1676382929
transform -1 0 34368 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__057_
timestamp 1676382929
transform 1 0 34272 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__058_
timestamp 1676382929
transform 1 0 35328 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__059_
timestamp 1676382929
transform 1 0 25344 0 1 2268
box -48 -56 336 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__060_
timestamp 1677577977
transform -1 0 21408 0 -1 2268
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__061_
timestamp 1683988354
transform 1 0 23520 0 1 3780
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_global_counter__062_
timestamp 1677175127
transform 1 0 21600 0 -1 5292
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__063_
timestamp 1676901763
transform -1 0 19968 0 1 3780
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__064_
timestamp 1685201930
transform 1 0 26208 0 -1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__065_
timestamp 1677516600
transform -1 0 20640 0 1 2268
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__066_
timestamp 1676627187
transform 1 0 28032 0 1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__067_
timestamp 1677516600
transform -1 0 29088 0 -1 5292
box -48 -56 816 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__068_
timestamp 1677577977
transform 1 0 29376 0 -1 6804
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__069_
timestamp 1685201930
transform -1 0 27744 0 -1 5292
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__070_
timestamp 1676627187
transform 1 0 25920 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__071_
timestamp 1683973020
transform -1 0 29376 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__072_
timestamp 1676627187
transform 1 0 28512 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__073_
timestamp 1677577977
transform 1 0 26784 0 -1 3780
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__074_
timestamp 1685201930
transform -1 0 27360 0 1 5292
box -48 -56 624 834
use sg13g2_nor3_2  u_ppwm_u_global_counter__075_
timestamp 1685180723
transform 1 0 26304 0 1 3780
box -48 -56 912 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__076_
timestamp 1683973020
transform -1 0 28320 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__077_
timestamp 1676627187
transform 1 0 26400 0 -1 3780
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__078_
timestamp 1677577977
transform -1 0 25536 0 -1 3780
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__079_
timestamp 1683988354
transform -1 0 26880 0 1 756
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_global_counter__080_
timestamp 1677175127
transform -1 0 26208 0 -1 3780
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__081_
timestamp 1676901763
transform 1 0 25920 0 1 756
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__082_
timestamp 1685201930
transform -1 0 25920 0 1 3780
box -48 -56 624 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__083_
timestamp 1677516600
transform -1 0 25920 0 1 756
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__084_
timestamp 1685201930
transform 1 0 25632 0 -1 6804
box -48 -56 624 834
use sg13g2_nor3_2  u_ppwm_u_global_counter__085_
timestamp 1685180723
transform -1 0 27168 0 -1 5292
box -48 -56 912 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__086_
timestamp 1685173987
transform 1 0 25056 0 -1 6804
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__087_
timestamp 1683973020
transform -1 0 34368 0 1 5292
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__088_
timestamp 1683988354
transform -1 0 34848 0 1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_global_counter__089_
timestamp 1685181386
transform 1 0 33408 0 1 5292
box -54 -56 528 834
use sg13g2_and3_2  u_ppwm_u_global_counter__090_
timestamp 1683976310
transform -1 0 35040 0 1 8316
box -48 -56 720 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__091_
timestamp 1685173987
transform -1 0 35424 0 1 5292
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__092_
timestamp 1683973020
transform -1 0 33888 0 -1 8316
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__093_
timestamp 1683988354
transform -1 0 34848 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_global_counter__094_
timestamp 1685181386
transform 1 0 33888 0 1 8316
box -54 -56 528 834
use sg13g2_and3_2  u_ppwm_u_global_counter__095_
timestamp 1683976310
transform -1 0 35520 0 -1 9828
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__096_
timestamp 1676901763
transform 1 0 35520 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__097_
timestamp 1683973020
transform -1 0 35712 0 1 8316
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__098_
timestamp 1683988354
transform -1 0 35712 0 1 9828
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__099_
timestamp 1677577977
transform 1 0 35712 0 1 9828
box -48 -56 816 834
use sg13g2_and2_1  u_ppwm_u_global_counter__100_
timestamp 1676901763
transform 1 0 34272 0 1 9828
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__101_
timestamp 1683988354
transform -1 0 35232 0 1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__102_
timestamp 1685173987
transform 1 0 34752 0 1 11340
box -48 -56 624 834
use sg13g2_and4_1  u_ppwm_u_global_counter__103_
timestamp 1676985977
transform 1 0 34560 0 -1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__104_
timestamp 1683973020
transform -1 0 36096 0 -1 12852
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__105_
timestamp 1677577977
transform -1 0 36864 0 -1 12852
box -48 -56 816 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__106_
timestamp 1746535184
transform 1 0 20832 0 1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__107_
timestamp 1746535184
transform 1 0 20832 0 1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__108_
timestamp 1746535184
transform 1 0 20544 0 -1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__109_
timestamp 1746535184
transform 1 0 29088 0 -1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__110_
timestamp 1746535184
transform 1 0 31008 0 -1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__111_
timestamp 1746535184
transform 1 0 30048 0 1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__112_
timestamp 1746535184
transform 1 0 27360 0 1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__113_
timestamp 1746535184
transform 1 0 29280 0 -1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__114_
timestamp 1746535184
transform 1 0 23520 0 -1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__115_
timestamp 1746535184
transform 1 0 26208 0 -1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__116_
timestamp 1746535184
transform -1 0 24480 0 1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__117_
timestamp 1746535184
transform -1 0 25824 0 -1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__118_
timestamp 1746535184
transform -1 0 36288 0 1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__119_
timestamp 1746535184
transform 1 0 35424 0 -1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__120_
timestamp 1746535184
transform 1 0 36480 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__121_
timestamp 1746535184
transform 1 0 36576 0 1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__122_
timestamp 1746535184
transform 1 0 37344 0 1 9828
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__123_
timestamp 1746535184
transform 1 0 35328 0 -1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__124_
timestamp 1746535184
transform 1 0 37056 0 1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__125_
timestamp 1746535184
transform 1 0 36864 0 1 12852
box -48 -56 2736 834
use sg13g2_inv_1  u_ppwm_u_mem__0613_
timestamp 1676382929
transform 1 0 11616 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0614_
timestamp 1676382929
transform 1 0 7776 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0615_
timestamp 1676382929
transform 1 0 16224 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0616_
timestamp 1676382929
transform -1 0 15840 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0617_
timestamp 1676382929
transform -1 0 5664 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0618_
timestamp 1676382929
transform 1 0 5664 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0619_
timestamp 1676382929
transform -1 0 5568 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0620_
timestamp 1676382929
transform -1 0 5664 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0621_
timestamp 1676382929
transform 1 0 10752 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0622_
timestamp 1676382929
transform -1 0 10560 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0623_
timestamp 1676382929
transform -1 0 9408 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0624_
timestamp 1676382929
transform -1 0 6240 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0625_
timestamp 1676382929
transform -1 0 2496 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0626_
timestamp 1676382929
transform 1 0 4800 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0627_
timestamp 1676382929
transform -1 0 6912 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0628_
timestamp 1676382929
transform 1 0 12576 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0629_
timestamp 1676382929
transform 1 0 18816 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0630_
timestamp 1676382929
transform 1 0 19872 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0631_
timestamp 1676382929
transform -1 0 21696 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0632_
timestamp 1676382929
transform 1 0 20448 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0633_
timestamp 1676382929
transform -1 0 10656 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0634_
timestamp 1676382929
transform -1 0 11328 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0635_
timestamp 1676382929
transform -1 0 13248 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0636_
timestamp 1676382929
transform 1 0 19104 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0637_
timestamp 1676382929
transform -1 0 19296 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0638_
timestamp 1676382929
transform -1 0 21216 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0639_
timestamp 1676382929
transform -1 0 19488 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0640_
timestamp 1676382929
transform -1 0 10272 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0641_
timestamp 1676382929
transform -1 0 6048 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0642_
timestamp 1676382929
transform -1 0 3456 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0643_
timestamp 1676382929
transform -1 0 3168 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0644_
timestamp 1676382929
transform -1 0 8064 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0645_
timestamp 1676382929
transform 1 0 13152 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0646_
timestamp 1676382929
transform 1 0 20256 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0647_
timestamp 1676382929
transform 1 0 21216 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0648_
timestamp 1676382929
transform -1 0 8832 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0649_
timestamp 1676382929
transform 1 0 7296 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0650_
timestamp 1676382929
transform -1 0 3936 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0651_
timestamp 1676382929
transform 1 0 7488 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0652_
timestamp 1676382929
transform 1 0 13728 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0653_
timestamp 1676382929
transform 1 0 14784 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0654_
timestamp 1676382929
transform -1 0 16320 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0655_
timestamp 1676382929
transform -1 0 13728 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0656_
timestamp 1676382929
transform -1 0 2880 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0657_
timestamp 1676382929
transform 1 0 4896 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0658_
timestamp 1676382929
transform -1 0 7776 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0659_
timestamp 1676382929
transform 1 0 10752 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0660_
timestamp 1676382929
transform 1 0 12384 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0661_
timestamp 1676382929
transform -1 0 14208 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0662_
timestamp 1676382929
transform -1 0 11328 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0663_
timestamp 1676382929
transform -1 0 10176 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0664_
timestamp 1676382929
transform -1 0 3648 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0665_
timestamp 1676382929
transform -1 0 4800 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0666_
timestamp 1676382929
transform 1 0 8736 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0667_
timestamp 1676382929
transform 1 0 14304 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0668_
timestamp 1676382929
transform 1 0 18240 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0669_
timestamp 1676382929
transform -1 0 21024 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0670_
timestamp 1676382929
transform -1 0 24288 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0671_
timestamp 1676382929
transform 1 0 28896 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0672_
timestamp 1676382929
transform -1 0 31104 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0673_
timestamp 1676382929
transform 1 0 37536 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0674_
timestamp 1676382929
transform -1 0 38688 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0675_
timestamp 1676382929
transform -1 0 39264 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0676_
timestamp 1676382929
transform -1 0 27744 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0677_
timestamp 1676382929
transform 1 0 25920 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0678_
timestamp 1676382929
transform 1 0 33024 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0679_
timestamp 1676382929
transform -1 0 34848 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0680_
timestamp 1676382929
transform 1 0 40032 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0681_
timestamp 1676382929
transform -1 0 43488 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0682_
timestamp 1676382929
transform -1 0 42336 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0683_
timestamp 1676382929
transform -1 0 31488 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0684_
timestamp 1676382929
transform -1 0 32640 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0685_
timestamp 1676382929
transform 1 0 28224 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0686_
timestamp 1676382929
transform 1 0 28320 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0687_
timestamp 1676382929
transform -1 0 31776 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0688_
timestamp 1676382929
transform -1 0 34464 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0689_
timestamp 1676382929
transform -1 0 33408 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0690_
timestamp 1676382929
transform -1 0 30048 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0691_
timestamp 1676382929
transform -1 0 28608 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0692_
timestamp 1676382929
transform -1 0 24288 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0693_
timestamp 1676382929
transform 1 0 27168 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0694_
timestamp 1676382929
transform -1 0 31008 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0695_
timestamp 1676382929
transform -1 0 36768 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0696_
timestamp 1676382929
transform -1 0 37920 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0697_
timestamp 1676382929
transform -1 0 33792 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0698_
timestamp 1676382929
transform 1 0 36000 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0699_
timestamp 1676382929
transform -1 0 39552 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0700_
timestamp 1676382929
transform 1 0 41856 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0701_
timestamp 1676382929
transform -1 0 43104 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0702_
timestamp 1676382929
transform -1 0 45984 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0703_
timestamp 1676382929
transform 1 0 45696 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0704_
timestamp 1676382929
transform -1 0 41568 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0705_
timestamp 1676382929
transform -1 0 38016 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0706_
timestamp 1676382929
transform -1 0 39264 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0707_
timestamp 1676382929
transform 1 0 45216 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0708_
timestamp 1676382929
transform -1 0 46656 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0709_
timestamp 1676382929
transform -1 0 46944 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0710_
timestamp 1676382929
transform -1 0 50016 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0711_
timestamp 1676382929
transform -1 0 42240 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0712_
timestamp 1676382929
transform -1 0 39168 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0713_
timestamp 1676382929
transform 1 0 40512 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0714_
timestamp 1676382929
transform 1 0 46848 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0715_
timestamp 1676382929
transform -1 0 46944 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0716_
timestamp 1676382929
transform 1 0 47136 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0717_
timestamp 1676382929
transform -1 0 49152 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0718_
timestamp 1676382929
transform -1 0 44640 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0719_
timestamp 1676382929
transform -1 0 37344 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0720_
timestamp 1676382929
transform 1 0 37056 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0721_
timestamp 1676382929
transform 1 0 46368 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0722_
timestamp 1676382929
transform -1 0 48576 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0723_
timestamp 1676382929
transform -1 0 43296 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0724_
timestamp 1676382929
transform -1 0 43008 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_mem__0725_
timestamp 1676382947
transform -1 0 8640 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_mem__0726_
timestamp 1676382929
transform -1 0 9216 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0727_
timestamp 1676382929
transform 1 0 38880 0 1 24948
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_mem__0728_
timestamp 1676382947
transform 1 0 25920 0 1 27972
box -48 -56 432 834
use sg13g2_inv_4  u_ppwm_u_mem__0729_
timestamp 1676383058
transform 1 0 24576 0 1 26460
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_mem__0730_
timestamp 1676639442
transform 1 0 8448 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__0731_
timestamp 1676627187
transform 1 0 8064 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0732_
timestamp 1683973020
transform -1 0 9216 0 1 14364
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_mem__0733_
timestamp 1683988354
transform 1 0 4224 0 -1 15876
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_mem__0734_
timestamp 1683988354
transform 1 0 4320 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__0735_
timestamp 1676639442
transform -1 0 7008 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_mem__0736_
timestamp 1676557249
transform -1 0 8640 0 -1 17388
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_mem__0737_
timestamp 1676643125
transform 1 0 6432 0 -1 15876
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_mem__0738_
timestamp 1677175127
transform 1 0 7104 0 -1 15876
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_mem__0739_
timestamp 1683988354
transform 1 0 7776 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0740_
timestamp 1685175443
transform 1 0 7776 0 -1 17388
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0741_
timestamp 1677247768
transform 1 0 13824 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0742_
timestamp 1677247768
transform -1 0 18240 0 -1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0743_
timestamp 1676557249
transform -1 0 17088 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0744_
timestamp 1683973020
transform -1 0 14976 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0745_
timestamp 1677247768
transform 1 0 11136 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0746_
timestamp 1676557249
transform 1 0 12192 0 1 27972
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0747_
timestamp 1677247768
transform 1 0 7584 0 -1 24948
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0748_
timestamp 1683973020
transform -1 0 12960 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0749_
timestamp 1685197497
transform 1 0 14208 0 -1 26460
box -48 -56 816 834
use sg13g2_mux4_1  u_ppwm_u_mem__0750_
timestamp 1677257233
transform -1 0 41760 0 -1 24948
box -48 -56 2064 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0751_
timestamp 1676567195
transform 1 0 40416 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0752_
timestamp 1677247768
transform 1 0 30816 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0753_
timestamp 1677247768
transform -1 0 32736 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0754_
timestamp 1676557249
transform 1 0 31872 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0755_
timestamp 1683973020
transform 1 0 30912 0 -1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0756_
timestamp 1683973020
transform 1 0 30816 0 1 26460
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0757_
timestamp 1683996397
transform 1 0 30432 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0758_
timestamp 1677247768
transform 1 0 4032 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0759_
timestamp 1677247768
transform -1 0 17760 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0760_
timestamp 1676557249
transform 1 0 17088 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0761_
timestamp 1683973020
transform -1 0 18048 0 1 24948
box -48 -56 528 834
use sg13g2_mux4_1  u_ppwm_u_mem__0762_
timestamp 1677257233
transform -1 0 19392 0 1 32508
box -48 -56 2064 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0763_
timestamp 1685175443
transform 1 0 17472 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0764_
timestamp 1683973020
transform -1 0 18528 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_mem__0765_
timestamp 1676557249
transform 1 0 36192 0 -1 27972
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0766_
timestamp 1685175443
transform 1 0 38112 0 -1 27972
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0767_
timestamp 1676557249
transform 1 0 40032 0 -1 35532
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0768_
timestamp 1685175443
transform -1 0 40704 0 1 34020
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0769_
timestamp 1676557249
transform 1 0 44640 0 -1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0770_
timestamp 1685175443
transform -1 0 44640 0 -1 26460
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0771_
timestamp 1676557249
transform 1 0 42240 0 1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0772_
timestamp 1685175443
transform -1 0 42624 0 -1 26460
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0773_
timestamp 1677257233
transform -1 0 41088 0 -1 26460
box -48 -56 2064 834
use sg13g2_a21o_2  u_ppwm_u_mem__0774_
timestamp 1683996397
transform 1 0 25344 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0775_
timestamp 1677247768
transform 1 0 4320 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0776_
timestamp 1676557249
transform 1 0 14976 0 -1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0777_
timestamp 1677247768
transform -1 0 20448 0 -1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0778_
timestamp 1683973020
transform 1 0 15936 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0779_
timestamp 1677247768
transform -1 0 14976 0 1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0780_
timestamp 1676557249
transform -1 0 13440 0 -1 30996
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0781_
timestamp 1677247768
transform 1 0 13344 0 1 34020
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0782_
timestamp 1683973020
transform -1 0 14496 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0783_
timestamp 1685197497
transform 1 0 14688 0 -1 27972
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_mem__0784_
timestamp 1676557249
transform -1 0 37344 0 -1 30996
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0785_
timestamp 1685175443
transform 1 0 37344 0 1 29484
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0786_
timestamp 1676557249
transform -1 0 40800 0 1 32508
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0787_
timestamp 1685175443
transform -1 0 42048 0 -1 30996
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0788_
timestamp 1676557249
transform 1 0 41568 0 -1 29484
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0789_
timestamp 1685175443
transform -1 0 43776 0 1 27972
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0790_
timestamp 1676557249
transform 1 0 44256 0 -1 27972
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0791_
timestamp 1685175443
transform 1 0 43584 0 -1 27972
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0792_
timestamp 1677257233
transform -1 0 41760 0 1 27972
box -48 -56 2064 834
use sg13g2_a21o_2  u_ppwm_u_mem__0793_
timestamp 1683996397
transform -1 0 25344 0 -1 27972
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0794_
timestamp 1677247768
transform 1 0 10464 0 1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0795_
timestamp 1676557249
transform 1 0 11808 0 1 27972
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0796_
timestamp 1677247768
transform -1 0 20160 0 1 26460
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0797_
timestamp 1683973020
transform 1 0 14976 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0798_
timestamp 1677247768
transform 1 0 12000 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0799_
timestamp 1676557249
transform 1 0 13920 0 1 29484
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0800_
timestamp 1677247768
transform 1 0 8448 0 -1 34020
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0801_
timestamp 1683973020
transform -1 0 13056 0 1 27972
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0802_
timestamp 1685197497
transform 1 0 13536 0 -1 27972
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0803_
timestamp 1677247768
transform 1 0 30720 0 -1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0804_
timestamp 1677247768
transform -1 0 37824 0 1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0805_
timestamp 1683973020
transform 1 0 31296 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0806_
timestamp 1685175443
transform 1 0 31392 0 -1 27972
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0807_
timestamp 1677257233
transform -1 0 45792 0 1 27972
box -48 -56 2064 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0808_
timestamp 1683973020
transform 1 0 30432 0 -1 27972
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0809_
timestamp 1683996397
transform 1 0 29856 0 1 26460
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0810_
timestamp 1685175443
transform 1 0 13920 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  u_ppwm_u_mem__0811_
timestamp 1677175127
transform -1 0 15168 0 1 24948
box -48 -56 720 834
use sg13g2_mux2_1  u_ppwm_u_mem__0812_
timestamp 1677247768
transform -1 0 18048 0 -1 24948
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0813_
timestamp 1683973020
transform -1 0 17568 0 1 24948
box -48 -56 528 834
use sg13g2_mux4_1  u_ppwm_u_mem__0814_
timestamp 1677257233
transform 1 0 6720 0 -1 30996
box -48 -56 2064 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0815_
timestamp 1685175443
transform 1 0 15840 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0816_
timestamp 1683973020
transform 1 0 16320 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0817_
timestamp 1677247768
transform -1 0 39648 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0818_
timestamp 1676557249
transform -1 0 29760 0 1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0819_
timestamp 1677247768
transform -1 0 42144 0 1 24948
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0820_
timestamp 1683973020
transform 1 0 29472 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0821_
timestamp 1685175443
transform -1 0 31008 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0822_
timestamp 1683973020
transform -1 0 30528 0 -1 29484
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0823_
timestamp 1677247768
transform 1 0 27360 0 -1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0824_
timestamp 1683973020
transform -1 0 29184 0 1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0825_
timestamp 1676567195
transform -1 0 28704 0 1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0826_
timestamp 1683973020
transform 1 0 28704 0 1 26460
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_mem__0827_
timestamp 1677175127
transform 1 0 27552 0 -1 24948
box -48 -56 720 834
use sg13g2_nor2b_1  u_ppwm_u_mem__0828_
timestamp 1685181386
transform 1 0 15168 0 -1 24948
box -54 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0829_
timestamp 1685175443
transform 1 0 14688 0 -1 24948
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0830_
timestamp 1676557249
transform 1 0 14592 0 1 23436
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0831_
timestamp 1676567195
transform 1 0 15552 0 1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0832_
timestamp 1683973020
transform -1 0 17088 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0833_
timestamp 1685175443
transform 1 0 15648 0 -1 24948
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0834_
timestamp 1677257233
transform 1 0 4416 0 1 29484
box -48 -56 2064 834
use sg13g2_nor2_1  u_ppwm_u_mem__0835_
timestamp 1676627187
transform -1 0 15744 0 -1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0836_
timestamp 1685175443
transform -1 0 16608 0 -1 24948
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0837_
timestamp 1677247768
transform 1 0 27168 0 -1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0838_
timestamp 1677247768
transform 1 0 27744 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0839_
timestamp 1677247768
transform -1 0 36192 0 1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0840_
timestamp 1677247768
transform -1 0 36384 0 -1 23436
box -48 -56 1008 834
use sg13g2_mux4_1  u_ppwm_u_mem__0841_
timestamp 1677257233
transform 1 0 27840 0 -1 27972
box -48 -56 2064 834
use sg13g2_nand2_1  u_ppwm_u_mem__0842_
timestamp 1676557249
transform -1 0 24576 0 1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0843_
timestamp 1685175443
transform 1 0 23616 0 -1 26460
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0844_
timestamp 1677247768
transform 1 0 7296 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0845_
timestamp 1676557249
transform 1 0 10176 0 -1 24948
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0846_
timestamp 1677247768
transform 1 0 12960 0 1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0847_
timestamp 1683973020
transform 1 0 13056 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0848_
timestamp 1677247768
transform 1 0 12096 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0849_
timestamp 1677247768
transform -1 0 12576 0 1 20412
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0850_
timestamp 1676557249
transform -1 0 11232 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0851_
timestamp 1683973020
transform -1 0 13536 0 -1 24948
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0852_
timestamp 1685197497
transform -1 0 14016 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0853_
timestamp 1677247768
transform -1 0 27840 0 1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0854_
timestamp 1677247768
transform 1 0 25440 0 -1 34020
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0855_
timestamp 1683973020
transform 1 0 26688 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0856_
timestamp 1685175443
transform -1 0 26784 0 1 27972
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0857_
timestamp 1677257233
transform 1 0 36576 0 -1 24948
box -48 -56 2064 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0858_
timestamp 1683973020
transform 1 0 28224 0 -1 24948
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0859_
timestamp 1683996397
transform 1 0 27072 0 -1 26460
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0860_
timestamp 1685175443
transform -1 0 44160 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0861_
timestamp 1683973020
transform -1 0 43488 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0862_
timestamp 1685175443
transform -1 0 43968 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0863_
timestamp 1683973020
transform -1 0 43584 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0864_
timestamp 1685175443
transform 1 0 47616 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0865_
timestamp 1683973020
transform 1 0 48192 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0866_
timestamp 1685175443
transform -1 0 49056 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0867_
timestamp 1683973020
transform -1 0 47424 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0868_
timestamp 1685175443
transform -1 0 41952 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0869_
timestamp 1683973020
transform -1 0 42048 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0870_
timestamp 1685175443
transform 1 0 34944 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0871_
timestamp 1683973020
transform 1 0 36384 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0872_
timestamp 1685175443
transform 1 0 44640 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0873_
timestamp 1683973020
transform 1 0 45120 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0874_
timestamp 1685175443
transform 1 0 47328 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0875_
timestamp 1683973020
transform 1 0 47904 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0876_
timestamp 1685175443
transform 1 0 47328 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0877_
timestamp 1683973020
transform 1 0 47808 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0878_
timestamp 1685175443
transform 1 0 45024 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0879_
timestamp 1683973020
transform 1 0 45888 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0880_
timestamp 1685175443
transform 1 0 47424 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0881_
timestamp 1683973020
transform -1 0 49440 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0882_
timestamp 1685175443
transform -1 0 42144 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0883_
timestamp 1683973020
transform -1 0 41664 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0884_
timestamp 1685175443
transform 1 0 37824 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0885_
timestamp 1683973020
transform -1 0 37824 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0886_
timestamp 1685175443
transform -1 0 40128 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0887_
timestamp 1683973020
transform -1 0 39360 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0888_
timestamp 1685175443
transform 1 0 47328 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0889_
timestamp 1683973020
transform 1 0 48384 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0890_
timestamp 1685175443
transform -1 0 48576 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0891_
timestamp 1683973020
transform -1 0 49056 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0892_
timestamp 1685175443
transform 1 0 48192 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0893_
timestamp 1683973020
transform -1 0 47424 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0894_
timestamp 1685175443
transform -1 0 45984 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0895_
timestamp 1683973020
transform -1 0 45216 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0896_
timestamp 1685175443
transform -1 0 39456 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0897_
timestamp 1683973020
transform -1 0 38496 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0898_
timestamp 1685175443
transform -1 0 35808 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0899_
timestamp 1683973020
transform 1 0 35808 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0900_
timestamp 1685175443
transform -1 0 38880 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0901_
timestamp 1683973020
transform 1 0 40128 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0902_
timestamp 1685175443
transform 1 0 44256 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0903_
timestamp 1683973020
transform -1 0 46464 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0904_
timestamp 1685175443
transform 1 0 43776 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0905_
timestamp 1683973020
transform 1 0 44256 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0906_
timestamp 1685175443
transform 1 0 43104 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0907_
timestamp 1683973020
transform 1 0 44736 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0908_
timestamp 1685175443
transform -1 0 43296 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0909_
timestamp 1683973020
transform -1 0 42816 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0910_
timestamp 1685175443
transform 1 0 38208 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0911_
timestamp 1683973020
transform 1 0 38496 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0912_
timestamp 1685175443
transform 1 0 34656 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0913_
timestamp 1683973020
transform 1 0 35520 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0914_
timestamp 1685175443
transform -1 0 34464 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0915_
timestamp 1683973020
transform -1 0 33120 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0916_
timestamp 1685175443
transform -1 0 34560 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0917_
timestamp 1683973020
transform -1 0 34272 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0918_
timestamp 1685175443
transform 1 0 37056 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0919_
timestamp 1683973020
transform -1 0 36384 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0920_
timestamp 1685175443
transform 1 0 32256 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0921_
timestamp 1683973020
transform -1 0 33696 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0922_
timestamp 1685175443
transform 1 0 27456 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0923_
timestamp 1683973020
transform -1 0 28224 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0924_
timestamp 1685175443
transform 1 0 27264 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0925_
timestamp 1683973020
transform 1 0 23424 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0926_
timestamp 1685175443
transform 1 0 26208 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0927_
timestamp 1683973020
transform 1 0 27168 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0928_
timestamp 1685175443
transform -1 0 28800 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0929_
timestamp 1683973020
transform 1 0 28992 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0930_
timestamp 1685175443
transform 1 0 30528 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0931_
timestamp 1683973020
transform 1 0 31392 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0932_
timestamp 1685175443
transform -1 0 34176 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0933_
timestamp 1683973020
transform 1 0 33408 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0934_
timestamp 1685175443
transform -1 0 35712 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0935_
timestamp 1683973020
transform -1 0 34656 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0936_
timestamp 1685175443
transform 1 0 30720 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0937_
timestamp 1683973020
transform -1 0 29472 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0938_
timestamp 1685175443
transform -1 0 26304 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0939_
timestamp 1683973020
transform 1 0 25824 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0940_
timestamp 1685175443
transform -1 0 25920 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0941_
timestamp 1683973020
transform 1 0 27840 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0942_
timestamp 1685175443
transform -1 0 32256 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0943_
timestamp 1683973020
transform -1 0 32064 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0944_
timestamp 1685175443
transform 1 0 39264 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0945_
timestamp 1683973020
transform 1 0 39744 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0946_
timestamp 1685175443
transform 1 0 42720 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0947_
timestamp 1683973020
transform -1 0 42336 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0948_
timestamp 1685175443
transform 1 0 41184 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0949_
timestamp 1683973020
transform 1 0 41568 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0950_
timestamp 1685175443
transform -1 0 36768 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0951_
timestamp 1683973020
transform -1 0 35712 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0952_
timestamp 1685175443
transform 1 0 29760 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0953_
timestamp 1683973020
transform 1 0 32160 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0954_
timestamp 1685175443
transform -1 0 27744 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0955_
timestamp 1683973020
transform -1 0 27168 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0956_
timestamp 1685175443
transform -1 0 25824 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0957_
timestamp 1683973020
transform 1 0 26208 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0958_
timestamp 1685175443
transform 1 0 35712 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0959_
timestamp 1683973020
transform 1 0 38304 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0960_
timestamp 1685175443
transform 1 0 38784 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0961_
timestamp 1683973020
transform 1 0 39264 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0962_
timestamp 1685175443
transform -1 0 39168 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0963_
timestamp 1683973020
transform -1 0 38400 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0964_
timestamp 1685175443
transform -1 0 34560 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0965_
timestamp 1683973020
transform -1 0 34080 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0966_
timestamp 1685175443
transform -1 0 30816 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0967_
timestamp 1683973020
transform -1 0 29952 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0968_
timestamp 1685175443
transform -1 0 26496 0 -1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0969_
timestamp 1683973020
transform -1 0 26016 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0970_
timestamp 1685175443
transform -1 0 21504 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0971_
timestamp 1683973020
transform -1 0 21984 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0972_
timestamp 1685175443
transform -1 0 19584 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0973_
timestamp 1683973020
transform -1 0 19008 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0974_
timestamp 1685175443
transform -1 0 17376 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0975_
timestamp 1683973020
transform -1 0 15072 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0976_
timestamp 1685175443
transform -1 0 11808 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0977_
timestamp 1683973020
transform -1 0 9504 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0978_
timestamp 1685175443
transform -1 0 6720 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0979_
timestamp 1683973020
transform -1 0 5760 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0980_
timestamp 1685175443
transform -1 0 2976 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0981_
timestamp 1683973020
transform -1 0 2496 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0982_
timestamp 1685175443
transform 1 0 3936 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0983_
timestamp 1683973020
transform 1 0 4416 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0984_
timestamp 1685175443
transform 1 0 12288 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0985_
timestamp 1683973020
transform -1 0 13920 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0986_
timestamp 1685175443
transform 1 0 14208 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0987_
timestamp 1683973020
transform 1 0 16416 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0988_
timestamp 1685175443
transform -1 0 13344 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0989_
timestamp 1683973020
transform -1 0 12960 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0990_
timestamp 1685175443
transform -1 0 12288 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0991_
timestamp 1683973020
transform -1 0 9216 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0992_
timestamp 1685175443
transform -1 0 5280 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0993_
timestamp 1683973020
transform 1 0 5760 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0994_
timestamp 1685175443
transform -1 0 6720 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0995_
timestamp 1683973020
transform -1 0 5664 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0996_
timestamp 1685175443
transform 1 0 3936 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0997_
timestamp 1683973020
transform 1 0 4416 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0998_
timestamp 1685175443
transform -1 0 11328 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0999_
timestamp 1683973020
transform 1 0 11520 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1000_
timestamp 1685175443
transform -1 0 14880 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1001_
timestamp 1683973020
transform -1 0 13920 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1002_
timestamp 1685175443
transform -1 0 15552 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1003_
timestamp 1683973020
transform 1 0 15072 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1004_
timestamp 1685175443
transform -1 0 13152 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1005_
timestamp 1683973020
transform 1 0 12192 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1006_
timestamp 1685175443
transform -1 0 8352 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1007_
timestamp 1683973020
transform -1 0 7200 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1008_
timestamp 1685175443
transform -1 0 3648 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1009_
timestamp 1683973020
transform 1 0 2688 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1010_
timestamp 1685175443
transform -1 0 4416 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1011_
timestamp 1683973020
transform 1 0 3936 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1012_
timestamp 1685175443
transform 1 0 6528 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1013_
timestamp 1683973020
transform 1 0 7008 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1014_
timestamp 1685175443
transform 1 0 18528 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1015_
timestamp 1683973020
transform 1 0 20736 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1016_
timestamp 1685175443
transform 1 0 17856 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1017_
timestamp 1683973020
transform 1 0 19392 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1018_
timestamp 1685175443
transform -1 0 16032 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1019_
timestamp 1683973020
transform -1 0 16896 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1020_
timestamp 1685175443
transform 1 0 7488 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1021_
timestamp 1683973020
transform -1 0 8928 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1022_
timestamp 1685175443
transform -1 0 5952 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1023_
timestamp 1683973020
transform -1 0 5472 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1024_
timestamp 1685175443
transform -1 0 4224 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1025_
timestamp 1683973020
transform -1 0 3936 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1026_
timestamp 1685175443
transform 1 0 3744 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1027_
timestamp 1683973020
transform 1 0 4224 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1028_
timestamp 1685175443
transform 1 0 7584 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1029_
timestamp 1683973020
transform 1 0 9024 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1030_
timestamp 1685175443
transform 1 0 18624 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1031_
timestamp 1683973020
transform 1 0 19968 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1032_
timestamp 1685175443
transform 1 0 19488 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1033_
timestamp 1683973020
transform 1 0 19968 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1034_
timestamp 1685175443
transform -1 0 19104 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1035_
timestamp 1683973020
transform 1 0 18528 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1036_
timestamp 1685175443
transform 1 0 16512 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1037_
timestamp 1683973020
transform -1 0 16512 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1038_
timestamp 1685175443
transform -1 0 15456 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1039_
timestamp 1683973020
transform -1 0 14016 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1040_
timestamp 1685175443
transform -1 0 14496 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1041_
timestamp 1683973020
transform -1 0 11040 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1042_
timestamp 1685175443
transform 1 0 12096 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1043_
timestamp 1683973020
transform -1 0 11136 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1044_
timestamp 1685175443
transform 1 0 19104 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1045_
timestamp 1683973020
transform 1 0 20448 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1046_
timestamp 1685175443
transform 1 0 20448 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1047_
timestamp 1683973020
transform 1 0 20928 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1048_
timestamp 1685175443
transform 1 0 19008 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1049_
timestamp 1683973020
transform 1 0 19488 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1050_
timestamp 1685175443
transform -1 0 18432 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1051_
timestamp 1683973020
transform -1 0 17088 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1052_
timestamp 1685175443
transform -1 0 13920 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1053_
timestamp 1683973020
transform -1 0 12672 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1054_
timestamp 1685175443
transform -1 0 8736 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1055_
timestamp 1683973020
transform -1 0 7392 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1056_
timestamp 1685175443
transform -1 0 5568 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1057_
timestamp 1683973020
transform -1 0 5376 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1058_
timestamp 1685175443
transform -1 0 3744 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1059_
timestamp 1683973020
transform -1 0 2976 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1060_
timestamp 1685175443
transform 1 0 5568 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1061_
timestamp 1683973020
transform 1 0 2976 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1062_
timestamp 1685175443
transform 1 0 6336 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1063_
timestamp 1683973020
transform 1 0 6720 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1064_
timestamp 1685175443
transform 1 0 9504 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1065_
timestamp 1683973020
transform 1 0 10272 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1066_
timestamp 1685175443
transform 1 0 11040 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1067_
timestamp 1683973020
transform 1 0 12000 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1068_
timestamp 1685175443
transform 1 0 5952 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1069_
timestamp 1683973020
transform 1 0 7584 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1070_
timestamp 1685175443
transform -1 0 5376 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1071_
timestamp 1683973020
transform 1 0 4416 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1072_
timestamp 1685175443
transform -1 0 4224 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1073_
timestamp 1683973020
transform 1 0 2592 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1074_
timestamp 1685175443
transform -1 0 4800 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1075_
timestamp 1683973020
transform 1 0 3840 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1076_
timestamp 1685175443
transform 1 0 9120 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1077_
timestamp 1683973020
transform 1 0 9600 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1078_
timestamp 1685175443
transform -1 0 16032 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1079_
timestamp 1683973020
transform 1 0 15072 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1080_
timestamp 1685175443
transform -1 0 15360 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1081_
timestamp 1683973020
transform -1 0 12384 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1082_
timestamp 1685175443
transform -1 0 10656 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1083_
timestamp 1683973020
transform -1 0 8832 0 1 17388
box -48 -56 528 834
use sg13g2_nand2b_2  u_ppwm_u_mem__1084_
timestamp 1685211885
transform -1 0 7680 0 1 15876
box -48 -56 816 834
use sg13g2_nand2_2  u_ppwm_u_mem__1085_
timestamp 1685180049
transform 1 0 6240 0 1 15876
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_mem__1086_
timestamp 1676627187
transform -1 0 5280 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1087_
timestamp 1676901763
transform -1 0 4512 0 -1 17388
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1088_
timestamp 1676639442
transform -1 0 4320 0 1 18900
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1089_
timestamp 1676627187
transform 1 0 3168 0 -1 17388
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1090_
timestamp 1676901763
transform 1 0 4704 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1091_
timestamp 1676639442
transform 1 0 3552 0 -1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1092_
timestamp 1683973020
transform 1 0 5376 0 1 15876
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_mem__1093_
timestamp 1676985977
transform 1 0 4512 0 -1 17388
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_mem__1094_
timestamp 1676639442
transform -1 0 6048 0 -1 17388
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1095_
timestamp 1676627187
transform 1 0 2976 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1096_
timestamp 1676901763
transform -1 0 4224 0 -1 15876
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1097_
timestamp 1676639442
transform 1 0 3360 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1098_
timestamp 1676627187
transform -1 0 4032 0 -1 12852
box -48 -56 432 834
use sg13g2_and3_1  u_ppwm_u_mem__1099_
timestamp 1676971669
transform -1 0 4032 0 1 14364
box -48 -56 720 834
use sg13g2_nor3_1  u_ppwm_u_mem__1100_
timestamp 1676639442
transform -1 0 3360 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1101_
timestamp 1676627187
transform -1 0 6240 0 1 15876
box -48 -56 432 834
use sg13g2_and4_1  u_ppwm_u_mem__1102_
timestamp 1676985977
transform 1 0 4032 0 1 14364
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_mem__1103_
timestamp 1676639442
transform 1 0 4128 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1104_
timestamp 1683973020
transform 1 0 5664 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1105_
timestamp 1683973020
transform -1 0 8352 0 1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_mem__1106_
timestamp 1685181386
transform 1 0 5088 0 -1 12852
box -54 -56 528 834
use sg13g2_tiehi  u_ppwm_u_mem__1107__173
timestamp 1680000651
transform 1 0 42048 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1107_
timestamp 1746535128
transform 1 0 41856 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1108__145
timestamp 1680000651
transform -1 0 42528 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1108_
timestamp 1746535128
transform 1 0 41664 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1109__143
timestamp 1680000651
transform 1 0 49728 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1109_
timestamp 1746535128
transform -1 0 51744 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1110_
timestamp 1746535128
transform 1 0 48096 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1110__141
timestamp 1680000651
transform -1 0 50496 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1111_
timestamp 1746535184
transform 1 0 42144 0 1 20412
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1111__139
timestamp 1680000651
transform -1 0 43104 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1112_
timestamp 1746535128
transform 1 0 34368 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1112__137
timestamp 1680000651
transform -1 0 35232 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1113_
timestamp 1746535128
transform -1 0 47520 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1113__135
timestamp 1680000651
transform 1 0 45888 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1114__133
timestamp 1680000651
transform 1 0 49248 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1114_
timestamp 1746535184
transform -1 0 51264 0 -1 23436
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1115__131
timestamp 1680000651
transform 1 0 48480 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1115_
timestamp 1746535128
transform 1 0 48672 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1116__129
timestamp 1680000651
transform -1 0 46752 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1116_
timestamp 1746535128
transform 1 0 45504 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1117__127
timestamp 1680000651
transform -1 0 51552 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1117_
timestamp 1746535128
transform -1 0 51744 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1118_
timestamp 1746535184
transform 1 0 42240 0 1 21924
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1118__125
timestamp 1680000651
transform 1 0 40800 0 -1 23436
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1119__123
timestamp 1680000651
transform -1 0 39168 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1119_
timestamp 1746535128
transform 1 0 38304 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1120__121
timestamp 1680000651
transform 1 0 39264 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1120_
timestamp 1746535128
transform 1 0 39168 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1121_
timestamp 1746535184
transform 1 0 49344 0 -1 24948
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1121__119
timestamp 1680000651
transform -1 0 50208 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1122_
timestamp 1746535128
transform 1 0 49536 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1122__117
timestamp 1680000651
transform -1 0 51168 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1123_
timestamp 1746535128
transform 1 0 47232 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1123__115
timestamp 1680000651
transform -1 0 48192 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1124_
timestamp 1746535128
transform 1 0 44640 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1124__113
timestamp 1680000651
transform 1 0 44544 0 1 32508
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1125__111
timestamp 1680000651
transform 1 0 38784 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1125_
timestamp 1746535128
transform 1 0 39264 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1126_
timestamp 1746535128
transform 1 0 36288 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1126__109
timestamp 1680000651
transform -1 0 37248 0 -1 27972
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1127__107
timestamp 1680000651
transform 1 0 37056 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1127_
timestamp 1746535128
transform -1 0 39456 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1128__105
timestamp 1680000651
transform -1 0 47904 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1128_
timestamp 1746535184
transform 1 0 46656 0 1 21924
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1129__103
timestamp 1680000651
transform -1 0 45600 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1129_
timestamp 1746535128
transform 1 0 44736 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1130_
timestamp 1746535128
transform 1 0 44448 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1130__101
timestamp 1680000651
transform -1 0 45600 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1131_
timestamp 1746535128
transform 1 0 42144 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1131__99
timestamp 1680000651
transform 1 0 42336 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1132__97
timestamp 1680000651
transform -1 0 41184 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1132_
timestamp 1746535128
transform 1 0 39648 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1133_
timestamp 1746535128
transform 1 0 36000 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1133__95
timestamp 1680000651
transform -1 0 37152 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1134_
timestamp 1746535128
transform 1 0 32736 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1134__93
timestamp 1680000651
transform 1 0 32256 0 1 24948
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1135__91
timestamp 1680000651
transform 1 0 32832 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1135_
timestamp 1746535128
transform -1 0 35328 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1136_
timestamp 1746535128
transform 1 0 35904 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1136__89
timestamp 1680000651
transform -1 0 36768 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1137_
timestamp 1746535128
transform 1 0 33600 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1137__87
timestamp 1680000651
transform -1 0 34944 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1138_
timestamp 1746535128
transform -1 0 30528 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1138__85
timestamp 1680000651
transform 1 0 28992 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1139__83
timestamp 1680000651
transform -1 0 24672 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1139_
timestamp 1746535128
transform 1 0 23232 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1140_
timestamp 1746535128
transform 1 0 22560 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1140__81
timestamp 1680000651
transform 1 0 22752 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1141_
timestamp 1746535128
transform 1 0 28800 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1141__79
timestamp 1680000651
transform 1 0 28512 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1142__77
timestamp 1680000651
transform 1 0 32736 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1142_
timestamp 1746535128
transform -1 0 33600 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1143_
timestamp 1746535128
transform 1 0 33120 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1143__75
timestamp 1680000651
transform 1 0 32832 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1144__73
timestamp 1680000651
transform 1 0 35136 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1144_
timestamp 1746535128
transform 1 0 34944 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1145__71
timestamp 1680000651
transform 1 0 28608 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1145_
timestamp 1746535128
transform 1 0 28896 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1146_
timestamp 1746535128
transform 1 0 24768 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1146__69
timestamp 1680000651
transform 1 0 24288 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1147_
timestamp 1746535128
transform -1 0 26688 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1147__67
timestamp 1680000651
transform 1 0 25152 0 -1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1148__65
timestamp 1680000651
transform 1 0 29952 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1148_
timestamp 1746535128
transform 1 0 31008 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1149_
timestamp 1746535184
transform 1 0 40800 0 -1 35532
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1149__63
timestamp 1680000651
transform 1 0 40416 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1150__61
timestamp 1680000651
transform 1 0 43392 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1150_
timestamp 1746535128
transform 1 0 43488 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1151_
timestamp 1746535128
transform 1 0 41664 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1151__59
timestamp 1680000651
transform 1 0 40800 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1152_
timestamp 1746535128
transform 1 0 35904 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1152__57
timestamp 1680000651
transform 1 0 34848 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1153_
timestamp 1746535184
transform 1 0 32640 0 1 35532
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1153__55
timestamp 1680000651
transform -1 0 33792 0 -1 37044
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1154__172
timestamp 1680000651
transform -1 0 28128 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1154_
timestamp 1746535128
transform 1 0 26976 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1155__170
timestamp 1680000651
transform -1 0 24192 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1155_
timestamp 1746535128
transform 1 0 23328 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1156_
timestamp 1746535184
transform -1 0 38112 0 1 35532
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1156__168
timestamp 1680000651
transform 1 0 36192 0 -1 37044
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1157__166
timestamp 1680000651
transform 1 0 38880 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1157_
timestamp 1746535128
transform 1 0 38976 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1158__164
timestamp 1680000651
transform -1 0 38688 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1158_
timestamp 1746535128
transform 1 0 37824 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1159__162
timestamp 1680000651
transform -1 0 34944 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1159_
timestamp 1746535128
transform 1 0 33312 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1160_
timestamp 1746535128
transform 1 0 29568 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1160__160
timestamp 1680000651
transform 1 0 29376 0 -1 37044
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1161__158
timestamp 1680000651
transform -1 0 25248 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1161_
timestamp 1746535128
transform 1 0 24384 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1162_
timestamp 1746535128
transform 1 0 21312 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1162__156
timestamp 1680000651
transform -1 0 22752 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1163__154
timestamp 1680000651
transform -1 0 20064 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1163_
timestamp 1746535128
transform 1 0 18720 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1164__152
timestamp 1680000651
transform -1 0 17760 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1164_
timestamp 1746535128
transform 1 0 15648 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1165_
timestamp 1746535128
transform 1 0 9216 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1165__150
timestamp 1680000651
transform -1 0 10752 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1166__148
timestamp 1680000651
transform -1 0 4800 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1166_
timestamp 1746535128
transform 1 0 3552 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1167__146
timestamp 1680000651
transform -1 0 2880 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1167_
timestamp 1746535128
transform 1 0 1920 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1168__142
timestamp 1680000651
transform -1 0 2016 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1168_
timestamp 1746535128
transform 1 0 1248 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1169__138
timestamp 1680000651
transform 1 0 11808 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1169_
timestamp 1746535128
transform -1 0 14304 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1170_
timestamp 1746535128
transform 1 0 15264 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1170__134
timestamp 1680000651
transform -1 0 16608 0 -1 37044
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1171__130
timestamp 1680000651
transform -1 0 14208 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1171_
timestamp 1746535128
transform 1 0 12672 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1172_
timestamp 1746535128
transform 1 0 9408 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1172__126
timestamp 1680000651
transform -1 0 10272 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1173_
timestamp 1746535128
transform 1 0 6144 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1173__122
timestamp 1680000651
transform -1 0 7488 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1174__118
timestamp 1680000651
transform 1 0 4896 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1174_
timestamp 1746535128
transform 1 0 4896 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1175_
timestamp 1746535128
transform 1 0 1152 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1175__114
timestamp 1680000651
transform 1 0 768 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1176__110
timestamp 1680000651
transform -1 0 11712 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1176_
timestamp 1746535128
transform 1 0 10848 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1177_
timestamp 1746535128
transform 1 0 14880 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1177__106
timestamp 1680000651
transform 1 0 14976 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1178_
timestamp 1746535128
transform 1 0 14784 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1178__102
timestamp 1680000651
transform 1 0 14400 0 -1 32508
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1179__98
timestamp 1680000651
transform 1 0 10176 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1179_
timestamp 1746535128
transform 1 0 11808 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1180__94
timestamp 1680000651
transform 1 0 8064 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1180_
timestamp 1746535128
transform 1 0 8352 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1181__90
timestamp 1680000651
transform -1 0 2208 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1181_
timestamp 1746535128
transform 1 0 1248 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1182_
timestamp 1746535128
transform 1 0 1248 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1182__86
timestamp 1680000651
transform -1 0 2112 0 -1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1183__82
timestamp 1680000651
transform 1 0 6144 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1183_
timestamp 1746535128
transform -1 0 7200 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1184_
timestamp 1746535184
transform 1 0 19872 0 -1 30996
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1184__78
timestamp 1680000651
transform 1 0 19488 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1185__74
timestamp 1680000651
transform 1 0 21120 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1185_
timestamp 1746535128
transform -1 0 22656 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1186_
timestamp 1746535128
transform 1 0 16896 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1186__70
timestamp 1680000651
transform -1 0 17760 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1187_
timestamp 1746535128
transform 1 0 8832 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1187__66
timestamp 1680000651
transform -1 0 10176 0 -1 30996
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1188__62
timestamp 1680000651
transform 1 0 7104 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1188_
timestamp 1746535128
transform -1 0 8544 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1189_
timestamp 1746535128
transform 1 0 1152 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1189__58
timestamp 1680000651
transform -1 0 2016 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1190_
timestamp 1746535128
transform 1 0 1152 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1190__54
timestamp 1680000651
transform 1 0 768 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1191__169
timestamp 1680000651
transform -1 0 10368 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1191_
timestamp 1746535128
transform 1 0 8928 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1192_
timestamp 1746535184
transform -1 0 19104 0 -1 29484
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1192__165
timestamp 1680000651
transform 1 0 16032 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1193_
timestamp 1746535128
transform -1 0 23040 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1193__161
timestamp 1680000651
transform 1 0 22080 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1194__157
timestamp 1680000651
transform 1 0 21120 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1194_
timestamp 1746535128
transform -1 0 21888 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1195__153
timestamp 1680000651
transform -1 0 18240 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1195_
timestamp 1746535128
transform 1 0 17280 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1196__149
timestamp 1680000651
transform -1 0 16032 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1196_
timestamp 1746535128
transform 1 0 13536 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1197__144
timestamp 1680000651
transform 1 0 9792 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1197_
timestamp 1746535128
transform 1 0 9984 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1198__136
timestamp 1680000651
transform 1 0 8640 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1198_
timestamp 1746535128
transform 1 0 9024 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1199_
timestamp 1746535184
transform -1 0 23424 0 -1 26460
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1199__128
timestamp 1680000651
transform 1 0 22080 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1200__120
timestamp 1680000651
transform -1 0 22656 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1200_
timestamp 1746535128
transform 1 0 21792 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1201__112
timestamp 1680000651
transform -1 0 21120 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1201_
timestamp 1746535128
transform 1 0 19968 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1202_
timestamp 1746535128
transform 1 0 17184 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1202__104
timestamp 1680000651
transform -1 0 18816 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1203_
timestamp 1746535128
transform 1 0 12960 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1203__96
timestamp 1680000651
transform -1 0 14304 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1204__88
timestamp 1680000651
transform 1 0 6048 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1204_
timestamp 1746535128
transform 1 0 7296 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1205_
timestamp 1746535128
transform 1 0 4992 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1205__80
timestamp 1680000651
transform -1 0 5952 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1206__72
timestamp 1680000651
transform -1 0 1920 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1206_
timestamp 1746535128
transform 1 0 1056 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1207_
timestamp 1746535128
transform 1 0 1152 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1207__64
timestamp 1680000651
transform -1 0 2016 0 1 23436
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1208__56
timestamp 1680000651
transform 1 0 6816 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1208_
timestamp 1746535128
transform 1 0 6528 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1209__167
timestamp 1680000651
transform -1 0 12096 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1209_
timestamp 1746535184
transform 1 0 10368 0 -1 20412
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1210__159
timestamp 1680000651
transform -1 0 14496 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1210_
timestamp 1746535184
transform 1 0 12480 0 1 17388
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1211_
timestamp 1746535128
transform 1 0 6432 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1211__151
timestamp 1680000651
transform 1 0 5568 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1212__140
timestamp 1680000651
transform 1 0 3456 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1212_
timestamp 1746535128
transform 1 0 4032 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1213__124
timestamp 1680000651
transform -1 0 2496 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1213_
timestamp 1746535128
transform 1 0 1632 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1214_
timestamp 1746535128
transform 1 0 1152 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1214__108
timestamp 1680000651
transform -1 0 2016 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1215__92
timestamp 1680000651
transform 1 0 10080 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1215_
timestamp 1746535128
transform -1 0 11712 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1216__76
timestamp 1680000651
transform -1 0 16416 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1216_
timestamp 1746535128
transform 1 0 14976 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1217_
timestamp 1746535128
transform 1 0 12384 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1217__60
timestamp 1680000651
transform -1 0 13536 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1218__163
timestamp 1680000651
transform -1 0 9696 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1218_
timestamp 1746535128
transform 1 0 8832 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1219_
timestamp 1746535128
transform 1 0 1248 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1219__147
timestamp 1680000651
transform 1 0 1056 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1220_
timestamp 1746535128
transform 1 0 1440 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1220__116
timestamp 1680000651
transform -1 0 2304 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1221_
timestamp 1746535128
transform 1 0 5664 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1221__84
timestamp 1680000651
transform 1 0 5472 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1222_
timestamp 1746535184
transform 1 0 864 0 -1 15876
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1222__171
timestamp 1680000651
transform -1 0 1728 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1223__132
timestamp 1680000651
transform -1 0 1824 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1223_
timestamp 1746535184
transform 1 0 960 0 -1 14364
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1224_
timestamp 1746535128
transform 1 0 3168 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1224__68
timestamp 1680000651
transform -1 0 4992 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1225_
timestamp 1746535128
transform 1 0 5568 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1225__174
timestamp 1680000651
transform -1 0 6528 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1226__175
timestamp 1680000651
transform -1 0 10464 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1226_
timestamp 1746535128
transform 1 0 9216 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1227__155
timestamp 1680000651
transform -1 0 8544 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1227_
timestamp 1746535184
transform 1 0 7104 0 1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1228_
timestamp 1746535128
transform 1 0 9312 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1228__100
timestamp 1680000651
transform -1 0 10176 0 -1 17388
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_pwm__124_
timestamp 1676382947
transform -1 0 15552 0 1 5292
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_pwm__125_
timestamp 1676382947
transform -1 0 16032 0 1 2268
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_pwm__126_
timestamp 1676382929
transform -1 0 10368 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__127_
timestamp 1676382929
transform -1 0 10080 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__128_
timestamp 1676382929
transform 1 0 7392 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__129_
timestamp 1676382929
transform -1 0 17088 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__130_
timestamp 1676382929
transform -1 0 16224 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__131_
timestamp 1676382929
transform 1 0 13344 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__132_
timestamp 1676382929
transform -1 0 13248 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__133_
timestamp 1676382929
transform -1 0 16416 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__134_
timestamp 1676382929
transform -1 0 17952 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__135_
timestamp 1676382929
transform -1 0 8352 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__136_
timestamp 1676382929
transform 1 0 10080 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__137_
timestamp 1676382929
transform 1 0 10272 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__138_
timestamp 1676382929
transform -1 0 7200 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__139_
timestamp 1676382929
transform -1 0 5952 0 1 5292
box -48 -56 336 834
use sg13g2_nor4_1  u_ppwm_u_pwm__140_
timestamp 1676643125
transform 1 0 9120 0 -1 6804
box -48 -56 624 834
use sg13g2_nor4_1  u_ppwm_u_pwm__141_
timestamp 1676643125
transform -1 0 12000 0 1 5292
box -48 -56 624 834
use sg13g2_nand4_1  u_ppwm_u_pwm__142_
timestamp 1685201930
transform 1 0 11616 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__143_
timestamp 1685175443
transform -1 0 11904 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__144_
timestamp 1683973020
transform -1 0 9888 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__145_
timestamp 1685175443
transform -1 0 11808 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__146_
timestamp 1683973020
transform -1 0 10272 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__147_
timestamp 1685175443
transform -1 0 15168 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__148_
timestamp 1683973020
transform -1 0 10752 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__149_
timestamp 1685175443
transform -1 0 14208 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__150_
timestamp 1683973020
transform -1 0 9696 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__151_
timestamp 1685175443
transform -1 0 14880 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__152_
timestamp 1683973020
transform -1 0 14688 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__153_
timestamp 1685175443
transform -1 0 14400 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__154_
timestamp 1683973020
transform 1 0 15168 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__155_
timestamp 1685175443
transform -1 0 13728 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__156_
timestamp 1683973020
transform 1 0 12768 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__157_
timestamp 1685175443
transform -1 0 11424 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__158_
timestamp 1683973020
transform -1 0 10464 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__159_
timestamp 1685175443
transform 1 0 15168 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__160_
timestamp 1683973020
transform -1 0 16704 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__161_
timestamp 1685175443
transform -1 0 15072 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__162_
timestamp 1683973020
transform 1 0 16128 0 -1 3780
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_pwm__163_
timestamp 1676901763
transform -1 0 6432 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__164_
timestamp 1685175443
transform -1 0 6048 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_pwm__165_
timestamp 1676627187
transform -1 0 6432 0 1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__166_
timestamp 1685175443
transform -1 0 5568 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__167_
timestamp 1683973020
transform 1 0 4608 0 -1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__168_
timestamp 1683973020
transform -1 0 6144 0 -1 5292
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_pwm__169_
timestamp 1676985977
transform -1 0 7968 0 -1 6804
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_pwm__170_
timestamp 1676639442
transform 1 0 4320 0 1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_pwm__171_
timestamp 1677516600
transform -1 0 7680 0 1 5292
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_pwm__172_
timestamp 1676627187
transform 1 0 5952 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__173_
timestamp 1683973020
transform -1 0 6816 0 1 2268
box -48 -56 528 834
use sg13g2_and3_1  u_ppwm_u_pwm__174_
timestamp 1676971669
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_nor3_1  u_ppwm_u_pwm__175_
timestamp 1676639442
transform 1 0 4128 0 -1 5292
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_pwm__176_
timestamp 1676985977
transform 1 0 7008 0 -1 5292
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__177_
timestamp 1685175443
transform 1 0 7680 0 1 5292
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_pwm__178_
timestamp 1676627187
transform 1 0 8352 0 1 2268
box -48 -56 432 834
use sg13g2_or2_1  u_ppwm_u_pwm__179_
timestamp 1684236171
transform 1 0 9024 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__180_
timestamp 1676557249
transform 1 0 7968 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  u_ppwm_u_pwm__181_
timestamp 1676971669
transform 1 0 9120 0 -1 3780
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_pwm__182_
timestamp 1683988354
transform 1 0 9312 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__183_
timestamp 1676557249
transform -1 0 10752 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__184_
timestamp 1683973020
transform -1 0 10080 0 -1 2268
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_pwm__185_
timestamp 1684236171
transform -1 0 11616 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__186_
timestamp 1676557249
transform -1 0 11328 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__187_
timestamp 1683973020
transform 1 0 12192 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__188_
timestamp 1685175443
transform -1 0 12096 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__189_
timestamp 1683973020
transform 1 0 13056 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_pwm__190_
timestamp 1683988354
transform -1 0 10752 0 -1 6804
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_pwm__191_
timestamp 1685201930
transform 1 0 14400 0 -1 5292
box -48 -56 624 834
use sg13g2_nand4_1  u_ppwm_u_pwm__192_
timestamp 1685201930
transform 1 0 9696 0 -1 6804
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_pwm__193_
timestamp 1676639442
transform 1 0 10464 0 1 5292
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__194_
timestamp 1676567195
transform 1 0 10176 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__195_
timestamp 1685181386
transform 1 0 8160 0 -1 6804
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__196_
timestamp 1676567195
transform -1 0 9120 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__197_
timestamp 1685181386
transform 1 0 7776 0 1 6804
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__198_
timestamp 1683973020
transform 1 0 8160 0 1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_pwm__199_
timestamp 1685197497
transform 1 0 9024 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__200_
timestamp 1676567195
transform 1 0 8256 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__201_
timestamp 1685181386
transform -1 0 8160 0 -1 8316
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_pwm__202_
timestamp 1685197497
transform 1 0 8736 0 1 6804
box -48 -56 816 834
use sg13g2_a21o_1  u_ppwm_u_pwm__203_
timestamp 1677175127
transform -1 0 10176 0 1 6804
box -48 -56 720 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__204_
timestamp 1676567195
transform 1 0 12096 0 1 5292
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__205_
timestamp 1676567195
transform -1 0 12768 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__206_
timestamp 1676557249
transform 1 0 11040 0 1 5292
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__207_
timestamp 1676567195
transform 1 0 11232 0 1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__208_
timestamp 1676567195
transform 1 0 11712 0 1 6804
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_pwm__209_
timestamp 1676627187
transform 1 0 13920 0 1 5292
box -48 -56 432 834
use sg13g2_nand4_1  u_ppwm_u_pwm__210_
timestamp 1685201930
transform 1 0 12768 0 -1 6804
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_pwm__211_
timestamp 1676627187
transform -1 0 14016 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__212_
timestamp 1685181386
transform 1 0 14688 0 1 6804
box -54 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_pwm__213_
timestamp 1677175127
transform 1 0 14496 0 -1 6804
box -48 -56 720 834
use sg13g2_nor2_1  u_ppwm_u_pwm__214_
timestamp 1676627187
transform 1 0 13536 0 1 5292
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_pwm__215_
timestamp 1676643125
transform 1 0 14112 0 1 6804
box -48 -56 624 834
use sg13g2_and2_1  u_ppwm_u_pwm__216_
timestamp 1676901763
transform 1 0 13440 0 1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_pwm__217_
timestamp 1685197497
transform 1 0 13632 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_pwm__218_
timestamp 1676557249
transform 1 0 14016 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_pwm__219_
timestamp 1676557249
transform -1 0 16416 0 1 2268
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_pwm__220_
timestamp 1685173987
transform 1 0 15360 0 -1 3780
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_pwm__221_
timestamp 1676557249
transform -1 0 16800 0 1 2268
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__222_
timestamp 1685181386
transform -1 0 16128 0 1 5292
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__223_
timestamp 1683973020
transform 1 0 14880 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__224_
timestamp 1685175443
transform 1 0 14688 0 1 3780
box -48 -56 538 834
use sg13g2_and2_1  u_ppwm_u_pwm__225_
timestamp 1676901763
transform 1 0 14400 0 -1 3780
box -48 -56 528 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__226_
timestamp 1746535128
transform 1 0 5952 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__226__190
timestamp 1680000651
transform -1 0 6912 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__227__187
timestamp 1680000651
transform 1 0 7200 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__227_
timestamp 1746535128
transform -1 0 9792 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__228_
timestamp 1746535128
transform 1 0 6624 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__228__185
timestamp 1680000651
transform 1 0 6528 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__229_
timestamp 1746535128
transform 1 0 5472 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__229__183
timestamp 1680000651
transform -1 0 6336 0 1 9828
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__230__181
timestamp 1680000651
transform -1 0 16800 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__230_
timestamp 1746535128
transform 1 0 14880 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__231_
timestamp 1746535128
transform 1 0 15648 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__231__179
timestamp 1680000651
transform 1 0 15168 0 1 6804
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__232__177
timestamp 1680000651
transform -1 0 11712 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__232_
timestamp 1746535128
transform 1 0 10944 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__233_
timestamp 1746535128
transform -1 0 12480 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__233__197
timestamp 1680000651
transform -1 0 12192 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__234__195
timestamp 1680000651
transform -1 0 17760 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__234_
timestamp 1746535128
transform 1 0 16896 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__235_
timestamp 1746535128
transform 1 0 16704 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__235__193
timestamp 1680000651
transform -1 0 17568 0 1 2268
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__236__191
timestamp 1680000651
transform -1 0 4224 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__236_
timestamp 1746535184
transform 1 0 3360 0 1 8316
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__237__189
timestamp 1680000651
transform -1 0 3168 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__237_
timestamp 1746535184
transform 1 0 2304 0 1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__238_
timestamp 1746535184
transform 1 0 3648 0 -1 6804
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__238__186
timestamp 1680000651
transform 1 0 3936 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__239_
timestamp 1746535128
transform 1 0 5376 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__239__182
timestamp 1680000651
transform -1 0 7200 0 1 2268
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__240__178
timestamp 1680000651
transform -1 0 4128 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__240_
timestamp 1746535184
transform 1 0 3264 0 1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__241_
timestamp 1746535184
transform 1 0 8640 0 -1 5292
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__241__196
timestamp 1680000651
transform 1 0 8928 0 1 3780
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__242__192
timestamp 1680000651
transform 1 0 10752 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__242_
timestamp 1746535184
transform 1 0 10656 0 -1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__243_
timestamp 1746535184
transform 1 0 9504 0 1 2268
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__243__188
timestamp 1680000651
transform -1 0 10464 0 -1 2268
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__244__180
timestamp 1680000651
transform -1 0 13056 0 -1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__244_
timestamp 1746535128
transform 1 0 12096 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__245_
timestamp 1746535128
transform 1 0 12768 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__245__194
timestamp 1680000651
transform -1 0 13632 0 -1 3780
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__246__184
timestamp 1680000651
transform -1 0 18720 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__246_
timestamp 1746535184
transform 1 0 17856 0 1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__247_
timestamp 1746535128
transform 1 0 14976 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__247__176
timestamp 1680000651
transform -1 0 15840 0 1 756
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel via3 78 36708 78 36708 0 clk
rlabel metal2 30576 28140 30576 28140 0 clknet_0_clk
rlabel metal3 9216 7140 9216 7140 0 clknet_4_0_0_clk
rlabel metal2 39120 16800 39120 16800 0 clknet_4_10_0_clk
rlabel metal2 40320 22428 40320 22428 0 clknet_4_11_0_clk
rlabel metal2 30048 31290 30048 31290 0 clknet_4_12_0_clk
rlabel metal2 30240 33810 30240 33810 0 clknet_4_13_0_clk
rlabel metal2 44160 30660 44160 30660 0 clknet_4_14_0_clk
rlabel metal2 40992 33012 40992 33012 0 clknet_4_15_0_clk
rlabel metal2 11424 13650 11424 13650 0 clknet_4_1_0_clk
rlabel metal3 18864 6468 18864 6468 0 clknet_4_2_0_clk
rlabel metal2 17184 14028 17184 14028 0 clknet_4_3_0_clk
rlabel metal3 5904 21588 5904 21588 0 clknet_4_4_0_clk
rlabel metal2 6192 31332 6192 31332 0 clknet_4_5_0_clk
rlabel metal3 14160 25284 14160 25284 0 clknet_4_6_0_clk
rlabel metal2 14976 31080 14976 31080 0 clknet_4_7_0_clk
rlabel metal3 31584 11676 31584 11676 0 clknet_4_8_0_clk
rlabel metal2 30384 22260 30384 22260 0 clknet_4_9_0_clk
rlabel metal3 5664 4116 5664 4116 0 clknet_5_0__leaf_clk
rlabel metal2 2496 27552 2496 27552 0 clknet_5_10__leaf_clk
rlabel metal2 4896 34188 4896 34188 0 clknet_5_11__leaf_clk
rlabel metal3 11184 29148 11184 29148 0 clknet_5_12__leaf_clk
rlabel metal2 11808 20076 11808 20076 0 clknet_5_13__leaf_clk
rlabel metal3 13488 33684 13488 33684 0 clknet_5_14__leaf_clk
rlabel metal3 16800 34356 16800 34356 0 clknet_5_15__leaf_clk
rlabel metal3 28128 1932 28128 1932 0 clknet_5_16__leaf_clk
rlabel metal3 31824 19236 31824 19236 0 clknet_5_17__leaf_clk
rlabel metal2 18624 21588 18624 21588 0 clknet_5_18__leaf_clk
rlabel metal2 34032 24612 34032 24612 0 clknet_5_19__leaf_clk
rlabel metal2 11952 1932 11952 1932 0 clknet_5_1__leaf_clk
rlabel metal2 37872 8652 37872 8652 0 clknet_5_20__leaf_clk
rlabel metal2 38352 21588 38352 21588 0 clknet_5_21__leaf_clk
rlabel metal3 36864 23016 36864 23016 0 clknet_5_22__leaf_clk
rlabel metal2 43584 22680 43584 22680 0 clknet_5_23__leaf_clk
rlabel metal2 23904 30450 23904 30450 0 clknet_5_24__leaf_clk
rlabel metal2 29472 31962 29472 31962 0 clknet_5_25__leaf_clk
rlabel metal2 20064 34776 20064 34776 0 clknet_5_26__leaf_clk
rlabel metal3 31296 32844 31296 32844 0 clknet_5_27__leaf_clk
rlabel metal2 45936 26628 45936 26628 0 clknet_5_28__leaf_clk
rlabel metal2 43056 26796 43056 26796 0 clknet_5_29__leaf_clk
rlabel metal2 2256 14028 2256 14028 0 clknet_5_2__leaf_clk
rlabel metal2 36288 31752 36288 31752 0 clknet_5_30__leaf_clk
rlabel metal2 40608 30576 40608 30576 0 clknet_5_31__leaf_clk
rlabel metal2 11808 14280 11808 14280 0 clknet_5_3__leaf_clk
rlabel metal2 16176 1932 16176 1932 0 clknet_5_4__leaf_clk
rlabel metal3 18672 5628 18672 5628 0 clknet_5_5__leaf_clk
rlabel metal2 16416 14238 16416 14238 0 clknet_5_6__leaf_clk
rlabel metal2 19200 11760 19200 11760 0 clknet_5_7__leaf_clk
rlabel metal2 2496 23856 2496 23856 0 clknet_5_8__leaf_clk
rlabel metal2 7008 18312 7008 18312 0 clknet_5_9__leaf_clk
rlabel metal2 864 19320 864 19320 0 net1
rlabel metal3 366 21588 366 21588 0 net10
rlabel metal2 9888 16548 9888 16548 0 net100
rlabel metal3 45120 30492 45120 30492 0 net101
rlabel metal2 14736 32004 14736 32004 0 net102
rlabel metal2 45312 25620 45312 25620 0 net103
rlabel metal3 18096 22428 18096 22428 0 net104
rlabel metal2 47136 22596 47136 22596 0 net105
rlabel metal2 15312 29820 15312 29820 0 net106
rlabel metal2 37344 22008 37344 22008 0 net107
rlabel metal2 1680 21420 1680 21420 0 net108
rlabel metal2 36960 27132 36960 27132 0 net109
rlabel metal3 366 8988 366 8988 0 net11
rlabel metal2 11424 28812 11424 28812 0 net110
rlabel metal2 39408 32004 39408 32004 0 net111
rlabel metal2 20832 24486 20832 24486 0 net112
rlabel metal2 44976 33012 44976 33012 0 net113
rlabel metal3 1344 29988 1344 29988 0 net114
rlabel metal2 47904 32592 47904 32592 0 net115
rlabel metal2 2016 18564 2016 18564 0 net116
rlabel metal2 50880 28140 50880 28140 0 net117
rlabel metal2 5184 32592 5184 32592 0 net118
rlabel metal2 49872 24612 49872 24612 0 net119
rlabel metal3 366 9828 366 9828 0 net12
rlabel metal2 22368 28056 22368 28056 0 net120
rlabel metal2 39600 20748 39600 20748 0 net121
rlabel metal2 7200 34692 7200 34692 0 net122
rlabel metal2 38784 23856 38784 23856 0 net123
rlabel metal2 2208 21084 2208 21084 0 net124
rlabel metal2 41088 22848 41088 22848 0 net125
rlabel metal2 9984 36204 9984 36204 0 net126
rlabel metal2 51264 28056 51264 28056 0 net127
rlabel metal3 22656 26124 22656 26124 0 net128
rlabel metal2 46464 27132 46464 27132 0 net129
rlabel metal3 366 10668 366 10668 0 net13
rlabel metal3 13536 36540 13536 36540 0 net130
rlabel metal3 48960 25956 48960 25956 0 net131
rlabel metal2 1488 14028 1488 14028 0 net132
rlabel metal2 50784 23520 50784 23520 0 net133
rlabel metal2 16320 36204 16320 36204 0 net134
rlabel metal2 46176 22554 46176 22554 0 net135
rlabel metal2 8928 25788 8928 25788 0 net136
rlabel metal2 34992 21420 34992 21420 0 net137
rlabel metal3 12912 35028 12912 35028 0 net138
rlabel metal2 42624 20454 42624 20454 0 net139
rlabel metal3 366 11508 366 11508 0 net14
rlabel metal3 4128 19404 4128 19404 0 net140
rlabel metal2 50208 30408 50208 30408 0 net141
rlabel metal2 1728 32592 1728 32592 0 net142
rlabel metal3 50640 30492 50640 30492 0 net143
rlabel metal3 10272 24444 10272 24444 0 net144
rlabel metal2 42240 27132 42240 27132 0 net145
rlabel metal2 2592 34104 2592 34104 0 net146
rlabel metal2 1392 17892 1392 17892 0 net147
rlabel metal2 4512 34692 4512 34692 0 net148
rlabel metal2 15744 22764 15744 22764 0 net149
rlabel metal3 366 12348 366 12348 0 net15
rlabel metal3 10080 34524 10080 34524 0 net150
rlabel metal3 6384 19404 6384 19404 0 net151
rlabel metal3 16800 35028 16800 35028 0 net152
rlabel metal2 17904 23940 17904 23940 0 net153
rlabel metal2 19584 36036 19584 36036 0 net154
rlabel metal2 7872 13188 7872 13188 0 net155
rlabel metal2 22464 34692 22464 34692 0 net156
rlabel metal2 21408 24864 21408 24864 0 net157
rlabel metal2 24960 36204 24960 36204 0 net158
rlabel metal2 12960 18060 12960 18060 0 net159
rlabel metal3 366 13188 366 13188 0 net16
rlabel metal2 29664 36582 29664 36582 0 net160
rlabel metal2 22368 29568 22368 29568 0 net161
rlabel metal2 34848 33516 34848 33516 0 net162
rlabel metal2 9408 18060 9408 18060 0 net163
rlabel metal2 38400 32424 38400 32424 0 net164
rlabel metal3 17472 29148 17472 29148 0 net165
rlabel metal2 39168 36582 39168 36582 0 net166
rlabel metal2 11808 20832 11808 20832 0 net167
rlabel metal2 37632 36204 37632 36204 0 net168
rlabel metal2 10080 27300 10080 27300 0 net169
rlabel metal3 510 14028 510 14028 0 net17
rlabel metal2 23856 36036 23856 36036 0 net170
rlabel metal2 1392 15540 1392 15540 0 net171
rlabel metal3 27648 37548 27648 37548 0 net172
rlabel metal2 42336 24108 42336 24108 0 net173
rlabel metal2 6240 13188 6240 13188 0 net174
rlabel metal2 10176 15204 10176 15204 0 net175
rlabel metal2 15504 1260 15504 1260 0 net176
rlabel metal2 11424 8232 11424 8232 0 net177
rlabel metal2 3792 4116 3792 4116 0 net178
rlabel metal2 15456 7056 15456 7056 0 net179
rlabel metal3 366 14868 366 14868 0 net18
rlabel metal2 12768 3696 12768 3696 0 net180
rlabel metal2 16512 7644 16512 7644 0 net181
rlabel metal3 6384 2772 6384 2772 0 net182
rlabel metal2 6048 9912 6048 9912 0 net183
rlabel metal2 18336 5754 18336 5754 0 net184
rlabel metal2 6816 10080 6816 10080 0 net185
rlabel metal2 4176 6468 4176 6468 0 net186
rlabel metal3 8400 11004 8400 11004 0 net187
rlabel metal2 10128 1764 10128 1764 0 net188
rlabel metal2 2832 7140 2832 7140 0 net189
rlabel metal3 366 3108 366 3108 0 net19
rlabel metal2 6624 12012 6624 12012 0 net190
rlabel metal2 3888 8652 3888 8652 0 net191
rlabel metal2 11040 1932 11040 1932 0 net192
rlabel metal2 17280 3108 17280 3108 0 net193
rlabel metal2 13344 2940 13344 2940 0 net194
rlabel metal2 17424 5796 17424 5796 0 net195
rlabel metal2 9168 4956 9168 4956 0 net196
rlabel metal2 11904 10500 11904 10500 0 net197
rlabel metal2 38208 9996 38208 9996 0 net198
rlabel metal2 37344 10164 37344 10164 0 net199
rlabel metal2 864 2184 864 2184 0 net2
rlabel metal3 366 3948 366 3948 0 net20
rlabel metal3 7872 12516 7872 12516 0 net200
rlabel metal3 6864 11676 6864 11676 0 net201
rlabel metal2 28032 4872 28032 4872 0 net202
rlabel metal2 27504 2604 27504 2604 0 net203
rlabel metal2 36768 13146 36768 13146 0 net204
rlabel metal2 36960 12936 36960 12936 0 net205
rlabel metal2 11664 18732 11664 18732 0 net206
rlabel metal2 12480 18942 12480 18942 0 net207
rlabel metal3 4560 31332 4560 31332 0 net208
rlabel metal2 4992 32508 4992 32508 0 net209
rlabel metal3 366 4788 366 4788 0 net21
rlabel metal3 13248 23940 13248 23940 0 net210
rlabel metal2 13680 23184 13680 23184 0 net211
rlabel metal3 4272 25284 4272 25284 0 net212
rlabel metal2 5136 24696 5136 24696 0 net213
rlabel metal3 17760 35196 17760 35196 0 net214
rlabel metal2 18864 35280 18864 35280 0 net215
rlabel metal2 27360 32844 27360 32844 0 net216
rlabel metal2 30432 33894 30432 33894 0 net217
rlabel metal2 10368 9744 10368 9744 0 net218
rlabel metal2 9840 11088 9840 11088 0 net219
rlabel metal3 366 5628 366 5628 0 net22
rlabel metal2 13344 7980 13344 7980 0 net220
rlabel metal2 11040 8946 11040 8946 0 net221
rlabel metal2 16320 5964 16320 5964 0 net222
rlabel metal3 16032 6552 16032 6552 0 net223
rlabel metal3 12384 34944 12384 34944 0 net224
rlabel metal2 3072 27678 3072 27678 0 net225
rlabel metal2 8448 29442 8448 29442 0 net226
rlabel metal2 25728 4200 25728 4200 0 net227
rlabel metal2 24384 1932 24384 1932 0 net228
rlabel metal3 19008 32172 19008 32172 0 net229
rlabel metal3 366 6468 366 6468 0 net23
rlabel metal2 19968 30912 19968 30912 0 net230
rlabel metal2 19392 28392 19392 28392 0 net231
rlabel metal2 19104 29148 19104 29148 0 net232
rlabel metal2 5952 21252 5952 21252 0 net233
rlabel metal2 4176 20160 4176 20160 0 net234
rlabel metal2 33888 27384 33888 27384 0 net235
rlabel metal2 32832 24780 32832 24780 0 net236
rlabel metal3 39552 33684 39552 33684 0 net237
rlabel metal2 39168 35868 39168 35868 0 net238
rlabel metal2 8064 30450 8064 30450 0 net239
rlabel metal3 366 7308 366 7308 0 net24
rlabel metal2 8928 30492 8928 30492 0 net240
rlabel metal3 45216 27678 45216 27678 0 net241
rlabel metal2 48672 25200 48672 25200 0 net242
rlabel metal2 7680 32424 7680 32424 0 net243
rlabel metal2 6288 34356 6288 34356 0 net244
rlabel metal2 19200 22386 19200 22386 0 net245
rlabel metal2 17376 23394 17376 23394 0 net246
rlabel metal2 26016 35826 26016 35826 0 net247
rlabel metal2 27264 35574 27264 35574 0 net248
rlabel metal2 13344 10164 13344 10164 0 net249
rlabel metal3 318 8148 318 8148 0 net25
rlabel metal2 12384 10458 12384 10458 0 net250
rlabel metal3 22128 3192 22128 3192 0 net251
rlabel metal2 20544 3444 20544 3444 0 net252
rlabel metal3 7104 34944 7104 34944 0 net253
rlabel metal2 36048 24612 36048 24612 0 net254
rlabel metal3 36384 25284 36384 25284 0 net255
rlabel metal3 27504 36708 27504 36708 0 net256
rlabel metal2 29712 35868 29712 35868 0 net257
rlabel metal2 19152 24780 19152 24780 0 net258
rlabel metal2 21792 25578 21792 25578 0 net259
rlabel metal2 18000 8820 18000 8820 0 net26
rlabel metal2 39168 35322 39168 35322 0 net260
rlabel metal2 38112 35868 38112 35868 0 net261
rlabel metal2 6816 23562 6816 23562 0 net262
rlabel metal2 7296 23688 7296 23688 0 net263
rlabel metal2 16128 4998 16128 4998 0 net264
rlabel metal2 16992 3990 16992 3990 0 net265
rlabel metal2 12384 25116 12384 25116 0 net266
rlabel metal2 10080 23898 10080 23898 0 net267
rlabel metal2 26592 6678 26592 6678 0 net268
rlabel metal2 20640 5376 20640 5376 0 net269
rlabel metal2 18624 19908 18624 19908 0 net27
rlabel metal2 12288 35616 12288 35616 0 net270
rlabel metal2 12864 35868 12864 35868 0 net271
rlabel metal3 25584 31164 25584 31164 0 net272
rlabel metal2 23328 33138 23328 33138 0 net273
rlabel metal2 20640 28224 20640 28224 0 net274
rlabel metal2 23328 26166 23328 26166 0 net275
rlabel metal3 15744 32172 15744 32172 0 net276
rlabel metal2 14976 30114 14976 30114 0 net277
rlabel metal3 13488 32676 13488 32676 0 net278
rlabel metal2 14880 33138 14880 33138 0 net279
rlabel metal2 18720 9744 18720 9744 0 net28
rlabel metal3 27408 33012 27408 33012 0 net280
rlabel metal2 28992 31626 28992 31626 0 net281
rlabel metal2 20928 34692 20928 34692 0 net282
rlabel metal2 21408 34650 21408 34650 0 net283
rlabel metal2 21216 27048 21216 27048 0 net284
rlabel metal3 22032 29232 22032 29232 0 net285
rlabel metal2 2400 23814 2400 23814 0 net286
rlabel metal3 3840 31920 3840 31920 0 net287
rlabel metal2 2016 33306 2016 33306 0 net288
rlabel metal2 30720 28644 30720 28644 0 net289
rlabel metal2 27264 18228 27264 18228 0 net29
rlabel metal2 28896 30114 28896 30114 0 net290
rlabel metal2 26496 1176 26496 1176 0 net291
rlabel metal3 24096 2688 24096 2688 0 net292
rlabel metal2 5952 30366 5952 30366 0 net293
rlabel metal2 8448 32508 8448 32508 0 net294
rlabel metal2 19968 22554 19968 22554 0 net295
rlabel metal2 20064 23814 20064 23814 0 net296
rlabel metal2 36576 33600 36576 33600 0 net297
rlabel metal2 41808 32844 41808 32844 0 net298
rlabel metal3 40368 29988 40368 29988 0 net299
rlabel metal3 366 15708 366 15708 0 net3
rlabel metal2 22176 11508 22176 11508 0 net30
rlabel metal2 42240 30954 42240 30954 0 net300
rlabel metal2 43776 31080 43776 31080 0 net301
rlabel metal2 44736 32466 44736 32466 0 net302
rlabel metal3 10560 34356 10560 34356 0 net303
rlabel metal2 17856 7812 17856 7812 0 net304
rlabel metal2 15072 8064 15072 8064 0 net305
rlabel metal3 35952 33600 35952 33600 0 net306
rlabel metal2 29280 18354 29280 18354 0 net307
rlabel metal2 35616 18144 35616 18144 0 net308
rlabel metal2 17568 14448 17568 14448 0 net309
rlabel metal2 40320 16716 40320 16716 0 net31
rlabel metal2 18432 12474 18432 12474 0 net310
rlabel metal2 17184 11424 17184 11424 0 net311
rlabel metal2 34944 18018 34944 18018 0 net312
rlabel metal2 16992 11508 16992 11508 0 net313
rlabel metal2 32448 17430 32448 17430 0 net314
rlabel metal3 17280 13230 17280 13230 0 net315
rlabel metal2 17664 14868 17664 14868 0 net316
rlabel metal2 31824 18564 31824 18564 0 net317
rlabel metal2 14016 14028 14016 14028 0 net318
rlabel metal3 15552 14700 15552 14700 0 net319
rlabel metal2 21216 11592 21216 11592 0 net32
rlabel metal3 26112 18564 26112 18564 0 net320
rlabel metal2 35904 15666 35904 15666 0 net321
rlabel metal2 29952 16254 29952 16254 0 net322
rlabel metal2 18912 16296 18912 16296 0 net323
rlabel metal2 26112 18144 26112 18144 0 net324
rlabel metal2 30624 15666 30624 15666 0 net325
rlabel metal2 24144 20076 24144 20076 0 net326
rlabel metal2 29760 15162 29760 15162 0 net327
rlabel metal2 11712 8736 11712 8736 0 net328
rlabel metal2 13536 9282 13536 9282 0 net329
rlabel metal2 18144 18060 18144 18060 0 net33
rlabel metal2 16320 4830 16320 4830 0 net330
rlabel metal2 35616 9492 35616 9492 0 net331
rlabel via2 39360 26121 39360 26121 0 net332
rlabel metal2 17952 25326 17952 25326 0 net333
rlabel metal2 14208 27006 14208 27006 0 net334
rlabel metal2 36672 24612 36672 24612 0 net335
rlabel metal3 21648 1932 21648 1932 0 net336
rlabel metal3 7296 4074 7296 4074 0 net337
rlabel metal2 7872 19194 7872 19194 0 net338
rlabel via2 12000 18648 12000 18648 0 net339
rlabel metal2 19776 8652 19776 8652 0 net34
rlabel metal2 4128 22218 4128 22218 0 net340
rlabel metal2 3648 25242 3648 25242 0 net341
rlabel metal3 12192 26754 12192 26754 0 net342
rlabel metal3 9168 20076 9168 20076 0 net343
rlabel metal2 16224 23646 16224 23646 0 net344
rlabel metal2 18336 21924 18336 21924 0 net345
rlabel metal2 4032 31416 4032 31416 0 net346
rlabel metal2 7584 29904 7584 29904 0 net347
rlabel metal2 8256 32508 8256 32508 0 net348
rlabel metal2 9216 34104 9216 34104 0 net349
rlabel metal2 34944 20916 34944 20916 0 net35
rlabel metal2 12384 34272 12384 34272 0 net350
rlabel metal3 14304 35070 14304 35070 0 net351
rlabel metal3 10800 32844 10800 32844 0 net352
rlabel metal2 19536 28308 19536 28308 0 net353
rlabel metal2 19008 26754 19008 26754 0 net354
rlabel metal2 15936 32088 15936 32088 0 net355
rlabel metal2 15456 32382 15456 32382 0 net356
rlabel metal2 19200 31080 19200 31080 0 net357
rlabel metal2 35040 23016 35040 23016 0 net358
rlabel metal3 35328 23604 35328 23604 0 net359
rlabel metal2 17568 16968 17568 16968 0 net36
rlabel metal2 46224 23772 46224 23772 0 net360
rlabel metal2 45696 26250 45696 26250 0 net361
rlabel metal2 41376 22890 41376 22890 0 net362
rlabel metal2 40416 22218 40416 22218 0 net363
rlabel metal2 30624 28602 30624 28602 0 net364
rlabel metal2 35616 29022 35616 29022 0 net365
rlabel metal2 29184 32886 29184 32886 0 net366
rlabel metal2 29664 35112 29664 35112 0 net367
rlabel metal3 35616 35196 35616 35196 0 net368
rlabel metal3 32352 34356 32352 34356 0 net369
rlabel metal3 23040 19236 23040 19236 0 net37
rlabel metal2 46176 27762 46176 27762 0 net370
rlabel metal2 45120 27468 45120 27468 0 net371
rlabel metal2 46272 30996 46272 30996 0 net372
rlabel metal2 41856 34062 41856 34062 0 net373
rlabel metal3 37236 33684 37236 33684 0 net374
rlabel metal2 32928 30198 32928 30198 0 net375
rlabel metal3 35520 21588 35520 21588 0 net376
rlabel metal3 21456 18900 21456 18900 0 net377
rlabel metal2 29184 13902 29184 13902 0 net378
rlabel metal2 36480 18228 36480 18228 0 net379
rlabel metal2 29040 20916 29040 20916 0 net38
rlabel metal3 36480 15162 36480 15162 0 net380
rlabel metal2 36288 14616 36288 14616 0 net381
rlabel metal2 34368 16044 34368 16044 0 net382
rlabel metal3 29760 16002 29760 16002 0 net383
rlabel metal2 25344 16548 25344 16548 0 net384
rlabel metal2 25056 15078 25056 15078 0 net385
rlabel metal2 17952 14784 17952 14784 0 net386
rlabel metal2 19776 12474 19776 12474 0 net387
rlabel metal4 11808 11634 11808 11634 0 net388
rlabel metal2 13824 13104 13824 13104 0 net389
rlabel metal2 39552 14280 39552 14280 0 net39
rlabel metal2 12672 10626 12672 10626 0 net390
rlabel metal3 18624 11508 18624 11508 0 net391
rlabel metal2 15216 11676 15216 11676 0 net392
rlabel metal2 29088 8106 29088 8106 0 net393
rlabel metal2 20064 13986 20064 13986 0 net394
rlabel metal2 29376 7728 29376 7728 0 net395
rlabel metal2 19584 13986 19584 13986 0 net396
rlabel metal2 25632 8526 25632 8526 0 net397
rlabel metal2 18576 16212 18576 16212 0 net398
rlabel metal2 25248 7098 25248 7098 0 net399
rlabel metal3 366 16548 366 16548 0 net4
rlabel metal2 28032 21462 28032 21462 0 net40
rlabel metal2 30912 23310 30912 23310 0 net400
rlabel metal2 30336 27426 30336 27426 0 net401
rlabel metal2 25728 28308 25728 28308 0 net402
rlabel metal2 17568 26586 17568 26586 0 net403
rlabel metal3 12384 26124 12384 26124 0 net404
rlabel metal2 14208 30114 14208 30114 0 net405
rlabel metal3 17088 30576 17088 30576 0 net406
rlabel metal2 29280 23604 29280 23604 0 net407
rlabel metal2 38963 25236 38963 25236 0 net408
rlabel metal2 29472 26628 29472 26628 0 net409
rlabel metal2 13056 15960 13056 15960 0 net41
rlabel metal2 12384 21714 12384 21714 0 net410
rlabel metal2 6912 31038 6912 31038 0 net411
rlabel metal2 17568 25620 17568 25620 0 net412
rlabel metal2 19200 33264 19200 33264 0 net413
rlabel metal2 12192 29946 12192 29946 0 net414
rlabel metal2 36192 23520 36192 23520 0 net415
rlabel metal2 31008 33894 31008 33894 0 net416
rlabel metal2 40704 26544 40704 26544 0 net417
rlabel metal3 39456 28434 39456 28434 0 net418
rlabel metal2 41856 30450 41856 30450 0 net419
rlabel metal2 25584 25284 25584 25284 0 net42
rlabel metal2 40128 27216 40128 27216 0 net420
rlabel metal3 37584 27636 37584 27636 0 net421
rlabel metal3 13008 16212 13008 16212 0 net422
rlabel metal2 12672 17346 12672 17346 0 net423
rlabel metal2 13920 9576 13920 9576 0 net424
rlabel metal2 14688 8652 14688 8652 0 net425
rlabel metal2 15744 13482 15744 13482 0 net426
rlabel metal2 15360 16044 15360 16044 0 net427
rlabel metal2 4032 25494 4032 25494 0 net428
rlabel metal2 6240 19698 6240 19698 0 net429
rlabel metal2 21600 22008 21600 22008 0 net43
rlabel metal2 6432 33726 6432 33726 0 net430
rlabel metal2 12864 31416 12864 31416 0 net431
rlabel metal2 11904 31080 11904 31080 0 net432
rlabel metal2 14208 24780 14208 24780 0 net433
rlabel metal2 17088 35028 17088 35028 0 net434
rlabel metal3 19872 30660 19872 30660 0 net435
rlabel metal2 12672 27510 12672 27510 0 net436
rlabel metal2 15936 17682 15936 17682 0 net437
rlabel metal2 29568 4788 29568 4788 0 net438
rlabel metal3 23250 1932 23250 1932 0 net439
rlabel metal2 29856 25032 29856 25032 0 net44
rlabel metal3 32112 12264 32112 12264 0 net440
rlabel metal2 32160 17472 32160 17472 0 net441
rlabel metal4 31968 17052 31968 17052 0 net442
rlabel metal2 35232 23520 35232 23520 0 net443
rlabel metal2 25536 34188 25536 34188 0 net444
rlabel metal2 33888 31248 33888 31248 0 net445
rlabel metal2 34176 25494 34176 25494 0 net446
rlabel metal2 45312 27006 45312 27006 0 net447
rlabel metal2 38592 22470 38592 22470 0 net448
rlabel metal2 37344 28476 37344 28476 0 net449
rlabel metal2 22896 13188 22896 13188 0 net45
rlabel metal2 47904 31080 47904 31080 0 net450
rlabel metal3 38880 23856 38880 23856 0 net451
rlabel metal2 33312 23772 33312 23772 0 net452
rlabel metal3 14448 31332 14448 31332 0 net453
rlabel metal2 10944 29820 10944 29820 0 net454
rlabel metal2 33120 35154 33120 35154 0 net455
rlabel metal2 32736 36330 32736 36330 0 net456
rlabel metal2 34752 35280 34752 35280 0 net457
rlabel metal2 21600 26208 21600 26208 0 net458
rlabel metal2 35520 30618 35520 30618 0 net459
rlabel metal3 33840 13860 33840 13860 0 net46
rlabel metal2 33216 30114 33216 30114 0 net460
rlabel metal2 30240 3864 30240 3864 0 net461
rlabel metal3 27600 3444 27600 3444 0 net462
rlabel metal2 29376 3864 29376 3864 0 net463
rlabel metal3 44160 23520 44160 23520 0 net464
rlabel metal2 51648 27930 51648 27930 0 net465
rlabel metal2 31680 30912 31680 30912 0 net466
rlabel metal2 14112 35028 14112 35028 0 net467
rlabel metal2 15408 35868 15408 35868 0 net468
rlabel metal2 41088 23562 41088 23562 0 net469
rlabel metal2 10080 13692 10080 13692 0 net47
rlabel metal2 42336 22470 42336 22470 0 net470
rlabel metal2 9696 20706 9696 20706 0 net471
rlabel metal2 6528 21588 6528 21588 0 net472
rlabel metal3 15264 22092 15264 22092 0 net473
rlabel metal3 17568 21672 17568 21672 0 net474
rlabel metal2 43440 29484 43440 29484 0 net475
rlabel metal2 44448 29736 44448 29736 0 net476
rlabel metal3 8400 19236 8400 19236 0 net477
rlabel metal3 12480 17724 12480 17724 0 net478
rlabel metal2 41472 22302 41472 22302 0 net479
rlabel metal2 39264 15372 39264 15372 0 net48
rlabel metal2 39408 21672 39408 21672 0 net480
rlabel metal2 44544 21630 44544 21630 0 net481
rlabel metal2 45792 22848 45792 22848 0 net482
rlabel metal2 46560 31668 46560 31668 0 net483
rlabel metal2 47376 31332 47376 31332 0 net484
rlabel metal3 11664 28308 11664 28308 0 net485
rlabel metal2 9216 27342 9216 27342 0 net486
rlabel metal2 15648 34650 15648 34650 0 net487
rlabel metal2 14304 33684 14304 33684 0 net488
rlabel metal3 12384 23268 12384 23268 0 net489
rlabel metal2 10848 12012 10848 12012 0 net49
rlabel metal2 13056 22260 13056 22260 0 net490
rlabel metal3 40224 21336 40224 21336 0 net491
rlabel metal2 38400 23478 38400 23478 0 net492
rlabel metal3 5040 33684 5040 33684 0 net493
rlabel metal2 33168 29148 33168 29148 0 net494
rlabel metal2 33360 28308 33360 28308 0 net495
rlabel metal2 8352 9492 8352 9492 0 net496
rlabel metal2 5568 9828 5568 9828 0 net497
rlabel metal2 10560 26880 10560 26880 0 net498
rlabel metal3 9600 25284 9600 25284 0 net499
rlabel metal3 366 17388 366 17388 0 net5
rlabel metal2 29952 19572 29952 19572 0 net50
rlabel metal3 46176 24948 46176 24948 0 net500
rlabel metal2 48480 28392 48480 28392 0 net501
rlabel metal2 51648 29820 51648 29820 0 net502
rlabel metal3 37632 27384 37632 27384 0 net503
rlabel metal2 39360 31206 39360 31206 0 net504
rlabel metal2 45888 29400 45888 29400 0 net505
rlabel metal3 44352 22512 44352 22512 0 net506
rlabel metal2 39264 21042 39264 21042 0 net507
rlabel metal2 13104 30828 13104 30828 0 net508
rlabel metal2 16992 31626 16992 31626 0 net509
rlabel metal2 32064 22596 32064 22596 0 net51
rlabel metal2 13824 31626 13824 31626 0 net510
rlabel metal2 43776 26376 43776 26376 0 net511
rlabel metal2 42336 25116 42336 25116 0 net512
rlabel metal3 9120 15582 9120 15582 0 net513
rlabel metal2 9312 15246 9312 15246 0 net514
rlabel metal3 29712 37380 29712 37380 0 net515
rlabel metal2 3792 26628 3792 26628 0 net516
rlabel metal2 30912 33138 30912 33138 0 net517
rlabel metal2 33744 32256 33744 32256 0 net518
rlabel metal2 42912 34650 42912 34650 0 net519
rlabel metal2 37728 19572 37728 19572 0 net52
rlabel metal3 41184 34608 41184 34608 0 net520
rlabel metal2 16224 18564 16224 18564 0 net521
rlabel metal2 15072 19530 15072 19530 0 net522
rlabel metal2 46848 28266 46848 28266 0 net523
rlabel metal2 3984 30828 3984 30828 0 net524
rlabel metal3 8736 29106 8736 29106 0 net525
rlabel metal2 7104 27258 7104 27258 0 net526
rlabel metal3 43632 22596 43632 22596 0 net527
rlabel metal2 29472 6510 29472 6510 0 net528
rlabel metal2 31008 6468 31008 6468 0 net529
rlabel metal2 19200 20748 19200 20748 0 net53
rlabel metal2 36720 32172 36720 32172 0 net530
rlabel metal2 36000 29442 36000 29442 0 net531
rlabel metal2 37152 23310 37152 23310 0 net532
rlabel metal2 42240 21042 42240 21042 0 net533
rlabel metal2 13344 18774 13344 18774 0 net534
rlabel metal2 7584 6426 7584 6426 0 net535
rlabel metal2 2400 7434 2400 7434 0 net536
rlabel metal2 37920 21420 37920 21420 0 net537
rlabel metal2 19104 32508 19104 32508 0 net538
rlabel metal2 31392 30576 31392 30576 0 net539
rlabel metal3 1344 25956 1344 25956 0 net54
rlabel metal2 31248 32844 31248 32844 0 net540
rlabel metal2 32544 31626 32544 31626 0 net541
rlabel metal3 27264 29736 27264 29736 0 net542
rlabel metal2 4992 23058 4992 23058 0 net543
rlabel metal2 7392 27888 7392 27888 0 net544
rlabel metal3 27696 31332 27696 31332 0 net545
rlabel metal2 28704 5208 28704 5208 0 net546
rlabel metal2 29184 5208 29184 5208 0 net547
rlabel metal2 43392 33936 43392 33936 0 net548
rlabel metal2 7104 14994 7104 14994 0 net549
rlabel metal2 33120 36246 33120 36246 0 net55
rlabel metal2 5472 12894 5472 12894 0 net550
rlabel metal2 5664 14700 5664 14700 0 net551
rlabel metal2 33792 8022 33792 8022 0 net552
rlabel metal3 34992 8148 34992 8148 0 net553
rlabel metal2 36576 8232 36576 8232 0 net554
rlabel metal2 34560 8148 34560 8148 0 net555
rlabel metal2 33792 5922 33792 5922 0 net556
rlabel metal3 35760 6636 35760 6636 0 net557
rlabel metal2 8736 22596 8736 22596 0 net558
rlabel metal2 24288 34356 24288 34356 0 net559
rlabel metal2 7056 22428 7056 22428 0 net56
rlabel metal2 49056 25242 49056 25242 0 net560
rlabel metal2 51168 23352 51168 23352 0 net561
rlabel metal2 10176 8232 10176 8232 0 net562
rlabel metal3 7488 8148 7488 8148 0 net563
rlabel metal2 35472 11928 35472 11928 0 net564
rlabel metal2 37056 11676 37056 11676 0 net565
rlabel metal3 5904 21000 5904 21000 0 net566
rlabel metal2 6816 18942 6816 18942 0 net567
rlabel metal2 16320 3024 16320 3024 0 net568
rlabel metal2 16800 3738 16800 3738 0 net569
rlabel metal3 35760 35028 35760 35028 0 net57
rlabel metal2 39600 27048 39600 27048 0 net570
rlabel metal2 39744 30114 39744 30114 0 net571
rlabel metal2 21216 18816 21216 18816 0 net572
rlabel metal2 19776 20202 19776 20202 0 net573
rlabel metal3 7056 27636 7056 27636 0 net574
rlabel metal2 37824 27888 37824 27888 0 net575
rlabel metal3 31344 36876 31344 36876 0 net576
rlabel metal3 36288 9492 36288 9492 0 net577
rlabel metal2 36576 8652 36576 8652 0 net578
rlabel metal2 6144 23142 6144 23142 0 net579
rlabel metal2 1728 27132 1728 27132 0 net58
rlabel metal2 10752 1260 10752 1260 0 net580
rlabel metal2 9696 2604 9696 2604 0 net581
rlabel metal2 5664 16296 5664 16296 0 net582
rlabel metal2 5760 17304 5760 17304 0 net583
rlabel metal2 5808 17724 5808 17724 0 net584
rlabel metal2 43200 28392 43200 28392 0 net585
rlabel metal3 31104 5922 31104 5922 0 net586
rlabel metal2 29280 5880 29280 5880 0 net587
rlabel metal2 30048 4116 30048 4116 0 net588
rlabel metal3 49152 26124 49152 26124 0 net589
rlabel metal3 41616 33012 41616 33012 0 net59
rlabel metal2 49440 25242 49440 25242 0 net590
rlabel metal2 46848 30702 46848 30702 0 net591
rlabel metal2 15600 20160 15600 20160 0 net592
rlabel metal2 10272 21882 10272 21882 0 net593
rlabel metal2 14784 4956 14784 4956 0 net594
rlabel metal3 12054 5544 12054 5544 0 net595
rlabel metal3 16512 5628 16512 5628 0 net596
rlabel metal2 4416 15582 4416 15582 0 net597
rlabel metal2 4416 12600 4416 12600 0 net598
rlabel metal2 3408 13188 3408 13188 0 net599
rlabel metal3 366 18228 366 18228 0 net6
rlabel metal2 13248 19572 13248 19572 0 net60
rlabel metal2 37248 23520 37248 23520 0 net600
rlabel metal2 34464 22764 34464 22764 0 net601
rlabel metal3 3888 14532 3888 14532 0 net602
rlabel metal3 7344 17052 7344 17052 0 net603
rlabel metal3 15120 3948 15120 3948 0 net604
rlabel metal2 12192 4410 12192 4410 0 net605
rlabel metal2 28512 29778 28512 29778 0 net606
rlabel metal3 21456 18564 21456 18564 0 net607
rlabel metal2 19440 18732 19440 18732 0 net608
rlabel metal3 25344 5796 25344 5796 0 net609
rlabel metal2 43680 34104 43680 34104 0 net61
rlabel metal2 25728 4998 25728 4998 0 net610
rlabel metal3 6576 6300 6576 6300 0 net611
rlabel metal3 5376 5628 5376 5628 0 net612
rlabel metal2 4896 6174 4896 6174 0 net613
rlabel metal2 35424 11424 35424 11424 0 net614
rlabel metal2 34752 8706 34752 8706 0 net615
rlabel metal2 35520 7098 35520 7098 0 net616
rlabel metal3 10512 31332 10512 31332 0 net617
rlabel metal3 4800 17724 4800 17724 0 net618
rlabel metal3 4032 17052 4032 17052 0 net619
rlabel metal2 7344 31500 7344 31500 0 net62
rlabel metal2 8976 29652 8976 29652 0 net620
rlabel metal2 6960 3948 6960 3948 0 net621
rlabel metal3 5328 4956 5328 4956 0 net622
rlabel metal2 3360 4158 3360 4158 0 net623
rlabel metal3 3552 16212 3552 16212 0 net624
rlabel metal3 8160 14196 8160 14196 0 net625
rlabel metal2 9552 4116 9552 4116 0 net626
rlabel metal2 30720 16968 30720 16968 0 net627
rlabel metal2 29088 15204 29088 15204 0 net628
rlabel metal2 28992 18438 28992 18438 0 net629
rlabel metal3 40992 35028 40992 35028 0 net63
rlabel metal2 6240 7350 6240 7350 0 net630
rlabel metal2 25632 23142 25632 23142 0 net631
rlabel metal3 26208 21588 26208 21588 0 net632
rlabel metal2 28176 21672 28176 21672 0 net633
rlabel metal2 22560 18228 22560 18228 0 net634
rlabel metal2 22176 19320 22176 19320 0 net635
rlabel metal3 34176 14196 34176 14196 0 net636
rlabel metal2 33792 13860 33792 13860 0 net637
rlabel metal2 24864 25578 24864 25578 0 net638
rlabel metal2 37344 16338 37344 16338 0 net639
rlabel metal2 1632 23520 1632 23520 0 net64
rlabel metal2 39936 17346 39936 17346 0 net640
rlabel metal2 24768 19404 24768 19404 0 net641
rlabel metal3 19296 17724 19296 17724 0 net642
rlabel metal2 7776 5334 7776 5334 0 net643
rlabel metal2 8640 3654 8640 3654 0 net644
rlabel metal2 8736 5208 8736 5208 0 net645
rlabel metal2 36384 18984 36384 18984 0 net646
rlabel metal2 34656 19488 34656 19488 0 net647
rlabel metal2 38880 18816 38880 18816 0 net648
rlabel metal2 19008 16548 19008 16548 0 net649
rlabel metal2 30288 35028 30288 35028 0 net65
rlabel metal2 17952 17094 17952 17094 0 net650
rlabel metal2 15552 13986 15552 13986 0 net651
rlabel metal2 12960 16170 12960 16170 0 net652
rlabel metal3 37524 17724 37524 17724 0 net653
rlabel metal3 22512 4956 22512 4956 0 net654
rlabel metal3 19920 4116 19920 4116 0 net655
rlabel metal2 21408 3066 21408 3066 0 net656
rlabel metal2 26640 1092 26640 1092 0 net657
rlabel metal2 30480 17052 30480 17052 0 net658
rlabel metal2 29760 17976 29760 17976 0 net659
rlabel metal2 9888 30156 9888 30156 0 net66
rlabel metal2 7872 4200 7872 4200 0 net660
rlabel metal2 20928 5040 20928 5040 0 net661
rlabel metal2 23712 9786 23712 9786 0 net662
rlabel metal3 38832 14028 38832 14028 0 net663
rlabel metal2 25056 11256 25056 11256 0 net664
rlabel metal3 22032 11676 22032 11676 0 net665
rlabel metal2 21072 9492 21072 9492 0 net666
rlabel metal2 17856 10080 17856 10080 0 net667
rlabel metal3 13728 11508 13728 11508 0 net668
rlabel metal2 12000 11970 12000 11970 0 net669
rlabel metal2 26208 29400 26208 29400 0 net67
rlabel metal2 22416 7140 22416 7140 0 net670
rlabel metal2 23424 16506 23424 16506 0 net671
rlabel metal2 33744 23100 33744 23100 0 net672
rlabel metal2 12480 13482 12480 13482 0 net673
rlabel metal3 11328 14112 11328 14112 0 net674
rlabel metal2 20976 8148 20976 8148 0 net675
rlabel metal2 25632 12768 25632 12768 0 net676
rlabel metal2 4704 12432 4704 12432 0 net68
rlabel metal3 24912 31500 24912 31500 0 net69
rlabel metal3 366 19068 366 19068 0 net7
rlabel metal2 17472 30912 17472 30912 0 net70
rlabel metal2 28992 33810 28992 33810 0 net71
rlabel metal2 1632 25032 1632 25032 0 net72
rlabel metal2 35424 29736 35424 29736 0 net73
rlabel metal3 21792 33012 21792 33012 0 net74
rlabel metal2 33120 30660 33120 30660 0 net75
rlabel metal2 15792 19236 15792 19236 0 net76
rlabel metal2 33072 28308 33072 28308 0 net77
rlabel metal2 20352 31080 20352 31080 0 net78
rlabel metal2 28800 30660 28800 30660 0 net79
rlabel metal3 366 19908 366 19908 0 net8
rlabel metal2 5664 25284 5664 25284 0 net80
rlabel metal2 23040 31080 23040 31080 0 net81
rlabel metal2 6432 27636 6432 27636 0 net82
rlabel metal3 24048 33516 24048 33516 0 net83
rlabel metal2 5760 18438 5760 18438 0 net84
rlabel metal2 29424 35028 29424 35028 0 net85
rlabel metal2 1824 28644 1824 28644 0 net86
rlabel metal2 34512 33012 34512 33012 0 net87
rlabel metal3 7056 23940 7056 23940 0 net88
rlabel metal2 36480 28728 36480 28728 0 net89
rlabel metal3 366 20748 366 20748 0 net9
rlabel metal2 1920 31080 1920 31080 0 net90
rlabel metal3 33984 27468 33984 27468 0 net91
rlabel metal2 10608 22932 10608 22932 0 net92
rlabel metal3 32928 25284 32928 25284 0 net93
rlabel metal3 8592 31500 8592 31500 0 net94
rlabel metal3 36672 25956 36672 25956 0 net95
rlabel metal3 13728 22428 13728 22428 0 net96
rlabel metal2 40896 29022 40896 29022 0 net97
rlabel metal2 12288 31962 12288 31962 0 net98
rlabel metal2 42624 32592 42624 32592 0 net99
rlabel metal3 174 37548 174 37548 0 rst_n
rlabel metal3 22032 6468 22032 6468 0 u_ppwm/global_counter_high\[0\]
rlabel metal3 22656 2688 22656 2688 0 u_ppwm/global_counter_high\[10\]
rlabel metal3 23808 5628 23808 5628 0 u_ppwm/global_counter_high\[11\]
rlabel metal3 33888 7392 33888 7392 0 u_ppwm/global_counter_high\[12\]
rlabel metal2 37920 6762 37920 6762 0 u_ppwm/global_counter_high\[13\]
rlabel metal2 38112 7182 38112 7182 0 u_ppwm/global_counter_high\[14\]
rlabel metal2 38016 9198 38016 9198 0 u_ppwm/global_counter_high\[15\]
rlabel metal2 38880 9786 38880 9786 0 u_ppwm/global_counter_high\[16\]
rlabel metal2 36096 11634 36096 11634 0 u_ppwm/global_counter_high\[17\]
rlabel metal3 39168 11676 39168 11676 0 u_ppwm/global_counter_high\[18\]
rlabel metal2 32832 13272 32832 13272 0 u_ppwm/global_counter_high\[19\]
rlabel metal2 26496 6678 26496 6678 0 u_ppwm/global_counter_high\[1\]
rlabel metal2 22272 6930 22272 6930 0 u_ppwm/global_counter_high\[2\]
rlabel metal2 31056 8652 31056 8652 0 u_ppwm/global_counter_high\[3\]
rlabel metal2 31296 7266 31296 7266 0 u_ppwm/global_counter_high\[4\]
rlabel metal2 31872 8526 31872 8526 0 u_ppwm/global_counter_high\[5\]
rlabel metal3 29664 2856 29664 2856 0 u_ppwm/global_counter_high\[6\]
rlabel metal2 31685 11130 31685 11130 0 u_ppwm/global_counter_high\[7\]
rlabel metal2 25968 1932 25968 1932 0 u_ppwm/global_counter_high\[8\]
rlabel metal2 27456 12474 27456 12474 0 u_ppwm/global_counter_high\[9\]
rlabel metal4 30624 24612 30624 24612 0 u_ppwm/instr\[0\]
rlabel metal2 28032 19614 28032 19614 0 u_ppwm/instr\[1\]
rlabel metal2 26784 18732 26784 18732 0 u_ppwm/instr\[2\]
rlabel metal2 29664 22680 29664 22680 0 u_ppwm/instr\[3\]
rlabel metal2 27648 24864 27648 24864 0 u_ppwm/instr\[4\]
rlabel metal2 24864 22134 24864 22134 0 u_ppwm/instr\[5\]
rlabel metal2 26976 23310 26976 23310 0 u_ppwm/instr\[6\]
rlabel metal2 9408 14868 9408 14868 0 u_ppwm/mem_write_done
rlabel metal3 33456 22512 33456 22512 0 u_ppwm/pc\[0\]
rlabel metal2 31776 25452 31776 25452 0 u_ppwm/pc\[1\]
rlabel metal2 29568 25830 29568 25830 0 u_ppwm/pc\[2\]
rlabel metal3 30624 23100 30624 23100 0 u_ppwm/pc\[3\]
rlabel metal2 34080 5586 34080 5586 0 u_ppwm/period_start
rlabel metal2 15456 16380 15456 16380 0 u_ppwm/pwm_value\[0\]
rlabel metal3 22368 6972 22368 6972 0 u_ppwm/pwm_value\[1\]
rlabel metal2 23328 10542 23328 10542 0 u_ppwm/pwm_value\[2\]
rlabel metal2 24384 11382 24384 11382 0 u_ppwm/pwm_value\[3\]
rlabel via2 21504 10248 21504 10248 0 u_ppwm/pwm_value\[4\]
rlabel metal2 19968 7938 19968 7938 0 u_ppwm/pwm_value\[5\]
rlabel metal3 12672 11676 12672 11676 0 u_ppwm/pwm_value\[6\]
rlabel metal3 11808 13860 11808 13860 0 u_ppwm/pwm_value\[7\]
rlabel metal3 29856 13230 29856 13230 0 u_ppwm/pwm_value\[8\]
rlabel metal2 15840 14532 15840 14532 0 u_ppwm/pwm_value\[9\]
rlabel metal2 20448 19992 20448 19992 0 u_ppwm/u_ex/_000_
rlabel metal2 18144 19026 18144 19026 0 u_ppwm/u_ex/_001_
rlabel metal2 21360 20160 21360 20160 0 u_ppwm/u_ex/_002_
rlabel metal2 31584 22554 31584 22554 0 u_ppwm/u_ex/_003_
rlabel metal2 29424 24024 29424 24024 0 u_ppwm/u_ex/_004_
rlabel metal3 25488 24780 25488 24780 0 u_ppwm/u_ex/_005_
rlabel metal3 26592 21756 26592 21756 0 u_ppwm/u_ex/_006_
rlabel metal2 28704 14742 28704 14742 0 u_ppwm/u_ex/_007_
rlabel metal2 20064 16968 20064 16968 0 u_ppwm/u_ex/_008_
rlabel metal3 18864 12264 18864 12264 0 u_ppwm/u_ex/_009_
rlabel metal2 20736 10458 20736 10458 0 u_ppwm/u_ex/_010_
rlabel metal2 21600 12558 21600 12558 0 u_ppwm/u_ex/_011_
rlabel metal2 17088 10248 17088 10248 0 u_ppwm/u_ex/_012_
rlabel metal2 17568 8652 17568 8652 0 u_ppwm/u_ex/_013_
rlabel metal3 13200 11928 13200 11928 0 u_ppwm/u_ex/_014_
rlabel metal2 13824 12642 13824 12642 0 u_ppwm/u_ex/_015_
rlabel metal3 22464 13146 22464 13146 0 u_ppwm/u_ex/_016_
rlabel metal3 15888 16380 15888 16380 0 u_ppwm/u_ex/_017_
rlabel metal4 23136 18270 23136 18270 0 u_ppwm/u_ex/_018_
rlabel metal2 21504 17808 21504 17808 0 u_ppwm/u_ex/_019_
rlabel metal3 26640 17976 26640 17976 0 u_ppwm/u_ex/_020_
rlabel metal2 29184 16254 29184 16254 0 u_ppwm/u_ex/_021_
rlabel metal2 33312 14532 33312 14532 0 u_ppwm/u_ex/_022_
rlabel metal3 35424 16212 35424 16212 0 u_ppwm/u_ex/_023_
rlabel metal2 38304 17556 38304 17556 0 u_ppwm/u_ex/_024_
rlabel metal2 38784 17808 38784 17808 0 u_ppwm/u_ex/_025_
rlabel metal2 33936 18396 33936 18396 0 u_ppwm/u_ex/_026_
rlabel metal2 36672 18102 36672 18102 0 u_ppwm/u_ex/_027_
rlabel metal2 20832 18774 20832 18774 0 u_ppwm/u_ex/_028_
rlabel metal2 29861 10332 29861 10332 0 u_ppwm/u_ex/_029_
rlabel metal2 31776 7854 31776 7854 0 u_ppwm/u_ex/_030_
rlabel metal2 28992 8442 28992 8442 0 u_ppwm/u_ex/_031_
rlabel metal2 28128 6888 28128 6888 0 u_ppwm/u_ex/_032_
rlabel metal2 26880 13020 26880 13020 0 u_ppwm/u_ex/_033_
rlabel metal3 26160 11676 26160 11676 0 u_ppwm/u_ex/_034_
rlabel metal2 26496 11088 26496 11088 0 u_ppwm/u_ex/_035_
rlabel metal2 26304 10248 26304 10248 0 u_ppwm/u_ex/_036_
rlabel metal2 31104 8232 31104 8232 0 u_ppwm/u_ex/_037_
rlabel metal3 31392 7980 31392 7980 0 u_ppwm/u_ex/_038_
rlabel metal2 24733 7231 24733 7231 0 u_ppwm/u_ex/_039_
rlabel metal4 25728 22890 25728 22890 0 u_ppwm/u_ex/_040_
rlabel metal2 23088 23100 23088 23100 0 u_ppwm/u_ex/_041_
rlabel metal2 19584 19698 19584 19698 0 u_ppwm/u_ex/_042_
rlabel metal3 21600 20748 21600 20748 0 u_ppwm/u_ex/_043_
rlabel metal2 31584 14070 31584 14070 0 u_ppwm/u_ex/_044_
rlabel metal2 25872 14196 25872 14196 0 u_ppwm/u_ex/_045_
rlabel metal2 26544 20076 26544 20076 0 u_ppwm/u_ex/_046_
rlabel metal2 22272 19488 22272 19488 0 u_ppwm/u_ex/_047_
rlabel metal2 19488 19992 19488 19992 0 u_ppwm/u_ex/_048_
rlabel metal3 20112 20076 20112 20076 0 u_ppwm/u_ex/_049_
rlabel metal3 21408 17220 21408 17220 0 u_ppwm/u_ex/_050_
rlabel metal3 22176 20580 22176 20580 0 u_ppwm/u_ex/_051_
rlabel metal3 20640 18564 20640 18564 0 u_ppwm/u_ex/_052_
rlabel metal2 27360 22428 27360 22428 0 u_ppwm/u_ex/_053_
rlabel metal2 24864 23730 24864 23730 0 u_ppwm/u_ex/_054_
rlabel metal2 31200 23016 31200 23016 0 u_ppwm/u_ex/_055_
rlabel metal2 31584 23352 31584 23352 0 u_ppwm/u_ex/_056_
rlabel metal2 26112 23520 26112 23520 0 u_ppwm/u_ex/_057_
rlabel metal2 29040 23856 29040 23856 0 u_ppwm/u_ex/_058_
rlabel metal3 29232 23604 29232 23604 0 u_ppwm/u_ex/_059_
rlabel metal3 28128 23058 28128 23058 0 u_ppwm/u_ex/_060_
rlabel metal2 29184 23142 29184 23142 0 u_ppwm/u_ex/_061_
rlabel metal2 28512 23352 28512 23352 0 u_ppwm/u_ex/_062_
rlabel metal2 29088 23310 29088 23310 0 u_ppwm/u_ex/_063_
rlabel metal2 29760 23520 29760 23520 0 u_ppwm/u_ex/_064_
rlabel metal3 29136 23772 29136 23772 0 u_ppwm/u_ex/_065_
rlabel metal2 25440 23604 25440 23604 0 u_ppwm/u_ex/_066_
rlabel metal3 25632 22092 25632 22092 0 u_ppwm/u_ex/_067_
rlabel metal2 25440 23226 25440 23226 0 u_ppwm/u_ex/_068_
rlabel metal2 26208 23352 26208 23352 0 u_ppwm/u_ex/_069_
rlabel metal2 23616 22512 23616 22512 0 u_ppwm/u_ex/_070_
rlabel metal2 24768 23058 24768 23058 0 u_ppwm/u_ex/_071_
rlabel metal4 25152 23142 25152 23142 0 u_ppwm/u_ex/_072_
rlabel metal3 25824 23016 25824 23016 0 u_ppwm/u_ex/_073_
rlabel metal2 25680 24612 25680 24612 0 u_ppwm/u_ex/_074_
rlabel metal2 25920 23604 25920 23604 0 u_ppwm/u_ex/_075_
rlabel metal2 23856 22260 23856 22260 0 u_ppwm/u_ex/_076_
rlabel metal2 23808 22596 23808 22596 0 u_ppwm/u_ex/_077_
rlabel metal2 24192 22932 24192 22932 0 u_ppwm/u_ex/_078_
rlabel metal2 24288 22932 24288 22932 0 u_ppwm/u_ex/_079_
rlabel metal2 23712 23016 23712 23016 0 u_ppwm/u_ex/_080_
rlabel metal2 23808 23394 23808 23394 0 u_ppwm/u_ex/_081_
rlabel metal2 24000 22680 24000 22680 0 u_ppwm/u_ex/_082_
rlabel metal3 24864 21588 24864 21588 0 u_ppwm/u_ex/_083_
rlabel metal3 26928 22260 26928 22260 0 u_ppwm/u_ex/_084_
rlabel metal3 32592 10164 32592 10164 0 u_ppwm/u_ex/_085_
rlabel metal2 31872 8148 31872 8148 0 u_ppwm/u_ex/_086_
rlabel metal2 24960 7182 24960 7182 0 u_ppwm/u_ex/_087_
rlabel metal2 24768 6552 24768 6552 0 u_ppwm/u_ex/_088_
rlabel metal2 30048 7896 30048 7896 0 u_ppwm/u_ex/_089_
rlabel metal3 30528 8022 30528 8022 0 u_ppwm/u_ex/_090_
rlabel metal2 24672 6216 24672 6216 0 u_ppwm/u_ex/_091_
rlabel metal4 30624 6930 30624 6930 0 u_ppwm/u_ex/_092_
rlabel metal3 29568 7308 29568 7308 0 u_ppwm/u_ex/_093_
rlabel metal2 29664 7602 29664 7602 0 u_ppwm/u_ex/_094_
rlabel metal2 30720 8064 30720 8064 0 u_ppwm/u_ex/_095_
rlabel metal2 30816 8442 30816 8442 0 u_ppwm/u_ex/_096_
rlabel metal2 32496 10164 32496 10164 0 u_ppwm/u_ex/_097_
rlabel metal4 33120 10038 33120 10038 0 u_ppwm/u_ex/_098_
rlabel metal2 33216 9996 33216 9996 0 u_ppwm/u_ex/_099_
rlabel metal2 32448 12264 32448 12264 0 u_ppwm/u_ex/_100_
rlabel metal3 33888 13188 33888 13188 0 u_ppwm/u_ex/_101_
rlabel metal2 34560 12600 34560 12600 0 u_ppwm/u_ex/_102_
rlabel metal2 33792 11760 33792 11760 0 u_ppwm/u_ex/_103_
rlabel metal2 33552 11676 33552 11676 0 u_ppwm/u_ex/_104_
rlabel metal2 33600 11823 33600 11823 0 u_ppwm/u_ex/_105_
rlabel metal2 33984 12180 33984 12180 0 u_ppwm/u_ex/_106_
rlabel metal2 33408 11508 33408 11508 0 u_ppwm/u_ex/_107_
rlabel metal2 31680 13146 31680 13146 0 u_ppwm/u_ex/_108_
rlabel metal2 32256 13272 32256 13272 0 u_ppwm/u_ex/_109_
rlabel metal2 32352 13608 32352 13608 0 u_ppwm/u_ex/_110_
rlabel metal2 29280 10941 29280 10941 0 u_ppwm/u_ex/_111_
rlabel metal2 29088 11088 29088 11088 0 u_ppwm/u_ex/_112_
rlabel metal3 23808 8148 23808 8148 0 u_ppwm/u_ex/_113_
rlabel metal2 24000 8568 24000 8568 0 u_ppwm/u_ex/_114_
rlabel metal2 24384 9996 24384 9996 0 u_ppwm/u_ex/_115_
rlabel metal2 24480 9492 24480 9492 0 u_ppwm/u_ex/_116_
rlabel metal2 23760 8652 23760 8652 0 u_ppwm/u_ex/_117_
rlabel metal2 24192 8946 24192 8946 0 u_ppwm/u_ex/_118_
rlabel metal2 24768 9366 24768 9366 0 u_ppwm/u_ex/_119_
rlabel metal3 29664 9534 29664 9534 0 u_ppwm/u_ex/_120_
rlabel metal2 28896 10122 28896 10122 0 u_ppwm/u_ex/_121_
rlabel metal2 29568 8946 29568 8946 0 u_ppwm/u_ex/_122_
rlabel metal2 29088 9828 29088 9828 0 u_ppwm/u_ex/_123_
rlabel via2 29275 9324 29275 9324 0 u_ppwm/u_ex/_124_
rlabel metal2 28224 9912 28224 9912 0 u_ppwm/u_ex/_125_
rlabel metal2 29472 9618 29472 9618 0 u_ppwm/u_ex/_126_
rlabel metal2 29760 9744 29760 9744 0 u_ppwm/u_ex/_127_
rlabel metal2 29568 10080 29568 10080 0 u_ppwm/u_ex/_128_
rlabel metal2 29376 11256 29376 11256 0 u_ppwm/u_ex/_129_
rlabel metal2 28992 13104 28992 13104 0 u_ppwm/u_ex/_130_
rlabel metal3 29424 13860 29424 13860 0 u_ppwm/u_ex/_131_
rlabel metal3 27072 14112 27072 14112 0 u_ppwm/u_ex/_132_
rlabel metal2 28704 13272 28704 13272 0 u_ppwm/u_ex/_133_
rlabel metal2 29664 14112 29664 14112 0 u_ppwm/u_ex/_134_
rlabel metal2 29568 14280 29568 14280 0 u_ppwm/u_ex/_135_
rlabel metal2 30048 14616 30048 14616 0 u_ppwm/u_ex/_136_
rlabel metal2 30240 14322 30240 14322 0 u_ppwm/u_ex/_137_
rlabel metal2 29664 14658 29664 14658 0 u_ppwm/u_ex/_138_
rlabel metal3 29226 14616 29226 14616 0 u_ppwm/u_ex/_139_
rlabel metal2 28128 15582 28128 15582 0 u_ppwm/u_ex/_140_
rlabel metal2 23232 7056 23232 7056 0 u_ppwm/u_ex/_141_
rlabel metal2 23040 7434 23040 7434 0 u_ppwm/u_ex/_142_
rlabel metal2 22944 7350 22944 7350 0 u_ppwm/u_ex/_143_
rlabel metal2 26208 6972 26208 6972 0 u_ppwm/u_ex/_144_
rlabel metal2 25728 7392 25728 7392 0 u_ppwm/u_ex/_145_
rlabel metal2 26304 7476 26304 7476 0 u_ppwm/u_ex/_146_
rlabel metal2 26592 8736 26592 8736 0 u_ppwm/u_ex/_147_
rlabel metal2 26592 8190 26592 8190 0 u_ppwm/u_ex/_148_
rlabel metal2 26928 8148 26928 8148 0 u_ppwm/u_ex/_149_
rlabel metal2 26448 7140 26448 7140 0 u_ppwm/u_ex/_150_
rlabel metal2 26544 6972 26544 6972 0 u_ppwm/u_ex/_151_
rlabel metal2 27168 9156 27168 9156 0 u_ppwm/u_ex/_152_
rlabel metal2 27360 9702 27360 9702 0 u_ppwm/u_ex/_153_
rlabel metal3 26304 11046 26304 11046 0 u_ppwm/u_ex/_154_
rlabel metal2 26112 10878 26112 10878 0 u_ppwm/u_ex/_155_
rlabel metal2 26592 10164 26592 10164 0 u_ppwm/u_ex/_156_
rlabel metal2 27024 11172 27024 11172 0 u_ppwm/u_ex/_157_
rlabel metal2 26208 10920 26208 10920 0 u_ppwm/u_ex/_158_
rlabel metal2 26304 11508 26304 11508 0 u_ppwm/u_ex/_159_
rlabel metal3 26784 11676 26784 11676 0 u_ppwm/u_ex/_160_
rlabel metal2 27264 11844 27264 11844 0 u_ppwm/u_ex/_161_
rlabel metal2 27360 12180 27360 12180 0 u_ppwm/u_ex/_162_
rlabel metal2 29376 13356 29376 13356 0 u_ppwm/u_ex/_163_
rlabel metal4 28032 13272 28032 13272 0 u_ppwm/u_ex/_164_
rlabel metal2 27744 13650 27744 13650 0 u_ppwm/u_ex/_165_
rlabel metal2 30144 9534 30144 9534 0 u_ppwm/u_ex/_166_
rlabel metal2 27072 6636 27072 6636 0 u_ppwm/u_ex/_167_
rlabel metal3 25344 6636 25344 6636 0 u_ppwm/u_ex/_168_
rlabel metal3 26064 7140 26064 7140 0 u_ppwm/u_ex/_169_
rlabel metal2 28128 7896 28128 7896 0 u_ppwm/u_ex/_170_
rlabel metal3 28368 6972 28368 6972 0 u_ppwm/u_ex/_171_
rlabel metal2 28320 7224 28320 7224 0 u_ppwm/u_ex/_172_
rlabel metal2 29280 7896 29280 7896 0 u_ppwm/u_ex/_173_
rlabel metal2 29472 10038 29472 10038 0 u_ppwm/u_ex/_174_
rlabel metal2 30624 9996 30624 9996 0 u_ppwm/u_ex/_175_
rlabel metal2 29280 11382 29280 11382 0 u_ppwm/u_ex/_176_
rlabel metal2 30048 10962 30048 10962 0 u_ppwm/u_ex/_177_
rlabel metal3 29424 11508 29424 11508 0 u_ppwm/u_ex/_178_
rlabel metal3 29808 12516 29808 12516 0 u_ppwm/u_ex/_179_
rlabel metal2 30144 12474 30144 12474 0 u_ppwm/u_ex/_180_
rlabel metal2 30000 11508 30000 11508 0 u_ppwm/u_ex/_181_
rlabel metal2 30000 13020 30000 13020 0 u_ppwm/u_ex/_182_
rlabel metal2 29088 11802 29088 11802 0 u_ppwm/u_ex/_183_
rlabel metal2 28992 12012 28992 12012 0 u_ppwm/u_ex/_184_
rlabel metal2 29472 11886 29472 11886 0 u_ppwm/u_ex/_185_
rlabel metal2 27552 13734 27552 13734 0 u_ppwm/u_ex/_186_
rlabel metal2 31104 10416 31104 10416 0 u_ppwm/u_ex/_187_
rlabel metal2 24480 6972 24480 6972 0 u_ppwm/u_ex/_188_
rlabel metal2 23808 6342 23808 6342 0 u_ppwm/u_ex/_189_
rlabel metal2 24144 7140 24144 7140 0 u_ppwm/u_ex/_190_
rlabel metal3 24720 7980 24720 7980 0 u_ppwm/u_ex/_191_
rlabel metal4 31872 8820 31872 8820 0 u_ppwm/u_ex/_192_
rlabel metal2 33216 8526 33216 8526 0 u_ppwm/u_ex/_193_
rlabel metal2 32160 8316 32160 8316 0 u_ppwm/u_ex/_194_
rlabel metal2 31296 7938 31296 7938 0 u_ppwm/u_ex/_195_
rlabel metal2 31488 8946 31488 8946 0 u_ppwm/u_ex/_196_
rlabel metal2 32640 8148 32640 8148 0 u_ppwm/u_ex/_197_
rlabel metal2 32112 8904 32112 8904 0 u_ppwm/u_ex/_198_
rlabel metal2 32112 9660 32112 9660 0 u_ppwm/u_ex/_199_
rlabel metal2 31296 10710 31296 10710 0 u_ppwm/u_ex/_200_
rlabel metal2 31488 11970 31488 11970 0 u_ppwm/u_ex/_201_
rlabel metal2 26784 11760 26784 11760 0 u_ppwm/u_ex/_202_
rlabel metal2 26640 12516 26640 12516 0 u_ppwm/u_ex/_203_
rlabel metal3 25440 13146 25440 13146 0 u_ppwm/u_ex/_204_
rlabel metal2 26784 12453 26784 12453 0 u_ppwm/u_ex/_205_
rlabel metal2 27072 12768 27072 12768 0 u_ppwm/u_ex/_206_
rlabel metal2 27168 13524 27168 13524 0 u_ppwm/u_ex/_207_
rlabel metal2 27072 13608 27072 13608 0 u_ppwm/u_ex/_208_
rlabel metal2 27264 14238 27264 14238 0 u_ppwm/u_ex/_209_
rlabel metal2 28416 15666 28416 15666 0 u_ppwm/u_ex/_210_
rlabel metal2 26256 20076 26256 20076 0 u_ppwm/u_ex/_211_
rlabel metal2 26592 17808 26592 17808 0 u_ppwm/u_ex/_212_
rlabel metal2 24288 14910 24288 14910 0 u_ppwm/u_ex/_213_
rlabel metal2 23040 14322 23040 14322 0 u_ppwm/u_ex/_214_
rlabel metal2 25152 18732 25152 18732 0 u_ppwm/u_ex/_215_
rlabel metal2 33408 17514 33408 17514 0 u_ppwm/u_ex/_216_
rlabel metal2 33216 19530 33216 19530 0 u_ppwm/u_ex/_217_
rlabel metal2 19584 15582 19584 15582 0 u_ppwm/u_ex/_218_
rlabel metal2 20640 15708 20640 15708 0 u_ppwm/u_ex/_219_
rlabel metal2 21024 16380 21024 16380 0 u_ppwm/u_ex/_220_
rlabel metal2 33216 17766 33216 17766 0 u_ppwm/u_ex/_221_
rlabel metal2 20640 16884 20640 16884 0 u_ppwm/u_ex/_222_
rlabel metal2 21024 15750 21024 15750 0 u_ppwm/u_ex/_223_
rlabel metal2 18912 15582 18912 15582 0 u_ppwm/u_ex/_224_
rlabel metal2 19104 16170 19104 16170 0 u_ppwm/u_ex/_225_
rlabel metal2 20448 16212 20448 16212 0 u_ppwm/u_ex/_226_
rlabel metal2 33792 16926 33792 16926 0 u_ppwm/u_ex/_227_
rlabel metal2 19008 12474 19008 12474 0 u_ppwm/u_ex/_228_
rlabel metal2 19104 12264 19104 12264 0 u_ppwm/u_ex/_229_
rlabel metal3 19440 12516 19440 12516 0 u_ppwm/u_ex/_230_
rlabel metal2 19968 14784 19968 14784 0 u_ppwm/u_ex/_231_
rlabel metal2 19872 14616 19872 14616 0 u_ppwm/u_ex/_232_
rlabel metal3 21072 15540 21072 15540 0 u_ppwm/u_ex/_233_
rlabel metal2 20352 14826 20352 14826 0 u_ppwm/u_ex/_234_
rlabel metal2 21600 14280 21600 14280 0 u_ppwm/u_ex/_235_
rlabel metal3 23328 15372 23328 15372 0 u_ppwm/u_ex/_236_
rlabel metal3 22752 15540 22752 15540 0 u_ppwm/u_ex/_237_
rlabel metal2 21696 14112 21696 14112 0 u_ppwm/u_ex/_238_
rlabel metal2 21936 11004 21936 11004 0 u_ppwm/u_ex/_239_
rlabel metal3 20736 13188 20736 13188 0 u_ppwm/u_ex/_240_
rlabel metal2 21024 14658 21024 14658 0 u_ppwm/u_ex/_241_
rlabel metal2 21312 13482 21312 13482 0 u_ppwm/u_ex/_242_
rlabel metal2 21312 12768 21312 12768 0 u_ppwm/u_ex/_243_
rlabel metal2 21408 12642 21408 12642 0 u_ppwm/u_ex/_244_
rlabel metal2 21024 12516 21024 12516 0 u_ppwm/u_ex/_245_
rlabel metal3 19968 13188 19968 13188 0 u_ppwm/u_ex/_246_
rlabel metal2 19680 13356 19680 13356 0 u_ppwm/u_ex/_247_
rlabel metal2 16128 13104 16128 13104 0 u_ppwm/u_ex/_248_
rlabel metal3 15984 8652 15984 8652 0 u_ppwm/u_ex/_249_
rlabel metal2 15552 12117 15552 12117 0 u_ppwm/u_ex/_250_
rlabel metal3 16608 11508 16608 11508 0 u_ppwm/u_ex/_251_
rlabel metal2 16128 10248 16128 10248 0 u_ppwm/u_ex/_252_
rlabel metal2 16800 9996 16800 9996 0 u_ppwm/u_ex/_253_
rlabel metal2 16896 10122 16896 10122 0 u_ppwm/u_ex/_254_
rlabel metal3 16320 9492 16320 9492 0 u_ppwm/u_ex/_255_
rlabel metal2 15984 8652 15984 8652 0 u_ppwm/u_ex/_256_
rlabel metal2 16320 8988 16320 8988 0 u_ppwm/u_ex/_257_
rlabel metal2 16224 9576 16224 9576 0 u_ppwm/u_ex/_258_
rlabel metal3 16848 9324 16848 9324 0 u_ppwm/u_ex/_259_
rlabel metal2 17280 10332 17280 10332 0 u_ppwm/u_ex/_260_
rlabel metal2 17040 8652 17040 8652 0 u_ppwm/u_ex/_261_
rlabel metal2 14400 13440 14400 13440 0 u_ppwm/u_ex/_262_
rlabel metal3 14304 12516 14304 12516 0 u_ppwm/u_ex/_263_
rlabel metal2 16608 12432 16608 12432 0 u_ppwm/u_ex/_264_
rlabel metal3 16224 12516 16224 12516 0 u_ppwm/u_ex/_265_
rlabel metal2 16080 12516 16080 12516 0 u_ppwm/u_ex/_266_
rlabel metal2 14400 12306 14400 12306 0 u_ppwm/u_ex/_267_
rlabel metal2 14304 13438 14304 13438 0 u_ppwm/u_ex/_268_
rlabel metal2 15312 13440 15312 13440 0 u_ppwm/u_ex/_269_
rlabel metal2 13920 12012 13920 12012 0 u_ppwm/u_ex/_270_
rlabel metal2 14016 11802 14016 11802 0 u_ppwm/u_ex/_271_
rlabel metal2 13632 11676 13632 11676 0 u_ppwm/u_ex/_272_
rlabel metal2 14496 13104 14496 13104 0 u_ppwm/u_ex/_273_
rlabel metal2 13344 13734 13344 13734 0 u_ppwm/u_ex/_274_
rlabel metal2 14688 13734 14688 13734 0 u_ppwm/u_ex/_275_
rlabel metal2 13920 12684 13920 12684 0 u_ppwm/u_ex/_276_
rlabel metal2 14016 12558 14016 12558 0 u_ppwm/u_ex/_277_
rlabel metal2 13680 12516 13680 12516 0 u_ppwm/u_ex/_278_
rlabel metal2 15168 12558 15168 12558 0 u_ppwm/u_ex/_279_
rlabel metal3 15168 12684 15168 12684 0 u_ppwm/u_ex/_280_
rlabel metal3 15936 13188 15936 13188 0 u_ppwm/u_ex/_281_
rlabel metal2 17280 14364 17280 14364 0 u_ppwm/u_ex/_282_
rlabel metal2 17856 14196 17856 14196 0 u_ppwm/u_ex/_283_
rlabel metal2 17376 14280 17376 14280 0 u_ppwm/u_ex/_284_
rlabel metal3 17328 13104 17328 13104 0 u_ppwm/u_ex/_285_
rlabel metal2 19296 13230 19296 13230 0 u_ppwm/u_ex/_286_
rlabel metal2 19392 12936 19392 12936 0 u_ppwm/u_ex/_287_
rlabel metal2 18624 12894 18624 12894 0 u_ppwm/u_ex/_288_
rlabel metal2 18672 14700 18672 14700 0 u_ppwm/u_ex/_289_
rlabel metal2 16032 15246 16032 15246 0 u_ppwm/u_ex/_290_
rlabel metal2 17856 14994 17856 14994 0 u_ppwm/u_ex/_291_
rlabel metal3 17136 16212 17136 16212 0 u_ppwm/u_ex/_292_
rlabel metal2 15792 14196 15792 14196 0 u_ppwm/u_ex/_293_
rlabel metal2 33120 18102 33120 18102 0 u_ppwm/u_ex/_294_
rlabel metal2 29280 17178 29280 17178 0 u_ppwm/u_ex/_295_
rlabel metal2 23616 16380 23616 16380 0 u_ppwm/u_ex/_296_
rlabel metal2 23520 17934 23520 17934 0 u_ppwm/u_ex/_297_
rlabel metal2 23376 17220 23376 17220 0 u_ppwm/u_ex/_298_
rlabel metal2 23040 18186 23040 18186 0 u_ppwm/u_ex/_299_
rlabel metal3 22704 17724 22704 17724 0 u_ppwm/u_ex/_300_
rlabel metal3 23232 17766 23232 17766 0 u_ppwm/u_ex/_301_
rlabel metal2 22848 16170 22848 16170 0 u_ppwm/u_ex/_302_
rlabel metal2 22272 16212 22272 16212 0 u_ppwm/u_ex/_303_
rlabel metal2 23424 17598 23424 17598 0 u_ppwm/u_ex/_304_
rlabel metal2 24624 17220 24624 17220 0 u_ppwm/u_ex/_305_
rlabel metal2 24384 17682 24384 17682 0 u_ppwm/u_ex/_306_
rlabel metal2 25440 17388 25440 17388 0 u_ppwm/u_ex/_307_
rlabel metal2 24192 17850 24192 17850 0 u_ppwm/u_ex/_308_
rlabel metal2 24192 17304 24192 17304 0 u_ppwm/u_ex/_309_
rlabel metal2 29280 15750 29280 15750 0 u_ppwm/u_ex/_310_
rlabel metal2 27840 16947 27840 16947 0 u_ppwm/u_ex/_311_
rlabel metal3 27312 16800 27312 16800 0 u_ppwm/u_ex/_312_
rlabel via2 27744 17291 27744 17291 0 u_ppwm/u_ex/_313_
rlabel metal2 26736 16464 26736 16464 0 u_ppwm/u_ex/_314_
rlabel metal3 25152 15540 25152 15540 0 u_ppwm/u_ex/_315_
rlabel metal2 25632 16044 25632 16044 0 u_ppwm/u_ex/_316_
rlabel metal2 26496 17220 26496 17220 0 u_ppwm/u_ex/_317_
rlabel metal2 26160 16212 26160 16212 0 u_ppwm/u_ex/_318_
rlabel metal2 27984 17052 27984 17052 0 u_ppwm/u_ex/_319_
rlabel metal2 28512 16128 28512 16128 0 u_ppwm/u_ex/_320_
rlabel metal2 28416 16506 28416 16506 0 u_ppwm/u_ex/_321_
rlabel metal2 29088 16128 29088 16128 0 u_ppwm/u_ex/_322_
rlabel metal2 28992 16506 28992 16506 0 u_ppwm/u_ex/_323_
rlabel metal2 29328 16212 29328 16212 0 u_ppwm/u_ex/_324_
rlabel metal2 29472 16254 29472 16254 0 u_ppwm/u_ex/_325_
rlabel metal2 29472 15624 29472 15624 0 u_ppwm/u_ex/_326_
rlabel metal2 33120 14910 33120 14910 0 u_ppwm/u_ex/_327_
rlabel metal3 34368 15540 34368 15540 0 u_ppwm/u_ex/_328_
rlabel metal2 35424 15498 35424 15498 0 u_ppwm/u_ex/_329_
rlabel metal2 34176 14616 34176 14616 0 u_ppwm/u_ex/_330_
rlabel metal2 32832 14490 32832 14490 0 u_ppwm/u_ex/_331_
rlabel via1 31968 14693 31968 14693 0 u_ppwm/u_ex/_332_
rlabel metal2 31872 14994 31872 14994 0 u_ppwm/u_ex/_333_
rlabel metal3 31776 14700 31776 14700 0 u_ppwm/u_ex/_334_
rlabel metal2 33696 15582 33696 15582 0 u_ppwm/u_ex/_335_
rlabel metal2 33408 15792 33408 15792 0 u_ppwm/u_ex/_336_
rlabel metal2 33600 16128 33600 16128 0 u_ppwm/u_ex/_337_
rlabel metal2 32928 16128 32928 16128 0 u_ppwm/u_ex/_338_
rlabel metal2 32784 15708 32784 15708 0 u_ppwm/u_ex/_339_
rlabel metal3 32736 16212 32736 16212 0 u_ppwm/u_ex/_340_
rlabel metal3 38784 16212 38784 16212 0 u_ppwm/u_ex/_341_
rlabel metal2 37584 15540 37584 15540 0 u_ppwm/u_ex/_342_
rlabel metal2 35760 15708 35760 15708 0 u_ppwm/u_ex/_343_
rlabel metal2 35712 15246 35712 15246 0 u_ppwm/u_ex/_344_
rlabel metal2 36288 15446 36288 15446 0 u_ppwm/u_ex/_345_
rlabel metal2 37536 15288 37536 15288 0 u_ppwm/u_ex/_346_
rlabel metal2 37152 16128 37152 16128 0 u_ppwm/u_ex/_347_
rlabel metal4 37152 15288 37152 15288 0 u_ppwm/u_ex/_348_
rlabel metal2 38400 16716 38400 16716 0 u_ppwm/u_ex/_349_
rlabel metal2 38496 16926 38496 16926 0 u_ppwm/u_ex/_350_
rlabel metal2 37680 16212 37680 16212 0 u_ppwm/u_ex/_351_
rlabel metal3 37056 15330 37056 15330 0 u_ppwm/u_ex/_352_
rlabel metal2 38880 15792 38880 15792 0 u_ppwm/u_ex/_353_
rlabel metal2 38976 15456 38976 15456 0 u_ppwm/u_ex/_354_
rlabel metal2 37728 17136 37728 17136 0 u_ppwm/u_ex/_355_
rlabel metal2 37440 17598 37440 17598 0 u_ppwm/u_ex/_356_
rlabel metal3 37344 17640 37344 17640 0 u_ppwm/u_ex/_357_
rlabel metal3 36480 15708 36480 15708 0 u_ppwm/u_ex/_358_
rlabel metal2 36240 16212 36240 16212 0 u_ppwm/u_ex/_359_
rlabel metal2 35808 16338 35808 16338 0 u_ppwm/u_ex/_360_
rlabel metal2 35616 20496 35616 20496 0 u_ppwm/u_ex/_361_
rlabel metal3 35184 17136 35184 17136 0 u_ppwm/u_ex/_362_
rlabel metal2 35136 19446 35136 19446 0 u_ppwm/u_ex/_363_
rlabel metal2 34176 18354 34176 18354 0 u_ppwm/u_ex/_364_
rlabel metal2 33744 18564 33744 18564 0 u_ppwm/u_ex/_365_
rlabel metal2 33600 18438 33600 18438 0 u_ppwm/u_ex/_366_
rlabel metal2 35424 18144 35424 18144 0 u_ppwm/u_ex/_367_
rlabel metal2 35328 20370 35328 20370 0 u_ppwm/u_ex/_368_
rlabel metal2 34656 18522 34656 18522 0 u_ppwm/u_ex/_369_
rlabel metal2 35904 18648 35904 18648 0 u_ppwm/u_ex/_370_
rlabel metal3 36384 17724 36384 17724 0 u_ppwm/u_ex/_371_
rlabel metal2 36768 17976 36768 17976 0 u_ppwm/u_ex/_372_
rlabel metal2 31584 11046 31584 11046 0 u_ppwm/u_ex/_373_
rlabel metal2 33024 10878 33024 10878 0 u_ppwm/u_ex/_374_
rlabel metal3 32352 8652 32352 8652 0 u_ppwm/u_ex/_375_
rlabel metal2 30144 8190 30144 8190 0 u_ppwm/u_ex/_376_
rlabel metal2 25056 8442 25056 8442 0 u_ppwm/u_ex/_377_
rlabel metal2 25344 7938 25344 7938 0 u_ppwm/u_ex/_378_
rlabel metal2 28416 13650 28416 13650 0 u_ppwm/u_ex/_379_
rlabel metal2 29280 12390 29280 12390 0 u_ppwm/u_ex/_380_
rlabel metal2 29952 9576 29952 9576 0 u_ppwm/u_ex/_381_
rlabel metal2 30240 9240 30240 9240 0 u_ppwm/u_ex/_382_
rlabel metal3 22944 11004 22944 11004 0 u_ppwm/u_ex/_383_
rlabel metal2 31104 23436 31104 23436 0 u_ppwm/u_ex/_384_
rlabel metal2 31440 17724 31440 17724 0 u_ppwm/u_ex/_385_
rlabel metal3 30960 15708 30960 15708 0 u_ppwm/u_ex/_386_
rlabel metal2 31104 19824 31104 19824 0 u_ppwm/u_ex/cmp_flag_q
rlabel metal2 23856 15708 23856 15708 0 u_ppwm/u_ex/reg_value_q\[0\]
rlabel metal2 21408 18270 21408 18270 0 u_ppwm/u_ex/reg_value_q\[1\]
rlabel metal2 30048 16926 30048 16926 0 u_ppwm/u_ex/reg_value_q\[2\]
rlabel metal2 31680 15708 31680 15708 0 u_ppwm/u_ex/reg_value_q\[3\]
rlabel metal2 36000 15120 36000 15120 0 u_ppwm/u_ex/reg_value_q\[4\]
rlabel metal2 37536 16792 37536 16792 0 u_ppwm/u_ex/reg_value_q\[5\]
rlabel metal3 37140 16212 37140 16212 0 u_ppwm/u_ex/reg_value_q\[6\]
rlabel metal2 32304 11676 32304 11676 0 u_ppwm/u_ex/reg_value_q\[7\]
rlabel metal2 36960 18564 36960 18564 0 u_ppwm/u_ex/reg_value_q\[8\]
rlabel metal2 39744 17556 39744 17556 0 u_ppwm/u_ex/reg_value_q\[9\]
rlabel metal2 22176 20790 22176 20790 0 u_ppwm/u_ex/state_q\[0\]
rlabel metal3 20928 19236 20928 19236 0 u_ppwm/u_ex/state_q\[1\]
rlabel metal2 23712 21924 23712 21924 0 u_ppwm/u_ex/state_q\[2\]
rlabel metal3 20448 2100 20448 2100 0 u_ppwm/u_global_counter/_000_
rlabel metal3 19872 3948 19872 3948 0 u_ppwm/u_global_counter/_001_
rlabel metal2 19968 3066 19968 3066 0 u_ppwm/u_global_counter/_002_
rlabel metal2 28464 5124 28464 5124 0 u_ppwm/u_global_counter/_003_
rlabel metal2 30240 6510 30240 6510 0 u_ppwm/u_global_counter/_004_
rlabel metal2 28800 5166 28800 5166 0 u_ppwm/u_global_counter/_005_
rlabel metal2 27360 3864 27360 3864 0 u_ppwm/u_global_counter/_006_
rlabel metal2 26592 3738 26592 3738 0 u_ppwm/u_global_counter/_007_
rlabel metal2 25104 2604 25104 2604 0 u_ppwm/u_global_counter/_008_
rlabel metal2 26304 1638 26304 1638 0 u_ppwm/u_global_counter/_009_
rlabel metal2 25056 1134 25056 1134 0 u_ppwm/u_global_counter/_010_
rlabel metal2 25632 5754 25632 5754 0 u_ppwm/u_global_counter/_011_
rlabel metal2 33792 5460 33792 5460 0 u_ppwm/u_global_counter/_012_
rlabel metal2 34992 7980 34992 7980 0 u_ppwm/u_global_counter/_013_
rlabel metal3 35232 8736 35232 8736 0 u_ppwm/u_global_counter/_014_
rlabel metal2 35808 8736 35808 8736 0 u_ppwm/u_global_counter/_015_
rlabel metal2 36288 10122 36288 10122 0 u_ppwm/u_global_counter/_016_
rlabel metal3 35232 11172 35232 11172 0 u_ppwm/u_global_counter/_017_
rlabel metal2 36288 11970 36288 11970 0 u_ppwm/u_global_counter/_018_
rlabel metal2 37632 12558 37632 12558 0 u_ppwm/u_global_counter/_019_
rlabel metal2 28032 5628 28032 5628 0 u_ppwm/u_global_counter/_020_
rlabel metal2 25248 5292 25248 5292 0 u_ppwm/u_global_counter/_021_
rlabel metal3 34272 5628 34272 5628 0 u_ppwm/u_global_counter/_022_
rlabel metal2 35424 8946 35424 8946 0 u_ppwm/u_global_counter/_023_
rlabel metal2 34656 11676 34656 11676 0 u_ppwm/u_global_counter/_024_
rlabel metal2 35808 12600 35808 12600 0 u_ppwm/u_global_counter/_025_
rlabel metal2 25536 2814 25536 2814 0 u_ppwm/u_global_counter/_026_
rlabel metal3 24960 3948 24960 3948 0 u_ppwm/u_global_counter/_027_
rlabel metal3 21216 4116 21216 4116 0 u_ppwm/u_global_counter/_028_
rlabel metal2 28272 5628 28272 5628 0 u_ppwm/u_global_counter/_029_
rlabel metal3 29760 6426 29760 6426 0 u_ppwm/u_global_counter/_030_
rlabel metal3 27168 4956 27168 4956 0 u_ppwm/u_global_counter/_031_
rlabel metal2 27936 5040 27936 5040 0 u_ppwm/u_global_counter/_032_
rlabel metal2 30048 5922 30048 5922 0 u_ppwm/u_global_counter/_033_
rlabel metal2 26832 4956 26832 4956 0 u_ppwm/u_global_counter/_034_
rlabel metal2 26784 1806 26784 1806 0 u_ppwm/u_global_counter/_035_
rlabel metal2 29184 3612 29184 3612 0 u_ppwm/u_global_counter/_036_
rlabel metal3 26256 924 26256 924 0 u_ppwm/u_global_counter/_037_
rlabel metal2 26112 2142 26112 2142 0 u_ppwm/u_global_counter/_038_
rlabel metal2 25536 5418 25536 5418 0 u_ppwm/u_global_counter/_039_
rlabel metal2 26496 5628 26496 5628 0 u_ppwm/u_global_counter/_040_
rlabel metal2 33504 8568 33504 8568 0 u_ppwm/u_global_counter/_041_
rlabel metal2 34368 5880 34368 5880 0 u_ppwm/u_global_counter/_042_
rlabel metal3 33984 5460 33984 5460 0 u_ppwm/u_global_counter/_043_
rlabel metal2 34416 8652 34416 8652 0 u_ppwm/u_global_counter/_044_
rlabel metal2 36384 7896 36384 7896 0 u_ppwm/u_global_counter/_045_
rlabel metal3 34656 8652 34656 8652 0 u_ppwm/u_global_counter/_046_
rlabel metal2 34992 10164 34992 10164 0 u_ppwm/u_global_counter/_047_
rlabel metal2 36096 10626 36096 10626 0 u_ppwm/u_global_counter/_048_
rlabel metal2 35328 10668 35328 10668 0 u_ppwm/u_global_counter/_049_
rlabel metal2 34992 11508 34992 11508 0 u_ppwm/u_global_counter/_050_
rlabel metal3 35376 10416 35376 10416 0 u_ppwm/u_global_counter/_051_
rlabel metal2 35952 12516 35952 12516 0 u_ppwm/u_global_counter/_052_
rlabel metal3 10224 22260 10224 22260 0 u_ppwm/u_mem/_0000_
rlabel metal2 16320 19782 16320 19782 0 u_ppwm/u_mem/_0001_
rlabel metal3 15024 19488 15024 19488 0 u_ppwm/u_mem/_0002_
rlabel metal2 12288 18270 12288 18270 0 u_ppwm/u_mem/_0003_
rlabel metal2 9984 14826 9984 14826 0 u_ppwm/u_mem/_0004_
rlabel metal2 7200 14238 7200 14238 0 u_ppwm/u_mem/_0005_
rlabel metal2 9408 16632 9408 16632 0 u_ppwm/u_mem/_0006_
rlabel metal2 43392 25578 43392 25578 0 u_ppwm/u_mem/_0007_
rlabel metal2 41760 27090 41760 27090 0 u_ppwm/u_mem/_0008_
rlabel metal2 48960 30576 48960 30576 0 u_ppwm/u_mem/_0009_
rlabel metal3 47760 29736 47760 29736 0 u_ppwm/u_mem/_0010_
rlabel metal2 42144 21504 42144 21504 0 u_ppwm/u_mem/_0011_
rlabel metal3 36144 23268 36144 23268 0 u_ppwm/u_mem/_0012_
rlabel metal2 45216 21756 45216 21756 0 u_ppwm/u_mem/_0013_
rlabel metal2 48432 23772 48432 23772 0 u_ppwm/u_mem/_0014_
rlabel metal2 47904 25578 47904 25578 0 u_ppwm/u_mem/_0015_
rlabel metal2 45600 27090 45600 27090 0 u_ppwm/u_mem/_0016_
rlabel metal2 49344 27678 49344 27678 0 u_ppwm/u_mem/_0017_
rlabel metal2 42240 23016 42240 23016 0 u_ppwm/u_mem/_0018_
rlabel metal2 39024 23100 39024 23100 0 u_ppwm/u_mem/_0019_
rlabel metal3 39744 21588 39744 21588 0 u_ppwm/u_mem/_0020_
rlabel metal2 48528 24444 48528 24444 0 u_ppwm/u_mem/_0021_
rlabel metal2 49632 26838 49632 26838 0 u_ppwm/u_mem/_0022_
rlabel metal2 47232 31500 47232 31500 0 u_ppwm/u_mem/_0023_
rlabel metal3 45408 31500 45408 31500 0 u_ppwm/u_mem/_0024_
rlabel metal2 38448 30408 38448 30408 0 u_ppwm/u_mem/_0025_
rlabel metal2 36384 26670 36384 26670 0 u_ppwm/u_mem/_0026_
rlabel metal2 40176 19908 40176 19908 0 u_ppwm/u_mem/_0027_
rlabel metal2 46752 24066 46752 24066 0 u_ppwm/u_mem/_0028_
rlabel metal2 44832 25368 44832 25368 0 u_ppwm/u_mem/_0029_
rlabel metal2 43680 30114 43680 30114 0 u_ppwm/u_mem/_0030_
rlabel metal2 42912 31626 42912 31626 0 u_ppwm/u_mem/_0031_
rlabel metal2 39552 30744 39552 30744 0 u_ppwm/u_mem/_0032_
rlabel metal2 35712 25452 35712 25452 0 u_ppwm/u_mem/_0033_
rlabel metal2 33888 25368 33888 25368 0 u_ppwm/u_mem/_0034_
rlabel metal3 34704 25956 34704 25956 0 u_ppwm/u_mem/_0035_
rlabel metal2 37152 29946 37152 29946 0 u_ppwm/u_mem/_0036_
rlabel metal2 33504 31332 33504 31332 0 u_ppwm/u_mem/_0037_
rlabel metal2 28032 31374 28032 31374 0 u_ppwm/u_mem/_0038_
rlabel metal2 23616 33012 23616 33012 0 u_ppwm/u_mem/_0039_
rlabel metal3 24912 30324 24912 30324 0 u_ppwm/u_mem/_0040_
rlabel metal2 29040 28980 29040 28980 0 u_ppwm/u_mem/_0041_
rlabel metal3 31344 29148 31344 29148 0 u_ppwm/u_mem/_0042_
rlabel metal2 33744 29316 33744 29316 0 u_ppwm/u_mem/_0043_
rlabel metal2 35040 31416 35040 31416 0 u_ppwm/u_mem/_0044_
rlabel metal2 29376 32424 29376 32424 0 u_ppwm/u_mem/_0045_
rlabel metal2 26016 31710 26016 31710 0 u_ppwm/u_mem/_0046_
rlabel metal3 28272 29064 28272 29064 0 u_ppwm/u_mem/_0047_
rlabel metal3 32016 33684 32016 33684 0 u_ppwm/u_mem/_0048_
rlabel metal2 40800 34314 40800 34314 0 u_ppwm/u_mem/_0049_
rlabel metal2 42144 32508 42144 32508 0 u_ppwm/u_mem/_0050_
rlabel metal2 41184 33936 41184 33936 0 u_ppwm/u_mem/_0051_
rlabel metal2 36000 34650 36000 34650 0 u_ppwm/u_mem/_0052_
rlabel metal2 32352 36120 32352 36120 0 u_ppwm/u_mem/_0053_
rlabel metal2 27936 35112 27936 35112 0 u_ppwm/u_mem/_0054_
rlabel metal3 24912 35280 24912 35280 0 u_ppwm/u_mem/_0055_
rlabel metal2 38496 35616 38496 35616 0 u_ppwm/u_mem/_0056_
rlabel metal2 39456 35322 39456 35322 0 u_ppwm/u_mem/_0057_
rlabel metal2 37920 33138 37920 33138 0 u_ppwm/u_mem/_0058_
rlabel metal2 33888 34188 33888 34188 0 u_ppwm/u_mem/_0059_
rlabel metal2 29760 35322 29760 35322 0 u_ppwm/u_mem/_0060_
rlabel metal2 24480 36204 24480 36204 0 u_ppwm/u_mem/_0061_
rlabel metal2 21744 33852 21744 33852 0 u_ppwm/u_mem/_0062_
rlabel metal2 18816 34230 18816 34230 0 u_ppwm/u_mem/_0063_
rlabel metal3 15312 34272 15312 34272 0 u_ppwm/u_mem/_0064_
rlabel metal2 9360 34608 9360 34608 0 u_ppwm/u_mem/_0065_
rlabel metal3 4656 34356 4656 34356 0 u_ppwm/u_mem/_0066_
rlabel metal2 3744 32928 3744 32928 0 u_ppwm/u_mem/_0067_
rlabel metal2 1344 32676 1344 32676 0 u_ppwm/u_mem/_0068_
rlabel metal3 14448 33096 14448 33096 0 u_ppwm/u_mem/_0069_
rlabel metal2 16464 34944 16464 34944 0 u_ppwm/u_mem/_0070_
rlabel metal2 13344 36708 13344 36708 0 u_ppwm/u_mem/_0071_
rlabel metal2 9024 35574 9024 35574 0 u_ppwm/u_mem/_0072_
rlabel metal2 7008 35238 7008 35238 0 u_ppwm/u_mem/_0073_
rlabel metal2 5568 32172 5568 32172 0 u_ppwm/u_mem/_0074_
rlabel metal2 1248 30492 1248 30492 0 u_ppwm/u_mem/_0075_
rlabel metal2 11616 30366 11616 30366 0 u_ppwm/u_mem/_0076_
rlabel metal2 14016 30576 14016 30576 0 u_ppwm/u_mem/_0077_
rlabel metal3 15600 33684 15600 33684 0 u_ppwm/u_mem/_0078_
rlabel metal2 12192 31584 12192 31584 0 u_ppwm/u_mem/_0079_
rlabel metal2 8160 32928 8160 32928 0 u_ppwm/u_mem/_0080_
rlabel metal2 1344 29820 1344 29820 0 u_ppwm/u_mem/_0081_
rlabel metal3 2736 28224 2736 28224 0 u_ppwm/u_mem/_0082_
rlabel metal2 8256 28266 8256 28266 0 u_ppwm/u_mem/_0083_
rlabel metal2 20640 31416 20640 31416 0 u_ppwm/u_mem/_0084_
rlabel metal2 22560 32466 22560 32466 0 u_ppwm/u_mem/_0085_
rlabel metal2 16800 31584 16800 31584 0 u_ppwm/u_mem/_0086_
rlabel metal2 9696 31290 9696 31290 0 u_ppwm/u_mem/_0087_
rlabel via1 5277 29232 5277 29232 0 u_ppwm/u_mem/_0088_
rlabel metal2 3840 27090 3840 27090 0 u_ppwm/u_mem/_0089_
rlabel metal3 2832 26208 2832 26208 0 u_ppwm/u_mem/_0090_
rlabel metal3 9552 26292 9552 26292 0 u_ppwm/u_mem/_0091_
rlabel metal2 19872 29064 19872 29064 0 u_ppwm/u_mem/_0092_
rlabel metal2 20064 28602 20064 28602 0 u_ppwm/u_mem/_0093_
rlabel metal2 18576 24444 18576 24444 0 u_ppwm/u_mem/_0094_
rlabel metal2 17088 23856 17088 23856 0 u_ppwm/u_mem/_0095_
rlabel metal2 14496 24066 14496 24066 0 u_ppwm/u_mem/_0096_
rlabel metal3 11808 24654 11808 24654 0 u_ppwm/u_mem/_0097_
rlabel metal2 10800 26124 10800 26124 0 u_ppwm/u_mem/_0098_
rlabel metal2 20496 26796 20496 26796 0 u_ppwm/u_mem/_0099_
rlabel metal3 21456 27468 21456 27468 0 u_ppwm/u_mem/_0100_
rlabel metal2 19584 24402 19584 24402 0 u_ppwm/u_mem/_0101_
rlabel metal2 16992 21630 16992 21630 0 u_ppwm/u_mem/_0102_
rlabel metal2 12768 23016 12768 23016 0 u_ppwm/u_mem/_0103_
rlabel metal3 6864 23268 6864 23268 0 u_ppwm/u_mem/_0104_
rlabel metal2 5856 25704 5856 25704 0 u_ppwm/u_mem/_0105_
rlabel metal2 2784 24150 2784 24150 0 u_ppwm/u_mem/_0106_
rlabel metal2 3168 23394 3168 23394 0 u_ppwm/u_mem/_0107_
rlabel metal3 6288 19908 6288 19908 0 u_ppwm/u_mem/_0108_
rlabel metal2 10464 20328 10464 20328 0 u_ppwm/u_mem/_0109_
rlabel metal2 12096 17052 12096 17052 0 u_ppwm/u_mem/_0110_
rlabel metal2 7488 18480 7488 18480 0 u_ppwm/u_mem/_0111_
rlabel metal2 5088 21000 5088 21000 0 u_ppwm/u_mem/_0112_
rlabel metal2 1776 20748 1776 20748 0 u_ppwm/u_mem/_0113_
rlabel metal2 1248 22554 1248 22554 0 u_ppwm/u_mem/_0114_
rlabel metal2 9648 22260 9648 22260 0 u_ppwm/u_mem/_0115_
rlabel metal3 15312 20076 15312 20076 0 u_ppwm/u_mem/_0116_
rlabel metal2 13152 18816 13152 18816 0 u_ppwm/u_mem/_0117_
rlabel metal2 8928 17808 8928 17808 0 u_ppwm/u_mem/_0118_
rlabel metal2 1344 18858 1344 18858 0 u_ppwm/u_mem/_0119_
rlabel metal2 1536 17430 1536 17430 0 u_ppwm/u_mem/_0120_
rlabel metal2 6624 18354 6624 18354 0 u_ppwm/u_mem/_0121_
rlabel metal2 3552 15792 3552 15792 0 u_ppwm/u_mem/_0122_
rlabel metal2 1056 14070 1056 14070 0 u_ppwm/u_mem/_0123_
rlabel metal2 4320 12642 4320 12642 0 u_ppwm/u_mem/_0124_
rlabel metal2 5376 14070 5376 14070 0 u_ppwm/u_mem/_0125_
rlabel metal3 11952 19236 11952 19236 0 u_ppwm/u_mem/_0126_
rlabel metal2 8544 15792 8544 15792 0 u_ppwm/u_mem/_0127_
rlabel metal2 16416 19656 16416 19656 0 u_ppwm/u_mem/_0128_
rlabel metal2 14688 24612 14688 24612 0 u_ppwm/u_mem/_0129_
rlabel metal3 4848 23100 4848 23100 0 u_ppwm/u_mem/_0130_
rlabel metal2 2976 21630 2976 21630 0 u_ppwm/u_mem/_0131_
rlabel metal2 5328 19488 5328 19488 0 u_ppwm/u_mem/_0132_
rlabel metal2 8016 18564 8016 18564 0 u_ppwm/u_mem/_0133_
rlabel metal2 10944 17262 10944 17262 0 u_ppwm/u_mem/_0134_
rlabel metal3 10512 19488 10512 19488 0 u_ppwm/u_mem/_0135_
rlabel metal3 8160 19908 8160 19908 0 u_ppwm/u_mem/_0136_
rlabel metal3 4704 23268 4704 23268 0 u_ppwm/u_mem/_0137_
rlabel metal3 2448 23772 2448 23772 0 u_ppwm/u_mem/_0138_
rlabel metal2 4992 24402 4992 24402 0 u_ppwm/u_mem/_0139_
rlabel metal3 6864 23100 6864 23100 0 u_ppwm/u_mem/_0140_
rlabel metal2 12288 23352 12288 23352 0 u_ppwm/u_mem/_0141_
rlabel metal3 17856 20748 17856 20748 0 u_ppwm/u_mem/_0142_
rlabel metal2 20064 22764 20064 22764 0 u_ppwm/u_mem/_0143_
rlabel metal2 21408 27636 21408 27636 0 u_ppwm/u_mem/_0144_
rlabel metal2 20736 26292 20736 26292 0 u_ppwm/u_mem/_0145_
rlabel metal2 10752 26712 10752 26712 0 u_ppwm/u_mem/_0146_
rlabel metal2 11136 23520 11136 23520 0 u_ppwm/u_mem/_0147_
rlabel metal2 13632 25242 13632 25242 0 u_ppwm/u_mem/_0148_
rlabel metal2 19296 22974 19296 22974 0 u_ppwm/u_mem/_0149_
rlabel metal2 18912 24864 18912 24864 0 u_ppwm/u_mem/_0150_
rlabel metal2 20352 28266 20352 28266 0 u_ppwm/u_mem/_0151_
rlabel metal3 19680 28476 19680 28476 0 u_ppwm/u_mem/_0152_
rlabel metal2 9408 26628 9408 26628 0 u_ppwm/u_mem/_0153_
rlabel metal2 4608 26208 4608 26208 0 u_ppwm/u_mem/_0154_
rlabel metal2 3552 27552 3552 27552 0 u_ppwm/u_mem/_0155_
rlabel metal3 4032 27384 4032 27384 0 u_ppwm/u_mem/_0156_
rlabel metal2 8544 31290 8544 31290 0 u_ppwm/u_mem/_0157_
rlabel metal2 16512 31374 16512 31374 0 u_ppwm/u_mem/_0158_
rlabel metal2 20448 33138 20448 33138 0 u_ppwm/u_mem/_0159_
rlabel metal2 21120 31248 21120 31248 0 u_ppwm/u_mem/_0160_
rlabel metal3 8016 29064 8016 29064 0 u_ppwm/u_mem/_0161_
rlabel metal2 7488 28056 7488 28056 0 u_ppwm/u_mem/_0162_
rlabel metal2 3072 29610 3072 29610 0 u_ppwm/u_mem/_0163_
rlabel metal3 7248 31500 7248 31500 0 u_ppwm/u_mem/_0164_
rlabel metal2 12576 31290 12576 31290 0 u_ppwm/u_mem/_0165_
rlabel metal2 14976 32550 14976 32550 0 u_ppwm/u_mem/_0166_
rlabel metal2 13536 30702 13536 30702 0 u_ppwm/u_mem/_0167_
rlabel metal2 11904 30030 11904 30030 0 u_ppwm/u_mem/_0168_
rlabel metal3 3744 31416 3744 31416 0 u_ppwm/u_mem/_0169_
rlabel metal2 5184 31332 5184 31332 0 u_ppwm/u_mem/_0170_
rlabel metal2 7584 32634 7584 32634 0 u_ppwm/u_mem/_0171_
rlabel metal2 10944 34902 10944 34902 0 u_ppwm/u_mem/_0172_
rlabel metal2 12576 36414 12576 36414 0 u_ppwm/u_mem/_0173_
rlabel metal2 16800 35238 16800 35238 0 u_ppwm/u_mem/_0174_
rlabel metal2 13536 32970 13536 32970 0 u_ppwm/u_mem/_0175_
rlabel metal2 9936 31500 9936 31500 0 u_ppwm/u_mem/_0176_
rlabel metal2 2112 32172 2112 32172 0 u_ppwm/u_mem/_0177_
rlabel metal2 4704 33852 4704 33852 0 u_ppwm/u_mem/_0178_
rlabel metal2 9024 34356 9024 34356 0 u_ppwm/u_mem/_0179_
rlabel metal2 14592 34356 14592 34356 0 u_ppwm/u_mem/_0180_
rlabel metal2 18624 33978 18624 33978 0 u_ppwm/u_mem/_0181_
rlabel metal2 21600 33642 21600 33642 0 u_ppwm/u_mem/_0182_
rlabel metal2 24096 35070 24096 35070 0 u_ppwm/u_mem/_0183_
rlabel metal2 29568 35826 29568 35826 0 u_ppwm/u_mem/_0184_
rlabel metal2 33696 33642 33696 33642 0 u_ppwm/u_mem/_0185_
rlabel metal2 37728 33012 37728 33012 0 u_ppwm/u_mem/_0186_
rlabel metal2 38496 34104 38496 34104 0 u_ppwm/u_mem/_0187_
rlabel metal2 38688 35238 38688 35238 0 u_ppwm/u_mem/_0188_
rlabel metal2 26592 36204 26592 36204 0 u_ppwm/u_mem/_0189_
rlabel metal3 26448 35196 26448 35196 0 u_ppwm/u_mem/_0190_
rlabel metal3 32880 35280 32880 35280 0 u_ppwm/u_mem/_0191_
rlabel metal2 35328 35238 35328 35238 0 u_ppwm/u_mem/_0192_
rlabel metal2 40224 32424 40224 32424 0 u_ppwm/u_mem/_0193_
rlabel metal2 41952 32256 41952 32256 0 u_ppwm/u_mem/_0194_
rlabel metal2 40608 34398 40608 34398 0 u_ppwm/u_mem/_0195_
rlabel metal2 31392 30828 31392 30828 0 u_ppwm/u_mem/_0196_
rlabel metal3 29856 29316 29856 29316 0 u_ppwm/u_mem/_0197_
rlabel metal2 26208 31290 26208 31290 0 u_ppwm/u_mem/_0198_
rlabel metal2 28512 32592 28512 32592 0 u_ppwm/u_mem/_0199_
rlabel metal2 31584 30912 31584 30912 0 u_ppwm/u_mem/_0200_
rlabel metal3 34032 29148 34032 29148 0 u_ppwm/u_mem/_0201_
rlabel metal3 32496 29316 32496 29316 0 u_ppwm/u_mem/_0202_
rlabel metal2 29616 29148 29616 29148 0 u_ppwm/u_mem/_0203_
rlabel metal3 27984 29148 27984 29148 0 u_ppwm/u_mem/_0204_
rlabel metal2 24096 31836 24096 31836 0 u_ppwm/u_mem/_0205_
rlabel metal2 27840 31416 27840 31416 0 u_ppwm/u_mem/_0206_
rlabel metal2 31200 31752 31200 31752 0 u_ppwm/u_mem/_0207_
rlabel metal2 36000 29862 36000 29862 0 u_ppwm/u_mem/_0208_
rlabel metal2 37728 27300 37728 27300 0 u_ppwm/u_mem/_0209_
rlabel metal2 32736 25578 32736 25578 0 u_ppwm/u_mem/_0210_
rlabel metal3 36768 24528 36768 24528 0 u_ppwm/u_mem/_0211_
rlabel metal3 39120 28560 39120 28560 0 u_ppwm/u_mem/_0212_
rlabel metal2 42192 31584 42192 31584 0 u_ppwm/u_mem/_0213_
rlabel metal2 45024 28056 45024 28056 0 u_ppwm/u_mem/_0214_
rlabel metal3 45216 25284 45216 25284 0 u_ppwm/u_mem/_0215_
rlabel metal2 46032 23940 46032 23940 0 u_ppwm/u_mem/_0216_
rlabel metal2 41040 21336 41040 21336 0 u_ppwm/u_mem/_0217_
rlabel metal2 37824 21630 37824 21630 0 u_ppwm/u_mem/_0218_
rlabel metal2 39072 28602 39072 28602 0 u_ppwm/u_mem/_0219_
rlabel metal2 44832 31290 44832 31290 0 u_ppwm/u_mem/_0220_
rlabel metal2 47040 30534 47040 30534 0 u_ppwm/u_mem/_0221_
rlabel metal3 43680 28266 43680 28266 0 u_ppwm/u_mem/_0222_
rlabel metal2 44544 26208 44544 26208 0 u_ppwm/u_mem/_0223_
rlabel metal3 40512 22260 40512 22260 0 u_ppwm/u_mem/_0224_
rlabel metal2 37440 23562 37440 23562 0 u_ppwm/u_mem/_0225_
rlabel metal2 40992 23100 40992 23100 0 u_ppwm/u_mem/_0226_
rlabel metal2 49056 27090 49056 27090 0 u_ppwm/u_mem/_0227_
rlabel metal2 44544 28224 44544 28224 0 u_ppwm/u_mem/_0228_
rlabel metal2 48192 26292 48192 26292 0 u_ppwm/u_mem/_0229_
rlabel metal2 48288 24654 48288 24654 0 u_ppwm/u_mem/_0230_
rlabel metal3 44976 21588 44976 21588 0 u_ppwm/u_mem/_0231_
rlabel metal2 36768 23352 36768 23352 0 u_ppwm/u_mem/_0232_
rlabel metal2 41664 21294 41664 21294 0 u_ppwm/u_mem/_0233_
rlabel metal3 46800 28308 46800 28308 0 u_ppwm/u_mem/_0234_
rlabel metal2 48384 28350 48384 28350 0 u_ppwm/u_mem/_0235_
rlabel metal2 43680 27720 43680 27720 0 u_ppwm/u_mem/_0236_
rlabel metal2 42672 26124 42672 26124 0 u_ppwm/u_mem/_0237_
rlabel metal3 7200 16464 7200 16464 0 u_ppwm/u_mem/_0238_
rlabel metal2 8976 14700 8976 14700 0 u_ppwm/u_mem/_0239_
rlabel metal2 39216 25284 39216 25284 0 u_ppwm/u_mem/_0240_
rlabel metal2 40032 28184 40032 28184 0 u_ppwm/u_mem/_0241_
rlabel via2 24288 26964 24288 26964 0 u_ppwm/u_mem/_0242_
rlabel metal3 9120 14784 9120 14784 0 u_ppwm/u_mem/_0243_
rlabel metal3 7968 15708 7968 15708 0 u_ppwm/u_mem/_0244_
rlabel metal2 6624 15498 6624 15498 0 u_ppwm/u_mem/_0245_
rlabel metal2 6720 16674 6720 16674 0 u_ppwm/u_mem/_0246_
rlabel metal3 6432 14868 6432 14868 0 u_ppwm/u_mem/_0247_
rlabel metal2 7968 16926 7968 16926 0 u_ppwm/u_mem/_0248_
rlabel metal2 7248 15540 7248 15540 0 u_ppwm/u_mem/_0249_
rlabel metal2 8112 16464 8112 16464 0 u_ppwm/u_mem/_0250_
rlabel metal2 14592 27300 14592 27300 0 u_ppwm/u_mem/_0251_
rlabel metal2 17280 33432 17280 33432 0 u_ppwm/u_mem/_0252_
rlabel metal2 14688 26292 14688 26292 0 u_ppwm/u_mem/_0253_
rlabel metal2 14784 26544 14784 26544 0 u_ppwm/u_mem/_0254_
rlabel metal2 12288 27678 12288 27678 0 u_ppwm/u_mem/_0255_
rlabel metal2 14592 26334 14592 26334 0 u_ppwm/u_mem/_0256_
rlabel metal2 12576 26040 12576 26040 0 u_ppwm/u_mem/_0257_
rlabel metal2 14400 26040 14400 26040 0 u_ppwm/u_mem/_0258_
rlabel metal2 30912 25872 30912 25872 0 u_ppwm/u_mem/_0259_
rlabel metal2 39888 24780 39888 24780 0 u_ppwm/u_mem/_0260_
rlabel metal3 34080 25914 34080 25914 0 u_ppwm/u_mem/_0261_
rlabel metal3 31728 27804 31728 27804 0 u_ppwm/u_mem/_0262_
rlabel metal2 31920 27636 31920 27636 0 u_ppwm/u_mem/_0263_
rlabel metal3 31536 26796 31536 26796 0 u_ppwm/u_mem/_0264_
rlabel metal2 31200 27048 31200 27048 0 u_ppwm/u_mem/_0265_
rlabel metal2 31104 26376 31104 26376 0 u_ppwm/u_mem/_0266_
rlabel metal3 14496 24486 14496 24486 0 u_ppwm/u_mem/_0267_
rlabel metal2 17136 26796 17136 26796 0 u_ppwm/u_mem/_0268_
rlabel metal2 18240 26166 18240 26166 0 u_ppwm/u_mem/_0269_
rlabel metal2 17952 25830 17952 25830 0 u_ppwm/u_mem/_0270_
rlabel metal2 17712 31500 17712 31500 0 u_ppwm/u_mem/_0271_
rlabel metal2 18432 26250 18432 26250 0 u_ppwm/u_mem/_0272_
rlabel metal2 25824 26040 25824 26040 0 u_ppwm/u_mem/_0273_
rlabel metal2 38400 27678 38400 27678 0 u_ppwm/u_mem/_0274_
rlabel metal2 40800 26208 40800 26208 0 u_ppwm/u_mem/_0275_
rlabel metal2 40416 34650 40416 34650 0 u_ppwm/u_mem/_0276_
rlabel metal2 40368 34188 40368 34188 0 u_ppwm/u_mem/_0277_
rlabel metal2 44352 26040 44352 26040 0 u_ppwm/u_mem/_0278_
rlabel metal3 39840 26166 39840 26166 0 u_ppwm/u_mem/_0279_
rlabel metal2 42384 25536 42384 25536 0 u_ppwm/u_mem/_0280_
rlabel metal3 41280 26124 41280 26124 0 u_ppwm/u_mem/_0281_
rlabel metal5 29512 26166 29512 26166 0 u_ppwm/u_mem/_0282_
rlabel metal2 14976 23898 14976 23898 0 u_ppwm/u_mem/_0283_
rlabel metal2 15168 26922 15168 26922 0 u_ppwm/u_mem/_0284_
rlabel metal3 17952 27636 17952 27636 0 u_ppwm/u_mem/_0285_
rlabel metal2 15325 27502 15325 27502 0 u_ppwm/u_mem/_0286_
rlabel metal2 13344 30744 13344 30744 0 u_ppwm/u_mem/_0287_
rlabel metal3 14160 29652 14160 29652 0 u_ppwm/u_mem/_0288_
rlabel metal2 14256 29652 14256 29652 0 u_ppwm/u_mem/_0289_
rlabel metal3 14640 27048 14640 27048 0 u_ppwm/u_mem/_0290_
rlabel metal3 14784 27342 14784 27342 0 u_ppwm/u_mem/_0291_
rlabel metal2 37632 30114 37632 30114 0 u_ppwm/u_mem/_0292_
rlabel metal2 41424 28308 41424 28308 0 u_ppwm/u_mem/_0293_
rlabel metal2 41760 30828 41760 30828 0 u_ppwm/u_mem/_0294_
rlabel metal3 41376 29736 41376 29736 0 u_ppwm/u_mem/_0295_
rlabel metal3 42624 29064 42624 29064 0 u_ppwm/u_mem/_0296_
rlabel metal3 41952 28308 41952 28308 0 u_ppwm/u_mem/_0297_
rlabel metal2 43872 27678 43872 27678 0 u_ppwm/u_mem/_0298_
rlabel metal2 40992 28014 40992 28014 0 u_ppwm/u_mem/_0299_
rlabel metal2 39840 27636 39840 27636 0 u_ppwm/u_mem/_0300_
rlabel metal3 11664 22512 11664 22512 0 u_ppwm/u_mem/_0301_
rlabel metal2 14016 27537 14016 27537 0 u_ppwm/u_mem/_0302_
rlabel metal3 17328 26796 17328 26796 0 u_ppwm/u_mem/_0303_
rlabel metal2 15024 27048 15024 27048 0 u_ppwm/u_mem/_0304_
rlabel metal3 13440 29820 13440 29820 0 u_ppwm/u_mem/_0305_
rlabel via1 13920 27634 13920 27634 0 u_ppwm/u_mem/_0306_
rlabel metal2 12768 32802 12768 32802 0 u_ppwm/u_mem/_0307_
rlabel metal3 13296 27636 13296 27636 0 u_ppwm/u_mem/_0308_
rlabel metal2 30336 26838 30336 26838 0 u_ppwm/u_mem/_0309_
rlabel metal2 31584 28182 31584 28182 0 u_ppwm/u_mem/_0310_
rlabel metal2 36864 27342 36864 27342 0 u_ppwm/u_mem/_0311_
rlabel metal2 31536 27048 31536 27048 0 u_ppwm/u_mem/_0312_
rlabel metal2 30432 27233 30432 27233 0 u_ppwm/u_mem/_0313_
rlabel metal2 30816 27468 30816 27468 0 u_ppwm/u_mem/_0314_
rlabel metal2 30528 27090 30528 27090 0 u_ppwm/u_mem/_0315_
rlabel metal2 14304 25368 14304 25368 0 u_ppwm/u_mem/_0316_
rlabel metal2 16608 26040 16608 26040 0 u_ppwm/u_mem/_0317_
rlabel metal2 17184 24864 17184 24864 0 u_ppwm/u_mem/_0318_
rlabel metal2 17472 25620 17472 25620 0 u_ppwm/u_mem/_0319_
rlabel metal2 16032 26250 16032 26250 0 u_ppwm/u_mem/_0320_
rlabel metal2 16320 26124 16320 26124 0 u_ppwm/u_mem/_0321_
rlabel metal2 16416 25326 16416 25326 0 u_ppwm/u_mem/_0322_
rlabel metal2 38688 27468 38688 27468 0 u_ppwm/u_mem/_0323_
rlabel metal3 29280 26796 29280 26796 0 u_ppwm/u_mem/_0324_
rlabel metal4 41280 25788 41280 25788 0 u_ppwm/u_mem/_0325_
rlabel metal2 29472 26292 29472 26292 0 u_ppwm/u_mem/_0326_
rlabel metal3 30528 29148 30528 29148 0 u_ppwm/u_mem/_0327_
rlabel metal2 30432 28602 30432 28602 0 u_ppwm/u_mem/_0328_
rlabel metal2 28272 30408 28272 30408 0 u_ppwm/u_mem/_0329_
rlabel metal3 28512 28182 28512 28182 0 u_ppwm/u_mem/_0330_
rlabel metal2 28320 27426 28320 27426 0 u_ppwm/u_mem/_0331_
rlabel via2 28128 24851 28128 24851 0 u_ppwm/u_mem/_0332_
rlabel metal2 15744 24528 15744 24528 0 u_ppwm/u_mem/_0333_
rlabel metal3 15456 24612 15456 24612 0 u_ppwm/u_mem/_0334_
rlabel metal2 14784 23604 14784 23604 0 u_ppwm/u_mem/_0335_
rlabel metal2 16704 24528 16704 24528 0 u_ppwm/u_mem/_0336_
rlabel metal2 16512 24696 16512 24696 0 u_ppwm/u_mem/_0337_
rlabel metal3 16224 24612 16224 24612 0 u_ppwm/u_mem/_0338_
rlabel metal2 15408 27720 15408 27720 0 u_ppwm/u_mem/_0339_
rlabel metal2 15456 25704 15456 25704 0 u_ppwm/u_mem/_0340_
rlabel metal2 16224 24822 16224 24822 0 u_ppwm/u_mem/_0341_
rlabel metal2 28032 29694 28032 29694 0 u_ppwm/u_mem/_0342_
rlabel metal3 28560 34020 28560 34020 0 u_ppwm/u_mem/_0343_
rlabel metal2 35328 28014 35328 28014 0 u_ppwm/u_mem/_0344_
rlabel metal4 28608 25200 28608 25200 0 u_ppwm/u_mem/_0345_
rlabel metal2 24480 27258 24480 27258 0 u_ppwm/u_mem/_0346_
rlabel metal2 23904 26418 23904 26418 0 u_ppwm/u_mem/_0347_
rlabel metal2 10272 24696 10272 24696 0 u_ppwm/u_mem/_0348_
rlabel metal2 13536 25494 13536 25494 0 u_ppwm/u_mem/_0349_
rlabel metal3 13632 28476 13632 28476 0 u_ppwm/u_mem/_0350_
rlabel via1 13378 26120 13378 26120 0 u_ppwm/u_mem/_0351_
rlabel metal2 13152 24486 13152 24486 0 u_ppwm/u_mem/_0352_
rlabel metal2 11616 25200 11616 25200 0 u_ppwm/u_mem/_0353_
rlabel metal3 13632 26082 13632 26082 0 u_ppwm/u_mem/_0354_
rlabel metal2 13344 25116 13344 25116 0 u_ppwm/u_mem/_0355_
rlabel metal3 17040 25872 17040 25872 0 u_ppwm/u_mem/_0356_
rlabel metal2 26928 29988 26928 29988 0 u_ppwm/u_mem/_0357_
rlabel metal2 27072 30114 27072 30114 0 u_ppwm/u_mem/_0358_
rlabel metal2 26496 28602 26496 28602 0 u_ppwm/u_mem/_0359_
rlabel metal2 27648 26163 27648 26163 0 u_ppwm/u_mem/_0360_
rlabel metal3 34080 24612 34080 24612 0 u_ppwm/u_mem/_0361_
rlabel metal2 28368 24780 28368 24780 0 u_ppwm/u_mem/_0362_
rlabel metal2 43680 25284 43680 25284 0 u_ppwm/u_mem/_0363_
rlabel metal2 43584 26964 43584 26964 0 u_ppwm/u_mem/_0364_
rlabel metal2 48144 30660 48144 30660 0 u_ppwm/u_mem/_0365_
rlabel metal3 48000 28140 48000 28140 0 u_ppwm/u_mem/_0366_
rlabel metal2 41952 21840 41952 21840 0 u_ppwm/u_mem/_0367_
rlabel metal3 35904 23100 35904 23100 0 u_ppwm/u_mem/_0368_
rlabel metal2 45120 21588 45120 21588 0 u_ppwm/u_mem/_0369_
rlabel metal2 47856 24612 47856 24612 0 u_ppwm/u_mem/_0370_
rlabel metal2 47808 26124 47808 26124 0 u_ppwm/u_mem/_0371_
rlabel metal3 45696 27636 45696 27636 0 u_ppwm/u_mem/_0372_
rlabel metal2 49344 26754 49344 26754 0 u_ppwm/u_mem/_0373_
rlabel metal2 41664 23100 41664 23100 0 u_ppwm/u_mem/_0374_
rlabel metal3 37968 23772 37968 23772 0 u_ppwm/u_mem/_0375_
rlabel metal2 39504 22260 39504 22260 0 u_ppwm/u_mem/_0376_
rlabel metal2 48480 24906 48480 24906 0 u_ppwm/u_mem/_0377_
rlabel metal3 48576 27636 48576 27636 0 u_ppwm/u_mem/_0378_
rlabel metal2 47424 30660 47424 30660 0 u_ppwm/u_mem/_0379_
rlabel metal3 45360 31332 45360 31332 0 u_ppwm/u_mem/_0380_
rlabel metal3 38736 30660 38736 30660 0 u_ppwm/u_mem/_0381_
rlabel metal3 35664 26628 35664 26628 0 u_ppwm/u_mem/_0382_
rlabel metal2 38592 21672 38592 21672 0 u_ppwm/u_mem/_0383_
rlabel metal2 44688 24780 44688 24780 0 u_ppwm/u_mem/_0384_
rlabel metal2 44160 25032 44160 25032 0 u_ppwm/u_mem/_0385_
rlabel metal2 43536 29652 43536 29652 0 u_ppwm/u_mem/_0386_
rlabel metal2 42816 32172 42816 32172 0 u_ppwm/u_mem/_0387_
rlabel metal2 38640 29820 38640 29820 0 u_ppwm/u_mem/_0388_
rlabel metal2 35616 24906 35616 24906 0 u_ppwm/u_mem/_0389_
rlabel metal3 33552 25284 33552 25284 0 u_ppwm/u_mem/_0390_
rlabel metal2 34176 26880 34176 26880 0 u_ppwm/u_mem/_0391_
rlabel metal2 37440 28518 37440 28518 0 u_ppwm/u_mem/_0392_
rlabel metal2 33600 31416 33600 31416 0 u_ppwm/u_mem/_0393_
rlabel metal2 28128 32004 28128 32004 0 u_ppwm/u_mem/_0394_
rlabel metal2 27648 31458 27648 31458 0 u_ppwm/u_mem/_0395_
rlabel metal3 26928 29148 26928 29148 0 u_ppwm/u_mem/_0396_
rlabel metal2 29184 29736 29184 29736 0 u_ppwm/u_mem/_0397_
rlabel metal3 31200 28308 31200 28308 0 u_ppwm/u_mem/_0398_
rlabel metal2 33504 29610 33504 29610 0 u_ppwm/u_mem/_0399_
rlabel metal3 34896 30660 34896 30660 0 u_ppwm/u_mem/_0400_
rlabel metal3 30336 30828 30336 30828 0 u_ppwm/u_mem/_0401_
rlabel metal2 25920 32004 25920 32004 0 u_ppwm/u_mem/_0402_
rlabel metal2 27936 29211 27936 29211 0 u_ppwm/u_mem/_0403_
rlabel metal2 31920 32340 31920 32340 0 u_ppwm/u_mem/_0404_
rlabel metal2 39744 34356 39744 34356 0 u_ppwm/u_mem/_0405_
rlabel metal2 42240 32634 42240 32634 0 u_ppwm/u_mem/_0406_
rlabel metal2 41568 33600 41568 33600 0 u_ppwm/u_mem/_0407_
rlabel metal2 36384 33894 36384 33894 0 u_ppwm/u_mem/_0408_
rlabel metal2 30144 34734 30144 34734 0 u_ppwm/u_mem/_0409_
rlabel metal2 27360 34776 27360 34776 0 u_ppwm/u_mem/_0410_
rlabel metal2 25440 34398 25440 34398 0 u_ppwm/u_mem/_0411_
rlabel metal2 38352 35280 38352 35280 0 u_ppwm/u_mem/_0412_
rlabel metal2 39216 34356 39216 34356 0 u_ppwm/u_mem/_0413_
rlabel metal2 38352 33684 38352 33684 0 u_ppwm/u_mem/_0414_
rlabel metal2 34080 33684 34080 33684 0 u_ppwm/u_mem/_0415_
rlabel metal3 30144 35196 30144 35196 0 u_ppwm/u_mem/_0416_
rlabel metal2 26016 36708 26016 36708 0 u_ppwm/u_mem/_0417_
rlabel metal3 21504 33684 21504 33684 0 u_ppwm/u_mem/_0418_
rlabel metal2 18912 33936 18912 33936 0 u_ppwm/u_mem/_0419_
rlabel metal2 14976 34440 14976 34440 0 u_ppwm/u_mem/_0420_
rlabel metal2 9408 34272 9408 34272 0 u_ppwm/u_mem/_0421_
rlabel metal2 6336 33936 6336 33936 0 u_ppwm/u_mem/_0422_
rlabel metal2 2496 32844 2496 32844 0 u_ppwm/u_mem/_0423_
rlabel metal2 4416 32844 4416 32844 0 u_ppwm/u_mem/_0424_
rlabel metal3 13248 32844 13248 32844 0 u_ppwm/u_mem/_0425_
rlabel metal3 15552 35196 15552 35196 0 u_ppwm/u_mem/_0426_
rlabel metal2 12960 34692 12960 34692 0 u_ppwm/u_mem/_0427_
rlabel metal2 11904 34482 11904 34482 0 u_ppwm/u_mem/_0428_
rlabel metal2 4896 33810 4896 33810 0 u_ppwm/u_mem/_0429_
rlabel metal2 5616 31332 5616 31332 0 u_ppwm/u_mem/_0430_
rlabel metal2 4416 31332 4416 31332 0 u_ppwm/u_mem/_0431_
rlabel metal2 11520 30240 11520 30240 0 u_ppwm/u_mem/_0432_
rlabel metal2 14496 30240 14496 30240 0 u_ppwm/u_mem/_0433_
rlabel metal2 15168 33348 15168 33348 0 u_ppwm/u_mem/_0434_
rlabel metal3 12528 31332 12528 31332 0 u_ppwm/u_mem/_0435_
rlabel metal2 8016 32340 8016 32340 0 u_ppwm/u_mem/_0436_
rlabel metal2 2784 29211 2784 29211 0 u_ppwm/u_mem/_0437_
rlabel metal2 4032 28980 4032 28980 0 u_ppwm/u_mem/_0438_
rlabel metal2 7008 28308 7008 28308 0 u_ppwm/u_mem/_0439_
rlabel metal2 20832 30576 20832 30576 0 u_ppwm/u_mem/_0440_
rlabel metal2 18240 32592 18240 32592 0 u_ppwm/u_mem/_0441_
rlabel metal2 16752 31332 16752 31332 0 u_ppwm/u_mem/_0442_
rlabel metal2 7872 30030 7872 30030 0 u_ppwm/u_mem/_0443_
rlabel metal2 5376 29232 5376 29232 0 u_ppwm/u_mem/_0444_
rlabel metal2 3840 26376 3840 26376 0 u_ppwm/u_mem/_0445_
rlabel metal2 4176 25284 4176 25284 0 u_ppwm/u_mem/_0446_
rlabel metal2 9120 26292 9120 26292 0 u_ppwm/u_mem/_0447_
rlabel metal2 19008 28602 19008 28602 0 u_ppwm/u_mem/_0448_
rlabel metal2 19968 28308 19968 28308 0 u_ppwm/u_mem/_0449_
rlabel metal2 18672 24612 18672 24612 0 u_ppwm/u_mem/_0450_
rlabel metal2 16704 23604 16704 23604 0 u_ppwm/u_mem/_0451_
rlabel metal3 14544 23688 14544 23688 0 u_ppwm/u_mem/_0452_
rlabel metal3 14112 24570 14112 24570 0 u_ppwm/u_mem/_0453_
rlabel metal2 12480 26838 12480 26838 0 u_ppwm/u_mem/_0454_
rlabel metal2 20352 26880 20352 26880 0 u_ppwm/u_mem/_0455_
rlabel metal2 20976 27636 20976 27636 0 u_ppwm/u_mem/_0456_
rlabel metal2 19488 23772 19488 23772 0 u_ppwm/u_mem/_0457_
rlabel metal2 17040 20748 17040 20748 0 u_ppwm/u_mem/_0458_
rlabel metal2 13536 22680 13536 22680 0 u_ppwm/u_mem/_0459_
rlabel metal3 7824 23100 7824 23100 0 u_ppwm/u_mem/_0460_
rlabel metal2 5184 24192 5184 24192 0 u_ppwm/u_mem/_0461_
rlabel metal2 2880 24444 2880 24444 0 u_ppwm/u_mem/_0462_
rlabel metal3 4512 23688 4512 23688 0 u_ppwm/u_mem/_0463_
rlabel metal2 6768 20076 6768 20076 0 u_ppwm/u_mem/_0464_
rlabel metal3 10128 20748 10128 20748 0 u_ppwm/u_mem/_0465_
rlabel metal2 12000 16212 12000 16212 0 u_ppwm/u_mem/_0466_
rlabel metal2 7680 18690 7680 18690 0 u_ppwm/u_mem/_0467_
rlabel metal2 4512 21672 4512 21672 0 u_ppwm/u_mem/_0468_
rlabel metal3 3264 21588 3264 21588 0 u_ppwm/u_mem/_0469_
rlabel metal2 3936 23310 3936 23310 0 u_ppwm/u_mem/_0470_
rlabel metal2 9600 23100 9600 23100 0 u_ppwm/u_mem/_0471_
rlabel metal3 15408 20748 15408 20748 0 u_ppwm/u_mem/_0472_
rlabel metal3 13632 18732 13632 18732 0 u_ppwm/u_mem/_0473_
rlabel metal3 9504 17724 9504 17724 0 u_ppwm/u_mem/_0474_
rlabel metal2 5808 16212 5808 16212 0 u_ppwm/u_mem/_0475_
rlabel metal3 3072 14700 3072 14700 0 u_ppwm/u_mem/_0476_
rlabel metal2 5184 16044 5184 16044 0 u_ppwm/u_mem/_0477_
rlabel metal3 3840 17136 3840 17136 0 u_ppwm/u_mem/_0478_
rlabel metal2 3840 17010 3840 17010 0 u_ppwm/u_mem/_0479_
rlabel metal2 3936 17262 3936 17262 0 u_ppwm/u_mem/_0480_
rlabel metal3 5040 16380 5040 16380 0 u_ppwm/u_mem/_0481_
rlabel metal3 5424 16800 5424 16800 0 u_ppwm/u_mem/_0482_
rlabel metal2 3648 16170 3648 16170 0 u_ppwm/u_mem/_0483_
rlabel metal2 3840 14826 3840 14826 0 u_ppwm/u_mem/_0484_
rlabel metal3 3408 12432 3408 12432 0 u_ppwm/u_mem/_0485_
rlabel metal3 4704 14868 4704 14868 0 u_ppwm/u_mem/_0486_
rlabel metal2 5568 14952 5568 14952 0 u_ppwm/u_mem/_0487_
rlabel metal3 6336 14952 6336 14952 0 u_ppwm/u_mem/_0488_
rlabel metal3 6144 12600 6144 12600 0 u_ppwm/u_mem/_0489_
rlabel metal2 5184 13524 5184 13524 0 u_ppwm/u_mem/_0490_
rlabel metal2 3744 18942 3744 18942 0 u_ppwm/u_mem/bit_count\[0\]
rlabel metal2 3936 18270 3936 18270 0 u_ppwm/u_mem/bit_count\[1\]
rlabel metal2 7680 17304 7680 17304 0 u_ppwm/u_mem/bit_count\[2\]
rlabel metal2 4416 14910 4416 14910 0 u_ppwm/u_mem/bit_count\[3\]
rlabel metal3 3936 14700 3936 14700 0 u_ppwm/u_mem/bit_count\[4\]
rlabel metal2 5616 13440 5616 13440 0 u_ppwm/u_mem/bit_count\[5\]
rlabel metal2 7920 14196 7920 14196 0 u_ppwm/u_mem/bit_count\[6\]
rlabel metal2 41472 24780 41472 24780 0 u_ppwm/u_mem/memory\[0\]
rlabel metal3 3936 23772 3936 23772 0 u_ppwm/u_mem/memory\[100\]
rlabel metal3 9984 21756 9984 21756 0 u_ppwm/u_mem/memory\[101\]
rlabel metal3 13440 21420 13440 21420 0 u_ppwm/u_mem/memory\[102\]
rlabel metal2 14016 18522 14016 18522 0 u_ppwm/u_mem/memory\[103\]
rlabel metal3 11760 20076 11760 20076 0 u_ppwm/u_mem/memory\[104\]
rlabel metal2 6864 20748 6864 20748 0 u_ppwm/u_mem/memory\[105\]
rlabel metal2 4176 21000 4176 21000 0 u_ppwm/u_mem/memory\[106\]
rlabel metal3 4608 22260 4608 22260 0 u_ppwm/u_mem/memory\[107\]
rlabel metal3 49968 27552 49968 27552 0 u_ppwm/u_mem/memory\[10\]
rlabel metal2 44736 23226 44736 23226 0 u_ppwm/u_mem/memory\[11\]
rlabel metal2 40800 23520 40800 23520 0 u_ppwm/u_mem/memory\[12\]
rlabel metal2 41568 21504 41568 21504 0 u_ppwm/u_mem/memory\[13\]
rlabel metal3 43806 24528 43806 24528 0 u_ppwm/u_mem/memory\[14\]
rlabel metal2 51648 26376 51648 26376 0 u_ppwm/u_mem/memory\[15\]
rlabel metal3 49104 32172 49104 32172 0 u_ppwm/u_mem/memory\[16\]
rlabel metal3 47424 32340 47424 32340 0 u_ppwm/u_mem/memory\[17\]
rlabel metal3 41040 31164 41040 31164 0 u_ppwm/u_mem/memory\[18\]
rlabel metal2 38976 27720 38976 27720 0 u_ppwm/u_mem/memory\[19\]
rlabel metal2 45024 26838 45024 26838 0 u_ppwm/u_mem/memory\[1\]
rlabel metal2 37536 22008 37536 22008 0 u_ppwm/u_mem/memory\[20\]
rlabel metal2 40512 24528 40512 24528 0 u_ppwm/u_mem/memory\[21\]
rlabel metal2 47232 25830 47232 25830 0 u_ppwm/u_mem/memory\[22\]
rlabel metal3 47376 29988 47376 29988 0 u_ppwm/u_mem/memory\[23\]
rlabel metal2 44640 31416 44640 31416 0 u_ppwm/u_mem/memory\[24\]
rlabel metal2 42144 29862 42144 29862 0 u_ppwm/u_mem/memory\[25\]
rlabel metal2 34848 25326 34848 25326 0 u_ppwm/u_mem/memory\[26\]
rlabel metal3 34752 25284 34752 25284 0 u_ppwm/u_mem/memory\[27\]
rlabel metal2 32832 27342 32832 27342 0 u_ppwm/u_mem/memory\[28\]
rlabel metal3 38064 28308 38064 28308 0 u_ppwm/u_mem/memory\[29\]
rlabel metal3 47952 30240 47952 30240 0 u_ppwm/u_mem/memory\[2\]
rlabel metal3 34272 32340 34272 32340 0 u_ppwm/u_mem/memory\[30\]
rlabel metal2 28032 33642 28032 33642 0 u_ppwm/u_mem/memory\[31\]
rlabel metal2 26400 32508 26400 32508 0 u_ppwm/u_mem/memory\[32\]
rlabel metal3 26352 30828 26352 30828 0 u_ppwm/u_mem/memory\[33\]
rlabel metal2 30624 30702 30624 30702 0 u_ppwm/u_mem/memory\[34\]
rlabel metal3 31872 28560 31872 28560 0 u_ppwm/u_mem/memory\[35\]
rlabel metal2 36048 28812 36048 28812 0 u_ppwm/u_mem/memory\[36\]
rlabel metal2 37056 30912 37056 30912 0 u_ppwm/u_mem/memory\[37\]
rlabel metal3 31152 31164 31152 31164 0 u_ppwm/u_mem/memory\[38\]
rlabel metal2 27984 32172 27984 32172 0 u_ppwm/u_mem/memory\[39\]
rlabel metal3 49824 29148 49824 29148 0 u_ppwm/u_mem/memory\[3\]
rlabel metal3 24960 30660 24960 30660 0 u_ppwm/u_mem/memory\[40\]
rlabel metal2 33504 32424 33504 32424 0 u_ppwm/u_mem/memory\[41\]
rlabel metal2 36960 35154 36960 35154 0 u_ppwm/u_mem/memory\[42\]
rlabel metal2 45984 34524 45984 34524 0 u_ppwm/u_mem/memory\[43\]
rlabel metal2 44160 33138 44160 33138 0 u_ppwm/u_mem/memory\[44\]
rlabel metal2 37344 33432 37344 33432 0 u_ppwm/u_mem/memory\[45\]
rlabel metal2 29952 34272 29952 34272 0 u_ppwm/u_mem/memory\[46\]
rlabel metal3 30144 36120 30144 36120 0 u_ppwm/u_mem/memory\[47\]
rlabel metal2 25824 35280 25824 35280 0 u_ppwm/u_mem/memory\[48\]
rlabel metal2 32256 37380 32256 37380 0 u_ppwm/u_mem/memory\[49\]
rlabel metal2 44592 22344 44592 22344 0 u_ppwm/u_mem/memory\[4\]
rlabel metal2 40320 35154 40320 35154 0 u_ppwm/u_mem/memory\[50\]
rlabel metal2 40512 32886 40512 32886 0 u_ppwm/u_mem/memory\[51\]
rlabel metal2 36864 33936 36864 33936 0 u_ppwm/u_mem/memory\[52\]
rlabel metal3 31344 35700 31344 35700 0 u_ppwm/u_mem/memory\[53\]
rlabel metal2 28032 35742 28032 35742 0 u_ppwm/u_mem/memory\[54\]
rlabel metal3 22560 34188 22560 34188 0 u_ppwm/u_mem/memory\[55\]
rlabel metal2 19392 34461 19392 34461 0 u_ppwm/u_mem/memory\[56\]
rlabel via2 19008 34343 19008 34343 0 u_ppwm/u_mem/memory\[57\]
rlabel metal2 13824 35154 13824 35154 0 u_ppwm/u_mem/memory\[58\]
rlabel metal2 8352 34902 8352 34902 0 u_ppwm/u_mem/memory\[59\]
rlabel metal2 36864 22806 36864 22806 0 u_ppwm/u_mem/memory\[5\]
rlabel metal2 6048 33642 6048 33642 0 u_ppwm/u_mem/memory\[60\]
rlabel via1 4800 32184 4800 32184 0 u_ppwm/u_mem/memory\[61\]
rlabel metal2 11808 31794 11808 31794 0 u_ppwm/u_mem/memory\[62\]
rlabel metal2 17712 35700 17712 35700 0 u_ppwm/u_mem/memory\[63\]
rlabel metal2 15456 34902 15456 34902 0 u_ppwm/u_mem/memory\[64\]
rlabel metal2 12960 35448 12960 35448 0 u_ppwm/u_mem/memory\[65\]
rlabel metal2 9024 33810 9024 33810 0 u_ppwm/u_mem/memory\[66\]
rlabel metal2 7440 31920 7440 31920 0 u_ppwm/u_mem/memory\[67\]
rlabel metal3 4368 29904 4368 29904 0 u_ppwm/u_mem/memory\[68\]
rlabel metal2 13536 30072 13536 30072 0 u_ppwm/u_mem/memory\[69\]
rlabel metal3 44400 22932 44400 22932 0 u_ppwm/u_mem/memory\[6\]
rlabel metal2 14688 29484 14688 29484 0 u_ppwm/u_mem/memory\[70\]
rlabel metal3 17952 32928 17952 32928 0 u_ppwm/u_mem/memory\[71\]
rlabel metal2 14304 32592 14304 32592 0 u_ppwm/u_mem/memory\[72\]
rlabel metal2 12384 30828 12384 30828 0 u_ppwm/u_mem/memory\[73\]
rlabel metal2 6624 30618 6624 30618 0 u_ppwm/u_mem/memory\[74\]
rlabel metal3 4512 29820 4512 29820 0 u_ppwm/u_mem/memory\[75\]
rlabel metal2 6720 28182 6720 28182 0 u_ppwm/u_mem/memory\[76\]
rlabel metal2 18720 29988 18720 29988 0 u_ppwm/u_mem/memory\[77\]
rlabel metal2 19344 32172 19344 32172 0 u_ppwm/u_mem/memory\[78\]
rlabel metal2 15840 32130 15840 32130 0 u_ppwm/u_mem/memory\[79\]
rlabel metal2 41088 24402 41088 24402 0 u_ppwm/u_mem/memory\[7\]
rlabel metal2 12576 29904 12576 29904 0 u_ppwm/u_mem/memory\[80\]
rlabel metal3 5904 29316 5904 29316 0 u_ppwm/u_mem/memory\[81\]
rlabel metal2 5184 27678 5184 27678 0 u_ppwm/u_mem/memory\[82\]
rlabel metal2 4656 26796 4656 26796 0 u_ppwm/u_mem/memory\[83\]
rlabel metal2 8736 27552 8736 27552 0 u_ppwm/u_mem/memory\[84\]
rlabel metal2 16608 28602 16608 28602 0 u_ppwm/u_mem/memory\[85\]
rlabel metal2 20064 27720 20064 27720 0 u_ppwm/u_mem/memory\[86\]
rlabel metal3 19296 26712 19296 26712 0 u_ppwm/u_mem/memory\[87\]
rlabel metal2 19728 24612 19728 24612 0 u_ppwm/u_mem/memory\[88\]
rlabel metal2 15744 23688 15744 23688 0 u_ppwm/u_mem/memory\[89\]
rlabel metal2 42528 25620 42528 25620 0 u_ppwm/u_mem/memory\[8\]
rlabel metal2 12528 24024 12528 24024 0 u_ppwm/u_mem/memory\[90\]
rlabel metal2 11712 25998 11712 25998 0 u_ppwm/u_mem/memory\[91\]
rlabel metal2 18720 26628 18720 26628 0 u_ppwm/u_mem/memory\[92\]
rlabel metal2 23424 28014 23424 28014 0 u_ppwm/u_mem/memory\[93\]
rlabel metal2 19488 26712 19488 26712 0 u_ppwm/u_mem/memory\[94\]
rlabel metal2 17472 23856 17472 23856 0 u_ppwm/u_mem/memory\[95\]
rlabel metal2 15552 21756 15552 21756 0 u_ppwm/u_mem/memory\[96\]
rlabel metal2 11424 23226 11424 23226 0 u_ppwm/u_mem/memory\[97\]
rlabel metal2 7488 24318 7488 24318 0 u_ppwm/u_mem/memory\[98\]
rlabel metal2 4512 24570 4512 24570 0 u_ppwm/u_mem/memory\[99\]
rlabel metal2 44544 27342 44544 27342 0 u_ppwm/u_mem/memory\[9\]
rlabel metal2 11712 16002 11712 16002 0 u_ppwm/u_mem/state_q\[0\]
rlabel metal2 11712 16464 11712 16464 0 u_ppwm/u_mem/state_q\[2\]
rlabel metal2 8352 12474 8352 12474 0 u_ppwm/u_pwm/_000_
rlabel metal2 10464 12516 10464 12516 0 u_ppwm/u_pwm/_001_
rlabel metal2 8928 8232 8928 8232 0 u_ppwm/u_pwm/_002_
rlabel metal2 9504 9912 9504 9912 0 u_ppwm/u_pwm/_003_
rlabel metal2 15840 8946 15840 8946 0 u_ppwm/u_pwm/_004_
rlabel metal3 15504 6636 15504 6636 0 u_ppwm/u_pwm/_005_
rlabel metal2 12672 9408 12672 9408 0 u_ppwm/u_pwm/_006_
rlabel metal2 10560 10920 10560 10920 0 u_ppwm/u_pwm/_007_
rlabel metal2 16800 4872 16800 4872 0 u_ppwm/u_pwm/_008_
rlabel metal2 16320 3864 16320 3864 0 u_ppwm/u_pwm/_009_
rlabel metal2 3456 8736 3456 8736 0 u_ppwm/u_pwm/_010_
rlabel metal2 4512 7896 4512 7896 0 u_ppwm/u_pwm/_011_
rlabel metal2 5568 5712 5568 5712 0 u_ppwm/u_pwm/_012_
rlabel metal3 5808 2688 5808 2688 0 u_ppwm/u_pwm/_013_
rlabel metal2 5376 4872 5376 4872 0 u_ppwm/u_pwm/_014_
rlabel metal2 8544 3486 8544 3486 0 u_ppwm/u_pwm/_015_
rlabel metal3 10128 1932 10128 1932 0 u_ppwm/u_pwm/_016_
rlabel metal3 10272 1764 10272 1764 0 u_ppwm/u_pwm/_017_
rlabel metal2 12384 4284 12384 4284 0 u_ppwm/u_pwm/_018_
rlabel metal2 12864 3654 12864 3654 0 u_ppwm/u_pwm/_019_
rlabel metal2 14400 5712 14400 5712 0 u_ppwm/u_pwm/_020_
rlabel metal2 15072 2268 15072 2268 0 u_ppwm/u_pwm/_021_
rlabel metal2 7200 5544 7200 5544 0 u_ppwm/u_pwm/_022_
rlabel metal2 6240 3276 6240 3276 0 u_ppwm/u_pwm/_023_
rlabel metal2 6768 2856 6768 2856 0 u_ppwm/u_pwm/_024_
rlabel metal3 6096 4368 6096 4368 0 u_ppwm/u_pwm/_025_
rlabel metal2 9312 4116 9312 4116 0 u_ppwm/u_pwm/_026_
rlabel metal2 7872 5208 7872 5208 0 u_ppwm/u_pwm/_027_
rlabel metal2 9408 3150 9408 3150 0 u_ppwm/u_pwm/_028_
rlabel metal3 9504 2436 9504 2436 0 u_ppwm/u_pwm/_029_
rlabel metal3 11952 4284 11952 4284 0 u_ppwm/u_pwm/_030_
rlabel metal2 9936 1932 9936 1932 0 u_ppwm/u_pwm/_031_
rlabel metal2 11904 4242 11904 4242 0 u_ppwm/u_pwm/_032_
rlabel metal2 11328 3318 11328 3318 0 u_ppwm/u_pwm/_033_
rlabel metal2 11712 4452 11712 4452 0 u_ppwm/u_pwm/_034_
rlabel metal2 10560 5922 10560 5922 0 u_ppwm/u_pwm/_035_
rlabel metal3 14160 5628 14160 5628 0 u_ppwm/u_pwm/_036_
rlabel metal2 10848 5670 10848 5670 0 u_ppwm/u_pwm/_037_
rlabel metal2 10512 6972 10512 6972 0 u_ppwm/u_pwm/_038_
rlabel metal3 8640 6636 8640 6636 0 u_ppwm/u_pwm/_039_
rlabel metal2 8640 5628 8640 5628 0 u_ppwm/u_pwm/_040_
rlabel metal3 8640 7392 8640 7392 0 u_ppwm/u_pwm/_041_
rlabel metal2 8304 5880 8304 5880 0 u_ppwm/u_pwm/_042_
rlabel metal2 9696 7266 9696 7266 0 u_ppwm/u_pwm/_043_
rlabel metal2 9120 7056 9120 7056 0 u_ppwm/u_pwm/_044_
rlabel metal2 8928 7434 8928 7434 0 u_ppwm/u_pwm/_045_
rlabel via1 9600 6970 9600 6970 0 u_ppwm/u_pwm/_046_
rlabel metal2 13824 6636 13824 6636 0 u_ppwm/u_pwm/_047_
rlabel metal2 13152 6048 13152 6048 0 u_ppwm/u_pwm/_048_
rlabel metal2 12384 6342 12384 6342 0 u_ppwm/u_pwm/_049_
rlabel metal2 11232 5922 11232 5922 0 u_ppwm/u_pwm/_050_
rlabel metal2 12960 6720 12960 6720 0 u_ppwm/u_pwm/_051_
rlabel metal3 12480 6468 12480 6468 0 u_ppwm/u_pwm/_052_
rlabel metal2 14112 5754 14112 5754 0 u_ppwm/u_pwm/_053_
rlabel metal2 13248 6888 13248 6888 0 u_ppwm/u_pwm/_054_
rlabel metal2 13824 5082 13824 5082 0 u_ppwm/u_pwm/_055_
rlabel metal2 14880 6720 14880 6720 0 u_ppwm/u_pwm/_056_
rlabel metal2 14496 6300 14496 6300 0 u_ppwm/u_pwm/_057_
rlabel metal2 13728 5754 13728 5754 0 u_ppwm/u_pwm/_058_
rlabel metal2 14016 6720 14016 6720 0 u_ppwm/u_pwm/_059_
rlabel metal2 13728 6720 13728 6720 0 u_ppwm/u_pwm/_060_
rlabel metal3 14592 4116 14592 4116 0 u_ppwm/u_pwm/_061_
rlabel metal2 15745 5678 15745 5678 0 u_ppwm/u_pwm/_062_
rlabel metal2 16224 2646 16224 2646 0 u_ppwm/u_pwm/_063_
rlabel metal2 16704 2940 16704 2940 0 u_ppwm/u_pwm/_064_
rlabel metal2 16608 3024 16608 3024 0 u_ppwm/u_pwm/_065_
rlabel metal2 14928 3444 14928 3444 0 u_ppwm/u_pwm/_066_
rlabel metal2 15024 3612 15024 3612 0 u_ppwm/u_pwm/_067_
rlabel metal2 14640 3444 14640 3444 0 u_ppwm/u_pwm/_068_
rlabel metal2 15456 3234 15456 3234 0 u_ppwm/u_pwm/_069_
rlabel metal2 15744 2982 15744 2982 0 u_ppwm/u_pwm/_070_
rlabel metal3 9984 1260 9984 1260 0 u_ppwm/u_pwm/_071_
rlabel metal2 9504 7896 9504 7896 0 u_ppwm/u_pwm/_072_
rlabel metal3 8400 7980 8400 7980 0 u_ppwm/u_pwm/_073_
rlabel metal2 16416 3150 16416 3150 0 u_ppwm/u_pwm/_074_
rlabel metal3 15072 4956 15072 4956 0 u_ppwm/u_pwm/_075_
rlabel metal2 10176 10710 10176 10710 0 u_ppwm/u_pwm/_076_
rlabel metal2 13056 8820 13056 8820 0 u_ppwm/u_pwm/_077_
rlabel metal3 15216 5460 15216 5460 0 u_ppwm/u_pwm/_078_
rlabel via2 15072 6707 15072 6707 0 u_ppwm/u_pwm/_079_
rlabel metal3 8784 9492 8784 9492 0 u_ppwm/u_pwm/_080_
rlabel metal3 9744 7728 9744 7728 0 u_ppwm/u_pwm/_081_
rlabel metal3 10224 9492 10224 9492 0 u_ppwm/u_pwm/_082_
rlabel metal2 9600 12432 9600 12432 0 u_ppwm/u_pwm/_083_
rlabel metal2 5760 5418 5760 5418 0 u_ppwm/u_pwm/_084_
rlabel metal2 11808 5040 11808 5040 0 u_ppwm/u_pwm/_085_
rlabel metal2 11712 5124 11712 5124 0 u_ppwm/u_pwm/_086_
rlabel metal2 12336 7140 12336 7140 0 u_ppwm/u_pwm/_087_
rlabel metal2 11520 10248 11520 10248 0 u_ppwm/u_pwm/_088_
rlabel metal2 11424 10542 11424 10542 0 u_ppwm/u_pwm/_089_
rlabel metal2 14784 9156 14784 9156 0 u_ppwm/u_pwm/_090_
rlabel metal3 9600 9534 9600 9534 0 u_ppwm/u_pwm/_091_
rlabel metal2 14496 8820 14496 8820 0 u_ppwm/u_pwm/_092_
rlabel metal2 15264 7014 15264 7014 0 u_ppwm/u_pwm/_093_
rlabel metal2 12864 9576 12864 9576 0 u_ppwm/u_pwm/_094_
rlabel metal2 11040 10332 11040 10332 0 u_ppwm/u_pwm/_095_
rlabel metal2 16608 6888 16608 6888 0 u_ppwm/u_pwm/_096_
rlabel metal2 16224 4326 16224 4326 0 u_ppwm/u_pwm/_097_
rlabel metal2 6000 6972 6000 6972 0 u_ppwm/u_pwm/_098_
rlabel metal2 5856 8148 5856 8148 0 u_ppwm/u_pwm/_099_
rlabel metal3 4944 7980 4944 7980 0 u_ppwm/u_pwm/_100_
rlabel metal3 6384 5040 6384 5040 0 u_ppwm/u_pwm/_101_
rlabel metal3 8880 11928 8880 11928 0 u_ppwm/u_pwm/cmp_value\[0\]
rlabel metal2 7872 10458 7872 10458 0 u_ppwm/u_pwm/cmp_value\[1\]
rlabel metal2 9659 8064 9659 8064 0 u_ppwm/u_pwm/cmp_value\[2\]
rlabel metal2 9120 9450 9120 9450 0 u_ppwm/u_pwm/cmp_value\[3\]
rlabel metal2 17280 8148 17280 8148 0 u_ppwm/u_pwm/cmp_value\[4\]
rlabel metal3 16320 7140 16320 7140 0 u_ppwm/u_pwm/cmp_value\[5\]
rlabel metal2 13440 8694 13440 8694 0 u_ppwm/u_pwm/cmp_value\[6\]
rlabel metal2 12576 10248 12576 10248 0 u_ppwm/u_pwm/cmp_value\[7\]
rlabel metal2 19392 4578 19392 4578 0 u_ppwm/u_pwm/cmp_value\[8\]
rlabel metal3 18960 2604 18960 2604 0 u_ppwm/u_pwm/cmp_value\[9\]
rlabel metal2 9504 6384 9504 6384 0 u_ppwm/u_pwm/counter\[0\]
rlabel metal2 8448 7014 8448 7014 0 u_ppwm/u_pwm/counter\[1\]
rlabel metal2 9312 6510 9312 6510 0 u_ppwm/u_pwm/counter\[2\]
rlabel metal2 8736 3402 8736 3402 0 u_ppwm/u_pwm/counter\[3\]
rlabel metal2 14496 4998 14496 4998 0 u_ppwm/u_pwm/counter\[4\]
rlabel metal2 14016 5502 14016 5502 0 u_ppwm/u_pwm/counter\[5\]
rlabel metal2 12096 3402 12096 3402 0 u_ppwm/u_pwm/counter\[6\]
rlabel metal2 12096 1848 12096 1848 0 u_ppwm/u_pwm/counter\[7\]
rlabel metal2 14544 4284 14544 4284 0 u_ppwm/u_pwm/counter\[8\]
rlabel metal2 15312 2856 15312 2856 0 u_ppwm/u_pwm/counter\[9\]
rlabel metal3 366 22428 366 22428 0 ui_in[0]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
