module tiny_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire clknet_leaf_0_clk;
 wire \ppwm_i.rst_n ;
 wire \ppwm_i.u_ppwm.data_o ;
 wire \ppwm_i.u_ppwm.global_counter[0] ;
 wire \ppwm_i.u_ppwm.global_counter[10] ;
 wire \ppwm_i.u_ppwm.global_counter[11] ;
 wire \ppwm_i.u_ppwm.global_counter[12] ;
 wire \ppwm_i.u_ppwm.global_counter[13] ;
 wire \ppwm_i.u_ppwm.global_counter[14] ;
 wire \ppwm_i.u_ppwm.global_counter[15] ;
 wire \ppwm_i.u_ppwm.global_counter[16] ;
 wire \ppwm_i.u_ppwm.global_counter[17] ;
 wire \ppwm_i.u_ppwm.global_counter[18] ;
 wire \ppwm_i.u_ppwm.global_counter[19] ;
 wire \ppwm_i.u_ppwm.global_counter[1] ;
 wire \ppwm_i.u_ppwm.global_counter[2] ;
 wire \ppwm_i.u_ppwm.global_counter[3] ;
 wire \ppwm_i.u_ppwm.global_counter[4] ;
 wire \ppwm_i.u_ppwm.global_counter[5] ;
 wire \ppwm_i.u_ppwm.global_counter[6] ;
 wire \ppwm_i.u_ppwm.global_counter[7] ;
 wire \ppwm_i.u_ppwm.global_counter[8] ;
 wire \ppwm_i.u_ppwm.global_counter[9] ;
 wire \ppwm_i.u_ppwm.mem_write_done ;
 wire \ppwm_i.u_ppwm.pc[0] ;
 wire \ppwm_i.u_ppwm.pc[1] ;
 wire \ppwm_i.u_ppwm.pc[2] ;
 wire \ppwm_i.u_ppwm.pc[3] ;
 wire \ppwm_i.u_ppwm.period_start ;
 wire \ppwm_i.u_ppwm.polarity ;
 wire \ppwm_i.u_ppwm.pwm_value[0] ;
 wire \ppwm_i.u_ppwm.pwm_value[1] ;
 wire \ppwm_i.u_ppwm.pwm_value[2] ;
 wire \ppwm_i.u_ppwm.pwm_value[3] ;
 wire \ppwm_i.u_ppwm.pwm_value[4] ;
 wire \ppwm_i.u_ppwm.pwm_value[5] ;
 wire \ppwm_i.u_ppwm.pwm_value[6] ;
 wire \ppwm_i.u_ppwm.pwm_value[7] ;
 wire \ppwm_i.u_ppwm.pwm_value[8] ;
 wire \ppwm_i.u_ppwm.pwm_value[9] ;
 wire \ppwm_i.u_ppwm.u_ex.cmp_flag_q ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[0] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[1] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[2] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[3] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[4] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[5] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[6] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[7] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[8] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[9] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[0] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[1] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[2] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[0] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[1] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[2] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[3] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[4] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[5] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[6] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[0] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[100] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[101] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[102] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[103] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[104] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[105] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[106] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[107] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[108] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[109] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[10] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[110] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[111] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[11] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[12] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[13] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[14] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[15] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[16] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[17] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[18] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[19] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[1] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[20] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[21] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[22] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[23] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[24] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[25] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[26] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[27] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[28] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[29] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[2] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[30] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[31] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[32] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[33] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[34] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[35] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[36] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[37] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[38] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[39] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[3] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[40] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[41] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[42] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[43] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[44] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[45] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[46] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[47] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[48] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[49] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[4] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[50] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[51] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[52] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[53] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[54] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[55] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[56] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[57] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[58] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[59] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[5] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[60] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[61] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[62] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[63] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[64] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[65] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[66] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[67] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[68] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[69] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[6] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[70] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[71] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[72] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[73] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[74] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[75] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[76] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[77] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[78] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[79] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[7] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[80] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[81] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[82] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[83] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[84] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[85] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[86] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[87] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[88] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[89] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[8] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[90] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[91] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[92] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[93] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[94] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[95] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[96] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[97] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[98] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[99] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[9] ;
 wire \ppwm_i.u_ppwm.u_mem.state_q[0] ;
 wire \ppwm_i.u_ppwm.u_mem.state_q[2] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[0] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[1] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[2] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[3] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[4] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[5] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[6] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[7] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[8] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[9] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[0] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[1] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[2] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[3] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[4] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[5] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[6] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[7] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[8] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[9] ;
 wire rst_n_sdr;
 wire \sdr_i.DP_1.matrix[0] ;
 wire \sdr_i.DP_1.matrix[10] ;
 wire \sdr_i.DP_1.matrix[18] ;
 wire \sdr_i.DP_1.matrix[19] ;
 wire \sdr_i.DP_1.matrix[1] ;
 wire \sdr_i.DP_1.matrix[27] ;
 wire \sdr_i.DP_1.matrix[28] ;
 wire \sdr_i.DP_1.matrix[36] ;
 wire \sdr_i.DP_1.matrix[37] ;
 wire \sdr_i.DP_1.matrix[45] ;
 wire \sdr_i.DP_1.matrix[46] ;
 wire \sdr_i.DP_1.matrix[54] ;
 wire \sdr_i.DP_1.matrix[55] ;
 wire \sdr_i.DP_1.matrix[63] ;
 wire \sdr_i.DP_1.matrix[64] ;
 wire \sdr_i.DP_1.matrix[72] ;
 wire \sdr_i.DP_1.matrix[73] ;
 wire \sdr_i.DP_1.matrix[9] ;
 wire \sdr_i.DP_2.matrix[0] ;
 wire \sdr_i.DP_2.matrix[10] ;
 wire \sdr_i.DP_2.matrix[18] ;
 wire \sdr_i.DP_2.matrix[19] ;
 wire \sdr_i.DP_2.matrix[1] ;
 wire \sdr_i.DP_2.matrix[27] ;
 wire \sdr_i.DP_2.matrix[28] ;
 wire \sdr_i.DP_2.matrix[36] ;
 wire \sdr_i.DP_2.matrix[37] ;
 wire \sdr_i.DP_2.matrix[45] ;
 wire \sdr_i.DP_2.matrix[46] ;
 wire \sdr_i.DP_2.matrix[54] ;
 wire \sdr_i.DP_2.matrix[55] ;
 wire \sdr_i.DP_2.matrix[63] ;
 wire \sdr_i.DP_2.matrix[64] ;
 wire \sdr_i.DP_2.matrix[72] ;
 wire \sdr_i.DP_2.matrix[73] ;
 wire \sdr_i.DP_2.matrix[9] ;
 wire \sdr_i.DP_3.matrix[0] ;
 wire \sdr_i.DP_3.matrix[10] ;
 wire \sdr_i.DP_3.matrix[18] ;
 wire \sdr_i.DP_3.matrix[19] ;
 wire \sdr_i.DP_3.matrix[1] ;
 wire \sdr_i.DP_3.matrix[27] ;
 wire \sdr_i.DP_3.matrix[28] ;
 wire \sdr_i.DP_3.matrix[36] ;
 wire \sdr_i.DP_3.matrix[37] ;
 wire \sdr_i.DP_3.matrix[45] ;
 wire \sdr_i.DP_3.matrix[46] ;
 wire \sdr_i.DP_3.matrix[54] ;
 wire \sdr_i.DP_3.matrix[55] ;
 wire \sdr_i.DP_3.matrix[63] ;
 wire \sdr_i.DP_3.matrix[64] ;
 wire \sdr_i.DP_3.matrix[72] ;
 wire \sdr_i.DP_3.matrix[73] ;
 wire \sdr_i.DP_3.matrix[9] ;
 wire \sdr_i.DP_4.matrix[0] ;
 wire \sdr_i.DP_4.matrix[10] ;
 wire \sdr_i.DP_4.matrix[18] ;
 wire \sdr_i.DP_4.matrix[19] ;
 wire \sdr_i.DP_4.matrix[1] ;
 wire \sdr_i.DP_4.matrix[27] ;
 wire \sdr_i.DP_4.matrix[28] ;
 wire \sdr_i.DP_4.matrix[36] ;
 wire \sdr_i.DP_4.matrix[37] ;
 wire \sdr_i.DP_4.matrix[45] ;
 wire \sdr_i.DP_4.matrix[46] ;
 wire \sdr_i.DP_4.matrix[54] ;
 wire \sdr_i.DP_4.matrix[55] ;
 wire \sdr_i.DP_4.matrix[63] ;
 wire \sdr_i.DP_4.matrix[64] ;
 wire \sdr_i.DP_4.matrix[72] ;
 wire \sdr_i.DP_4.matrix[73] ;
 wire \sdr_i.DP_4.matrix[9] ;
 wire \sdr_i.mac1.products_ff[0] ;
 wire \sdr_i.mac1.products_ff[102] ;
 wire \sdr_i.mac1.products_ff[103] ;
 wire \sdr_i.mac1.products_ff[119] ;
 wire \sdr_i.mac1.products_ff[120] ;
 wire \sdr_i.mac1.products_ff[136] ;
 wire \sdr_i.mac1.products_ff[137] ;
 wire \sdr_i.mac1.products_ff[17] ;
 wire \sdr_i.mac1.products_ff[18] ;
 wire \sdr_i.mac1.products_ff[1] ;
 wire \sdr_i.mac1.products_ff[34] ;
 wire \sdr_i.mac1.products_ff[35] ;
 wire \sdr_i.mac1.products_ff[51] ;
 wire \sdr_i.mac1.products_ff[52] ;
 wire \sdr_i.mac1.products_ff[68] ;
 wire \sdr_i.mac1.products_ff[69] ;
 wire \sdr_i.mac1.products_ff[85] ;
 wire \sdr_i.mac1.products_ff[86] ;
 wire \sdr_i.mac1.sum_lvl1_ff[0] ;
 wire \sdr_i.mac1.sum_lvl1_ff[16] ;
 wire \sdr_i.mac1.sum_lvl1_ff[17] ;
 wire \sdr_i.mac1.sum_lvl1_ff[1] ;
 wire \sdr_i.mac1.sum_lvl1_ff[24] ;
 wire \sdr_i.mac1.sum_lvl1_ff[25] ;
 wire \sdr_i.mac1.sum_lvl1_ff[32] ;
 wire \sdr_i.mac1.sum_lvl1_ff[33] ;
 wire \sdr_i.mac1.sum_lvl1_ff[8] ;
 wire \sdr_i.mac1.sum_lvl1_ff[9] ;
 wire \sdr_i.mac1.sum_lvl2_ff[0] ;
 wire \sdr_i.mac1.sum_lvl2_ff[1] ;
 wire \sdr_i.mac1.sum_lvl2_ff[4] ;
 wire \sdr_i.mac1.sum_lvl2_ff[5] ;
 wire \sdr_i.mac1.sum_lvl2_ff[8] ;
 wire \sdr_i.mac1.sum_lvl2_ff[9] ;
 wire \sdr_i.mac1.sum_lvl3_ff[0] ;
 wire \sdr_i.mac1.sum_lvl3_ff[1] ;
 wire \sdr_i.mac1.sum_lvl3_ff[2] ;
 wire \sdr_i.mac1.sum_lvl3_ff[3] ;
 wire \sdr_i.mac1.total_sum[0] ;
 wire \sdr_i.mac1.total_sum[1] ;
 wire \sdr_i.mac2.products_ff[0] ;
 wire \sdr_i.mac2.products_ff[102] ;
 wire \sdr_i.mac2.products_ff[103] ;
 wire \sdr_i.mac2.products_ff[119] ;
 wire \sdr_i.mac2.products_ff[120] ;
 wire \sdr_i.mac2.products_ff[136] ;
 wire \sdr_i.mac2.products_ff[137] ;
 wire \sdr_i.mac2.products_ff[17] ;
 wire \sdr_i.mac2.products_ff[18] ;
 wire \sdr_i.mac2.products_ff[1] ;
 wire \sdr_i.mac2.products_ff[34] ;
 wire \sdr_i.mac2.products_ff[35] ;
 wire \sdr_i.mac2.products_ff[51] ;
 wire \sdr_i.mac2.products_ff[52] ;
 wire \sdr_i.mac2.products_ff[68] ;
 wire \sdr_i.mac2.products_ff[69] ;
 wire \sdr_i.mac2.products_ff[85] ;
 wire \sdr_i.mac2.products_ff[86] ;
 wire \sdr_i.mac2.sum_lvl1_ff[0] ;
 wire \sdr_i.mac2.sum_lvl1_ff[16] ;
 wire \sdr_i.mac2.sum_lvl1_ff[17] ;
 wire \sdr_i.mac2.sum_lvl1_ff[1] ;
 wire \sdr_i.mac2.sum_lvl1_ff[24] ;
 wire \sdr_i.mac2.sum_lvl1_ff[25] ;
 wire \sdr_i.mac2.sum_lvl1_ff[32] ;
 wire \sdr_i.mac2.sum_lvl1_ff[33] ;
 wire \sdr_i.mac2.sum_lvl1_ff[8] ;
 wire \sdr_i.mac2.sum_lvl1_ff[9] ;
 wire \sdr_i.mac2.sum_lvl2_ff[0] ;
 wire \sdr_i.mac2.sum_lvl2_ff[1] ;
 wire \sdr_i.mac2.sum_lvl2_ff[4] ;
 wire \sdr_i.mac2.sum_lvl2_ff[5] ;
 wire \sdr_i.mac2.sum_lvl2_ff[8] ;
 wire \sdr_i.mac2.sum_lvl2_ff[9] ;
 wire \sdr_i.mac2.sum_lvl3_ff[0] ;
 wire \sdr_i.mac2.sum_lvl3_ff[1] ;
 wire \sdr_i.mac2.sum_lvl3_ff[2] ;
 wire \sdr_i.mac2.sum_lvl3_ff[3] ;
 wire \sdr_i.mac2.total_sum[0] ;
 wire \sdr_i.mac2.total_sum[1] ;
 wire \sdr_i.mac2.total_sum[2] ;
 wire \sdr_i.total_sum1[2] ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net1;
 wire net2;
 wire net3;
 wire net16;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;

 sg13g2_inv_1 _1526_ (.Y(_1097_),
    .A(net582));
 sg13g2_inv_1 _1527_ (.Y(_1098_),
    .A(net3));
 sg13g2_inv_1 _1528_ (.Y(_1099_),
    .A(net604));
 sg13g2_inv_1 _1529_ (.Y(_1100_),
    .A(net627));
 sg13g2_inv_1 _1530_ (.Y(_1101_),
    .A(net616));
 sg13g2_inv_1 _1531_ (.Y(_1102_),
    .A(net612));
 sg13g2_inv_1 _1532_ (.Y(_1103_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[106] ));
 sg13g2_inv_1 _1533_ (.Y(_1104_),
    .A(net749));
 sg13g2_inv_1 _1534_ (.Y(_1105_),
    .A(net645));
 sg13g2_inv_1 _1535_ (.Y(_1106_),
    .A(net594));
 sg13g2_inv_1 _1536_ (.Y(_1107_),
    .A(net625));
 sg13g2_inv_1 _1537_ (.Y(_1108_),
    .A(net649));
 sg13g2_inv_1 _1538_ (.Y(_1109_),
    .A(net362));
 sg13g2_inv_1 _1539_ (.Y(_1110_),
    .A(net555));
 sg13g2_inv_1 _1540_ (.Y(_1111_),
    .A(net773));
 sg13g2_inv_1 _1541_ (.Y(_1112_),
    .A(net680));
 sg13g2_inv_1 _1542_ (.Y(_1113_),
    .A(net635));
 sg13g2_inv_1 _1543_ (.Y(_1114_),
    .A(net597));
 sg13g2_inv_1 _1544_ (.Y(_1115_),
    .A(net640));
 sg13g2_inv_1 _1545_ (.Y(_1116_),
    .A(net672));
 sg13g2_inv_1 _1546_ (.Y(_1117_),
    .A(net568));
 sg13g2_inv_1 _1547_ (.Y(_1118_),
    .A(net727));
 sg13g2_inv_1 _1548_ (.Y(_1119_),
    .A(net614));
 sg13g2_inv_1 _1549_ (.Y(_1120_),
    .A(net687));
 sg13g2_inv_1 _1550_ (.Y(_1121_),
    .A(net354));
 sg13g2_inv_1 _1551_ (.Y(_1122_),
    .A(net368));
 sg13g2_inv_1 _1552_ (.Y(_1123_),
    .A(net634));
 sg13g2_inv_1 _1553_ (.Y(_1124_),
    .A(net358));
 sg13g2_inv_1 _1554_ (.Y(_1125_),
    .A(net681));
 sg13g2_inv_1 _1555_ (.Y(_1126_),
    .A(net678));
 sg13g2_inv_1 _1556_ (.Y(_1127_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[82] ));
 sg13g2_inv_1 _1557_ (.Y(_1128_),
    .A(net700));
 sg13g2_inv_1 _1558_ (.Y(_1129_),
    .A(net706));
 sg13g2_inv_1 _1559_ (.Y(_1130_),
    .A(net364));
 sg13g2_inv_1 _1560_ (.Y(_1131_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[78] ));
 sg13g2_inv_1 _1561_ (.Y(_1132_),
    .A(net652));
 sg13g2_inv_1 _1562_ (.Y(_1133_),
    .A(net677));
 sg13g2_inv_1 _1563_ (.Y(_1134_),
    .A(net607));
 sg13g2_inv_1 _1564_ (.Y(_1135_),
    .A(net630));
 sg13g2_inv_1 _1565_ (.Y(_1136_),
    .A(net704));
 sg13g2_inv_1 _1566_ (.Y(_1137_),
    .A(net559));
 sg13g2_inv_1 _1567_ (.Y(_1138_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[71] ));
 sg13g2_inv_1 _1568_ (.Y(_1139_),
    .A(net667));
 sg13g2_inv_1 _1569_ (.Y(_1140_),
    .A(net637));
 sg13g2_inv_1 _1570_ (.Y(_1141_),
    .A(net574));
 sg13g2_inv_1 _1571_ (.Y(_1142_),
    .A(net671));
 sg13g2_inv_1 _1572_ (.Y(_1143_),
    .A(net659));
 sg13g2_inv_1 _1573_ (.Y(_1144_),
    .A(net347));
 sg13g2_inv_1 _1574_ (.Y(_1145_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[64] ));
 sg13g2_inv_1 _1575_ (.Y(_1146_),
    .A(net650));
 sg13g2_inv_1 _1576_ (.Y(_1147_),
    .A(net660));
 sg13g2_inv_1 _1577_ (.Y(_1148_),
    .A(net590));
 sg13g2_inv_1 _1578_ (.Y(_1149_),
    .A(net619));
 sg13g2_inv_1 _1579_ (.Y(_1150_),
    .A(net728));
 sg13g2_inv_1 _1580_ (.Y(_1151_),
    .A(net563));
 sg13g2_inv_1 _1581_ (.Y(_1152_),
    .A(net632));
 sg13g2_inv_2 _1582_ (.Y(_1153_),
    .A(net673));
 sg13g2_inv_1 _1583_ (.Y(_1154_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[55] ));
 sg13g2_inv_1 _1584_ (.Y(_1155_),
    .A(net669));
 sg13g2_inv_1 _1585_ (.Y(_1156_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[53] ));
 sg13g2_inv_1 _1586_ (.Y(_1157_),
    .A(net657));
 sg13g2_inv_1 _1587_ (.Y(_1158_),
    .A(net366));
 sg13g2_inv_1 _1588_ (.Y(_1159_),
    .A(net639));
 sg13g2_inv_1 _1589_ (.Y(_1160_),
    .A(net638));
 sg13g2_inv_1 _1590_ (.Y(_1161_),
    .A(net570));
 sg13g2_inv_2 _1591_ (.Y(_1162_),
    .A(net703));
 sg13g2_inv_1 _1592_ (.Y(_1163_),
    .A(net592));
 sg13g2_inv_1 _1593_ (.Y(_1164_),
    .A(net611));
 sg13g2_inv_1 _1594_ (.Y(_1165_),
    .A(net356));
 sg13g2_inv_1 _1595_ (.Y(_1166_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[43] ));
 sg13g2_inv_1 _1596_ (.Y(_1167_),
    .A(net682));
 sg13g2_inv_1 _1597_ (.Y(_1168_),
    .A(net702));
 sg13g2_inv_1 _1598_ (.Y(_1169_),
    .A(net699));
 sg13g2_inv_1 _1599_ (.Y(_1170_),
    .A(net698));
 sg13g2_inv_1 _1600_ (.Y(_1171_),
    .A(net643));
 sg13g2_inv_1 _1601_ (.Y(_1172_),
    .A(net606));
 sg13g2_inv_1 _1602_ (.Y(_1173_),
    .A(net584));
 sg13g2_inv_1 _1603_ (.Y(_1174_),
    .A(net714));
 sg13g2_inv_1 _1604_ (.Y(_1175_),
    .A(net675));
 sg13g2_inv_1 _1605_ (.Y(_1176_),
    .A(net688));
 sg13g2_inv_1 _1606_ (.Y(_1177_),
    .A(net345));
 sg13g2_inv_1 _1607_ (.Y(_1178_),
    .A(net360));
 sg13g2_inv_1 _1608_ (.Y(_1179_),
    .A(net576));
 sg13g2_inv_1 _1609_ (.Y(_1180_),
    .A(net636));
 sg13g2_inv_1 _1610_ (.Y(_1181_),
    .A(net596));
 sg13g2_inv_1 _1611_ (.Y(_1182_),
    .A(net550));
 sg13g2_inv_2 _1612_ (.Y(_1183_),
    .A(net691));
 sg13g2_inv_1 _1613_ (.Y(_1184_),
    .A(net586));
 sg13g2_inv_1 _1614_ (.Y(_1185_),
    .A(net599));
 sg13g2_inv_1 _1615_ (.Y(_1186_),
    .A(net617));
 sg13g2_inv_1 _1616_ (.Y(_1187_),
    .A(net621));
 sg13g2_inv_1 _1617_ (.Y(_1188_),
    .A(net733));
 sg13g2_inv_1 _1618_ (.Y(_1189_),
    .A(net623));
 sg13g2_inv_1 _1619_ (.Y(_1190_),
    .A(net705));
 sg13g2_inv_1 _1620_ (.Y(_1191_),
    .A(net697));
 sg13g2_inv_1 _1621_ (.Y(_1192_),
    .A(net352));
 sg13g2_inv_1 _1622_ (.Y(_1193_),
    .A(net646));
 sg13g2_inv_1 _1623_ (.Y(_1194_),
    .A(net588));
 sg13g2_inv_1 _1624_ (.Y(_1195_),
    .A(net666));
 sg13g2_inv_1 _1625_ (.Y(_1196_),
    .A(net609));
 sg13g2_inv_1 _1626_ (.Y(_1197_),
    .A(net686));
 sg13g2_inv_1 _1627_ (.Y(_1198_),
    .A(net647));
 sg13g2_inv_1 _1628_ (.Y(_1199_),
    .A(net642));
 sg13g2_inv_1 _1629_ (.Y(_1200_),
    .A(net561));
 sg13g2_inv_1 _1630_ (.Y(_1201_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[8] ));
 sg13g2_inv_1 _1631_ (.Y(_1202_),
    .A(net692));
 sg13g2_inv_1 _1632_ (.Y(_1203_),
    .A(net628));
 sg13g2_inv_1 _1633_ (.Y(_1204_),
    .A(net684));
 sg13g2_inv_1 _1634_ (.Y(_1205_),
    .A(net656));
 sg13g2_inv_1 _1635_ (.Y(_1206_),
    .A(net342));
 sg13g2_inv_1 _1636_ (.Y(_1207_),
    .A(net337));
 sg13g2_inv_1 _1637_ (.Y(_1208_),
    .A(net343));
 sg13g2_inv_1 _1638_ (.Y(_1209_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[0] ));
 sg13g2_inv_2 _1639_ (.Y(_1210_),
    .A(net805));
 sg13g2_inv_2 _1640_ (.Y(_1211_),
    .A(net809));
 sg13g2_inv_2 _1641_ (.Y(_1212_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ));
 sg13g2_inv_1 _1642_ (.Y(_1213_),
    .A(net502));
 sg13g2_inv_2 _1643_ (.Y(_1214_),
    .A(net821));
 sg13g2_inv_4 _1644_ (.A(net818),
    .Y(_1215_));
 sg13g2_inv_2 _1645_ (.Y(_1216_),
    .A(net816));
 sg13g2_inv_2 _1646_ (.Y(_1217_),
    .A(net811));
 sg13g2_inv_2 _1647_ (.Y(_1218_),
    .A(net826));
 sg13g2_inv_2 _1648_ (.Y(_1219_),
    .A(net812));
 sg13g2_inv_4 _1649_ (.A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .Y(_1220_));
 sg13g2_inv_2 _1650_ (.Y(_1221_),
    .A(\ppwm_i.u_ppwm.pwm_value[8] ));
 sg13g2_inv_2 _1651_ (.Y(_1222_),
    .A(net503));
 sg13g2_inv_2 _1652_ (.Y(_1223_),
    .A(net504));
 sg13g2_inv_4 _1653_ (.A(\ppwm_i.u_ppwm.pwm_value[5] ),
    .Y(_1224_));
 sg13g2_inv_4 _1654_ (.A(net505),
    .Y(_1225_));
 sg13g2_inv_2 _1655_ (.Y(_1226_),
    .A(net506));
 sg13g2_inv_2 _1656_ (.Y(_1227_),
    .A(\ppwm_i.u_ppwm.pwm_value[2] ));
 sg13g2_inv_2 _1657_ (.Y(_1228_),
    .A(net507));
 sg13g2_inv_4 _1658_ (.A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .Y(_1229_));
 sg13g2_inv_1 _1659_ (.Y(_1230_),
    .A(net712));
 sg13g2_inv_4 _1660_ (.A(net508),
    .Y(_1231_));
 sg13g2_inv_2 _1661_ (.Y(_1232_),
    .A(net768));
 sg13g2_inv_1 _1662_ (.Y(_1233_),
    .A(net512));
 sg13g2_inv_1 _1663_ (.Y(_1234_),
    .A(net752));
 sg13g2_inv_1 _1664_ (.Y(_1235_),
    .A(net715));
 sg13g2_inv_1 _1665_ (.Y(_1236_),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[8] ));
 sg13g2_inv_1 _1666_ (.Y(_1237_),
    .A(net819));
 sg13g2_inv_1 _1667_ (.Y(_1238_),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[6] ));
 sg13g2_inv_1 _1668_ (.Y(_1239_),
    .A(net520));
 sg13g2_inv_1 _1669_ (.Y(_1240_),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[1] ));
 sg13g2_inv_1 _1670_ (.Y(_1241_),
    .A(net725));
 sg13g2_inv_1 _1671_ (.Y(_1242_),
    .A(net802));
 sg13g2_inv_1 _1672_ (.Y(_1243_),
    .A(net791));
 sg13g2_inv_1 _1673_ (.Y(_1244_),
    .A(net796));
 sg13g2_inv_1 _1674_ (.Y(_1245_),
    .A(\ppwm_i.u_ppwm.u_pwm.cmp_value[3] ));
 sg13g2_inv_1 _1675_ (.Y(_1246_),
    .A(\ppwm_i.u_ppwm.u_pwm.cmp_value[2] ));
 sg13g2_inv_1 _1676_ (.Y(_1247_),
    .A(net322));
 sg13g2_inv_1 _1677_ (.Y(_1248_),
    .A(net548));
 sg13g2_inv_1 _1678_ (.Y(_1249_),
    .A(net326));
 sg13g2_inv_1 _1679_ (.Y(_1250_),
    .A(\ppwm_i.u_ppwm.data_o ));
 sg13g2_inv_1 _1680_ (.Y(_1251_),
    .A(\ppwm_i.u_ppwm.global_counter[19] ));
 sg13g2_inv_1 _1681_ (.Y(_1252_),
    .A(\ppwm_i.u_ppwm.global_counter[18] ));
 sg13g2_inv_1 _1682_ (.Y(_1253_),
    .A(net798));
 sg13g2_inv_2 _1683_ (.Y(_1254_),
    .A(net780));
 sg13g2_inv_1 _1684_ (.Y(_1255_),
    .A(net572));
 sg13g2_inv_2 _1685_ (.Y(_1256_),
    .A(net776));
 sg13g2_inv_1 _1686_ (.Y(_1257_),
    .A(\ppwm_i.u_ppwm.global_counter[12] ));
 sg13g2_inv_2 _1687_ (.Y(_1258_),
    .A(net787));
 sg13g2_inv_2 _1688_ (.Y(_1259_),
    .A(net335));
 sg13g2_inv_1 _1689_ (.Y(_1260_),
    .A(\ppwm_i.u_ppwm.global_counter[8] ));
 sg13g2_inv_2 _1690_ (.Y(_1261_),
    .A(net320));
 sg13g2_inv_1 _1691_ (.Y(_1262_),
    .A(\ppwm_i.u_ppwm.global_counter[5] ));
 sg13g2_inv_1 _1692_ (.Y(_1263_),
    .A(\ppwm_i.u_ppwm.global_counter[4] ));
 sg13g2_inv_2 _1693_ (.Y(_1264_),
    .A(net789));
 sg13g2_inv_1 _1694_ (.Y(_1265_),
    .A(\ppwm_i.u_ppwm.global_counter[2] ));
 sg13g2_nand2_1 _1695_ (.Y(_1266_),
    .A(net2),
    .B(_1248_));
 sg13g2_inv_4 _1696_ (.A(net457),
    .Y(\ppwm_i.rst_n ));
 sg13g2_nor2_1 _1697_ (.A(_1098_),
    .B(net457),
    .Y(_1267_));
 sg13g2_nor3_1 _1698_ (.A(net3),
    .B(net324),
    .C(net457),
    .Y(_1268_));
 sg13g2_a21oi_1 _1699_ (.A1(_1235_),
    .A2(_1267_),
    .Y(_0003_),
    .B1(_1268_));
 sg13g2_nand2_1 _1700_ (.Y(_1269_),
    .A(net694),
    .B(net330));
 sg13g2_nand4_1 _1701_ (.B(net716),
    .C(net339),
    .A(net661),
    .Y(_1270_),
    .D(net751));
 sg13g2_nor3_1 _1702_ (.A(net748),
    .B(_1269_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_nand2_1 _1703_ (.Y(_1272_),
    .A(net471),
    .B(net421));
 sg13g2_nand3_1 _1704_ (.B(net421),
    .C(_1271_),
    .A(net471),
    .Y(_1273_));
 sg13g2_nand3_1 _1705_ (.B(net715),
    .C(net421),
    .A(_1098_),
    .Y(_1274_));
 sg13g2_nand2_1 _1706_ (.Y(_0004_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_nand2_1 _1707_ (.Y(_1275_),
    .A(net324),
    .B(_1267_));
 sg13g2_o21ai_1 _1708_ (.B1(_1275_),
    .Y(_0005_),
    .A1(_1271_),
    .A2(_1272_));
 sg13g2_and2_1 _1709_ (.A(net514),
    .B(net517),
    .X(_1276_));
 sg13g2_and3_1 _1710_ (.X(_1277_),
    .A(net508),
    .B(net510),
    .C(net450));
 sg13g2_nand3_1 _1711_ (.B(net510),
    .C(net450),
    .A(net508),
    .Y(_1278_));
 sg13g2_nand2_1 _1712_ (.Y(_1279_),
    .A(net768),
    .B(net419));
 sg13g2_nor2_1 _1713_ (.A(net514),
    .B(net517),
    .Y(_1280_));
 sg13g2_nor3_1 _1714_ (.A(\ppwm_i.u_ppwm.u_mem.memory[87] ),
    .B(net515),
    .C(net518),
    .Y(_1281_));
 sg13g2_nor2b_2 _1715_ (.A(net514),
    .B_N(net517),
    .Y(_1282_));
 sg13g2_nor2b_2 _1716_ (.A(net517),
    .B_N(net514),
    .Y(_1283_));
 sg13g2_a21oi_1 _1717_ (.A1(_1115_),
    .A2(net443),
    .Y(_1284_),
    .B1(net460));
 sg13g2_a221oi_1 _1718_ (.B2(_1108_),
    .C1(_1281_),
    .B1(net439),
    .A1(_1101_),
    .Y(_1285_),
    .A2(net451));
 sg13g2_a22oi_1 _1719_ (.Y(_1286_),
    .B1(net439),
    .B2(_1136_),
    .A2(net443),
    .A1(_1143_));
 sg13g2_a221oi_1 _1720_ (.B2(_1150_),
    .C1(net510),
    .B1(net447),
    .A1(_1129_),
    .Y(_1287_),
    .A2(net451));
 sg13g2_a221oi_1 _1721_ (.B2(_1287_),
    .C1(_1231_),
    .B1(_1286_),
    .A1(_1284_),
    .Y(_1288_),
    .A2(_1285_));
 sg13g2_nor3_1 _1722_ (.A(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .B(net516),
    .C(net519),
    .Y(_1289_));
 sg13g2_a21oi_1 _1723_ (.A1(_1192_),
    .A2(net441),
    .Y(_1290_),
    .B1(net512));
 sg13g2_a221oi_1 _1724_ (.B2(_1199_),
    .C1(_1289_),
    .B1(net444),
    .A1(_1185_),
    .Y(_1291_),
    .A2(net453));
 sg13g2_a22oi_1 _1725_ (.Y(_1292_),
    .B1(net441),
    .B2(_1164_),
    .A2(net448),
    .A1(_1178_));
 sg13g2_a221oi_1 _1726_ (.B2(_1171_),
    .C1(net460),
    .B1(net446),
    .A1(_1157_),
    .Y(_1293_),
    .A2(net454));
 sg13g2_a221oi_1 _1727_ (.B2(_1293_),
    .C1(net509),
    .B1(_1292_),
    .A1(_1290_),
    .Y(_1294_),
    .A2(_1291_));
 sg13g2_nor2_2 _1728_ (.A(_1288_),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_or2_1 _1729_ (.X(_1296_),
    .B(_1294_),
    .A(_1288_));
 sg13g2_a21oi_1 _1730_ (.A1(_1114_),
    .A2(net442),
    .Y(_1297_),
    .B1(net460));
 sg13g2_nor3_1 _1731_ (.A(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .B(net515),
    .C(net518),
    .Y(_1298_));
 sg13g2_a221oi_1 _1732_ (.B2(_1107_),
    .C1(_1298_),
    .B1(net438),
    .A1(_1100_),
    .Y(_1299_),
    .A2(net450));
 sg13g2_a22oi_1 _1733_ (.Y(_1300_),
    .B1(net442),
    .B2(_1142_),
    .A2(net450),
    .A1(_1128_));
 sg13g2_a221oi_1 _1734_ (.B2(_1135_),
    .C1(net510),
    .B1(net438),
    .A1(_1149_),
    .Y(_1301_),
    .A2(net447));
 sg13g2_a22oi_1 _1735_ (.Y(_1302_),
    .B1(_1300_),
    .B2(_1301_),
    .A2(_1299_),
    .A1(_1297_));
 sg13g2_nand2_1 _1736_ (.Y(_1303_),
    .A(_1177_),
    .B(net448));
 sg13g2_nand2_1 _1737_ (.Y(_1304_),
    .A(_1163_),
    .B(net441));
 sg13g2_a22oi_1 _1738_ (.Y(_1305_),
    .B1(net446),
    .B2(_1170_),
    .A2(net454),
    .A1(_1156_));
 sg13g2_nand4_1 _1739_ (.B(_1303_),
    .C(_1304_),
    .A(net512),
    .Y(_1306_),
    .D(_1305_));
 sg13g2_a22oi_1 _1740_ (.Y(_1307_),
    .B1(net440),
    .B2(_1191_),
    .A2(net453),
    .A1(_1184_));
 sg13g2_a221oi_1 _1741_ (.B2(_1198_),
    .C1(net512),
    .B1(net444),
    .A1(_1205_),
    .Y(_1308_),
    .A2(net448));
 sg13g2_a21oi_2 _1742_ (.B1(net509),
    .Y(_1309_),
    .A2(_1308_),
    .A1(_1307_));
 sg13g2_a22oi_1 _1743_ (.Y(_1310_),
    .B1(_1306_),
    .B2(_1309_),
    .A2(_1302_),
    .A1(net508));
 sg13g2_inv_4 _1744_ (.A(net397),
    .Y(_1311_));
 sg13g2_nand2_2 _1745_ (.Y(_1312_),
    .A(net404),
    .B(_1311_));
 sg13g2_nor3_1 _1746_ (.A(\ppwm_i.u_ppwm.u_mem.memory[84] ),
    .B(net515),
    .C(net518),
    .Y(_1313_));
 sg13g2_a21oi_1 _1747_ (.A1(_1111_),
    .A2(net438),
    .Y(_1314_),
    .B1(net460));
 sg13g2_a221oi_1 _1748_ (.B2(_1118_),
    .C1(_1313_),
    .B1(net442),
    .A1(_1104_),
    .Y(_1315_),
    .A2(net450));
 sg13g2_a22oi_1 _1749_ (.Y(_1316_),
    .B1(net438),
    .B2(_1139_),
    .A2(net442),
    .A1(_1146_));
 sg13g2_a221oi_1 _1750_ (.B2(_1153_),
    .C1(net510),
    .B1(net447),
    .A1(_1132_),
    .Y(_1317_),
    .A2(net450));
 sg13g2_a221oi_1 _1751_ (.B2(_1317_),
    .C1(_1231_),
    .B1(_1316_),
    .A1(_1314_),
    .Y(_1318_),
    .A2(_1315_));
 sg13g2_a21oi_1 _1752_ (.A1(_1167_),
    .A2(net440),
    .Y(_1319_),
    .B1(net461));
 sg13g2_nor3_1 _1753_ (.A(\ppwm_i.u_ppwm.u_mem.memory[28] ),
    .B(net514),
    .C(net517),
    .Y(_1320_));
 sg13g2_a221oi_1 _1754_ (.B2(_1174_),
    .C1(_1320_),
    .B1(net444),
    .A1(_1160_),
    .Y(_1321_),
    .A2(net453));
 sg13g2_a22oi_1 _1755_ (.Y(_1322_),
    .B1(net448),
    .B2(_1209_),
    .A2(net453),
    .A1(_1188_));
 sg13g2_a221oi_1 _1756_ (.B2(_1195_),
    .C1(net512),
    .B1(net440),
    .A1(_1202_),
    .Y(_1323_),
    .A2(net445));
 sg13g2_a22oi_1 _1757_ (.Y(_1324_),
    .B1(_1322_),
    .B2(_1323_),
    .A2(_1321_),
    .A1(_1319_));
 sg13g2_a21o_2 _1758_ (.A2(_1324_),
    .A1(_1231_),
    .B1(_1318_),
    .X(_1325_));
 sg13g2_a21oi_1 _1759_ (.A1(_1103_),
    .A2(net451),
    .Y(_1326_),
    .B1(net460));
 sg13g2_nor3_1 _1760_ (.A(\ppwm_i.u_ppwm.u_mem.memory[85] ),
    .B(net515),
    .C(net518),
    .Y(_1327_));
 sg13g2_a221oi_1 _1761_ (.B2(_1110_),
    .C1(_1327_),
    .B1(net439),
    .A1(_1117_),
    .Y(_1328_),
    .A2(net443));
 sg13g2_a22oi_1 _1762_ (.Y(_1329_),
    .B1(net439),
    .B2(_1138_),
    .A2(net447),
    .A1(_1152_));
 sg13g2_a221oi_1 _1763_ (.B2(_1145_),
    .C1(net510),
    .B1(net443),
    .A1(_1131_),
    .Y(_1330_),
    .A2(net451));
 sg13g2_a22oi_1 _1764_ (.Y(_1331_),
    .B1(_1329_),
    .B2(_1330_),
    .A2(_1328_),
    .A1(_1326_));
 sg13g2_nor3_1 _1765_ (.A(\ppwm_i.u_ppwm.u_mem.memory[1] ),
    .B(net514),
    .C(net517),
    .Y(_1332_));
 sg13g2_a21oi_1 _1766_ (.A1(_1187_),
    .A2(net453),
    .Y(_1333_),
    .B1(net512));
 sg13g2_a221oi_1 _1767_ (.B2(_1194_),
    .C1(_1332_),
    .B1(net440),
    .A1(_1201_),
    .Y(_1334_),
    .A2(net444));
 sg13g2_a22oi_1 _1768_ (.Y(_1335_),
    .B1(net448),
    .B2(_1180_),
    .A2(net453),
    .A1(_1159_));
 sg13g2_a221oi_1 _1769_ (.B2(_1166_),
    .C1(net461),
    .B1(net440),
    .A1(_1173_),
    .Y(_1336_),
    .A2(net444));
 sg13g2_a221oi_1 _1770_ (.B2(_1336_),
    .C1(net509),
    .B1(_1335_),
    .A1(_1333_),
    .Y(_1337_),
    .A2(_1334_));
 sg13g2_a21o_2 _1771_ (.A2(_1331_),
    .A1(net509),
    .B1(_1337_),
    .X(_1338_));
 sg13g2_nand2_1 _1772_ (.Y(_1339_),
    .A(_1325_),
    .B(net394));
 sg13g2_a21oi_1 _1773_ (.A1(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .A2(net445),
    .Y(_1340_),
    .B1(net513));
 sg13g2_and3_1 _1774_ (.X(_1341_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .B(net514),
    .C(net517));
 sg13g2_a221oi_1 _1775_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .C1(_1341_),
    .B1(net440),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .Y(_1342_),
    .A2(net449));
 sg13g2_a21oi_1 _1776_ (.A1(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .A2(net448),
    .Y(_1343_),
    .B1(net461));
 sg13g2_and3_1 _1777_ (.X(_1344_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[55] ),
    .B(net514),
    .C(net517));
 sg13g2_a221oi_1 _1778_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .C1(_1344_),
    .B1(net440),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .Y(_1345_),
    .A2(net444));
 sg13g2_a221oi_1 _1779_ (.B2(_1345_),
    .C1(net509),
    .B1(_1343_),
    .A1(_1340_),
    .Y(_1346_),
    .A2(_1342_));
 sg13g2_a22oi_1 _1780_ (.Y(_1347_),
    .B1(net442),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .A2(net450),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[83] ));
 sg13g2_a221oi_1 _1781_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .C1(net510),
    .B1(net438),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .Y(_1348_),
    .A2(net447));
 sg13g2_a21oi_1 _1782_ (.A1(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .A2(net447),
    .Y(_1349_),
    .B1(net460));
 sg13g2_and3_1 _1783_ (.X(_1350_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .B(net515),
    .C(net518));
 sg13g2_a221oi_1 _1784_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .C1(_1350_),
    .B1(net438),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .Y(_1351_),
    .A2(net442));
 sg13g2_a221oi_1 _1785_ (.B2(_1351_),
    .C1(_1231_),
    .B1(_1349_),
    .A1(_1347_),
    .Y(_1352_),
    .A2(_1348_));
 sg13g2_nor2_2 _1786_ (.A(net407),
    .B(net406),
    .Y(_0335_));
 sg13g2_or2_1 _1787_ (.X(_0336_),
    .B(net406),
    .A(net407));
 sg13g2_a22oi_1 _1788_ (.Y(_0337_),
    .B1(net438),
    .B2(_1106_),
    .A2(net452),
    .A1(_1099_));
 sg13g2_a221oi_1 _1789_ (.B2(_1113_),
    .C1(net460),
    .B1(net442),
    .A1(_1120_),
    .Y(_0338_),
    .A2(net447));
 sg13g2_a22oi_1 _1790_ (.Y(_0339_),
    .B1(net438),
    .B2(_1134_),
    .A2(net447),
    .A1(_1148_));
 sg13g2_a221oi_1 _1791_ (.B2(_1141_),
    .C1(net510),
    .B1(net442),
    .A1(_1127_),
    .Y(_0340_),
    .A2(net450));
 sg13g2_a221oi_1 _1792_ (.B2(_0340_),
    .C1(_1231_),
    .B1(_0339_),
    .A1(_0337_),
    .Y(_0341_),
    .A2(_0338_));
 sg13g2_a22oi_1 _1793_ (.Y(_0342_),
    .B1(net441),
    .B2(_1162_),
    .A2(net448),
    .A1(_1176_));
 sg13g2_a221oi_1 _1794_ (.B2(_1169_),
    .C1(net461),
    .B1(net444),
    .A1(_1155_),
    .Y(_0343_),
    .A2(net453));
 sg13g2_nor3_1 _1795_ (.A(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .B(net516),
    .C(net519),
    .Y(_0344_));
 sg13g2_a221oi_1 _1796_ (.B2(_1190_),
    .C1(_0344_),
    .B1(net441),
    .A1(_1197_),
    .Y(_0345_),
    .A2(net445));
 sg13g2_a21oi_1 _1797_ (.A1(_1183_),
    .A2(net453),
    .Y(_0346_),
    .B1(net512));
 sg13g2_a221oi_1 _1798_ (.B2(_0346_),
    .C1(net509),
    .B1(_0345_),
    .A1(_0342_),
    .Y(_0347_),
    .A2(_0343_));
 sg13g2_nor2_1 _1799_ (.A(_0341_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_or2_1 _1800_ (.X(_0349_),
    .B(_0347_),
    .A(_0341_));
 sg13g2_nor2_2 _1801_ (.A(net390),
    .B(net387),
    .Y(_0350_));
 sg13g2_nand2_2 _1802_ (.Y(_0351_),
    .A(net392),
    .B(net385));
 sg13g2_a22oi_1 _1803_ (.Y(_0352_),
    .B1(net439),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .A2(net443),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[93] ));
 sg13g2_a221oi_1 _1804_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .C1(net460),
    .B1(net449),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .Y(_0353_),
    .A2(net452));
 sg13g2_nand2_1 _1805_ (.Y(_0354_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .B(net439));
 sg13g2_a21oi_1 _1806_ (.A1(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .A2(net443),
    .Y(_0355_),
    .B1(net511));
 sg13g2_a22oi_1 _1807_ (.Y(_0356_),
    .B1(net449),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .A2(net451),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[79] ));
 sg13g2_nand3_1 _1808_ (.B(_0355_),
    .C(_0356_),
    .A(_0354_),
    .Y(_0357_));
 sg13g2_a21oi_1 _1809_ (.A1(_0352_),
    .A2(_0353_),
    .Y(_0358_),
    .B1(_1231_));
 sg13g2_a22oi_1 _1810_ (.Y(_0359_),
    .B1(net441),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .A2(net448),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[2] ));
 sg13g2_a221oi_1 _1811_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .C1(net513),
    .B1(net445),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .Y(_0360_),
    .A2(net454));
 sg13g2_a21oi_1 _1812_ (.A1(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .A2(net449),
    .Y(_0361_),
    .B1(net461));
 sg13g2_and3_1 _1813_ (.X(_0362_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .B(net516),
    .C(net519));
 sg13g2_a221oi_1 _1814_ (.B2(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .C1(_0362_),
    .B1(net440),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .Y(_0363_),
    .A2(net444));
 sg13g2_a221oi_1 _1815_ (.B2(_0363_),
    .C1(net509),
    .B1(_0361_),
    .A1(_0359_),
    .Y(_0364_),
    .A2(_0360_));
 sg13g2_a21o_2 _1816_ (.A2(_0358_),
    .A1(_0357_),
    .B1(_0364_),
    .X(_0365_));
 sg13g2_nor3_1 _1817_ (.A(_1339_),
    .B(_0351_),
    .C(_0365_),
    .Y(_0366_));
 sg13g2_nand2b_1 _1818_ (.Y(_0367_),
    .B(_0366_),
    .A_N(_1312_));
 sg13g2_nand2b_1 _1819_ (.Y(_0368_),
    .B(_0367_),
    .A_N(_1279_));
 sg13g2_nor2_1 _1820_ (.A(_1249_),
    .B(net457),
    .Y(_0369_));
 sg13g2_a21oi_1 _1821_ (.A1(_1249_),
    .A2(net759),
    .Y(_0370_),
    .B1(net457));
 sg13g2_o21ai_1 _1822_ (.B1(_0370_),
    .Y(_0000_),
    .A1(_1278_),
    .A2(_0368_));
 sg13g2_o21ai_1 _1823_ (.B1(_0369_),
    .Y(_0371_),
    .A1(net759),
    .A2(net317));
 sg13g2_o21ai_1 _1824_ (.B1(_0371_),
    .Y(_0002_),
    .A1(_1277_),
    .A2(_0368_));
 sg13g2_nand3_1 _1825_ (.B(net317),
    .C(net414),
    .A(_1249_),
    .Y(_0372_));
 sg13g2_o21ai_1 _1826_ (.B1(net318),
    .Y(_0001_),
    .A1(_1279_),
    .A2(_0367_));
 sg13g2_or2_1 _1827_ (.X(_0373_),
    .B(\sdr_i.mac2.total_sum[0] ),
    .A(\sdr_i.mac1.total_sum[0] ));
 sg13g2_nand2_1 _1828_ (.Y(_0374_),
    .A(\sdr_i.mac1.total_sum[0] ),
    .B(\sdr_i.mac2.total_sum[0] ));
 sg13g2_nand3_1 _1829_ (.B(_0373_),
    .C(_0374_),
    .A(net548),
    .Y(_0375_));
 sg13g2_o21ai_1 _1830_ (.B1(_0375_),
    .Y(net12),
    .A1(net548),
    .A2(_1250_));
 sg13g2_nand2_1 _1831_ (.Y(_0376_),
    .A(\sdr_i.mac1.total_sum[1] ),
    .B(\sdr_i.mac2.total_sum[1] ));
 sg13g2_xnor2_1 _1832_ (.Y(_0377_),
    .A(\sdr_i.mac1.total_sum[1] ),
    .B(\sdr_i.mac2.total_sum[1] ));
 sg13g2_or2_1 _1833_ (.X(_0378_),
    .B(_0377_),
    .A(_0374_));
 sg13g2_nand2_1 _1834_ (.Y(_0379_),
    .A(net548),
    .B(_0378_));
 sg13g2_a21oi_2 _1835_ (.B1(_0379_),
    .Y(net13),
    .A2(_0377_),
    .A1(_0374_));
 sg13g2_nand2_1 _1836_ (.Y(_0380_),
    .A(\sdr_i.total_sum1[2] ),
    .B(\sdr_i.mac2.total_sum[2] ));
 sg13g2_xnor2_1 _1837_ (.Y(_0381_),
    .A(\sdr_i.total_sum1[2] ),
    .B(\sdr_i.mac2.total_sum[2] ));
 sg13g2_nand3_1 _1838_ (.B(_0378_),
    .C(_0381_),
    .A(_0376_),
    .Y(_0382_));
 sg13g2_a21o_1 _1839_ (.A2(_0378_),
    .A1(_0376_),
    .B1(_0381_),
    .X(_0383_));
 sg13g2_and3_2 _1840_ (.X(net14),
    .A(net548),
    .B(_0382_),
    .C(_0383_));
 sg13g2_a21oi_2 _1841_ (.B1(_1248_),
    .Y(net15),
    .A2(_0383_),
    .A1(_0380_));
 sg13g2_nand2_1 _1842_ (.Y(_0384_),
    .A(net286),
    .B(net221));
 sg13g2_nand2_1 _1843_ (.Y(_0385_),
    .A(net289),
    .B(net233));
 sg13g2_xor2_1 _1844_ (.B(_0385_),
    .A(_0384_),
    .X(_0053_));
 sg13g2_nand2_1 _1845_ (.Y(_0386_),
    .A(net274),
    .B(net220));
 sg13g2_nand2_1 _1846_ (.Y(_0387_),
    .A(net285),
    .B(net237));
 sg13g2_xor2_1 _1847_ (.B(_0387_),
    .A(_0386_),
    .X(_0055_));
 sg13g2_nand2_1 _1848_ (.Y(_0388_),
    .A(net280),
    .B(net223));
 sg13g2_nand2_1 _1849_ (.Y(_0389_),
    .A(net288),
    .B(net247));
 sg13g2_xor2_1 _1850_ (.B(_0389_),
    .A(_0388_),
    .X(_0057_));
 sg13g2_nand2_1 _1851_ (.Y(_0390_),
    .A(net312),
    .B(net263));
 sg13g2_nand2_1 _1852_ (.Y(_0391_),
    .A(net295),
    .B(net249));
 sg13g2_xor2_1 _1853_ (.B(_0391_),
    .A(_0390_),
    .X(_0059_));
 sg13g2_nand2_1 _1854_ (.Y(_0392_),
    .A(net294),
    .B(net245));
 sg13g2_nand2_1 _1855_ (.Y(_0393_),
    .A(net293),
    .B(net234));
 sg13g2_xor2_1 _1856_ (.B(_0393_),
    .A(_0392_),
    .X(_0063_));
 sg13g2_nand2_1 _1857_ (.Y(_0394_),
    .A(net301),
    .B(net236));
 sg13g2_nand2_1 _1858_ (.Y(_0395_),
    .A(net278),
    .B(net228));
 sg13g2_xor2_1 _1859_ (.B(_0395_),
    .A(_0394_),
    .X(_0065_));
 sg13g2_nand2_1 _1860_ (.Y(_0396_),
    .A(net300),
    .B(net243));
 sg13g2_nand2_1 _1861_ (.Y(_0397_),
    .A(net309),
    .B(net239));
 sg13g2_xor2_1 _1862_ (.B(_0397_),
    .A(_0396_),
    .X(_0067_));
 sg13g2_nand2_1 _1863_ (.Y(_0398_),
    .A(net302),
    .B(net250));
 sg13g2_nand2_1 _1864_ (.Y(_0399_),
    .A(net271),
    .B(net253));
 sg13g2_xor2_1 _1865_ (.B(_0399_),
    .A(_0398_),
    .X(_0069_));
 sg13g2_nand2_1 _1866_ (.Y(_0400_),
    .A(net315),
    .B(net238));
 sg13g2_nand2_1 _1867_ (.Y(_0401_),
    .A(net316),
    .B(net246));
 sg13g2_xor2_1 _1868_ (.B(_0401_),
    .A(_0400_),
    .X(_0071_));
 sg13g2_nand2_1 _1869_ (.Y(_0402_),
    .A(net284),
    .B(net232));
 sg13g2_nand2_1 _1870_ (.Y(_0403_),
    .A(net272),
    .B(net224));
 sg13g2_xor2_1 _1871_ (.B(_0403_),
    .A(_0402_),
    .X(_0073_));
 sg13g2_nand2_1 _1872_ (.Y(_0404_),
    .A(net287),
    .B(net229));
 sg13g2_nand2_1 _1873_ (.Y(_0405_),
    .A(net276),
    .B(net252));
 sg13g2_xor2_1 _1874_ (.B(_0405_),
    .A(_0404_),
    .X(_0075_));
 sg13g2_and2_1 _1875_ (.A(net2),
    .B(net1),
    .X(rst_n_sdr));
 sg13g2_and2_1 _1876_ (.A(net273),
    .B(net281),
    .X(_0040_));
 sg13g2_and2_1 _1877_ (.A(net304),
    .B(net275),
    .X(_0042_));
 sg13g2_and2_1 _1878_ (.A(net282),
    .B(net283),
    .X(_0044_));
 sg13g2_and2_1 _1879_ (.A(net299),
    .B(net277),
    .X(_0046_));
 sg13g2_and2_1 _1880_ (.A(net279),
    .B(net311),
    .X(_0048_));
 sg13g2_and2_1 _1881_ (.A(net303),
    .B(net310),
    .X(_0050_));
 sg13g2_and2_1 _1882_ (.A(net289),
    .B(net286),
    .X(_0052_));
 sg13g2_nand2_1 _1883_ (.Y(_0406_),
    .A(net734),
    .B(net217));
 sg13g2_xor2_1 _1884_ (.B(net217),
    .A(\sdr_i.mac1.products_ff[0] ),
    .X(_0015_));
 sg13g2_and2_1 _1885_ (.A(net285),
    .B(net274),
    .X(_0054_));
 sg13g2_xor2_1 _1886_ (.B(\sdr_i.mac1.products_ff[18] ),
    .A(\sdr_i.mac1.products_ff[1] ),
    .X(_0407_));
 sg13g2_xnor2_1 _1887_ (.Y(_0016_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_and2_1 _1888_ (.A(net288),
    .B(net280),
    .X(_0056_));
 sg13g2_and2_1 _1889_ (.A(net295),
    .B(net312),
    .X(_0058_));
 sg13g2_nand2_1 _1890_ (.Y(_0408_),
    .A(\sdr_i.mac2.products_ff[85] ),
    .B(net265));
 sg13g2_xor2_1 _1891_ (.B(net265),
    .A(\sdr_i.mac2.products_ff[85] ),
    .X(_0036_));
 sg13g2_xor2_1 _1892_ (.B(net754),
    .A(\sdr_i.mac2.products_ff[86] ),
    .X(_0409_));
 sg13g2_xnor2_1 _1893_ (.Y(_0037_),
    .A(_0408_),
    .B(net755));
 sg13g2_nand2_1 _1894_ (.Y(_0410_),
    .A(net757),
    .B(net254));
 sg13g2_xor2_1 _1895_ (.B(net254),
    .A(\sdr_i.mac2.products_ff[17] ),
    .X(_0032_));
 sg13g2_xor2_1 _1896_ (.B(\sdr_i.mac2.products_ff[1] ),
    .A(\sdr_i.mac2.products_ff[18] ),
    .X(_0411_));
 sg13g2_xnor2_1 _1897_ (.Y(_0033_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_and2_1 _1898_ (.A(net290),
    .B(net296),
    .X(_0060_));
 sg13g2_and2_1 _1899_ (.A(net293),
    .B(net294),
    .X(_0062_));
 sg13g2_and2_1 _1900_ (.A(net278),
    .B(net301),
    .X(_0064_));
 sg13g2_and2_1 _1901_ (.A(net309),
    .B(net300),
    .X(_0066_));
 sg13g2_and2_1 _1902_ (.A(net271),
    .B(net302),
    .X(_0068_));
 sg13g2_and2_1 _1903_ (.A(net316),
    .B(net315),
    .X(_0070_));
 sg13g2_and2_1 _1904_ (.A(net272),
    .B(net284),
    .X(_0072_));
 sg13g2_nand2_1 _1905_ (.Y(_0412_),
    .A(net774),
    .B(net261));
 sg13g2_xor2_1 _1906_ (.B(net261),
    .A(\sdr_i.mac1.sum_lvl3_ff[2] ),
    .X(_0030_));
 sg13g2_nand2_1 _1907_ (.Y(_0413_),
    .A(net552),
    .B(\sdr_i.mac1.sum_lvl3_ff[1] ));
 sg13g2_nor2_1 _1908_ (.A(net552),
    .B(\sdr_i.mac1.sum_lvl3_ff[1] ),
    .Y(_0414_));
 sg13g2_xor2_1 _1909_ (.B(\sdr_i.mac1.sum_lvl3_ff[1] ),
    .A(net552),
    .X(_0415_));
 sg13g2_xnor2_1 _1910_ (.Y(_0031_),
    .A(_0412_),
    .B(_0415_));
 sg13g2_and2_1 _1911_ (.A(net276),
    .B(net287),
    .X(_0074_));
 sg13g2_nand2_1 _1912_ (.Y(_0416_),
    .A(\sdr_i.mac2.sum_lvl3_ff[2] ),
    .B(net259));
 sg13g2_xor2_1 _1913_ (.B(net259),
    .A(\sdr_i.mac2.sum_lvl3_ff[2] ),
    .X(_0007_));
 sg13g2_nand2_1 _1914_ (.Y(_0417_),
    .A(net601),
    .B(\sdr_i.mac2.sum_lvl3_ff[1] ));
 sg13g2_nor2_1 _1915_ (.A(net601),
    .B(\sdr_i.mac2.sum_lvl3_ff[1] ),
    .Y(_0418_));
 sg13g2_xor2_1 _1916_ (.B(net782),
    .A(net601),
    .X(_0419_));
 sg13g2_xnor2_1 _1917_ (.Y(_0008_),
    .A(_0416_),
    .B(_0419_));
 sg13g2_nand2_1 _1918_ (.Y(_0420_),
    .A(net764),
    .B(net297));
 sg13g2_xor2_1 _1919_ (.B(net297),
    .A(\sdr_i.mac2.sum_lvl2_ff[4] ),
    .X(_0009_));
 sg13g2_xor2_1 _1920_ (.B(\sdr_i.mac2.sum_lvl2_ff[1] ),
    .A(\sdr_i.mac2.sum_lvl2_ff[5] ),
    .X(_0421_));
 sg13g2_xnor2_1 _1921_ (.Y(_0010_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_nand2_1 _1922_ (.Y(_0422_),
    .A(net731),
    .B(net291));
 sg13g2_xor2_1 _1923_ (.B(net291),
    .A(\sdr_i.mac2.sum_lvl1_ff[8] ),
    .X(_0013_));
 sg13g2_xor2_1 _1924_ (.B(\sdr_i.mac2.sum_lvl1_ff[1] ),
    .A(\sdr_i.mac2.sum_lvl1_ff[9] ),
    .X(_0423_));
 sg13g2_xnor2_1 _1925_ (.Y(_0014_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_nand2_1 _1926_ (.Y(_0424_),
    .A(net778),
    .B(net313));
 sg13g2_xor2_1 _1927_ (.B(net313),
    .A(\sdr_i.mac1.products_ff[51] ),
    .X(_0017_));
 sg13g2_xor2_1 _1928_ (.B(\sdr_i.mac1.products_ff[35] ),
    .A(\sdr_i.mac1.products_ff[52] ),
    .X(_0425_));
 sg13g2_xnor2_1 _1929_ (.Y(_0018_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_nand2_1 _1930_ (.Y(_0426_),
    .A(net741),
    .B(net307));
 sg13g2_xor2_1 _1931_ (.B(net307),
    .A(\sdr_i.mac1.products_ff[68] ),
    .X(_0019_));
 sg13g2_xor2_1 _1932_ (.B(\sdr_i.mac1.products_ff[86] ),
    .A(\sdr_i.mac1.products_ff[69] ),
    .X(_0427_));
 sg13g2_xnor2_1 _1933_ (.Y(_0020_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_nand2_1 _1934_ (.Y(_0428_),
    .A(\sdr_i.mac1.products_ff[119] ),
    .B(net230));
 sg13g2_xor2_1 _1935_ (.B(net230),
    .A(\sdr_i.mac1.products_ff[119] ),
    .X(_0021_));
 sg13g2_xor2_1 _1936_ (.B(net761),
    .A(\sdr_i.mac1.products_ff[120] ),
    .X(_0429_));
 sg13g2_xnor2_1 _1937_ (.Y(_0022_),
    .A(_0428_),
    .B(net762));
 sg13g2_nand2_1 _1938_ (.Y(_0430_),
    .A(\sdr_i.mac1.sum_lvl1_ff[8] ),
    .B(net215));
 sg13g2_xor2_1 _1939_ (.B(net215),
    .A(\sdr_i.mac1.sum_lvl1_ff[8] ),
    .X(_0023_));
 sg13g2_xor2_1 _1940_ (.B(net736),
    .A(\sdr_i.mac1.sum_lvl1_ff[9] ),
    .X(_0431_));
 sg13g2_xnor2_1 _1941_ (.Y(_0024_),
    .A(_0430_),
    .B(net737));
 sg13g2_nand2_1 _1942_ (.Y(_0432_),
    .A(net746),
    .B(net267));
 sg13g2_xor2_1 _1943_ (.B(net267),
    .A(\sdr_i.mac1.sum_lvl1_ff[24] ),
    .X(_0025_));
 sg13g2_xor2_1 _1944_ (.B(\sdr_i.mac1.sum_lvl1_ff[17] ),
    .A(\sdr_i.mac1.sum_lvl1_ff[25] ),
    .X(_0433_));
 sg13g2_xnor2_1 _1945_ (.Y(_0026_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_nand2_1 _1946_ (.Y(_0434_),
    .A(\sdr_i.mac1.sum_lvl2_ff[4] ),
    .B(net305));
 sg13g2_xor2_1 _1947_ (.B(net305),
    .A(\sdr_i.mac1.sum_lvl2_ff[4] ),
    .X(_0027_));
 sg13g2_xor2_1 _1948_ (.B(net743),
    .A(\sdr_i.mac1.sum_lvl2_ff[5] ),
    .X(_0435_));
 sg13g2_xnor2_1 _1949_ (.Y(_0028_),
    .A(_0434_),
    .B(net744));
 sg13g2_nand2_1 _1950_ (.Y(_0436_),
    .A(net729),
    .B(net213));
 sg13g2_xor2_1 _1951_ (.B(net213),
    .A(\sdr_i.mac2.products_ff[34] ),
    .X(_0034_));
 sg13g2_xor2_1 _1952_ (.B(\sdr_i.mac2.products_ff[52] ),
    .A(\sdr_i.mac2.products_ff[35] ),
    .X(_0437_));
 sg13g2_xnor2_1 _1953_ (.Y(_0035_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_nand2_1 _1954_ (.Y(_0438_),
    .A(net739),
    .B(net257));
 sg13g2_xor2_1 _1955_ (.B(net257),
    .A(\sdr_i.mac2.products_ff[102] ),
    .X(_0038_));
 sg13g2_xor2_1 _1956_ (.B(\sdr_i.mac2.products_ff[120] ),
    .A(\sdr_i.mac2.products_ff[103] ),
    .X(_0439_));
 sg13g2_xnor2_1 _1957_ (.Y(_0039_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nand2_1 _1958_ (.Y(_0440_),
    .A(net269),
    .B(\sdr_i.mac2.sum_lvl1_ff[16] ));
 sg13g2_xor2_1 _1959_ (.B(\sdr_i.mac2.sum_lvl1_ff[16] ),
    .A(net269),
    .X(_0011_));
 sg13g2_xor2_1 _1960_ (.B(net722),
    .A(\sdr_i.mac2.sum_lvl1_ff[25] ),
    .X(_0441_));
 sg13g2_xnor2_1 _1961_ (.Y(_0012_),
    .A(_0440_),
    .B(net723));
 sg13g2_nand2_1 _1962_ (.Y(_0442_),
    .A(net290),
    .B(net222));
 sg13g2_nand2_1 _1963_ (.Y(_0443_),
    .A(net296),
    .B(net219));
 sg13g2_xor2_1 _1964_ (.B(_0443_),
    .A(_0442_),
    .X(_0061_));
 sg13g2_o21ai_1 _1965_ (.B1(net553),
    .Y(_0029_),
    .A1(_0412_),
    .A2(_0414_));
 sg13g2_nand2_1 _1966_ (.Y(_0444_),
    .A(net273),
    .B(net241));
 sg13g2_nand2_1 _1967_ (.Y(_0445_),
    .A(net281),
    .B(net240));
 sg13g2_xor2_1 _1968_ (.B(_0445_),
    .A(_0444_),
    .X(_0041_));
 sg13g2_nand2_1 _1969_ (.Y(_0446_),
    .A(net304),
    .B(net226));
 sg13g2_nand2_1 _1970_ (.Y(_0447_),
    .A(net275),
    .B(net235));
 sg13g2_xor2_1 _1971_ (.B(_0447_),
    .A(_0446_),
    .X(_0043_));
 sg13g2_o21ai_1 _1972_ (.B1(net602),
    .Y(_0006_),
    .A1(_0416_),
    .A2(_0418_));
 sg13g2_nand2_1 _1973_ (.Y(_0448_),
    .A(net283),
    .B(net242));
 sg13g2_nand2_1 _1974_ (.Y(_0449_),
    .A(net282),
    .B(net227));
 sg13g2_xor2_1 _1975_ (.B(_0449_),
    .A(_0448_),
    .X(_0045_));
 sg13g2_nand2_1 _1976_ (.Y(_0450_),
    .A(net299),
    .B(net251));
 sg13g2_nand2_1 _1977_ (.Y(_0451_),
    .A(net277),
    .B(net256));
 sg13g2_xor2_1 _1978_ (.B(_0451_),
    .A(_0450_),
    .X(_0047_));
 sg13g2_nand2_1 _1979_ (.Y(_0452_),
    .A(net279),
    .B(net248));
 sg13g2_nand2_1 _1980_ (.Y(_0453_),
    .A(net311),
    .B(net244));
 sg13g2_xor2_1 _1981_ (.B(_0453_),
    .A(_0452_),
    .X(_0049_));
 sg13g2_nand2_1 _1982_ (.Y(_0454_),
    .A(net310),
    .B(net264));
 sg13g2_nand2_1 _1983_ (.Y(_0455_),
    .A(net303),
    .B(net225));
 sg13g2_xor2_1 _1984_ (.B(_0455_),
    .A(_0454_),
    .X(_0051_));
 sg13g2_xor2_1 _1985_ (.B(\ppwm_i.u_ppwm.global_counter[0] ),
    .A(net326),
    .X(_0148_));
 sg13g2_nand3_1 _1986_ (.B(net822),
    .C(\ppwm_i.u_ppwm.global_counter[0] ),
    .A(net326),
    .Y(_0456_));
 sg13g2_a21o_1 _1987_ (.A2(\ppwm_i.u_ppwm.global_counter[0] ),
    .A1(net326),
    .B1(net822),
    .X(_0457_));
 sg13g2_and2_1 _1988_ (.A(_0456_),
    .B(net823),
    .X(_0149_));
 sg13g2_and4_1 _1989_ (.A(net326),
    .B(net710),
    .C(\ppwm_i.u_ppwm.global_counter[1] ),
    .D(\ppwm_i.u_ppwm.global_counter[0] ),
    .X(_0458_));
 sg13g2_xnor2_1 _1990_ (.Y(_0150_),
    .A(net710),
    .B(_0456_));
 sg13g2_xnor2_1 _1991_ (.Y(_0151_),
    .A(_1264_),
    .B(_0458_));
 sg13g2_nand3_1 _1992_ (.B(net789),
    .C(_0458_),
    .A(net806),
    .Y(_0459_));
 sg13g2_a21o_1 _1993_ (.A2(_0458_),
    .A1(net789),
    .B1(net806),
    .X(_0460_));
 sg13g2_and2_1 _1994_ (.A(_0459_),
    .B(_0460_),
    .X(_0152_));
 sg13g2_nand4_1 _1995_ (.B(\ppwm_i.u_ppwm.global_counter[4] ),
    .C(\ppwm_i.u_ppwm.global_counter[3] ),
    .A(net333),
    .Y(_0461_),
    .D(_0458_));
 sg13g2_xnor2_1 _1996_ (.Y(_0153_),
    .A(net333),
    .B(_0459_));
 sg13g2_nor2_1 _1997_ (.A(_1261_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_xnor2_1 _1998_ (.Y(_0154_),
    .A(net320),
    .B(_0461_));
 sg13g2_xor2_1 _1999_ (.B(_0462_),
    .A(net654),
    .X(_0155_));
 sg13g2_nand3_1 _2000_ (.B(net654),
    .C(_0462_),
    .A(net807),
    .Y(_0463_));
 sg13g2_a21o_1 _2001_ (.A2(_0462_),
    .A1(net654),
    .B1(net807),
    .X(_0464_));
 sg13g2_and2_1 _2002_ (.A(_0463_),
    .B(_0464_),
    .X(_0156_));
 sg13g2_nor2_2 _2003_ (.A(_1259_),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_xnor2_1 _2004_ (.Y(_0157_),
    .A(net335),
    .B(_0463_));
 sg13g2_and2_1 _2005_ (.A(net557),
    .B(_0465_),
    .X(_0466_));
 sg13g2_xor2_1 _2006_ (.B(_0465_),
    .A(net557),
    .X(_0158_));
 sg13g2_xnor2_1 _2007_ (.Y(_0159_),
    .A(_1258_),
    .B(_0466_));
 sg13g2_and3_2 _2008_ (.X(_0467_),
    .A(net719),
    .B(net787),
    .C(_0466_));
 sg13g2_a21oi_1 _2009_ (.A1(\ppwm_i.u_ppwm.global_counter[11] ),
    .A2(_0466_),
    .Y(_0468_),
    .B1(net719));
 sg13g2_nor2_1 _2010_ (.A(_0467_),
    .B(net720),
    .Y(_0160_));
 sg13g2_xnor2_1 _2011_ (.Y(_0161_),
    .A(_1256_),
    .B(_0467_));
 sg13g2_nand3_1 _2012_ (.B(net776),
    .C(_0467_),
    .A(net813),
    .Y(_0469_));
 sg13g2_a21o_1 _2013_ (.A2(_0467_),
    .A1(net776),
    .B1(net813),
    .X(_0470_));
 sg13g2_and2_1 _2014_ (.A(_0469_),
    .B(_0470_),
    .X(_0162_));
 sg13g2_nor2_1 _2015_ (.A(_1255_),
    .B(_0469_),
    .Y(_0471_));
 sg13g2_xnor2_1 _2016_ (.Y(_0163_),
    .A(net572),
    .B(_0469_));
 sg13g2_nor3_2 _2017_ (.A(_1254_),
    .B(_1255_),
    .C(_0469_),
    .Y(_0472_));
 sg13g2_xnor2_1 _2018_ (.Y(_0164_),
    .A(_1254_),
    .B(_0471_));
 sg13g2_xnor2_1 _2019_ (.Y(_0165_),
    .A(_1253_),
    .B(_0472_));
 sg13g2_nand3_1 _2020_ (.B(net798),
    .C(_0472_),
    .A(net804),
    .Y(_0473_));
 sg13g2_a21o_1 _2021_ (.A2(_0472_),
    .A1(net798),
    .B1(net804),
    .X(_0474_));
 sg13g2_and2_1 _2022_ (.A(_0473_),
    .B(_0474_),
    .X(_0166_));
 sg13g2_xnor2_1 _2023_ (.Y(_0167_),
    .A(net328),
    .B(_0473_));
 sg13g2_nor4_1 _2024_ (.A(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .Y(_0475_));
 sg13g2_nor4_1 _2025_ (.A(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .C(net520),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .Y(_0476_));
 sg13g2_nand4_1 _2026_ (.B(_1236_),
    .C(_0475_),
    .A(_1234_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_o21ai_1 _2027_ (.B1(net421),
    .Y(_0478_),
    .A1(\ppwm_i.u_ppwm.pwm_value[0] ),
    .A2(net409));
 sg13g2_a21oi_1 _2028_ (.A1(_1247_),
    .A2(net409),
    .Y(_0168_),
    .B1(_0478_));
 sg13g2_nor2_1 _2029_ (.A(net507),
    .B(net409),
    .Y(_0479_));
 sg13g2_nor2b_1 _2030_ (.A(net578),
    .B_N(net409),
    .Y(_0480_));
 sg13g2_nor3_1 _2031_ (.A(net457),
    .B(_0479_),
    .C(_0480_),
    .Y(_0169_));
 sg13g2_nor2_1 _2032_ (.A(net794),
    .B(net409),
    .Y(_0481_));
 sg13g2_a21oi_1 _2033_ (.A1(_1246_),
    .A2(net409),
    .Y(_0482_),
    .B1(net456));
 sg13g2_nor2b_1 _2034_ (.A(_0481_),
    .B_N(_0482_),
    .Y(_0170_));
 sg13g2_nor2_1 _2035_ (.A(net770),
    .B(net411),
    .Y(_0483_));
 sg13g2_a21oi_1 _2036_ (.A1(_1245_),
    .A2(net409),
    .Y(_0484_),
    .B1(net456));
 sg13g2_nor2b_1 _2037_ (.A(net771),
    .B_N(_0484_),
    .Y(_0171_));
 sg13g2_nand2_1 _2038_ (.Y(_0485_),
    .A(_1244_),
    .B(net410));
 sg13g2_o21ai_1 _2039_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net505),
    .A2(net409));
 sg13g2_nor2_1 _2040_ (.A(net456),
    .B(net797),
    .Y(_0172_));
 sg13g2_nand2_1 _2041_ (.Y(_0487_),
    .A(_1243_),
    .B(net410));
 sg13g2_o21ai_1 _2042_ (.B1(_0487_),
    .Y(_0488_),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ),
    .A2(net410));
 sg13g2_nor2_1 _2043_ (.A(net455),
    .B(net792),
    .Y(_0173_));
 sg13g2_nor2_1 _2044_ (.A(net504),
    .B(net411),
    .Y(_0489_));
 sg13g2_nor2b_1 _2045_ (.A(net664),
    .B_N(net410),
    .Y(_0490_));
 sg13g2_nor3_1 _2046_ (.A(net456),
    .B(_0489_),
    .C(_0490_),
    .Y(_0174_));
 sg13g2_nor2_1 _2047_ (.A(net503),
    .B(net410),
    .Y(_0491_));
 sg13g2_nor2b_1 _2048_ (.A(net580),
    .B_N(net411),
    .Y(_0492_));
 sg13g2_nor3_1 _2049_ (.A(net455),
    .B(_0491_),
    .C(_0492_),
    .Y(_0175_));
 sg13g2_nand2_1 _2050_ (.Y(_0493_),
    .A(_1242_),
    .B(net410));
 sg13g2_o21ai_1 _2051_ (.B1(_0493_),
    .Y(_0494_),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .A2(net410));
 sg13g2_nor2_1 _2052_ (.A(net456),
    .B(net803),
    .Y(_0176_));
 sg13g2_nand2_1 _2053_ (.Y(_0495_),
    .A(_1241_),
    .B(net410));
 sg13g2_o21ai_1 _2054_ (.B1(_0495_),
    .Y(_0496_),
    .A1(net793),
    .A2(net411));
 sg13g2_nor2_1 _2055_ (.A(net455),
    .B(_0496_),
    .Y(_0177_));
 sg13g2_xnor2_1 _2056_ (.Y(_0497_),
    .A(net715),
    .B(net769));
 sg13g2_nor2_1 _2057_ (.A(net455),
    .B(_0497_),
    .Y(_0178_));
 sg13g2_a21oi_1 _2058_ (.A1(\ppwm_i.u_ppwm.mem_write_done ),
    .A2(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .Y(_0498_),
    .B1(net707));
 sg13g2_and3_1 _2059_ (.X(_0499_),
    .A(net715),
    .B(net707),
    .C(net769));
 sg13g2_nor3_1 _2060_ (.A(net455),
    .B(net708),
    .C(_0499_),
    .Y(_0179_));
 sg13g2_and2_1 _2061_ (.A(net784),
    .B(_0499_),
    .X(_0500_));
 sg13g2_o21ai_1 _2062_ (.B1(net422),
    .Y(_0501_),
    .A1(net784),
    .A2(_0499_));
 sg13g2_nor2_1 _2063_ (.A(_0500_),
    .B(_0501_),
    .Y(_0180_));
 sg13g2_and2_1 _2064_ (.A(net786),
    .B(_0500_),
    .X(_0502_));
 sg13g2_o21ai_1 _2065_ (.B1(net422),
    .Y(_0503_),
    .A1(net786),
    .A2(_0500_));
 sg13g2_nor2_1 _2066_ (.A(_0502_),
    .B(_0503_),
    .Y(_0181_));
 sg13g2_and2_1 _2067_ (.A(net785),
    .B(_0502_),
    .X(_0504_));
 sg13g2_o21ai_1 _2068_ (.B1(net422),
    .Y(_0505_),
    .A1(net785),
    .A2(_0502_));
 sg13g2_nor2_1 _2069_ (.A(_0504_),
    .B(_0505_),
    .Y(_0182_));
 sg13g2_nand4_1 _2070_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .A(net565),
    .Y(_0506_),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[2] ));
 sg13g2_o21ai_1 _2071_ (.B1(net422),
    .Y(_0507_),
    .A1(net520),
    .A2(_0504_));
 sg13g2_a21oi_1 _2072_ (.A1(net520),
    .A2(_0504_),
    .Y(_0183_),
    .B1(_0507_));
 sg13g2_a21o_1 _2073_ (.A2(_0504_),
    .A1(net520),
    .B1(net808),
    .X(_0508_));
 sg13g2_nand3_1 _2074_ (.B(net520),
    .C(_0504_),
    .A(net808),
    .Y(_0509_));
 sg13g2_and3_1 _2075_ (.X(_0184_),
    .A(net422),
    .B(_0508_),
    .C(_0509_));
 sg13g2_and2_1 _2076_ (.A(_1237_),
    .B(_0509_),
    .X(_0510_));
 sg13g2_and4_1 _2077_ (.A(net819),
    .B(net808),
    .C(net520),
    .D(_0504_),
    .X(_0511_));
 sg13g2_nor3_1 _2078_ (.A(net455),
    .B(_0510_),
    .C(_0511_),
    .Y(_0185_));
 sg13g2_nor2_1 _2079_ (.A(net766),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_and2_1 _2080_ (.A(net766),
    .B(_0511_),
    .X(_0513_));
 sg13g2_nor3_1 _2081_ (.A(net455),
    .B(net767),
    .C(_0513_),
    .Y(_0186_));
 sg13g2_xnor2_1 _2082_ (.Y(_0514_),
    .A(net752),
    .B(_0513_));
 sg13g2_nor2_1 _2083_ (.A(net455),
    .B(net753),
    .Y(_0187_));
 sg13g2_nand3_1 _2084_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .C(net423),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .Y(_0515_));
 sg13g2_nand4_1 _2085_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .Y(_0516_),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[0] ));
 sg13g2_nor3_1 _2086_ (.A(net566),
    .B(_0515_),
    .C(_0516_),
    .Y(_0188_));
 sg13g2_nor2b_1 _2087_ (.A(net395),
    .B_N(_0365_),
    .Y(_0517_));
 sg13g2_o21ai_1 _2088_ (.B1(_0517_),
    .Y(_0518_),
    .A1(\ppwm_i.u_ppwm.u_ex.cmp_flag_q ),
    .A2(net394));
 sg13g2_nor2_1 _2089_ (.A(net401),
    .B(_0518_),
    .Y(_0519_));
 sg13g2_nor2_1 _2090_ (.A(_1232_),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_o21ai_1 _2091_ (.B1(net427),
    .Y(_0521_),
    .A1(net518),
    .A2(_0520_));
 sg13g2_a21oi_1 _2092_ (.A1(net518),
    .A2(_0520_),
    .Y(_0189_),
    .B1(_0521_));
 sg13g2_and2_1 _2093_ (.A(net518),
    .B(net401),
    .X(_0522_));
 sg13g2_and2_1 _2094_ (.A(net515),
    .B(net396),
    .X(_0523_));
 sg13g2_xor2_1 _2095_ (.B(net397),
    .A(net515),
    .X(_0524_));
 sg13g2_nand2_1 _2096_ (.Y(_0525_),
    .A(_1232_),
    .B(net515));
 sg13g2_o21ai_1 _2097_ (.B1(_0518_),
    .Y(_0526_),
    .A1(net451),
    .A2(net449));
 sg13g2_xor2_1 _2098_ (.B(_0524_),
    .A(_0522_),
    .X(_0527_));
 sg13g2_o21ai_1 _2099_ (.B1(net768),
    .Y(_0528_),
    .A1(_0518_),
    .A2(_0527_));
 sg13g2_nand2b_1 _2100_ (.Y(_0529_),
    .B(_0526_),
    .A_N(_0528_));
 sg13g2_a21oi_1 _2101_ (.A1(_0525_),
    .A2(_0529_),
    .Y(_0190_),
    .B1(net458));
 sg13g2_a21oi_1 _2102_ (.A1(_0522_),
    .A2(_0524_),
    .Y(_0530_),
    .B1(_0523_));
 sg13g2_nand2_1 _2103_ (.Y(_0531_),
    .A(net511),
    .B(net389));
 sg13g2_xnor2_1 _2104_ (.Y(_0532_),
    .A(net511),
    .B(net389));
 sg13g2_xnor2_1 _2105_ (.Y(_0533_),
    .A(net511),
    .B(net451));
 sg13g2_nand2_1 _2106_ (.Y(_0534_),
    .A(_1232_),
    .B(net512));
 sg13g2_xor2_1 _2107_ (.B(_0532_),
    .A(_0530_),
    .X(_0535_));
 sg13g2_a21oi_1 _2108_ (.A1(_0518_),
    .A2(_0533_),
    .Y(_0536_),
    .B1(_1232_));
 sg13g2_o21ai_1 _2109_ (.B1(_0536_),
    .Y(_0537_),
    .A1(_0518_),
    .A2(_0535_));
 sg13g2_a21oi_1 _2110_ (.A1(_0534_),
    .A2(_0537_),
    .Y(_0191_),
    .B1(net458));
 sg13g2_nor2_1 _2111_ (.A(_1231_),
    .B(net406),
    .Y(_0538_));
 sg13g2_nor2_1 _2112_ (.A(net408),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_o21ai_1 _2113_ (.B1(_0531_),
    .Y(_0540_),
    .A1(_0530_),
    .A2(_0532_));
 sg13g2_a21oi_1 _2114_ (.A1(_0539_),
    .A2(_0540_),
    .Y(_0541_),
    .B1(_0518_));
 sg13g2_o21ai_1 _2115_ (.B1(_0541_),
    .Y(_0542_),
    .A1(_0539_),
    .A2(_0540_));
 sg13g2_a21oi_1 _2116_ (.A1(net511),
    .A2(net451),
    .Y(_0543_),
    .B1(net508));
 sg13g2_o21ai_1 _2117_ (.B1(_0518_),
    .Y(_0544_),
    .A1(_1277_),
    .A2(_0543_));
 sg13g2_and2_1 _2118_ (.A(net768),
    .B(_0544_),
    .X(_0545_));
 sg13g2_a22oi_1 _2119_ (.Y(_0546_),
    .B1(_0542_),
    .B2(_0545_),
    .A2(_1232_),
    .A1(net508));
 sg13g2_nor2_1 _2120_ (.A(net458),
    .B(_0546_),
    .Y(_0192_));
 sg13g2_and2_1 _2121_ (.A(net395),
    .B(_0365_),
    .X(_0547_));
 sg13g2_nand2_1 _2122_ (.Y(_0548_),
    .A(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .B(_0547_));
 sg13g2_nor2_1 _2123_ (.A(net394),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_o21ai_1 _2124_ (.B1(net349),
    .Y(_0550_),
    .A1(net394),
    .A2(_0548_));
 sg13g2_nand2_2 _2125_ (.Y(_0551_),
    .A(_1311_),
    .B(net388));
 sg13g2_a22oi_1 _2126_ (.Y(_0552_),
    .B1(\ppwm_i.u_ppwm.global_counter[18] ),
    .B2(_1221_),
    .A2(\ppwm_i.u_ppwm.global_counter[19] ),
    .A1(_1220_));
 sg13g2_nor2_1 _2127_ (.A(\ppwm_i.u_ppwm.pwm_value[3] ),
    .B(_1256_),
    .Y(_0553_));
 sg13g2_nand2b_1 _2128_ (.Y(_0554_),
    .B(net507),
    .A_N(\ppwm_i.u_ppwm.global_counter[11] ));
 sg13g2_nor2b_1 _2129_ (.A(net507),
    .B_N(\ppwm_i.u_ppwm.global_counter[11] ),
    .Y(_0555_));
 sg13g2_nand2b_1 _2130_ (.Y(_0556_),
    .B(\ppwm_i.u_ppwm.pwm_value[0] ),
    .A_N(\ppwm_i.u_ppwm.global_counter[10] ));
 sg13g2_a221oi_1 _2131_ (.B2(_0556_),
    .C1(_0555_),
    .B1(_0554_),
    .A1(_1227_),
    .Y(_0557_),
    .A2(\ppwm_i.u_ppwm.global_counter[12] ));
 sg13g2_nand2b_1 _2132_ (.Y(_0558_),
    .B(net505),
    .A_N(\ppwm_i.u_ppwm.global_counter[14] ));
 sg13g2_a221oi_1 _2133_ (.B2(\ppwm_i.u_ppwm.pwm_value[2] ),
    .C1(_0557_),
    .B1(_1257_),
    .A1(net506),
    .Y(_0559_),
    .A2(_1256_));
 sg13g2_o21ai_1 _2134_ (.B1(_0558_),
    .Y(_0560_),
    .A1(_0553_),
    .A2(_0559_));
 sg13g2_a22oi_1 _2135_ (.Y(_0561_),
    .B1(\ppwm_i.u_ppwm.global_counter[14] ),
    .B2(_1225_),
    .A2(\ppwm_i.u_ppwm.global_counter[15] ),
    .A1(_1224_));
 sg13g2_nor2_1 _2136_ (.A(_1224_),
    .B(\ppwm_i.u_ppwm.global_counter[15] ),
    .Y(_0562_));
 sg13g2_a221oi_1 _2137_ (.B2(_0561_),
    .C1(_0562_),
    .B1(_0560_),
    .A1(net504),
    .Y(_0563_),
    .A2(_1254_));
 sg13g2_nand2_1 _2138_ (.Y(_0564_),
    .A(_1222_),
    .B(\ppwm_i.u_ppwm.global_counter[17] ));
 sg13g2_o21ai_1 _2139_ (.B1(_0564_),
    .Y(_0565_),
    .A1(net504),
    .A2(_1254_));
 sg13g2_a22oi_1 _2140_ (.Y(_0566_),
    .B1(_1253_),
    .B2(net503),
    .A2(_1252_),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ));
 sg13g2_o21ai_1 _2141_ (.B1(_0566_),
    .Y(_0567_),
    .A1(_0563_),
    .A2(_0565_));
 sg13g2_a22oi_1 _2142_ (.Y(_0568_),
    .B1(_0552_),
    .B2(_0567_),
    .A2(_1251_),
    .A1(\ppwm_i.u_ppwm.pwm_value[9] ));
 sg13g2_nand2_1 _2143_ (.Y(_0569_),
    .A(_1211_),
    .B(\ppwm_i.u_ppwm.global_counter[18] ));
 sg13g2_nor2b_1 _2144_ (.A(\ppwm_i.u_ppwm.global_counter[10] ),
    .B_N(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .Y(_0570_));
 sg13g2_o21ai_1 _2145_ (.B1(_0570_),
    .Y(_0571_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(_1258_));
 sg13g2_a22oi_1 _2146_ (.Y(_0572_),
    .B1(_1258_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(_1257_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ));
 sg13g2_nor2_1 _2147_ (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .B(_1256_),
    .Y(_0573_));
 sg13g2_a221oi_1 _2148_ (.B2(_0572_),
    .C1(_0573_),
    .B1(_0571_),
    .A1(_1217_),
    .Y(_0574_),
    .A2(\ppwm_i.u_ppwm.global_counter[12] ));
 sg13g2_nand2_1 _2149_ (.Y(_0575_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .B(_1256_));
 sg13g2_o21ai_1 _2150_ (.B1(_0575_),
    .Y(_0576_),
    .A1(_1215_),
    .A2(\ppwm_i.u_ppwm.global_counter[14] ));
 sg13g2_a22oi_1 _2151_ (.Y(_0577_),
    .B1(\ppwm_i.u_ppwm.global_counter[14] ),
    .B2(_1215_),
    .A2(\ppwm_i.u_ppwm.global_counter[15] ),
    .A1(_1214_));
 sg13g2_o21ai_1 _2152_ (.B1(_0577_),
    .Y(_0578_),
    .A1(_0574_),
    .A2(_0576_));
 sg13g2_a22oi_1 _2153_ (.Y(_0579_),
    .B1(_1255_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A2(_1254_),
    .A1(net502));
 sg13g2_nor2b_1 _2154_ (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .B_N(\ppwm_i.u_ppwm.global_counter[17] ),
    .Y(_0580_));
 sg13g2_a221oi_1 _2155_ (.B2(_0579_),
    .C1(_0580_),
    .B1(_0578_),
    .A1(_1213_),
    .Y(_0581_),
    .A2(\ppwm_i.u_ppwm.global_counter[16] ));
 sg13g2_nor2_1 _2156_ (.A(_1212_),
    .B(\ppwm_i.u_ppwm.global_counter[17] ),
    .Y(_0582_));
 sg13g2_o21ai_1 _2157_ (.B1(_0569_),
    .Y(_0583_),
    .A1(_0581_),
    .A2(_0582_));
 sg13g2_a22oi_1 _2158_ (.Y(_0584_),
    .B1(_1252_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .A2(_1251_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ));
 sg13g2_nand2_2 _2159_ (.Y(_0585_),
    .A(net398),
    .B(_1311_));
 sg13g2_nand2_1 _2160_ (.Y(_0586_),
    .A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .B(_1259_));
 sg13g2_a22oi_1 _2161_ (.Y(_0587_),
    .B1(\ppwm_i.u_ppwm.global_counter[8] ),
    .B2(_1221_),
    .A2(\ppwm_i.u_ppwm.global_counter[9] ),
    .A1(_1220_));
 sg13g2_nand2_1 _2162_ (.Y(_0588_),
    .A(_1227_),
    .B(\ppwm_i.u_ppwm.global_counter[2] ));
 sg13g2_nor2b_1 _2163_ (.A(\ppwm_i.u_ppwm.pwm_value[1] ),
    .B_N(\ppwm_i.u_ppwm.global_counter[1] ),
    .Y(_0589_));
 sg13g2_nand2b_1 _2164_ (.Y(_0590_),
    .B(\ppwm_i.u_ppwm.pwm_value[0] ),
    .A_N(\ppwm_i.u_ppwm.global_counter[0] ));
 sg13g2_nand2b_1 _2165_ (.Y(_0591_),
    .B(\ppwm_i.u_ppwm.pwm_value[1] ),
    .A_N(\ppwm_i.u_ppwm.global_counter[1] ));
 sg13g2_o21ai_1 _2166_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0589_),
    .A2(_0590_));
 sg13g2_nor2_1 _2167_ (.A(_1227_),
    .B(\ppwm_i.u_ppwm.global_counter[2] ),
    .Y(_0593_));
 sg13g2_a221oi_1 _2168_ (.B2(_0592_),
    .C1(_0593_),
    .B1(_0588_),
    .A1(net506),
    .Y(_0594_),
    .A2(_1264_));
 sg13g2_nand2_1 _2169_ (.Y(_0595_),
    .A(_1226_),
    .B(\ppwm_i.u_ppwm.global_counter[3] ));
 sg13g2_o21ai_1 _2170_ (.B1(_0595_),
    .Y(_0596_),
    .A1(net505),
    .A2(_1263_));
 sg13g2_a22oi_1 _2171_ (.Y(_0597_),
    .B1(_1263_),
    .B2(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A2(_1262_),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ));
 sg13g2_o21ai_1 _2172_ (.B1(_0597_),
    .Y(_0598_),
    .A1(_0594_),
    .A2(_0596_));
 sg13g2_nand2_1 _2173_ (.Y(_0599_),
    .A(_1224_),
    .B(\ppwm_i.u_ppwm.global_counter[5] ));
 sg13g2_a22oi_1 _2174_ (.Y(_0600_),
    .B1(_0598_),
    .B2(_0599_),
    .A2(_1261_),
    .A1(net504));
 sg13g2_a221oi_1 _2175_ (.B2(_1223_),
    .C1(_0600_),
    .B1(\ppwm_i.u_ppwm.global_counter[6] ),
    .A1(_1222_),
    .Y(_0601_),
    .A2(\ppwm_i.u_ppwm.global_counter[7] ));
 sg13g2_nand2b_1 _2176_ (.Y(_0602_),
    .B(net503),
    .A_N(\ppwm_i.u_ppwm.global_counter[7] ));
 sg13g2_o21ai_1 _2177_ (.B1(_0602_),
    .Y(_0603_),
    .A1(_1221_),
    .A2(\ppwm_i.u_ppwm.global_counter[8] ));
 sg13g2_o21ai_1 _2178_ (.B1(_0587_),
    .Y(_0604_),
    .A1(_0601_),
    .A2(_0603_));
 sg13g2_a21oi_1 _2179_ (.A1(_0586_),
    .A2(_0604_),
    .Y(_0605_),
    .B1(_0585_));
 sg13g2_nor2_1 _2180_ (.A(_1212_),
    .B(\ppwm_i.u_ppwm.global_counter[7] ),
    .Y(_0606_));
 sg13g2_nand2_1 _2181_ (.Y(_0607_),
    .A(_1218_),
    .B(\ppwm_i.u_ppwm.global_counter[1] ));
 sg13g2_nor2_1 _2182_ (.A(_1219_),
    .B(\ppwm_i.u_ppwm.global_counter[0] ),
    .Y(_0608_));
 sg13g2_nor2_1 _2183_ (.A(_1218_),
    .B(\ppwm_i.u_ppwm.global_counter[1] ),
    .Y(_0609_));
 sg13g2_a221oi_1 _2184_ (.B2(_0608_),
    .C1(_0609_),
    .B1(_0607_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .Y(_0610_),
    .A2(_1265_));
 sg13g2_a221oi_1 _2185_ (.B2(_1217_),
    .C1(_0610_),
    .B1(\ppwm_i.u_ppwm.global_counter[2] ),
    .A1(_1216_),
    .Y(_0611_),
    .A2(\ppwm_i.u_ppwm.global_counter[3] ));
 sg13g2_nand2_1 _2186_ (.Y(_0612_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .B(_1264_));
 sg13g2_o21ai_1 _2187_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_1215_),
    .A2(\ppwm_i.u_ppwm.global_counter[4] ));
 sg13g2_a22oi_1 _2188_ (.Y(_0614_),
    .B1(\ppwm_i.u_ppwm.global_counter[4] ),
    .B2(_1215_),
    .A2(\ppwm_i.u_ppwm.global_counter[5] ),
    .A1(_1214_));
 sg13g2_o21ai_1 _2189_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0611_),
    .A2(_0613_));
 sg13g2_a22oi_1 _2190_ (.Y(_0616_),
    .B1(_1262_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A2(_1261_),
    .A1(net502));
 sg13g2_nor2_1 _2191_ (.A(net502),
    .B(_1261_),
    .Y(_0617_));
 sg13g2_a221oi_1 _2192_ (.B2(_0616_),
    .C1(_0617_),
    .B1(_0615_),
    .A1(_1212_),
    .Y(_0618_),
    .A2(\ppwm_i.u_ppwm.global_counter[7] ));
 sg13g2_nand2_1 _2193_ (.Y(_0619_),
    .A(_1211_),
    .B(\ppwm_i.u_ppwm.global_counter[8] ));
 sg13g2_o21ai_1 _2194_ (.B1(_0619_),
    .Y(_0620_),
    .A1(_0606_),
    .A2(_0618_));
 sg13g2_a22oi_1 _2195_ (.Y(_0621_),
    .B1(_1260_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .A2(_1259_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ));
 sg13g2_a221oi_1 _2196_ (.B2(_0621_),
    .C1(_1312_),
    .B1(_0620_),
    .A1(_1210_),
    .Y(_0622_),
    .A2(\ppwm_i.u_ppwm.global_counter[9] ));
 sg13g2_o21ai_1 _2197_ (.B1(net385),
    .Y(_0623_),
    .A1(_0605_),
    .A2(_0622_));
 sg13g2_nand2b_1 _2198_ (.Y(_0624_),
    .B(net507),
    .A_N(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ));
 sg13g2_nand3_1 _2199_ (.B(_1229_),
    .C(_0624_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .Y(_0625_));
 sg13g2_nor2_1 _2200_ (.A(_1216_),
    .B(net506),
    .Y(_0626_));
 sg13g2_a22oi_1 _2201_ (.Y(_0627_),
    .B1(_1228_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(_1227_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ));
 sg13g2_a22oi_1 _2202_ (.Y(_0628_),
    .B1(_0625_),
    .B2(_0627_),
    .A2(\ppwm_i.u_ppwm.pwm_value[2] ),
    .A1(_1217_));
 sg13g2_a22oi_1 _2203_ (.Y(_0629_),
    .B1(net506),
    .B2(_1216_),
    .A2(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A1(_1215_));
 sg13g2_o21ai_1 _2204_ (.B1(_0629_),
    .Y(_0630_),
    .A1(_0626_),
    .A2(_0628_));
 sg13g2_a22oi_1 _2205_ (.Y(_0631_),
    .B1(_1225_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .A2(_1224_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ));
 sg13g2_nor2_1 _2206_ (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .B(_1223_),
    .Y(_0632_));
 sg13g2_a221oi_1 _2207_ (.B2(_0631_),
    .C1(_0632_),
    .B1(_0630_),
    .A1(_1214_),
    .Y(_0633_),
    .A2(\ppwm_i.u_ppwm.pwm_value[5] ));
 sg13g2_a221oi_1 _2208_ (.B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .C1(_0633_),
    .B1(_1223_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .Y(_0634_),
    .A2(_1222_));
 sg13g2_nand2_1 _2209_ (.Y(_0635_),
    .A(_1212_),
    .B(net503));
 sg13g2_o21ai_1 _2210_ (.B1(_0635_),
    .Y(_0636_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .A2(_1221_));
 sg13g2_a22oi_1 _2211_ (.Y(_0637_),
    .B1(_1221_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .A2(_1220_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ));
 sg13g2_o21ai_1 _2212_ (.B1(_0637_),
    .Y(_0638_),
    .A1(_0634_),
    .A2(_0636_));
 sg13g2_nand2_2 _2213_ (.Y(_0639_),
    .A(net397),
    .B(net385));
 sg13g2_a221oi_1 _2214_ (.B2(_0584_),
    .C1(_0551_),
    .B1(_0583_),
    .A1(_1210_),
    .Y(_0640_),
    .A2(\ppwm_i.u_ppwm.global_counter[19] ));
 sg13g2_nand2b_1 _2215_ (.Y(_0641_),
    .B(net402),
    .A_N(_0640_));
 sg13g2_a21oi_1 _2216_ (.A1(net399),
    .A2(_0568_),
    .Y(_0642_),
    .B1(_0551_));
 sg13g2_a21oi_1 _2217_ (.A1(_1210_),
    .A2(\ppwm_i.u_ppwm.pwm_value[9] ),
    .Y(_0643_),
    .B1(net381));
 sg13g2_and2_1 _2218_ (.A(_0638_),
    .B(_0643_),
    .X(_0644_));
 sg13g2_o21ai_1 _2219_ (.B1(_0641_),
    .Y(_0645_),
    .A1(_0642_),
    .A2(_0644_));
 sg13g2_o21ai_1 _2220_ (.B1(net396),
    .Y(_0646_),
    .A1(net401),
    .A2(net389));
 sg13g2_nand2_1 _2221_ (.Y(_0647_),
    .A(_0549_),
    .B(_0646_));
 sg13g2_a21o_1 _2222_ (.A2(_0645_),
    .A1(_0623_),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_a21oi_1 _2223_ (.A1(net350),
    .A2(_0648_),
    .Y(_0193_),
    .B1(net458));
 sg13g2_nand3_1 _2224_ (.B(net396),
    .C(_0366_),
    .A(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .Y(_0649_));
 sg13g2_o21ai_1 _2225_ (.B1(net419),
    .Y(_0650_),
    .A1(net401),
    .A2(_0649_));
 sg13g2_a21oi_1 _2226_ (.A1(_1230_),
    .A2(_0649_),
    .Y(_0194_),
    .B1(_0650_));
 sg13g2_or2_1 _2227_ (.X(_0651_),
    .B(_0365_),
    .A(net394));
 sg13g2_nor3_1 _2228_ (.A(_1325_),
    .B(net394),
    .C(_0365_),
    .Y(_0652_));
 sg13g2_nor4_2 _2229_ (.A(net396),
    .B(net395),
    .C(net390),
    .Y(_0653_),
    .D(_0651_));
 sg13g2_nor2_1 _2230_ (.A(_1218_),
    .B(net398),
    .Y(_0654_));
 sg13g2_a21oi_2 _2231_ (.B1(_0654_),
    .Y(_0655_),
    .A2(net400),
    .A1(net507));
 sg13g2_mux2_1 _2232_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .A1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .S(net398),
    .X(_0656_));
 sg13g2_nor2_1 _2233_ (.A(net384),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_a21oi_1 _2234_ (.A1(net384),
    .A2(_0655_),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_nor4_2 _2235_ (.A(net396),
    .B(net395),
    .C(net392),
    .Y(_0659_),
    .D(_0651_));
 sg13g2_nor2_1 _2236_ (.A(_1215_),
    .B(net399),
    .Y(_0660_));
 sg13g2_a21oi_1 _2237_ (.A1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A2(net399),
    .Y(_0661_),
    .B1(_0660_));
 sg13g2_mux2_1 _2238_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .A1(net505),
    .S(net399),
    .X(_0662_));
 sg13g2_nor2_1 _2239_ (.A(net384),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_nor2_1 _2240_ (.A(_1216_),
    .B(net398),
    .Y(_0664_));
 sg13g2_nor2_1 _2241_ (.A(_1226_),
    .B(net403),
    .Y(_0665_));
 sg13g2_nor2_1 _2242_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nor3_1 _2243_ (.A(net388),
    .B(_0664_),
    .C(_0665_),
    .Y(_0667_));
 sg13g2_nor2_1 _2244_ (.A(_0663_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_a22oi_1 _2245_ (.Y(_0669_),
    .B1(_0659_),
    .B2(_0668_),
    .A2(_0658_),
    .A1(net379));
 sg13g2_mux2_1 _2246_ (.A0(\ppwm_i.u_ppwm.global_counter[10] ),
    .A1(\ppwm_i.u_ppwm.global_counter[0] ),
    .S(net398),
    .X(_0670_));
 sg13g2_and3_2 _2247_ (.X(_0671_),
    .A(net395),
    .B(net394),
    .C(_0365_));
 sg13g2_nand2_2 _2248_ (.Y(_0672_),
    .A(net394),
    .B(_0547_));
 sg13g2_nor2_2 _2249_ (.A(_0551_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_nand2_1 _2250_ (.Y(_0674_),
    .A(_0651_),
    .B(_0672_));
 sg13g2_nor2_1 _2251_ (.A(_1311_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_and2_1 _2252_ (.A(_0551_),
    .B(net380),
    .X(_0676_));
 sg13g2_a221oi_1 _2253_ (.B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .C1(_0675_),
    .B1(net375),
    .A1(_0670_),
    .Y(_0677_),
    .A2(net376));
 sg13g2_nand2_1 _2254_ (.Y(_0678_),
    .A(_1229_),
    .B(_1311_));
 sg13g2_o21ai_1 _2255_ (.B1(net385),
    .Y(_0679_),
    .A1(net401),
    .A2(net397));
 sg13g2_a21oi_1 _2256_ (.A1(net395),
    .A2(_1338_),
    .Y(_0680_),
    .B1(_0365_));
 sg13g2_a22oi_1 _2257_ (.Y(_0681_),
    .B1(_0680_),
    .B2(net398),
    .A2(_0679_),
    .A1(net380));
 sg13g2_nand2b_1 _2258_ (.Y(_0682_),
    .B(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .A_N(_0681_));
 sg13g2_a21oi_2 _2259_ (.B1(_0682_),
    .Y(_0683_),
    .A2(net375),
    .A1(_0585_));
 sg13g2_nor2b_2 _2260_ (.A(_0651_),
    .B_N(net395),
    .Y(_0684_));
 sg13g2_nand2b_2 _2261_ (.Y(_0685_),
    .B(net395),
    .A_N(_0651_));
 sg13g2_a221oi_1 _2262_ (.B2(_1309_),
    .C1(_1229_),
    .B1(_1306_),
    .A1(net508),
    .Y(_0686_),
    .A2(_1302_));
 sg13g2_nand2_1 _2263_ (.Y(_0687_),
    .A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .B(net396));
 sg13g2_nor2_1 _2264_ (.A(net800),
    .B(net371),
    .Y(_0688_));
 sg13g2_nand3_1 _2265_ (.B(net377),
    .C(_0687_),
    .A(_0678_),
    .Y(_0689_));
 sg13g2_and4_1 _2266_ (.A(_0669_),
    .B(_0677_),
    .C(net371),
    .D(_0689_),
    .X(_0690_));
 sg13g2_nor3_1 _2267_ (.A(net457),
    .B(_0688_),
    .C(_0690_),
    .Y(_0195_));
 sg13g2_and2_1 _2268_ (.A(net396),
    .B(_0652_),
    .X(_0691_));
 sg13g2_nand2_2 _2269_ (.Y(_0692_),
    .A(net396),
    .B(_0652_));
 sg13g2_nand2_1 _2270_ (.Y(_0693_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .B(net401));
 sg13g2_o21ai_1 _2271_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_1229_),
    .A2(net401));
 sg13g2_inv_1 _2272_ (.Y(_0695_),
    .A(_0694_));
 sg13g2_nor3_1 _2273_ (.A(_0351_),
    .B(_0692_),
    .C(_0695_),
    .Y(_0696_));
 sg13g2_mux2_1 _2274_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ),
    .S(net399),
    .X(_0697_));
 sg13g2_mux2_1 _2275_ (.A0(_0662_),
    .A1(_0697_),
    .S(net387),
    .X(_0698_));
 sg13g2_nor2_1 _2276_ (.A(net386),
    .B(_0656_),
    .Y(_0699_));
 sg13g2_a21oi_1 _2277_ (.A1(net386),
    .A2(_0666_),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_a221oi_1 _2278_ (.B2(net379),
    .C1(_0696_),
    .B1(_0700_),
    .A1(_0659_),
    .Y(_0701_),
    .A2(_0698_));
 sg13g2_o21ai_1 _2279_ (.B1(_1228_),
    .Y(_0702_),
    .A1(_0341_),
    .A2(_0347_));
 sg13g2_nor3_1 _2280_ (.A(_1228_),
    .B(_0341_),
    .C(_0347_),
    .Y(_0703_));
 sg13g2_xnor2_1 _2281_ (.Y(_0704_),
    .A(net507),
    .B(net386));
 sg13g2_a21oi_1 _2282_ (.A1(_0687_),
    .A2(_0704_),
    .Y(_0705_),
    .B1(_0685_));
 sg13g2_o21ai_1 _2283_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0687_),
    .A2(_0704_));
 sg13g2_nor2_1 _2284_ (.A(net385),
    .B(_0674_),
    .Y(_0707_));
 sg13g2_nand2_1 _2285_ (.Y(_0708_),
    .A(\ppwm_i.u_ppwm.global_counter[1] ),
    .B(net398));
 sg13g2_o21ai_1 _2286_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_1258_),
    .A2(net398));
 sg13g2_a221oi_1 _2287_ (.B2(net376),
    .C1(_0707_),
    .B1(_0709_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .Y(_0710_),
    .A2(net375));
 sg13g2_nand4_1 _2288_ (.B(_0701_),
    .C(_0706_),
    .A(net371),
    .Y(_0711_),
    .D(_0710_));
 sg13g2_o21ai_1 _2289_ (.B1(net424),
    .Y(_0712_),
    .A1(net507),
    .A2(net371));
 sg13g2_nor2b_1 _2290_ (.A(_0712_),
    .B_N(_0711_),
    .Y(_0196_));
 sg13g2_a21o_2 _2291_ (.A2(_0702_),
    .A1(_0686_),
    .B1(_0703_),
    .X(_0713_));
 sg13g2_or3_1 _2292_ (.A(\ppwm_i.u_ppwm.pwm_value[2] ),
    .B(net407),
    .C(net405),
    .X(_0714_));
 sg13g2_nor2_1 _2293_ (.A(_1227_),
    .B(net393),
    .Y(_0715_));
 sg13g2_o21ai_1 _2294_ (.B1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .Y(_0716_),
    .A1(net407),
    .A2(net405));
 sg13g2_and2_1 _2295_ (.A(_0714_),
    .B(_0716_),
    .X(_0717_));
 sg13g2_xnor2_1 _2296_ (.Y(_0718_),
    .A(_0713_),
    .B(_0717_));
 sg13g2_or2_1 _2297_ (.X(_0719_),
    .B(_0718_),
    .A(_0685_));
 sg13g2_nand2_1 _2298_ (.Y(_0720_),
    .A(net392),
    .B(_0691_));
 sg13g2_a221oi_1 _2299_ (.B2(net386),
    .C1(_0720_),
    .B1(_0695_),
    .A1(_0350_),
    .Y(_0721_),
    .A2(_0655_));
 sg13g2_mux2_1 _2300_ (.A0(net502),
    .A1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .S(net399),
    .X(_0722_));
 sg13g2_inv_1 _2301_ (.Y(_0723_),
    .A(_0722_));
 sg13g2_nor2_1 _2302_ (.A(net387),
    .B(_0697_),
    .Y(_0724_));
 sg13g2_a21oi_1 _2303_ (.A1(net387),
    .A2(_0723_),
    .Y(_0725_),
    .B1(_0724_));
 sg13g2_a221oi_1 _2304_ (.B2(_0659_),
    .C1(_0721_),
    .B1(_0725_),
    .A1(net379),
    .Y(_0726_),
    .A2(_0668_));
 sg13g2_nor2_1 _2305_ (.A(net393),
    .B(_0674_),
    .Y(_0727_));
 sg13g2_nand2_1 _2306_ (.Y(_0728_),
    .A(\ppwm_i.u_ppwm.global_counter[12] ),
    .B(net401));
 sg13g2_o21ai_1 _2307_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_1265_),
    .A2(_1295_));
 sg13g2_a221oi_1 _2308_ (.B2(net376),
    .C1(_0727_),
    .B1(_0729_),
    .A1(net820),
    .Y(_0730_),
    .A2(net375));
 sg13g2_nand4_1 _2309_ (.B(_0719_),
    .C(_0726_),
    .A(net373),
    .Y(_0731_),
    .D(_0730_));
 sg13g2_o21ai_1 _2310_ (.B1(net435),
    .Y(_0732_),
    .A1(net794),
    .A2(net373));
 sg13g2_nor2b_1 _2311_ (.A(_0732_),
    .B_N(_0731_),
    .Y(_0197_));
 sg13g2_o21ai_1 _2312_ (.B1(net506),
    .Y(_0733_),
    .A1(net408),
    .A2(net405));
 sg13g2_or3_1 _2313_ (.A(net506),
    .B(net408),
    .C(net405),
    .X(_0734_));
 sg13g2_nand2_1 _2314_ (.Y(_0735_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_a21oi_1 _2315_ (.A1(_0713_),
    .A2(_0717_),
    .Y(_0736_),
    .B1(_0715_));
 sg13g2_o21ai_1 _2316_ (.B1(net378),
    .Y(_0737_),
    .A1(_0735_),
    .A2(_0736_));
 sg13g2_a21o_1 _2317_ (.A2(_0736_),
    .A1(_0735_),
    .B1(_0737_),
    .X(_0738_));
 sg13g2_nor2_2 _2318_ (.A(net392),
    .B(net384),
    .Y(_0739_));
 sg13g2_nand2_1 _2319_ (.Y(_0740_),
    .A(net390),
    .B(net386));
 sg13g2_o21ai_1 _2320_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0351_),
    .A2(_0656_));
 sg13g2_a221oi_1 _2321_ (.B2(net390),
    .C1(_0741_),
    .B1(_0695_),
    .A1(net386),
    .Y(_0742_),
    .A2(_0655_));
 sg13g2_mux2_1 _2322_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .A1(\ppwm_i.u_ppwm.pwm_value[7] ),
    .S(net400),
    .X(_0743_));
 sg13g2_inv_2 _2323_ (.Y(_0744_),
    .A(_0743_));
 sg13g2_nor2_1 _2324_ (.A(net387),
    .B(_0722_),
    .Y(_0745_));
 sg13g2_a21oi_1 _2325_ (.A1(net387),
    .A2(_0744_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_and2_1 _2326_ (.A(_0659_),
    .B(_0746_),
    .X(_0747_));
 sg13g2_a221oi_1 _2327_ (.B2(_0691_),
    .C1(_0747_),
    .B1(_0742_),
    .A1(net379),
    .Y(_0748_),
    .A2(_0698_));
 sg13g2_nand2_1 _2328_ (.Y(_0749_),
    .A(\ppwm_i.u_ppwm.global_counter[13] ),
    .B(net403));
 sg13g2_o21ai_1 _2329_ (.B1(_0749_),
    .Y(_0750_),
    .A1(_1264_),
    .A2(net403));
 sg13g2_a22oi_1 _2330_ (.Y(_0751_),
    .B1(_0750_),
    .B2(net376),
    .A2(net375),
    .A1(net816));
 sg13g2_nand4_1 _2331_ (.B(_0738_),
    .C(_0748_),
    .A(net373),
    .Y(_0752_),
    .D(_0751_));
 sg13g2_o21ai_1 _2332_ (.B1(net435),
    .Y(_0753_),
    .A1(net506),
    .A2(net373));
 sg13g2_nor2b_1 _2333_ (.A(_0753_),
    .B_N(_0752_),
    .Y(_0198_));
 sg13g2_nor2_1 _2334_ (.A(_1225_),
    .B(net391),
    .Y(_0754_));
 sg13g2_xnor2_1 _2335_ (.Y(_0755_),
    .A(net505),
    .B(net391));
 sg13g2_and4_1 _2336_ (.A(_0714_),
    .B(_0716_),
    .C(_0733_),
    .D(_0734_),
    .X(_0756_));
 sg13g2_nand2_1 _2337_ (.Y(_0757_),
    .A(_0716_),
    .B(_0733_));
 sg13g2_a21o_2 _2338_ (.A2(_0756_),
    .A1(_0713_),
    .B1(_0757_),
    .X(_0758_));
 sg13g2_o21ai_1 _2339_ (.B1(net377),
    .Y(_0759_),
    .A1(_0755_),
    .A2(_0758_));
 sg13g2_a21oi_1 _2340_ (.A1(_0755_),
    .A2(_0758_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_o21ai_1 _2341_ (.B1(_0691_),
    .Y(_0761_),
    .A1(_0694_),
    .A2(_0740_));
 sg13g2_nand2_1 _2342_ (.Y(_0762_),
    .A(_0350_),
    .B(_0666_));
 sg13g2_nor2_2 _2343_ (.A(_0350_),
    .B(_0739_),
    .Y(_0763_));
 sg13g2_nand2_2 _2344_ (.Y(_0764_),
    .A(_0351_),
    .B(_0740_));
 sg13g2_o21ai_1 _2345_ (.B1(_0762_),
    .Y(_0765_),
    .A1(_0658_),
    .A2(_0764_));
 sg13g2_mux2_1 _2346_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .S(net399),
    .X(_0766_));
 sg13g2_nor2_1 _2347_ (.A(net384),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_a21oi_1 _2348_ (.A1(net384),
    .A2(_0744_),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_a22oi_1 _2349_ (.Y(_0769_),
    .B1(_0768_),
    .B2(_0659_),
    .A2(_0725_),
    .A1(net379));
 sg13g2_o21ai_1 _2350_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_0761_),
    .A2(_0765_));
 sg13g2_nand2_1 _2351_ (.Y(_0771_),
    .A(\ppwm_i.u_ppwm.global_counter[14] ),
    .B(net403));
 sg13g2_o21ai_1 _2352_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_1263_),
    .A2(net403));
 sg13g2_a22oi_1 _2353_ (.Y(_0773_),
    .B1(_0772_),
    .B2(net376),
    .A2(net375),
    .A1(net818));
 sg13g2_nand2_1 _2354_ (.Y(_0774_),
    .A(net373),
    .B(_0773_));
 sg13g2_nor3_1 _2355_ (.A(_0760_),
    .B(_0770_),
    .C(_0774_),
    .Y(_0775_));
 sg13g2_o21ai_1 _2356_ (.B1(net421),
    .Y(_0776_),
    .A1(net505),
    .A2(net371));
 sg13g2_nor2_1 _2357_ (.A(_0775_),
    .B(_0776_),
    .Y(_0199_));
 sg13g2_a21oi_1 _2358_ (.A1(_0755_),
    .A2(_0758_),
    .Y(_0777_),
    .B1(_0754_));
 sg13g2_xnor2_1 _2359_ (.Y(_0778_),
    .A(\ppwm_i.u_ppwm.pwm_value[5] ),
    .B(net391));
 sg13g2_nand2b_1 _2360_ (.Y(_0779_),
    .B(_0777_),
    .A_N(_0778_));
 sg13g2_nand2b_1 _2361_ (.Y(_0780_),
    .B(_0778_),
    .A_N(_0777_));
 sg13g2_nand3_1 _2362_ (.B(_0779_),
    .C(_0780_),
    .A(net377),
    .Y(_0781_));
 sg13g2_nand2b_1 _2363_ (.Y(_0782_),
    .B(_0763_),
    .A_N(_0700_));
 sg13g2_a221oi_1 _2364_ (.B2(_0655_),
    .C1(_0692_),
    .B1(_0739_),
    .A1(_0350_),
    .Y(_0783_),
    .A2(_0661_));
 sg13g2_nand2_1 _2365_ (.Y(_0784_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .B(net404));
 sg13g2_o21ai_1 _2366_ (.B1(_0784_),
    .Y(_0785_),
    .A1(_1220_),
    .A2(net404));
 sg13g2_nor2_1 _2367_ (.A(net386),
    .B(_0766_),
    .Y(_0786_));
 sg13g2_mux2_1 _2368_ (.A0(_0766_),
    .A1(_0785_),
    .S(net386),
    .X(_0787_));
 sg13g2_and2_1 _2369_ (.A(_0659_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_a221oi_1 _2370_ (.B2(_0783_),
    .C1(_0788_),
    .B1(_0782_),
    .A1(net379),
    .Y(_0789_),
    .A2(_0746_));
 sg13g2_nand2_1 _2371_ (.Y(_0790_),
    .A(\ppwm_i.u_ppwm.global_counter[15] ),
    .B(net402));
 sg13g2_o21ai_1 _2372_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_1262_),
    .A2(net402));
 sg13g2_a22oi_1 _2373_ (.Y(_0792_),
    .B1(_0791_),
    .B2(net376),
    .A2(net375),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ));
 sg13g2_nand4_1 _2374_ (.B(_0781_),
    .C(_0789_),
    .A(net371),
    .Y(_0793_),
    .D(_0792_));
 sg13g2_o21ai_1 _2375_ (.B1(net422),
    .Y(_0794_),
    .A1(net828),
    .A2(net371));
 sg13g2_nor2b_1 _2376_ (.A(_0794_),
    .B_N(_0793_),
    .Y(_0200_));
 sg13g2_nor2_1 _2377_ (.A(_1223_),
    .B(net391),
    .Y(_0795_));
 sg13g2_xnor2_1 _2378_ (.Y(_0796_),
    .A(net504),
    .B(net391));
 sg13g2_o21ai_1 _2379_ (.B1(net390),
    .Y(_0797_),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ),
    .A2(net505));
 sg13g2_a21oi_1 _2380_ (.A1(_1224_),
    .A2(_1225_),
    .Y(_0798_),
    .B1(net392));
 sg13g2_and2_1 _2381_ (.A(_0755_),
    .B(_0778_),
    .X(_0799_));
 sg13g2_a21o_1 _2382_ (.A2(_0799_),
    .A1(_0758_),
    .B1(_0798_),
    .X(_0800_));
 sg13g2_o21ai_1 _2383_ (.B1(net377),
    .Y(_0801_),
    .A1(_0796_),
    .A2(_0800_));
 sg13g2_a21oi_1 _2384_ (.A1(_0796_),
    .A2(_0800_),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_o21ai_1 _2385_ (.B1(_0764_),
    .Y(_0803_),
    .A1(_0657_),
    .A2(_0724_));
 sg13g2_o21ai_1 _2386_ (.B1(_0763_),
    .Y(_0804_),
    .A1(_0663_),
    .A2(_0667_));
 sg13g2_nand3_1 _2387_ (.B(_0803_),
    .C(_0804_),
    .A(_0691_),
    .Y(_0805_));
 sg13g2_and2_1 _2388_ (.A(net384),
    .B(_0785_),
    .X(_0806_));
 sg13g2_a22oi_1 _2389_ (.Y(_0807_),
    .B1(_0806_),
    .B2(_0659_),
    .A2(_0768_),
    .A1(net379));
 sg13g2_nand2_1 _2390_ (.Y(_0808_),
    .A(\ppwm_i.u_ppwm.global_counter[16] ),
    .B(net403));
 sg13g2_o21ai_1 _2391_ (.B1(_0808_),
    .Y(_0809_),
    .A1(_1261_),
    .A2(net402));
 sg13g2_a22oi_1 _2392_ (.Y(_0810_),
    .B1(_0809_),
    .B2(net376),
    .A2(net375),
    .A1(net502));
 sg13g2_nand4_1 _2393_ (.B(_0805_),
    .C(_0807_),
    .A(_0683_),
    .Y(_0811_),
    .D(_0810_));
 sg13g2_nor2_1 _2394_ (.A(net504),
    .B(net371),
    .Y(_0812_));
 sg13g2_o21ai_1 _2395_ (.B1(net423),
    .Y(_0813_),
    .A1(_0802_),
    .A2(_0811_));
 sg13g2_nor2_1 _2396_ (.A(_0812_),
    .B(_0813_),
    .Y(_0201_));
 sg13g2_a21oi_1 _2397_ (.A1(_0796_),
    .A2(_0800_),
    .Y(_0814_),
    .B1(_0795_));
 sg13g2_xnor2_1 _2398_ (.Y(_0815_),
    .A(net503),
    .B(net391));
 sg13g2_inv_1 _2399_ (.Y(_0816_),
    .A(_0815_));
 sg13g2_nand2b_1 _2400_ (.Y(_0817_),
    .B(_0815_),
    .A_N(_0814_));
 sg13g2_a21oi_1 _2401_ (.A1(_0814_),
    .A2(_0816_),
    .Y(_0818_),
    .B1(_0685_));
 sg13g2_nand2b_1 _2402_ (.Y(_0819_),
    .B(_0763_),
    .A_N(_0698_));
 sg13g2_a221oi_1 _2403_ (.B2(_0666_),
    .C1(_0692_),
    .B1(_0739_),
    .A1(_0350_),
    .Y(_0820_),
    .A2(_0723_));
 sg13g2_a22oi_1 _2404_ (.Y(_0821_),
    .B1(_0819_),
    .B2(_0820_),
    .A2(_0787_),
    .A1(net379));
 sg13g2_mux2_1 _2405_ (.A0(\ppwm_i.u_ppwm.global_counter[17] ),
    .A1(\ppwm_i.u_ppwm.global_counter[7] ),
    .S(net399),
    .X(_0822_));
 sg13g2_a22oi_1 _2406_ (.Y(_0823_),
    .B1(_0822_),
    .B2(net376),
    .A2(_0676_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ));
 sg13g2_nand3_1 _2407_ (.B(_0821_),
    .C(_0823_),
    .A(_0683_),
    .Y(_0824_));
 sg13g2_a21oi_1 _2408_ (.A1(_0817_),
    .A2(_0818_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_o21ai_1 _2409_ (.B1(net423),
    .Y(_0826_),
    .A1(net503),
    .A2(net372));
 sg13g2_nor2_1 _2410_ (.A(_0825_),
    .B(_0826_),
    .Y(_0202_));
 sg13g2_and4_1 _2411_ (.A(_0755_),
    .B(_0778_),
    .C(_0796_),
    .D(_0815_),
    .X(_0827_));
 sg13g2_o21ai_1 _2412_ (.B1(_0336_),
    .Y(_0828_),
    .A1(net503),
    .A2(net504));
 sg13g2_nand2_1 _2413_ (.Y(_0829_),
    .A(_0797_),
    .B(_0828_));
 sg13g2_a21oi_1 _2414_ (.A1(_0758_),
    .A2(_0827_),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_nand2_1 _2415_ (.Y(_0831_),
    .A(net814),
    .B(_0336_));
 sg13g2_xnor2_1 _2416_ (.Y(_0832_),
    .A(\ppwm_i.u_ppwm.pwm_value[8] ),
    .B(net391));
 sg13g2_nand2b_1 _2417_ (.Y(_0833_),
    .B(_0830_),
    .A_N(_0832_));
 sg13g2_nand2b_1 _2418_ (.Y(_0834_),
    .B(_0832_),
    .A_N(_0830_));
 sg13g2_nand3_1 _2419_ (.B(_0833_),
    .C(_0834_),
    .A(net377),
    .Y(_0835_));
 sg13g2_nand2b_1 _2420_ (.Y(_0836_),
    .B(_0763_),
    .A_N(_0725_));
 sg13g2_a221oi_1 _2421_ (.B2(_0350_),
    .C1(_0692_),
    .B1(_0744_),
    .A1(_0661_),
    .Y(_0837_),
    .A2(_0739_));
 sg13g2_a22oi_1 _2422_ (.Y(_0838_),
    .B1(_0836_),
    .B2(_0837_),
    .A2(_0806_),
    .A1(_0653_));
 sg13g2_nand2_1 _2423_ (.Y(_0839_),
    .A(\ppwm_i.u_ppwm.global_counter[18] ),
    .B(net402));
 sg13g2_o21ai_1 _2424_ (.B1(_0839_),
    .Y(_0840_),
    .A1(_1260_),
    .A2(net402));
 sg13g2_a22oi_1 _2425_ (.Y(_0841_),
    .B1(_0840_),
    .B2(_0673_),
    .A2(_0676_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ));
 sg13g2_nand4_1 _2426_ (.B(_0835_),
    .C(_0838_),
    .A(net372),
    .Y(_0842_),
    .D(_0841_));
 sg13g2_o21ai_1 _2427_ (.B1(net424),
    .Y(_0843_),
    .A1(net814),
    .A2(net372));
 sg13g2_nor2b_1 _2428_ (.A(_0843_),
    .B_N(_0842_),
    .Y(_0203_));
 sg13g2_xnor2_1 _2429_ (.Y(_0844_),
    .A(_1220_),
    .B(net391));
 sg13g2_nand3_1 _2430_ (.B(_0834_),
    .C(_0844_),
    .A(_0831_),
    .Y(_0845_));
 sg13g2_a21o_1 _2431_ (.A2(_0834_),
    .A1(_0831_),
    .B1(_0844_),
    .X(_0846_));
 sg13g2_nand3_1 _2432_ (.B(_0845_),
    .C(_0846_),
    .A(net377),
    .Y(_0847_));
 sg13g2_o21ai_1 _2433_ (.B1(_0764_),
    .Y(_0848_),
    .A1(net384),
    .A2(_0697_));
 sg13g2_nand2_1 _2434_ (.Y(_0849_),
    .A(_0746_),
    .B(_0763_));
 sg13g2_o21ai_1 _2435_ (.B1(_0849_),
    .Y(_0850_),
    .A1(_0786_),
    .A2(_0848_));
 sg13g2_nand2_1 _2436_ (.Y(_0851_),
    .A(\ppwm_i.u_ppwm.global_counter[19] ),
    .B(net402));
 sg13g2_o21ai_1 _2437_ (.B1(_0851_),
    .Y(_0852_),
    .A1(_1259_),
    .A2(net402));
 sg13g2_a22oi_1 _2438_ (.Y(_0853_),
    .B1(_0852_),
    .B2(_0673_),
    .A2(_0676_),
    .A1(net805));
 sg13g2_nand2_1 _2439_ (.Y(_0854_),
    .A(net373),
    .B(_0853_));
 sg13g2_a21oi_1 _2440_ (.A1(_0691_),
    .A2(_0850_),
    .Y(_0855_),
    .B1(_0854_));
 sg13g2_o21ai_1 _2441_ (.B1(net423),
    .Y(_0856_),
    .A1(net793),
    .A2(net372));
 sg13g2_a21oi_1 _2442_ (.A1(_0847_),
    .A2(_0855_),
    .Y(_0204_),
    .B1(_0856_));
 sg13g2_nor2_1 _2443_ (.A(net383),
    .B(_0670_),
    .Y(_0857_));
 sg13g2_a21oi_1 _2444_ (.A1(_1229_),
    .A2(net383),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_or2_1 _2445_ (.X(_0859_),
    .B(_0680_),
    .A(net380));
 sg13g2_and3_2 _2446_ (.X(_0860_),
    .A(net768),
    .B(_0681_),
    .C(_0859_));
 sg13g2_inv_2 _2447_ (.Y(_0861_),
    .A(net374));
 sg13g2_a221oi_1 _2448_ (.B2(_1309_),
    .C1(_1219_),
    .B1(_1306_),
    .A1(net508),
    .Y(_0862_),
    .A2(_1302_));
 sg13g2_nand2_1 _2449_ (.Y(_0863_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .B(net397));
 sg13g2_xnor2_1 _2450_ (.Y(_0864_),
    .A(_1219_),
    .B(net397));
 sg13g2_a221oi_1 _2451_ (.B2(net377),
    .C1(_0675_),
    .B1(_0864_),
    .A1(net380),
    .Y(_0865_),
    .A2(_0858_));
 sg13g2_and2_1 _2452_ (.A(net374),
    .B(_0865_),
    .X(_0866_));
 sg13g2_a221oi_1 _2453_ (.B2(_0669_),
    .C1(net458),
    .B1(_0866_),
    .A1(_1219_),
    .Y(_0205_),
    .A2(net370));
 sg13g2_o21ai_1 _2454_ (.B1(_1218_),
    .Y(_0867_),
    .A1(_0341_),
    .A2(_0347_));
 sg13g2_nor3_1 _2455_ (.A(_1218_),
    .B(_0341_),
    .C(_0347_),
    .Y(_0868_));
 sg13g2_xnor2_1 _2456_ (.Y(_0869_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .B(net389));
 sg13g2_o21ai_1 _2457_ (.B1(net377),
    .Y(_0870_),
    .A1(_0863_),
    .A2(_0869_));
 sg13g2_a21oi_1 _2458_ (.A1(_0863_),
    .A2(_0869_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_o21ai_1 _2459_ (.B1(net380),
    .Y(_0872_),
    .A1(net383),
    .A2(_0709_));
 sg13g2_a21oi_1 _2460_ (.A1(_1228_),
    .A2(net383),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_nor4_1 _2461_ (.A(_0707_),
    .B(net370),
    .C(_0871_),
    .D(_0873_),
    .Y(_0874_));
 sg13g2_a221oi_1 _2462_ (.B2(_0701_),
    .C1(net458),
    .B1(_0874_),
    .A1(_1218_),
    .Y(_0206_),
    .A2(net370));
 sg13g2_a21o_2 _2463_ (.A2(_0867_),
    .A1(_0862_),
    .B1(_0868_),
    .X(_0875_));
 sg13g2_or3_1 _2464_ (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .B(net407),
    .C(net405),
    .X(_0876_));
 sg13g2_o21ai_1 _2465_ (.B1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .Y(_0877_),
    .A1(net407),
    .A2(net405));
 sg13g2_and2_1 _2466_ (.A(_0876_),
    .B(_0877_),
    .X(_0878_));
 sg13g2_nand2_1 _2467_ (.Y(_0879_),
    .A(_0875_),
    .B(_0878_));
 sg13g2_or2_1 _2468_ (.X(_0880_),
    .B(_0878_),
    .A(_0875_));
 sg13g2_nand3_1 _2469_ (.B(_0879_),
    .C(_0880_),
    .A(net378),
    .Y(_0881_));
 sg13g2_nor2_1 _2470_ (.A(net383),
    .B(_0729_),
    .Y(_0882_));
 sg13g2_a21oi_1 _2471_ (.A1(_1227_),
    .A2(net383),
    .Y(_0883_),
    .B1(_0882_));
 sg13g2_a21oi_1 _2472_ (.A1(net380),
    .A2(_0883_),
    .Y(_0884_),
    .B1(_0727_));
 sg13g2_and3_1 _2473_ (.X(_0885_),
    .A(_0726_),
    .B(net374),
    .C(_0884_));
 sg13g2_a221oi_1 _2474_ (.B2(_0885_),
    .C1(net458),
    .B1(_0881_),
    .A1(_1217_),
    .Y(_0207_),
    .A2(net370));
 sg13g2_o21ai_1 _2475_ (.B1(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .Y(_0886_),
    .A1(net407),
    .A2(net405));
 sg13g2_or3_1 _2476_ (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .B(net407),
    .C(net405),
    .X(_0887_));
 sg13g2_nand2_1 _2477_ (.Y(_0888_),
    .A(_0886_),
    .B(_0887_));
 sg13g2_a21o_1 _2478_ (.A2(_0879_),
    .A1(_0877_),
    .B1(_0888_),
    .X(_0889_));
 sg13g2_nand3_1 _2479_ (.B(_0879_),
    .C(_0888_),
    .A(_0877_),
    .Y(_0890_));
 sg13g2_nand3_1 _2480_ (.B(_0889_),
    .C(_0890_),
    .A(net378),
    .Y(_0891_));
 sg13g2_a21oi_1 _2481_ (.A1(_1226_),
    .A2(net383),
    .Y(_0892_),
    .B1(_0672_));
 sg13g2_o21ai_1 _2482_ (.B1(_0892_),
    .Y(_0893_),
    .A1(net383),
    .A2(_0750_));
 sg13g2_and3_1 _2483_ (.X(_0894_),
    .A(_0748_),
    .B(net374),
    .C(_0893_));
 sg13g2_a221oi_1 _2484_ (.B2(_0894_),
    .C1(net458),
    .B1(_0891_),
    .A1(_1216_),
    .Y(_0208_),
    .A2(net370));
 sg13g2_nor2_1 _2485_ (.A(_1215_),
    .B(net393),
    .Y(_0895_));
 sg13g2_xnor2_1 _2486_ (.Y(_0896_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .B(net393));
 sg13g2_and4_1 _2487_ (.A(_0876_),
    .B(_0877_),
    .C(_0886_),
    .D(_0887_),
    .X(_0897_));
 sg13g2_nand2_1 _2488_ (.Y(_0898_),
    .A(_0877_),
    .B(_0886_));
 sg13g2_a21oi_1 _2489_ (.A1(_0875_),
    .A2(_0897_),
    .Y(_0899_),
    .B1(_0898_));
 sg13g2_a21o_2 _2490_ (.A2(_0897_),
    .A1(_0875_),
    .B1(_0898_),
    .X(_0900_));
 sg13g2_and2_1 _2491_ (.A(_0896_),
    .B(_0900_),
    .X(_0901_));
 sg13g2_o21ai_1 _2492_ (.B1(net378),
    .Y(_0902_),
    .A1(_0896_),
    .A2(_0900_));
 sg13g2_o21ai_1 _2493_ (.B1(net380),
    .Y(_0903_),
    .A1(net382),
    .A2(_0772_));
 sg13g2_a21oi_1 _2494_ (.A1(_1225_),
    .A2(net382),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_o21ai_1 _2495_ (.B1(net374),
    .Y(_0905_),
    .A1(_0901_),
    .A2(_0902_));
 sg13g2_nor3_1 _2496_ (.A(_0770_),
    .B(_0904_),
    .C(_0905_),
    .Y(_0906_));
 sg13g2_o21ai_1 _2497_ (.B1(net423),
    .Y(_0907_),
    .A1(net818),
    .A2(net374));
 sg13g2_nor2_1 _2498_ (.A(_0906_),
    .B(_0907_),
    .Y(_0209_));
 sg13g2_xnor2_1 _2499_ (.Y(_0908_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .B(net393));
 sg13g2_o21ai_1 _2500_ (.B1(_0908_),
    .Y(_0909_),
    .A1(_0895_),
    .A2(_0901_));
 sg13g2_or3_1 _2501_ (.A(_0895_),
    .B(_0901_),
    .C(_0908_),
    .X(_0910_));
 sg13g2_nand3_1 _2502_ (.B(_0909_),
    .C(_0910_),
    .A(net378),
    .Y(_0911_));
 sg13g2_a21oi_1 _2503_ (.A1(_1224_),
    .A2(net382),
    .Y(_0912_),
    .B1(_0672_));
 sg13g2_o21ai_1 _2504_ (.B1(_0912_),
    .Y(_0913_),
    .A1(net382),
    .A2(_0791_));
 sg13g2_and3_1 _2505_ (.X(_0914_),
    .A(_0789_),
    .B(net374),
    .C(_0913_));
 sg13g2_a221oi_1 _2506_ (.B2(_0914_),
    .C1(net459),
    .B1(_0911_),
    .A1(_1214_),
    .Y(_0210_),
    .A2(net370));
 sg13g2_nor2_1 _2507_ (.A(_1213_),
    .B(net393),
    .Y(_0915_));
 sg13g2_xnor2_1 _2508_ (.Y(_0916_),
    .A(net502),
    .B(net393));
 sg13g2_o21ai_1 _2509_ (.B1(net390),
    .Y(_0917_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A2(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ));
 sg13g2_nand2_1 _2510_ (.Y(_0918_),
    .A(_0896_),
    .B(_0908_));
 sg13g2_o21ai_1 _2511_ (.B1(_0917_),
    .Y(_0919_),
    .A1(_0899_),
    .A2(_0918_));
 sg13g2_o21ai_1 _2512_ (.B1(net378),
    .Y(_0920_),
    .A1(_0916_),
    .A2(_0919_));
 sg13g2_a21oi_1 _2513_ (.A1(_0916_),
    .A2(_0919_),
    .Y(_0921_),
    .B1(_0920_));
 sg13g2_a21oi_1 _2514_ (.A1(_1223_),
    .A2(net381),
    .Y(_0922_),
    .B1(_0672_));
 sg13g2_o21ai_1 _2515_ (.B1(_0922_),
    .Y(_0923_),
    .A1(net381),
    .A2(_0809_));
 sg13g2_nand4_1 _2516_ (.B(_0807_),
    .C(net374),
    .A(_0805_),
    .Y(_0924_),
    .D(_0923_));
 sg13g2_o21ai_1 _2517_ (.B1(net436),
    .Y(_0925_),
    .A1(_0921_),
    .A2(_0924_));
 sg13g2_a21oi_1 _2518_ (.A1(_1213_),
    .A2(net370),
    .Y(_0211_),
    .B1(_0925_));
 sg13g2_a21oi_1 _2519_ (.A1(_0916_),
    .A2(_0919_),
    .Y(_0926_),
    .B1(_0915_));
 sg13g2_xnor2_1 _2520_ (.Y(_0927_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .B(net393));
 sg13g2_inv_1 _2521_ (.Y(_0928_),
    .A(_0927_));
 sg13g2_nand2b_1 _2522_ (.Y(_0929_),
    .B(_0927_),
    .A_N(_0926_));
 sg13g2_a21oi_1 _2523_ (.A1(_0926_),
    .A2(_0928_),
    .Y(_0930_),
    .B1(_0685_));
 sg13g2_nor2_1 _2524_ (.A(net381),
    .B(_0822_),
    .Y(_0931_));
 sg13g2_a21oi_1 _2525_ (.A1(_1222_),
    .A2(net382),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_nand2_1 _2526_ (.Y(_0933_),
    .A(_0821_),
    .B(_0860_));
 sg13g2_a221oi_1 _2527_ (.B2(net380),
    .C1(_0933_),
    .B1(_0932_),
    .A1(_0929_),
    .Y(_0934_),
    .A2(_0930_));
 sg13g2_o21ai_1 _2528_ (.B1(net423),
    .Y(_0935_),
    .A1(net817),
    .A2(_0860_));
 sg13g2_nor2_1 _2529_ (.A(_0934_),
    .B(_0935_),
    .Y(_0212_));
 sg13g2_and4_1 _2530_ (.A(_0896_),
    .B(_0908_),
    .C(_0916_),
    .D(_0927_),
    .X(_0936_));
 sg13g2_o21ai_1 _2531_ (.B1(net390),
    .Y(_0937_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .A2(net502));
 sg13g2_nand2_1 _2532_ (.Y(_0938_),
    .A(_0917_),
    .B(_0937_));
 sg13g2_a21oi_1 _2533_ (.A1(_0900_),
    .A2(_0936_),
    .Y(_0939_),
    .B1(_0938_));
 sg13g2_nand2_1 _2534_ (.Y(_0940_),
    .A(net841),
    .B(net390));
 sg13g2_xnor2_1 _2535_ (.Y(_0941_),
    .A(_1211_),
    .B(_0335_));
 sg13g2_a21oi_1 _2536_ (.A1(_0939_),
    .A2(_0941_),
    .Y(_0942_),
    .B1(_0685_));
 sg13g2_o21ai_1 _2537_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0939_),
    .A2(_0941_));
 sg13g2_a21oi_1 _2538_ (.A1(_1221_),
    .A2(net381),
    .Y(_0944_),
    .B1(_0672_));
 sg13g2_o21ai_1 _2539_ (.B1(_0944_),
    .Y(_0945_),
    .A1(net381),
    .A2(_0840_));
 sg13g2_and3_1 _2540_ (.X(_0946_),
    .A(_0838_),
    .B(_0860_),
    .C(_0945_));
 sg13g2_a221oi_1 _2541_ (.B2(_0946_),
    .C1(net459),
    .B1(_0943_),
    .A1(_1211_),
    .Y(_0213_),
    .A2(net370));
 sg13g2_o21ai_1 _2542_ (.B1(_0940_),
    .Y(_0947_),
    .A1(_0939_),
    .A2(_0941_));
 sg13g2_xnor2_1 _2543_ (.Y(_0948_),
    .A(net805),
    .B(net392));
 sg13g2_a21oi_1 _2544_ (.A1(_0947_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(_0685_));
 sg13g2_o21ai_1 _2545_ (.B1(_0949_),
    .Y(_0950_),
    .A1(_0947_),
    .A2(_0948_));
 sg13g2_nor2_1 _2546_ (.A(net381),
    .B(_0852_),
    .Y(_0951_));
 sg13g2_a21oi_1 _2547_ (.A1(_1220_),
    .A2(net381),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_a221oi_1 _2548_ (.B2(_0671_),
    .C1(_0861_),
    .B1(_0952_),
    .A1(_0691_),
    .Y(_0953_),
    .A2(_0850_));
 sg13g2_a221oi_1 _2549_ (.B2(_0953_),
    .C1(net459),
    .B1(_0950_),
    .A1(_1210_),
    .Y(_0214_),
    .A2(_0861_));
 sg13g2_o21ai_1 _2550_ (.B1(net429),
    .Y(_0954_),
    .A1(net495),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[0] ));
 sg13g2_a21oi_1 _2551_ (.A1(net495),
    .A2(_1208_),
    .Y(_0215_),
    .B1(_0954_));
 sg13g2_o21ai_1 _2552_ (.B1(net430),
    .Y(_0955_),
    .A1(net490),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[1] ));
 sg13g2_a21oi_1 _2553_ (.A1(net490),
    .A2(_1207_),
    .Y(_0216_),
    .B1(_0955_));
 sg13g2_o21ai_1 _2554_ (.B1(net431),
    .Y(_0956_),
    .A1(net489),
    .A2(net337));
 sg13g2_a21oi_1 _2555_ (.A1(net489),
    .A2(_1206_),
    .Y(_0217_),
    .B1(_0956_));
 sg13g2_o21ai_1 _2556_ (.B1(net431),
    .Y(_0957_),
    .A1(net497),
    .A2(net342));
 sg13g2_a21oi_1 _2557_ (.A1(net497),
    .A2(_1205_),
    .Y(_0218_),
    .B1(_0957_));
 sg13g2_o21ai_1 _2558_ (.B1(net433),
    .Y(_0958_),
    .A1(net498),
    .A2(net656));
 sg13g2_a21oi_1 _2559_ (.A1(net498),
    .A2(_1204_),
    .Y(_0219_),
    .B1(_0958_));
 sg13g2_o21ai_1 _2560_ (.B1(net433),
    .Y(_0959_),
    .A1(net499),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[5] ));
 sg13g2_a21oi_1 _2561_ (.A1(net499),
    .A2(_1203_),
    .Y(_0220_),
    .B1(_0959_));
 sg13g2_o21ai_1 _2562_ (.B1(net432),
    .Y(_0960_),
    .A1(net494),
    .A2(net628));
 sg13g2_a21oi_1 _2563_ (.A1(net494),
    .A2(_1202_),
    .Y(_0221_),
    .B1(_0960_));
 sg13g2_o21ai_1 _2564_ (.B1(net432),
    .Y(_0961_),
    .A1(net494),
    .A2(net692));
 sg13g2_a21oi_1 _2565_ (.A1(net494),
    .A2(_1201_),
    .Y(_0222_),
    .B1(_0961_));
 sg13g2_o21ai_1 _2566_ (.B1(net432),
    .Y(_0962_),
    .A1(net495),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[8] ));
 sg13g2_a21oi_1 _2567_ (.A1(net495),
    .A2(_1200_),
    .Y(_0223_),
    .B1(_0962_));
 sg13g2_o21ai_1 _2568_ (.B1(net431),
    .Y(_0963_),
    .A1(net489),
    .A2(net561));
 sg13g2_a21oi_1 _2569_ (.A1(net497),
    .A2(_1199_),
    .Y(_0224_),
    .B1(_0963_));
 sg13g2_o21ai_1 _2570_ (.B1(net431),
    .Y(_0964_),
    .A1(net497),
    .A2(net642));
 sg13g2_a21oi_1 _2571_ (.A1(net498),
    .A2(_1198_),
    .Y(_0225_),
    .B1(_0964_));
 sg13g2_o21ai_1 _2572_ (.B1(net433),
    .Y(_0965_),
    .A1(net498),
    .A2(net647));
 sg13g2_a21oi_1 _2573_ (.A1(net499),
    .A2(_1197_),
    .Y(_0226_),
    .B1(_0965_));
 sg13g2_o21ai_1 _2574_ (.B1(net433),
    .Y(_0966_),
    .A1(net499),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[12] ));
 sg13g2_a21oi_1 _2575_ (.A1(net499),
    .A2(_1196_),
    .Y(_0227_),
    .B1(_0966_));
 sg13g2_o21ai_1 _2576_ (.B1(net432),
    .Y(_0967_),
    .A1(net499),
    .A2(net609));
 sg13g2_a21oi_1 _2577_ (.A1(net495),
    .A2(_1195_),
    .Y(_0228_),
    .B1(_0967_));
 sg13g2_o21ai_1 _2578_ (.B1(net432),
    .Y(_0968_),
    .A1(net495),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[14] ));
 sg13g2_a21oi_1 _2579_ (.A1(net495),
    .A2(_1194_),
    .Y(_0229_),
    .B1(_0968_));
 sg13g2_o21ai_1 _2580_ (.B1(net431),
    .Y(_0969_),
    .A1(net489),
    .A2(net588));
 sg13g2_a21oi_1 _2581_ (.A1(net489),
    .A2(_1193_),
    .Y(_0230_),
    .B1(_0969_));
 sg13g2_o21ai_1 _2582_ (.B1(net427),
    .Y(_0970_),
    .A1(net484),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[16] ));
 sg13g2_a21oi_1 _2583_ (.A1(net484),
    .A2(_1192_),
    .Y(_0231_),
    .B1(_0970_));
 sg13g2_o21ai_1 _2584_ (.B1(net427),
    .Y(_0971_),
    .A1(net486),
    .A2(net352));
 sg13g2_a21oi_1 _2585_ (.A1(net486),
    .A2(_1191_),
    .Y(_0232_),
    .B1(_0971_));
 sg13g2_o21ai_1 _2586_ (.B1(net433),
    .Y(_0972_),
    .A1(net498),
    .A2(net697));
 sg13g2_a21oi_1 _2587_ (.A1(net498),
    .A2(_1190_),
    .Y(_0233_),
    .B1(_0972_));
 sg13g2_o21ai_1 _2588_ (.B1(net432),
    .Y(_0973_),
    .A1(net499),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[19] ));
 sg13g2_a21oi_1 _2589_ (.A1(net499),
    .A2(_1189_),
    .Y(_0234_),
    .B1(_0973_));
 sg13g2_o21ai_1 _2590_ (.B1(net432),
    .Y(_0974_),
    .A1(net493),
    .A2(net623));
 sg13g2_a21oi_1 _2591_ (.A1(net493),
    .A2(_1188_),
    .Y(_0235_),
    .B1(_0974_));
 sg13g2_o21ai_1 _2592_ (.B1(net428),
    .Y(_0975_),
    .A1(net493),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[21] ));
 sg13g2_a21oi_1 _2593_ (.A1(net493),
    .A2(_1187_),
    .Y(_0236_),
    .B1(_0975_));
 sg13g2_o21ai_1 _2594_ (.B1(net429),
    .Y(_0976_),
    .A1(net493),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[22] ));
 sg13g2_a21oi_1 _2595_ (.A1(net495),
    .A2(_1186_),
    .Y(_0237_),
    .B1(_0976_));
 sg13g2_o21ai_1 _2596_ (.B1(net431),
    .Y(_0977_),
    .A1(net490),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[23] ));
 sg13g2_a21oi_1 _2597_ (.A1(net489),
    .A2(_1185_),
    .Y(_0238_),
    .B1(_0977_));
 sg13g2_o21ai_1 _2598_ (.B1(net431),
    .Y(_0978_),
    .A1(net497),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[24] ));
 sg13g2_a21oi_1 _2599_ (.A1(net497),
    .A2(_1184_),
    .Y(_0239_),
    .B1(_0978_));
 sg13g2_o21ai_1 _2600_ (.B1(net433),
    .Y(_0979_),
    .A1(net497),
    .A2(net586));
 sg13g2_a21oi_1 _2601_ (.A1(net497),
    .A2(_1183_),
    .Y(_0240_),
    .B1(_0979_));
 sg13g2_o21ai_1 _2602_ (.B1(net432),
    .Y(_0980_),
    .A1(net500),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[26] ));
 sg13g2_a21oi_1 _2603_ (.A1(net493),
    .A2(_1182_),
    .Y(_0241_),
    .B1(_0980_));
 sg13g2_o21ai_1 _2604_ (.B1(net429),
    .Y(_0981_),
    .A1(net493),
    .A2(net550));
 sg13g2_a21oi_1 _2605_ (.A1(net493),
    .A2(_1181_),
    .Y(_0242_),
    .B1(_0981_));
 sg13g2_o21ai_1 _2606_ (.B1(net429),
    .Y(_0982_),
    .A1(net491),
    .A2(net596));
 sg13g2_a21oi_1 _2607_ (.A1(net492),
    .A2(_1180_),
    .Y(_0243_),
    .B1(_0982_));
 sg13g2_o21ai_1 _2608_ (.B1(net430),
    .Y(_0983_),
    .A1(net487),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[29] ));
 sg13g2_a21oi_1 _2609_ (.A1(net487),
    .A2(_1179_),
    .Y(_0244_),
    .B1(_0983_));
 sg13g2_o21ai_1 _2610_ (.B1(net425),
    .Y(_0984_),
    .A1(net484),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[30] ));
 sg13g2_a21oi_1 _2611_ (.A1(net484),
    .A2(_1178_),
    .Y(_0245_),
    .B1(_0984_));
 sg13g2_o21ai_1 _2612_ (.B1(net426),
    .Y(_0985_),
    .A1(net483),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[31] ));
 sg13g2_a21oi_1 _2613_ (.A1(net483),
    .A2(_1177_),
    .Y(_0246_),
    .B1(_0985_));
 sg13g2_o21ai_1 _2614_ (.B1(net427),
    .Y(_0986_),
    .A1(net483),
    .A2(net345));
 sg13g2_a21oi_1 _2615_ (.A1(net483),
    .A2(_1176_),
    .Y(_0247_),
    .B1(_0986_));
 sg13g2_o21ai_1 _2616_ (.B1(net431),
    .Y(_0987_),
    .A1(net484),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[33] ));
 sg13g2_a21oi_1 _2617_ (.A1(net489),
    .A2(_1175_),
    .Y(_0248_),
    .B1(_0987_));
 sg13g2_o21ai_1 _2618_ (.B1(net430),
    .Y(_0988_),
    .A1(net489),
    .A2(net675));
 sg13g2_a21oi_1 _2619_ (.A1(net487),
    .A2(_1174_),
    .Y(_0249_),
    .B1(_0988_));
 sg13g2_o21ai_1 _2620_ (.B1(net428),
    .Y(_0989_),
    .A1(net491),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[35] ));
 sg13g2_a21oi_1 _2621_ (.A1(net491),
    .A2(_1173_),
    .Y(_0250_),
    .B1(_0989_));
 sg13g2_o21ai_1 _2622_ (.B1(net430),
    .Y(_0990_),
    .A1(net487),
    .A2(net584));
 sg13g2_a21oi_1 _2623_ (.A1(net487),
    .A2(_1172_),
    .Y(_0251_),
    .B1(_0990_));
 sg13g2_o21ai_1 _2624_ (.B1(net425),
    .Y(_0991_),
    .A1(net482),
    .A2(net606));
 sg13g2_a21oi_1 _2625_ (.A1(net482),
    .A2(_1171_),
    .Y(_0252_),
    .B1(_0991_));
 sg13g2_o21ai_1 _2626_ (.B1(net425),
    .Y(_0992_),
    .A1(net482),
    .A2(net643));
 sg13g2_a21oi_1 _2627_ (.A1(net482),
    .A2(_1170_),
    .Y(_0253_),
    .B1(_0992_));
 sg13g2_o21ai_1 _2628_ (.B1(net425),
    .Y(_0993_),
    .A1(net481),
    .A2(net698));
 sg13g2_a21oi_1 _2629_ (.A1(net481),
    .A2(_1169_),
    .Y(_0254_),
    .B1(_0993_));
 sg13g2_o21ai_1 _2630_ (.B1(net430),
    .Y(_0994_),
    .A1(net488),
    .A2(net699));
 sg13g2_a21oi_1 _2631_ (.A1(net487),
    .A2(_1168_),
    .Y(_0255_),
    .B1(_0994_));
 sg13g2_o21ai_1 _2632_ (.B1(net428),
    .Y(_0995_),
    .A1(net487),
    .A2(net702));
 sg13g2_a21oi_1 _2633_ (.A1(net491),
    .A2(_1167_),
    .Y(_0256_),
    .B1(_0995_));
 sg13g2_o21ai_1 _2634_ (.B1(net428),
    .Y(_0996_),
    .A1(net491),
    .A2(net682));
 sg13g2_a21oi_1 _2635_ (.A1(net491),
    .A2(_1166_),
    .Y(_0257_),
    .B1(_0996_));
 sg13g2_o21ai_1 _2636_ (.B1(net430),
    .Y(_0997_),
    .A1(net488),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[43] ));
 sg13g2_a21oi_1 _2637_ (.A1(net488),
    .A2(_1165_),
    .Y(_0258_),
    .B1(_0997_));
 sg13g2_o21ai_1 _2638_ (.B1(net426),
    .Y(_0998_),
    .A1(net481),
    .A2(net356));
 sg13g2_a21oi_1 _2639_ (.A1(net481),
    .A2(_1164_),
    .Y(_0259_),
    .B1(_0998_));
 sg13g2_o21ai_1 _2640_ (.B1(net426),
    .Y(_0999_),
    .A1(net483),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[45] ));
 sg13g2_a21oi_1 _2641_ (.A1(net483),
    .A2(_1163_),
    .Y(_0260_),
    .B1(_0999_));
 sg13g2_o21ai_1 _2642_ (.B1(net425),
    .Y(_1000_),
    .A1(net483),
    .A2(net592));
 sg13g2_a21oi_1 _2643_ (.A1(net483),
    .A2(_1162_),
    .Y(_0261_),
    .B1(_1000_));
 sg13g2_o21ai_1 _2644_ (.B1(net428),
    .Y(_1001_),
    .A1(net492),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[47] ));
 sg13g2_a21oi_1 _2645_ (.A1(net492),
    .A2(_1161_),
    .Y(_0262_),
    .B1(_1001_));
 sg13g2_o21ai_1 _2646_ (.B1(net428),
    .Y(_1002_),
    .A1(net492),
    .A2(net570));
 sg13g2_a21oi_1 _2647_ (.A1(net492),
    .A2(_1160_),
    .Y(_0263_),
    .B1(_1002_));
 sg13g2_o21ai_1 _2648_ (.B1(net428),
    .Y(_1003_),
    .A1(net492),
    .A2(net638));
 sg13g2_a21oi_1 _2649_ (.A1(net491),
    .A2(_1159_),
    .Y(_0264_),
    .B1(_1003_));
 sg13g2_o21ai_1 _2650_ (.B1(net428),
    .Y(_1004_),
    .A1(net491),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[50] ));
 sg13g2_a21oi_1 _2651_ (.A1(net487),
    .A2(_1158_),
    .Y(_0265_),
    .B1(_1004_));
 sg13g2_o21ai_1 _2652_ (.B1(net430),
    .Y(_1005_),
    .A1(net488),
    .A2(net366));
 sg13g2_a21oi_1 _2653_ (.A1(net481),
    .A2(_1157_),
    .Y(_0266_),
    .B1(_1005_));
 sg13g2_o21ai_1 _2654_ (.B1(net425),
    .Y(_1006_),
    .A1(net482),
    .A2(net657));
 sg13g2_a21oi_1 _2655_ (.A1(net482),
    .A2(_1156_),
    .Y(_0267_),
    .B1(_1006_));
 sg13g2_o21ai_1 _2656_ (.B1(net425),
    .Y(_1007_),
    .A1(net482),
    .A2(net726));
 sg13g2_a21oi_1 _2657_ (.A1(net481),
    .A2(_1155_),
    .Y(_0268_),
    .B1(_1007_));
 sg13g2_o21ai_1 _2658_ (.B1(net425),
    .Y(_1008_),
    .A1(net481),
    .A2(net669));
 sg13g2_a21oi_1 _2659_ (.A1(net481),
    .A2(_1154_),
    .Y(_0269_),
    .B1(_1008_));
 sg13g2_o21ai_1 _2660_ (.B1(net426),
    .Y(_1009_),
    .A1(net485),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[55] ));
 sg13g2_a21oi_1 _2661_ (.A1(net485),
    .A2(_1153_),
    .Y(_0270_),
    .B1(_1009_));
 sg13g2_o21ai_1 _2662_ (.B1(net426),
    .Y(_1010_),
    .A1(net485),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[56] ));
 sg13g2_a21oi_1 _2663_ (.A1(net485),
    .A2(_1152_),
    .Y(_0271_),
    .B1(_1010_));
 sg13g2_o21ai_1 _2664_ (.B1(net426),
    .Y(_1011_),
    .A1(net485),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[57] ));
 sg13g2_a21oi_1 _2665_ (.A1(net485),
    .A2(_1151_),
    .Y(_0272_),
    .B1(_1011_));
 sg13g2_o21ai_1 _2666_ (.B1(net417),
    .Y(_1012_),
    .A1(net479),
    .A2(net563));
 sg13g2_a21oi_1 _2667_ (.A1(net479),
    .A2(_1150_),
    .Y(_0273_),
    .B1(_1012_));
 sg13g2_o21ai_1 _2668_ (.B1(net416),
    .Y(_1013_),
    .A1(net474),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[59] ));
 sg13g2_a21oi_1 _2669_ (.A1(net466),
    .A2(_1149_),
    .Y(_0274_),
    .B1(_1013_));
 sg13g2_o21ai_1 _2670_ (.B1(net412),
    .Y(_1014_),
    .A1(net465),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[60] ));
 sg13g2_a21oi_1 _2671_ (.A1(net465),
    .A2(_1148_),
    .Y(_0275_),
    .B1(_1014_));
 sg13g2_o21ai_1 _2672_ (.B1(net413),
    .Y(_1015_),
    .A1(net462),
    .A2(net590));
 sg13g2_a21oi_1 _2673_ (.A1(net462),
    .A2(_1147_),
    .Y(_0276_),
    .B1(_1015_));
 sg13g2_o21ai_1 _2674_ (.B1(net412),
    .Y(_1016_),
    .A1(net466),
    .A2(net660));
 sg13g2_a21oi_1 _2675_ (.A1(net466),
    .A2(_1146_),
    .Y(_0277_),
    .B1(_1016_));
 sg13g2_o21ai_1 _2676_ (.B1(net416),
    .Y(_1017_),
    .A1(net473),
    .A2(net650));
 sg13g2_a21oi_1 _2677_ (.A1(net473),
    .A2(_1145_),
    .Y(_0278_),
    .B1(_1017_));
 sg13g2_o21ai_1 _2678_ (.B1(net417),
    .Y(_1018_),
    .A1(net477),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[64] ));
 sg13g2_a21oi_1 _2679_ (.A1(net477),
    .A2(_1144_),
    .Y(_0279_),
    .B1(_1018_));
 sg13g2_o21ai_1 _2680_ (.B1(net417),
    .Y(_1019_),
    .A1(net477),
    .A2(net347));
 sg13g2_a21oi_1 _2681_ (.A1(net478),
    .A2(_1143_),
    .Y(_0280_),
    .B1(_1019_));
 sg13g2_o21ai_1 _2682_ (.B1(net418),
    .Y(_1020_),
    .A1(net473),
    .A2(net659));
 sg13g2_a21oi_1 _2683_ (.A1(net466),
    .A2(_1142_),
    .Y(_0281_),
    .B1(_1020_));
 sg13g2_o21ai_1 _2684_ (.B1(net412),
    .Y(_1021_),
    .A1(net465),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[67] ));
 sg13g2_a21oi_1 _2685_ (.A1(net467),
    .A2(_1141_),
    .Y(_0282_),
    .B1(_1021_));
 sg13g2_o21ai_1 _2686_ (.B1(net413),
    .Y(_1022_),
    .A1(net463),
    .A2(net574));
 sg13g2_a21oi_1 _2687_ (.A1(net463),
    .A2(_1140_),
    .Y(_0283_),
    .B1(_1022_));
 sg13g2_o21ai_1 _2688_ (.B1(net413),
    .Y(_1023_),
    .A1(net462),
    .A2(net637));
 sg13g2_a21oi_1 _2689_ (.A1(net462),
    .A2(_1139_),
    .Y(_0284_),
    .B1(_1023_));
 sg13g2_o21ai_1 _2690_ (.B1(net416),
    .Y(_1024_),
    .A1(net473),
    .A2(net667));
 sg13g2_a21oi_1 _2691_ (.A1(net473),
    .A2(_1138_),
    .Y(_0285_),
    .B1(_1024_));
 sg13g2_o21ai_1 _2692_ (.B1(net426),
    .Y(_1025_),
    .A1(net485),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[71] ));
 sg13g2_a21oi_1 _2693_ (.A1(net485),
    .A2(_1137_),
    .Y(_0286_),
    .B1(_1025_));
 sg13g2_o21ai_1 _2694_ (.B1(net417),
    .Y(_1026_),
    .A1(net477),
    .A2(net559));
 sg13g2_a21oi_1 _2695_ (.A1(net479),
    .A2(_1136_),
    .Y(_0287_),
    .B1(_1026_));
 sg13g2_o21ai_1 _2696_ (.B1(net416),
    .Y(_1027_),
    .A1(net473),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[73] ));
 sg13g2_a21oi_1 _2697_ (.A1(net466),
    .A2(_1135_),
    .Y(_0288_),
    .B1(_1027_));
 sg13g2_o21ai_1 _2698_ (.B1(net412),
    .Y(_1028_),
    .A1(net465),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[74] ));
 sg13g2_a21oi_1 _2699_ (.A1(net465),
    .A2(_1134_),
    .Y(_0289_),
    .B1(_1028_));
 sg13g2_o21ai_1 _2700_ (.B1(net413),
    .Y(_1029_),
    .A1(net462),
    .A2(net607));
 sg13g2_a21oi_1 _2701_ (.A1(net465),
    .A2(_1133_),
    .Y(_0290_),
    .B1(_1029_));
 sg13g2_o21ai_1 _2702_ (.B1(net412),
    .Y(_1030_),
    .A1(net466),
    .A2(net677));
 sg13g2_a21oi_1 _2703_ (.A1(net466),
    .A2(_1132_),
    .Y(_0291_),
    .B1(_1030_));
 sg13g2_o21ai_1 _2704_ (.B1(net417),
    .Y(_1031_),
    .A1(net478),
    .A2(net652));
 sg13g2_a21oi_1 _2705_ (.A1(net478),
    .A2(_1131_),
    .Y(_0292_),
    .B1(_1031_));
 sg13g2_o21ai_1 _2706_ (.B1(net417),
    .Y(_1032_),
    .A1(net477),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[78] ));
 sg13g2_a21oi_1 _2707_ (.A1(net477),
    .A2(_1130_),
    .Y(_0293_),
    .B1(_1032_));
 sg13g2_o21ai_1 _2708_ (.B1(net418),
    .Y(_1033_),
    .A1(net477),
    .A2(net364));
 sg13g2_a21oi_1 _2709_ (.A1(net477),
    .A2(_1129_),
    .Y(_0294_),
    .B1(_1033_));
 sg13g2_o21ai_1 _2710_ (.B1(net412),
    .Y(_1034_),
    .A1(net469),
    .A2(net706));
 sg13g2_a21oi_1 _2711_ (.A1(net469),
    .A2(_1128_),
    .Y(_0295_),
    .B1(_1034_));
 sg13g2_o21ai_1 _2712_ (.B1(net413),
    .Y(_1035_),
    .A1(net462),
    .A2(net700));
 sg13g2_a21oi_1 _2713_ (.A1(net463),
    .A2(_1127_),
    .Y(_0296_),
    .B1(_1035_));
 sg13g2_o21ai_1 _2714_ (.B1(net413),
    .Y(_1036_),
    .A1(net462),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[82] ));
 sg13g2_a21oi_1 _2715_ (.A1(net462),
    .A2(_1126_),
    .Y(_0297_),
    .B1(_1036_));
 sg13g2_o21ai_1 _2716_ (.B1(net413),
    .Y(_1037_),
    .A1(net463),
    .A2(net678));
 sg13g2_a21oi_1 _2717_ (.A1(net463),
    .A2(_1125_),
    .Y(_0298_),
    .B1(_1037_));
 sg13g2_o21ai_1 _2718_ (.B1(net412),
    .Y(_1038_),
    .A1(net466),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[84] ));
 sg13g2_a21oi_1 _2719_ (.A1(net467),
    .A2(_1124_),
    .Y(_0299_),
    .B1(_1038_));
 sg13g2_o21ai_1 _2720_ (.B1(net418),
    .Y(_1039_),
    .A1(net476),
    .A2(net358));
 sg13g2_a21oi_1 _2721_ (.A1(net475),
    .A2(_1123_),
    .Y(_0300_),
    .B1(_1039_));
 sg13g2_o21ai_1 _2722_ (.B1(net419),
    .Y(_1040_),
    .A1(net475),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[86] ));
 sg13g2_a21oi_1 _2723_ (.A1(net475),
    .A2(_1122_),
    .Y(_0301_),
    .B1(_1040_));
 sg13g2_o21ai_1 _2724_ (.B1(net419),
    .Y(_1041_),
    .A1(net474),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[87] ));
 sg13g2_a21oi_1 _2725_ (.A1(net474),
    .A2(_1121_),
    .Y(_0302_),
    .B1(_1041_));
 sg13g2_o21ai_1 _2726_ (.B1(net414),
    .Y(_1042_),
    .A1(net469),
    .A2(net354));
 sg13g2_a21oi_1 _2727_ (.A1(net468),
    .A2(_1120_),
    .Y(_0303_),
    .B1(_1042_));
 sg13g2_o21ai_1 _2728_ (.B1(net413),
    .Y(_1043_),
    .A1(net464),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[89] ));
 sg13g2_a21oi_1 _2729_ (.A1(net464),
    .A2(_1119_),
    .Y(_0304_),
    .B1(_1043_));
 sg13g2_o21ai_1 _2730_ (.B1(net415),
    .Y(_1044_),
    .A1(net465),
    .A2(net614));
 sg13g2_a21oi_1 _2731_ (.A1(net465),
    .A2(_1118_),
    .Y(_0305_),
    .B1(_1044_));
 sg13g2_o21ai_1 _2732_ (.B1(net416),
    .Y(_1045_),
    .A1(net473),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[91] ));
 sg13g2_a21oi_1 _2733_ (.A1(net473),
    .A2(_1117_),
    .Y(_0306_),
    .B1(_1045_));
 sg13g2_o21ai_1 _2734_ (.B1(net416),
    .Y(_1046_),
    .A1(net478),
    .A2(net568));
 sg13g2_a21oi_1 _2735_ (.A1(net478),
    .A2(_1116_),
    .Y(_0307_),
    .B1(_1046_));
 sg13g2_o21ai_1 _2736_ (.B1(net417),
    .Y(_1047_),
    .A1(net479),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[93] ));
 sg13g2_a21oi_1 _2737_ (.A1(net474),
    .A2(_1115_),
    .Y(_0308_),
    .B1(_1047_));
 sg13g2_o21ai_1 _2738_ (.B1(net419),
    .Y(_1048_),
    .A1(net474),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[94] ));
 sg13g2_a21oi_1 _2739_ (.A1(net468),
    .A2(_1114_),
    .Y(_0309_),
    .B1(_1048_));
 sg13g2_o21ai_1 _2740_ (.B1(net414),
    .Y(_1049_),
    .A1(net468),
    .A2(net597));
 sg13g2_a21oi_1 _2741_ (.A1(net468),
    .A2(_1113_),
    .Y(_0310_),
    .B1(_1049_));
 sg13g2_o21ai_1 _2742_ (.B1(net414),
    .Y(_1050_),
    .A1(net464),
    .A2(net635));
 sg13g2_a21oi_1 _2743_ (.A1(net464),
    .A2(_1112_),
    .Y(_0311_),
    .B1(_1050_));
 sg13g2_o21ai_1 _2744_ (.B1(net412),
    .Y(_1051_),
    .A1(net468),
    .A2(net680));
 sg13g2_a21oi_1 _2745_ (.A1(net468),
    .A2(_1111_),
    .Y(_0312_),
    .B1(_1051_));
 sg13g2_o21ai_1 _2746_ (.B1(net416),
    .Y(_1052_),
    .A1(net476),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[98] ));
 sg13g2_a21oi_1 _2747_ (.A1(net476),
    .A2(_1110_),
    .Y(_0313_),
    .B1(_1052_));
 sg13g2_o21ai_1 _2748_ (.B1(net418),
    .Y(_1053_),
    .A1(net478),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[99] ));
 sg13g2_a21oi_1 _2749_ (.A1(net478),
    .A2(_1109_),
    .Y(_0314_),
    .B1(_1053_));
 sg13g2_o21ai_1 _2750_ (.B1(net419),
    .Y(_1054_),
    .A1(net475),
    .A2(net362));
 sg13g2_a21oi_1 _2751_ (.A1(net475),
    .A2(_1108_),
    .Y(_0315_),
    .B1(_1054_));
 sg13g2_o21ai_1 _2752_ (.B1(net419),
    .Y(_1055_),
    .A1(net474),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[101] ));
 sg13g2_a21oi_1 _2753_ (.A1(net474),
    .A2(_1107_),
    .Y(_0316_),
    .B1(_1055_));
 sg13g2_o21ai_1 _2754_ (.B1(net415),
    .Y(_1056_),
    .A1(net472),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[102] ));
 sg13g2_a21oi_1 _2755_ (.A1(net472),
    .A2(_1106_),
    .Y(_0317_),
    .B1(_1056_));
 sg13g2_o21ai_1 _2756_ (.B1(net414),
    .Y(_1057_),
    .A1(net464),
    .A2(net594));
 sg13g2_a21oi_1 _2757_ (.A1(net464),
    .A2(_1105_),
    .Y(_0318_),
    .B1(_1057_));
 sg13g2_o21ai_1 _2758_ (.B1(net415),
    .Y(_1058_),
    .A1(net468),
    .A2(net645));
 sg13g2_a21oi_1 _2759_ (.A1(net468),
    .A2(_1104_),
    .Y(_0319_),
    .B1(_1058_));
 sg13g2_o21ai_1 _2760_ (.B1(net416),
    .Y(_1059_),
    .A1(net475),
    .A2(net749));
 sg13g2_a21oi_1 _2761_ (.A1(net479),
    .A2(_1103_),
    .Y(_0320_),
    .B1(_1059_));
 sg13g2_o21ai_1 _2762_ (.B1(net417),
    .Y(_1060_),
    .A1(net480),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[106] ));
 sg13g2_a21oi_1 _2763_ (.A1(net480),
    .A2(_1102_),
    .Y(_0321_),
    .B1(_1060_));
 sg13g2_o21ai_1 _2764_ (.B1(net420),
    .Y(_1061_),
    .A1(net479),
    .A2(net612));
 sg13g2_a21oi_1 _2765_ (.A1(net479),
    .A2(_1101_),
    .Y(_0322_),
    .B1(_1061_));
 sg13g2_o21ai_1 _2766_ (.B1(net419),
    .Y(_1062_),
    .A1(net474),
    .A2(net616));
 sg13g2_a21oi_1 _2767_ (.A1(net469),
    .A2(_1100_),
    .Y(_0323_),
    .B1(_1062_));
 sg13g2_o21ai_1 _2768_ (.B1(net415),
    .Y(_1063_),
    .A1(net472),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[109] ));
 sg13g2_a21oi_1 _2769_ (.A1(net472),
    .A2(_1099_),
    .Y(_0324_),
    .B1(_1063_));
 sg13g2_o21ai_1 _2770_ (.B1(net414),
    .Y(_1064_),
    .A1(net471),
    .A2(\ppwm_i.u_ppwm.u_mem.memory[110] ));
 sg13g2_a21oi_1 _2771_ (.A1(_1097_),
    .A2(net471),
    .Y(_0325_),
    .B1(_1064_));
 sg13g2_o21ai_1 _2772_ (.B1(net414),
    .Y(_1065_),
    .A1(net582),
    .A2(net471));
 sg13g2_a21oi_1 _2773_ (.A1(_1098_),
    .A2(net471),
    .Y(_0326_),
    .B1(_1065_));
 sg13g2_nand2b_1 _2774_ (.Y(_1066_),
    .B(net324),
    .A_N(net471));
 sg13g2_nand2_2 _2775_ (.Y(_1067_),
    .A(net421),
    .B(_1066_));
 sg13g2_xnor2_1 _2776_ (.Y(_1068_),
    .A(net751),
    .B(net471));
 sg13g2_nor2_1 _2777_ (.A(_1067_),
    .B(_1068_),
    .Y(_0327_));
 sg13g2_a21oi_1 _2778_ (.A1(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .A2(net472),
    .Y(_1069_),
    .B1(net339));
 sg13g2_and3_1 _2779_ (.X(_1070_),
    .A(net339),
    .B(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .C(net472));
 sg13g2_nor3_1 _2780_ (.A(_1067_),
    .B(net340),
    .C(_1070_),
    .Y(_0328_));
 sg13g2_nor2_1 _2781_ (.A(net716),
    .B(_1070_),
    .Y(_1071_));
 sg13g2_and2_1 _2782_ (.A(net716),
    .B(_1070_),
    .X(_1072_));
 sg13g2_nor3_1 _2783_ (.A(_1067_),
    .B(net717),
    .C(_1072_),
    .Y(_0329_));
 sg13g2_and2_1 _2784_ (.A(net661),
    .B(_1072_),
    .X(_1073_));
 sg13g2_nor2_1 _2785_ (.A(net661),
    .B(_1072_),
    .Y(_1074_));
 sg13g2_nor3_1 _2786_ (.A(_1067_),
    .B(_1073_),
    .C(net662),
    .Y(_0330_));
 sg13g2_xnor2_1 _2787_ (.Y(_1075_),
    .A(net748),
    .B(_1073_));
 sg13g2_nor2_1 _2788_ (.A(_1067_),
    .B(_1075_),
    .Y(_0331_));
 sg13g2_a21oi_1 _2789_ (.A1(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .A2(_1073_),
    .Y(_1076_),
    .B1(net330));
 sg13g2_and3_1 _2790_ (.X(_1077_),
    .A(net330),
    .B(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .C(_1073_));
 sg13g2_nor3_1 _2791_ (.A(_1067_),
    .B(net331),
    .C(_1077_),
    .Y(_0332_));
 sg13g2_and2_1 _2792_ (.A(net694),
    .B(_1077_),
    .X(_1078_));
 sg13g2_a21oi_1 _2793_ (.A1(net694),
    .A2(_1066_),
    .Y(_1079_),
    .B1(_1077_));
 sg13g2_nor3_1 _2794_ (.A(net457),
    .B(_1078_),
    .C(net695),
    .Y(_0333_));
 sg13g2_nand2b_1 _2795_ (.Y(_1080_),
    .B(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .A_N(\ppwm_i.u_ppwm.u_pwm.counter[1] ));
 sg13g2_o21ai_1 _2796_ (.B1(_1080_),
    .Y(_1081_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .A2(_1247_));
 sg13g2_o21ai_1 _2797_ (.B1(_1081_),
    .Y(_1082_),
    .A1(_1240_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ));
 sg13g2_o21ai_1 _2798_ (.B1(_1082_),
    .Y(_1083_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .A2(_1246_));
 sg13g2_a22oi_1 _2799_ (.Y(_1084_),
    .B1(_1246_),
    .B2(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .A2(_1245_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[3] ));
 sg13g2_nand2b_1 _2800_ (.Y(_1085_),
    .B(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .A_N(\ppwm_i.u_ppwm.u_pwm.counter[4] ));
 sg13g2_o21ai_1 _2801_ (.B1(_1085_),
    .Y(_1086_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .A2(_1245_));
 sg13g2_a21oi_1 _2802_ (.A1(_1083_),
    .A2(_1084_),
    .Y(_1087_),
    .B1(_1086_));
 sg13g2_a221oi_1 _2803_ (.B2(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .C1(_1087_),
    .B1(_1244_),
    .A1(net520),
    .Y(_1088_),
    .A2(_1243_));
 sg13g2_a221oi_1 _2804_ (.B2(_1239_),
    .C1(_1088_),
    .B1(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .A1(_1238_),
    .Y(_1089_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ));
 sg13g2_nand2b_1 _2805_ (.Y(_1090_),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .A_N(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ));
 sg13g2_o21ai_1 _2806_ (.B1(_1090_),
    .Y(_1091_),
    .A1(_1238_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ));
 sg13g2_a22oi_1 _2807_ (.Y(_1092_),
    .B1(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ),
    .B2(_1237_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .A1(_1236_));
 sg13g2_o21ai_1 _2808_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_1089_),
    .A2(_1091_));
 sg13g2_a22oi_1 _2809_ (.Y(_1094_),
    .B1(_1242_),
    .B2(net839),
    .A2(_1241_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[9] ));
 sg13g2_a22oi_1 _2810_ (.Y(_1095_),
    .B1(_1093_),
    .B2(net840),
    .A2(net725),
    .A1(_1234_));
 sg13g2_o21ai_1 _2811_ (.B1(net414),
    .Y(_1096_),
    .A1(net712),
    .A2(_1095_));
 sg13g2_a21oi_1 _2812_ (.A1(net712),
    .A2(_1095_),
    .Y(_0334_),
    .B1(_1096_));
 sg13g2_buf_1 _2813_ (.A(net276),
    .X(_0076_));
 sg13g2_buf_1 _2814_ (.A(net229),
    .X(_0077_));
 sg13g2_buf_1 _2815_ (.A(net285),
    .X(_0078_));
 sg13g2_buf_1 _2816_ (.A(net220),
    .X(_0079_));
 sg13g2_buf_1 _2817_ (.A(net273),
    .X(_0080_));
 sg13g2_buf_1 _2818_ (.A(net240),
    .X(_0081_));
 sg13g2_buf_1 _2819_ (.A(net304),
    .X(_0082_));
 sg13g2_buf_1 _2820_ (.A(net235),
    .X(_0083_));
 sg13g2_buf_1 _2821_ (.A(net295),
    .X(_0084_));
 sg13g2_buf_1 _2822_ (.A(net263),
    .X(_0085_));
 sg13g2_buf_1 _2823_ (.A(net279),
    .X(_0086_));
 sg13g2_buf_1 _2824_ (.A(net244),
    .X(_0087_));
 sg13g2_buf_1 _2825_ (.A(net303),
    .X(_0088_));
 sg13g2_buf_1 _2826_ (.A(net264),
    .X(_0089_));
 sg13g2_buf_1 _2827_ (.A(net289),
    .X(_0090_));
 sg13g2_buf_1 _2828_ (.A(net221),
    .X(_0091_));
 sg13g2_buf_1 _2829_ (.A(net272),
    .X(_0092_));
 sg13g2_buf_1 _2830_ (.A(net232),
    .X(_0093_));
 sg13g2_buf_1 _2831_ (.A(net287),
    .X(_0094_));
 sg13g2_buf_1 _2832_ (.A(net252),
    .X(_0095_));
 sg13g2_buf_1 _2833_ (.A(net274),
    .X(_0096_));
 sg13g2_buf_1 _2834_ (.A(net237),
    .X(_0097_));
 sg13g2_buf_1 _2835_ (.A(net281),
    .X(_0098_));
 sg13g2_buf_1 _2836_ (.A(net241),
    .X(_0099_));
 sg13g2_buf_1 _2837_ (.A(net275),
    .X(_0100_));
 sg13g2_buf_1 _2838_ (.A(net226),
    .X(_0101_));
 sg13g2_buf_1 _2839_ (.A(net312),
    .X(_0102_));
 sg13g2_buf_1 _2840_ (.A(net249),
    .X(_0103_));
 sg13g2_buf_1 _2841_ (.A(net311),
    .X(_0104_));
 sg13g2_buf_1 _2842_ (.A(net248),
    .X(_0105_));
 sg13g2_buf_1 _2843_ (.A(net310),
    .X(_0106_));
 sg13g2_buf_1 _2844_ (.A(net225),
    .X(_0107_));
 sg13g2_buf_1 _2845_ (.A(net286),
    .X(_0108_));
 sg13g2_buf_1 _2846_ (.A(net233),
    .X(_0109_));
 sg13g2_buf_1 _2847_ (.A(net284),
    .X(_0110_));
 sg13g2_buf_1 _2848_ (.A(net224),
    .X(_0111_));
 sg13g2_buf_1 _2849_ (.A(net288),
    .X(_0112_));
 sg13g2_buf_1 _2850_ (.A(net223),
    .X(_0113_));
 sg13g2_buf_1 _2851_ (.A(net290),
    .X(_0114_));
 sg13g2_buf_1 _2852_ (.A(net219),
    .X(_0115_));
 sg13g2_buf_1 _2853_ (.A(net293),
    .X(_0116_));
 sg13g2_buf_1 _2854_ (.A(net245),
    .X(_0117_));
 sg13g2_buf_1 _2855_ (.A(net278),
    .X(_0118_));
 sg13g2_buf_1 _2856_ (.A(net236),
    .X(_0119_));
 sg13g2_buf_1 _2857_ (.A(net299),
    .X(_0120_));
 sg13g2_buf_1 _2858_ (.A(net256),
    .X(_0121_));
 sg13g2_buf_1 _2859_ (.A(net309),
    .X(_0122_));
 sg13g2_buf_1 _2860_ (.A(net243),
    .X(_0123_));
 sg13g2_buf_1 _2861_ (.A(net282),
    .X(_0124_));
 sg13g2_buf_1 _2862_ (.A(net242),
    .X(_0125_));
 sg13g2_buf_1 _2863_ (.A(net271),
    .X(_0126_));
 sg13g2_buf_1 _2864_ (.A(net250),
    .X(_0127_));
 sg13g2_buf_1 _2865_ (.A(net316),
    .X(_0128_));
 sg13g2_buf_1 _2866_ (.A(net238),
    .X(_0129_));
 sg13g2_buf_1 _2867_ (.A(net280),
    .X(_0130_));
 sg13g2_buf_1 _2868_ (.A(net247),
    .X(_0131_));
 sg13g2_buf_1 _2869_ (.A(net296),
    .X(_0132_));
 sg13g2_buf_1 _2870_ (.A(net222),
    .X(_0133_));
 sg13g2_buf_1 _2871_ (.A(net294),
    .X(_0134_));
 sg13g2_buf_1 _2872_ (.A(net234),
    .X(_0135_));
 sg13g2_buf_1 _2873_ (.A(net301),
    .X(_0136_));
 sg13g2_buf_1 _2874_ (.A(net228),
    .X(_0137_));
 sg13g2_buf_1 _2875_ (.A(net277),
    .X(_0138_));
 sg13g2_buf_1 _2876_ (.A(net251),
    .X(_0139_));
 sg13g2_buf_1 _2877_ (.A(net300),
    .X(_0140_));
 sg13g2_buf_1 _2878_ (.A(net239),
    .X(_0141_));
 sg13g2_buf_1 _2879_ (.A(net283),
    .X(_0142_));
 sg13g2_buf_1 _2880_ (.A(net227),
    .X(_0143_));
 sg13g2_buf_1 _2881_ (.A(net302),
    .X(_0144_));
 sg13g2_buf_1 _2882_ (.A(net253),
    .X(_0145_));
 sg13g2_buf_1 _2883_ (.A(net315),
    .X(_0146_));
 sg13g2_buf_1 _2884_ (.A(net246),
    .X(_0147_));
 sg13g2_dfrbpq_1 _2885_ (.RESET_B(net523),
    .D(_0076_),
    .Q(\sdr_i.DP_1.matrix[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2886_ (.RESET_B(net523),
    .D(_0077_),
    .Q(\sdr_i.DP_1.matrix[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2887_ (.RESET_B(net521),
    .D(_0078_),
    .Q(\sdr_i.DP_1.matrix[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2888_ (.RESET_B(net521),
    .D(_0079_),
    .Q(\sdr_i.DP_1.matrix[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2889_ (.RESET_B(net527),
    .D(_0080_),
    .Q(\sdr_i.DP_1.matrix[18] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2890_ (.RESET_B(net525),
    .D(_0081_),
    .Q(\sdr_i.DP_1.matrix[19] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2891_ (.RESET_B(net535),
    .D(_0082_),
    .Q(\sdr_i.DP_1.matrix[27] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2892_ (.RESET_B(net535),
    .D(_0083_),
    .Q(\sdr_i.DP_1.matrix[28] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2893_ (.RESET_B(net529),
    .D(_0084_),
    .Q(\sdr_i.DP_1.matrix[36] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2894_ (.RESET_B(net529),
    .D(_0085_),
    .Q(\sdr_i.DP_1.matrix[37] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2895_ (.RESET_B(net531),
    .D(_0086_),
    .Q(\sdr_i.DP_1.matrix[45] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2896_ (.RESET_B(net531),
    .D(_0087_),
    .Q(\sdr_i.DP_1.matrix[46] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2897_ (.RESET_B(net528),
    .D(_0088_),
    .Q(\sdr_i.DP_1.matrix[54] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2898_ (.RESET_B(net529),
    .D(_0089_),
    .Q(\sdr_i.DP_1.matrix[55] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2899_ (.RESET_B(net528),
    .D(_0090_),
    .Q(\sdr_i.DP_1.matrix[63] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2900_ (.RESET_B(net528),
    .D(_0091_),
    .Q(\sdr_i.DP_1.matrix[64] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2901_ (.RESET_B(net521),
    .D(_0092_),
    .Q(\sdr_i.DP_1.matrix[72] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2902_ (.RESET_B(net521),
    .D(_0093_),
    .Q(\sdr_i.DP_1.matrix[73] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2903_ (.RESET_B(net523),
    .D(_0094_),
    .Q(\sdr_i.DP_2.matrix[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2904_ (.RESET_B(net523),
    .D(_0095_),
    .Q(\sdr_i.DP_2.matrix[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2905_ (.RESET_B(net521),
    .D(_0096_),
    .Q(\sdr_i.DP_2.matrix[9] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2906_ (.RESET_B(net521),
    .D(_0097_),
    .Q(\sdr_i.DP_2.matrix[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2907_ (.RESET_B(net525),
    .D(_0098_),
    .Q(\sdr_i.DP_2.matrix[18] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2908_ (.RESET_B(net527),
    .D(_0099_),
    .Q(\sdr_i.DP_2.matrix[19] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2909_ (.RESET_B(net535),
    .D(_0100_),
    .Q(\sdr_i.DP_2.matrix[27] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2910_ (.RESET_B(net535),
    .D(_0101_),
    .Q(\sdr_i.DP_2.matrix[28] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2911_ (.RESET_B(net529),
    .D(_0102_),
    .Q(\sdr_i.DP_2.matrix[36] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2912_ (.RESET_B(net529),
    .D(_0103_),
    .Q(\sdr_i.DP_2.matrix[37] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2913_ (.RESET_B(net532),
    .D(_0104_),
    .Q(\sdr_i.DP_2.matrix[45] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2914_ (.RESET_B(net532),
    .D(_0105_),
    .Q(\sdr_i.DP_2.matrix[46] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2915_ (.RESET_B(net528),
    .D(_0106_),
    .Q(\sdr_i.DP_2.matrix[54] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2916_ (.RESET_B(net528),
    .D(_0107_),
    .Q(\sdr_i.DP_2.matrix[55] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2917_ (.RESET_B(net530),
    .D(_0108_),
    .Q(\sdr_i.DP_2.matrix[63] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2918_ (.RESET_B(net528),
    .D(_0109_),
    .Q(\sdr_i.DP_2.matrix[64] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2919_ (.RESET_B(net521),
    .D(_0110_),
    .Q(\sdr_i.DP_2.matrix[72] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2920_ (.RESET_B(net521),
    .D(_0111_),
    .Q(\sdr_i.DP_2.matrix[73] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2921_ (.RESET_B(net544),
    .D(_0112_),
    .Q(\sdr_i.DP_3.matrix[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2922_ (.RESET_B(net545),
    .D(_0113_),
    .Q(\sdr_i.DP_3.matrix[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2923_ (.RESET_B(net546),
    .D(_0114_),
    .Q(\sdr_i.DP_3.matrix[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2924_ (.RESET_B(net546),
    .D(_0115_),
    .Q(\sdr_i.DP_3.matrix[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2925_ (.RESET_B(net538),
    .D(_0116_),
    .Q(\sdr_i.DP_3.matrix[18] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2926_ (.RESET_B(net538),
    .D(_0117_),
    .Q(\sdr_i.DP_3.matrix[19] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2927_ (.RESET_B(net540),
    .D(_0118_),
    .Q(\sdr_i.DP_3.matrix[27] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2928_ (.RESET_B(net539),
    .D(_0119_),
    .Q(\sdr_i.DP_3.matrix[28] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2929_ (.RESET_B(net537),
    .D(_0120_),
    .Q(\sdr_i.DP_3.matrix[36] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2930_ (.RESET_B(net536),
    .D(_0121_),
    .Q(\sdr_i.DP_3.matrix[37] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2931_ (.RESET_B(net542),
    .D(_0122_),
    .Q(\sdr_i.DP_3.matrix[45] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2932_ (.RESET_B(net543),
    .D(_0123_),
    .Q(\sdr_i.DP_3.matrix[46] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2933_ (.RESET_B(net535),
    .D(_0124_),
    .Q(\sdr_i.DP_3.matrix[54] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2934_ (.RESET_B(net535),
    .D(_0125_),
    .Q(\sdr_i.DP_3.matrix[55] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2935_ (.RESET_B(net538),
    .D(_0126_),
    .Q(\sdr_i.DP_3.matrix[63] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2936_ (.RESET_B(net538),
    .D(_0127_),
    .Q(\sdr_i.DP_3.matrix[64] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2937_ (.RESET_B(net533),
    .D(_0128_),
    .Q(\sdr_i.DP_3.matrix[72] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2938_ (.RESET_B(net527),
    .D(_0129_),
    .Q(\sdr_i.DP_3.matrix[73] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2939_ (.RESET_B(net545),
    .D(_0130_),
    .Q(\sdr_i.DP_4.matrix[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2940_ (.RESET_B(net545),
    .D(_0131_),
    .Q(\sdr_i.DP_4.matrix[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2941_ (.RESET_B(net546),
    .D(_0132_),
    .Q(\sdr_i.DP_4.matrix[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2942_ (.RESET_B(net546),
    .D(_0133_),
    .Q(\sdr_i.DP_4.matrix[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2943_ (.RESET_B(net539),
    .D(_0134_),
    .Q(\sdr_i.DP_4.matrix[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2944_ (.RESET_B(net539),
    .D(_0135_),
    .Q(\sdr_i.DP_4.matrix[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2945_ (.RESET_B(net539),
    .D(_0136_),
    .Q(\sdr_i.DP_4.matrix[27] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2946_ (.RESET_B(net540),
    .D(_0137_),
    .Q(\sdr_i.DP_4.matrix[28] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2947_ (.RESET_B(net536),
    .D(_0138_),
    .Q(\sdr_i.DP_4.matrix[36] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2948_ (.RESET_B(net536),
    .D(_0139_),
    .Q(\sdr_i.DP_4.matrix[37] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2949_ (.RESET_B(net542),
    .D(_0140_),
    .Q(\sdr_i.DP_4.matrix[45] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2950_ (.RESET_B(net542),
    .D(_0141_),
    .Q(\sdr_i.DP_4.matrix[46] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2951_ (.RESET_B(net535),
    .D(_0142_),
    .Q(\sdr_i.DP_4.matrix[54] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2952_ (.RESET_B(net537),
    .D(_0143_),
    .Q(\sdr_i.DP_4.matrix[55] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2953_ (.RESET_B(net538),
    .D(_0144_),
    .Q(\sdr_i.DP_4.matrix[63] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2954_ (.RESET_B(net538),
    .D(_0145_),
    .Q(\sdr_i.DP_4.matrix[64] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2955_ (.RESET_B(net533),
    .D(_0146_),
    .Q(\sdr_i.DP_4.matrix[72] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2956_ (.RESET_B(net533),
    .D(_0147_),
    .Q(\sdr_i.DP_4.matrix[73] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _2957_ (.RESET_B(net421),
    .D(net327),
    .Q(\ppwm_i.u_ppwm.global_counter[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _2958_ (.RESET_B(net421),
    .D(net824),
    .Q(\ppwm_i.u_ppwm.global_counter[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _2959_ (.RESET_B(net422),
    .D(net711),
    .Q(\ppwm_i.u_ppwm.global_counter[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _2960_ (.RESET_B(net435),
    .D(net790),
    .Q(\ppwm_i.u_ppwm.global_counter[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2961_ (.RESET_B(net435),
    .D(_0152_),
    .Q(\ppwm_i.u_ppwm.global_counter[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2962_ (.RESET_B(net435),
    .D(net334),
    .Q(\ppwm_i.u_ppwm.global_counter[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2963_ (.RESET_B(net436),
    .D(net321),
    .Q(\ppwm_i.u_ppwm.global_counter[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2964_ (.RESET_B(net436),
    .D(net655),
    .Q(\ppwm_i.u_ppwm.global_counter[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2965_ (.RESET_B(net436),
    .D(_0156_),
    .Q(\ppwm_i.u_ppwm.global_counter[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2966_ (.RESET_B(net437),
    .D(net336),
    .Q(\ppwm_i.u_ppwm.global_counter[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2967_ (.RESET_B(net435),
    .D(net558),
    .Q(\ppwm_i.u_ppwm.global_counter[10] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2968_ (.RESET_B(net435),
    .D(_0159_),
    .Q(\ppwm_i.u_ppwm.global_counter[11] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2969_ (.RESET_B(net435),
    .D(net721),
    .Q(\ppwm_i.u_ppwm.global_counter[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2970_ (.RESET_B(net437),
    .D(net777),
    .Q(\ppwm_i.u_ppwm.global_counter[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2971_ (.RESET_B(net437),
    .D(_0162_),
    .Q(\ppwm_i.u_ppwm.global_counter[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2972_ (.RESET_B(net436),
    .D(net573),
    .Q(\ppwm_i.u_ppwm.global_counter[15] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2973_ (.RESET_B(net436),
    .D(net781),
    .Q(\ppwm_i.u_ppwm.global_counter[16] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2974_ (.RESET_B(net436),
    .D(net799),
    .Q(\ppwm_i.u_ppwm.global_counter[17] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2975_ (.RESET_B(net436),
    .D(_0166_),
    .Q(\ppwm_i.u_ppwm.global_counter[18] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2976_ (.RESET_B(net423),
    .D(net329),
    .Q(\ppwm_i.u_ppwm.global_counter[19] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2977_ (.RESET_B(net192),
    .D(net323),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2978_ (.RESET_B(net190),
    .D(net579),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2979_ (.RESET_B(net188),
    .D(net795),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2980_ (.RESET_B(net186),
    .D(net772),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2981_ (.RESET_B(net184),
    .D(_0172_),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2982_ (.RESET_B(net182),
    .D(_0173_),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2983_ (.RESET_B(net180),
    .D(net665),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2984_ (.RESET_B(net179),
    .D(net581),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2985_ (.RESET_B(net177),
    .D(_0176_),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2986_ (.RESET_B(net175),
    .D(_0177_),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[9] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2987_ (.RESET_B(net173),
    .D(_0178_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2988_ (.RESET_B(net171),
    .D(net709),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2989_ (.RESET_B(net169),
    .D(_0180_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2990_ (.RESET_B(net167),
    .D(_0181_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2991_ (.RESET_B(net165),
    .D(_0182_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2992_ (.RESET_B(net163),
    .D(_0183_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2993_ (.RESET_B(net161),
    .D(_0184_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2994_ (.RESET_B(net159),
    .D(_0185_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2995_ (.RESET_B(net157),
    .D(_0186_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2996_ (.RESET_B(net155),
    .D(_0187_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2997_ (.RESET_B(net153),
    .D(net567),
    .Q(\ppwm_i.u_ppwm.period_start ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2998_ (.RESET_B(net152),
    .D(_0189_),
    .Q(\ppwm_i.u_ppwm.pc[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2999_ (.RESET_B(net150),
    .D(_0190_),
    .Q(\ppwm_i.u_ppwm.pc[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3000_ (.RESET_B(net148),
    .D(_0191_),
    .Q(\ppwm_i.u_ppwm.pc[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3001_ (.RESET_B(net146),
    .D(_0192_),
    .Q(\ppwm_i.u_ppwm.pc[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3002_ (.RESET_B(net144),
    .D(net351),
    .Q(\ppwm_i.u_ppwm.u_ex.cmp_flag_q ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3003_ (.RESET_B(net142),
    .D(net713),
    .Q(\ppwm_i.u_ppwm.polarity ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3004_ (.RESET_B(net140),
    .D(net801),
    .Q(\ppwm_i.u_ppwm.pwm_value[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _3005_ (.RESET_B(net138),
    .D(net832),
    .Q(\ppwm_i.u_ppwm.pwm_value[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _3006_ (.RESET_B(net136),
    .D(_0197_),
    .Q(\ppwm_i.u_ppwm.pwm_value[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3007_ (.RESET_B(net134),
    .D(_0198_),
    .Q(\ppwm_i.u_ppwm.pwm_value[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3008_ (.RESET_B(net132),
    .D(_0199_),
    .Q(\ppwm_i.u_ppwm.pwm_value[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _3009_ (.RESET_B(net130),
    .D(net829),
    .Q(\ppwm_i.u_ppwm.pwm_value[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _3010_ (.RESET_B(net128),
    .D(_0201_),
    .Q(\ppwm_i.u_ppwm.pwm_value[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3011_ (.RESET_B(net126),
    .D(net834),
    .Q(\ppwm_i.u_ppwm.pwm_value[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _3012_ (.RESET_B(net124),
    .D(net815),
    .Q(\ppwm_i.u_ppwm.pwm_value[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _3013_ (.RESET_B(net122),
    .D(_0204_),
    .Q(\ppwm_i.u_ppwm.pwm_value[9] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _3014_ (.RESET_B(net120),
    .D(_0205_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _3015_ (.RESET_B(net118),
    .D(_0206_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _3016_ (.RESET_B(net116),
    .D(_0207_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3017_ (.RESET_B(net115),
    .D(_0208_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3018_ (.RESET_B(net113),
    .D(_0209_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _3019_ (.RESET_B(net111),
    .D(_0210_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3020_ (.RESET_B(net109),
    .D(net837),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _3021_ (.RESET_B(net107),
    .D(_0212_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _3022_ (.RESET_B(net105),
    .D(net810),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _3023_ (.RESET_B(net103),
    .D(_0214_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3024_ (.RESET_B(net101),
    .D(net344),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3025_ (.RESET_B(net99),
    .D(net338),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3026_ (.RESET_B(net97),
    .D(_0217_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3027_ (.RESET_B(net95),
    .D(_0218_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3028_ (.RESET_B(net93),
    .D(net685),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3029_ (.RESET_B(net91),
    .D(net629),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3030_ (.RESET_B(net89),
    .D(_0221_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3031_ (.RESET_B(net87),
    .D(net693),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3032_ (.RESET_B(net85),
    .D(net562),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[8] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3033_ (.RESET_B(net83),
    .D(_0224_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3034_ (.RESET_B(net81),
    .D(net648),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[10] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3035_ (.RESET_B(net79),
    .D(_0226_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3036_ (.RESET_B(net77),
    .D(net610),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[12] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3037_ (.RESET_B(net75),
    .D(_0228_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3038_ (.RESET_B(net73),
    .D(net589),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[14] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3039_ (.RESET_B(net71),
    .D(_0230_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[15] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(net69),
    .D(net353),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(net67),
    .D(_0232_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[17] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(net65),
    .D(_0233_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[18] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3043_ (.RESET_B(net63),
    .D(net624),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[19] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3044_ (.RESET_B(net61),
    .D(_0235_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3045_ (.RESET_B(net59),
    .D(net622),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[21] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3046_ (.RESET_B(net57),
    .D(net618),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3047_ (.RESET_B(net55),
    .D(net600),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3048_ (.RESET_B(net53),
    .D(net587),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[24] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3049_ (.RESET_B(net52),
    .D(_0240_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[25] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3050_ (.RESET_B(net50),
    .D(net551),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[26] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3051_ (.RESET_B(net48),
    .D(_0242_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3052_ (.RESET_B(net46),
    .D(_0243_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[28] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3053_ (.RESET_B(net44),
    .D(net577),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[29] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3054_ (.RESET_B(net42),
    .D(net361),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3055_ (.RESET_B(net40),
    .D(net346),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[31] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3056_ (.RESET_B(net38),
    .D(net689),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[32] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3057_ (.RESET_B(net36),
    .D(net676),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[33] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3058_ (.RESET_B(net34),
    .D(_0249_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3059_ (.RESET_B(net32),
    .D(net585),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[35] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3060_ (.RESET_B(net30),
    .D(_0251_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3061_ (.RESET_B(net28),
    .D(net644),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3062_ (.RESET_B(net189),
    .D(_0253_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3063_ (.RESET_B(net185),
    .D(_0254_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[39] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3064_ (.RESET_B(net181),
    .D(_0255_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[40] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3065_ (.RESET_B(net178),
    .D(_0256_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3066_ (.RESET_B(net174),
    .D(net683),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[42] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3067_ (.RESET_B(net170),
    .D(net357),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[43] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3068_ (.RESET_B(net166),
    .D(_0259_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3069_ (.RESET_B(net162),
    .D(net593),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[45] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3070_ (.RESET_B(net158),
    .D(_0261_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[46] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3071_ (.RESET_B(net154),
    .D(net571),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[47] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _3072_ (.RESET_B(net149),
    .D(_0263_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3073_ (.RESET_B(net145),
    .D(_0264_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[49] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3074_ (.RESET_B(net141),
    .D(net367),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[50] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3075_ (.RESET_B(net137),
    .D(_0266_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3076_ (.RESET_B(net133),
    .D(net658),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[52] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3077_ (.RESET_B(net129),
    .D(_0268_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[53] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3078_ (.RESET_B(net125),
    .D(net670),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[54] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3079_ (.RESET_B(net121),
    .D(net674),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[55] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3080_ (.RESET_B(net117),
    .D(net633),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[56] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3081_ (.RESET_B(net114),
    .D(net564),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3082_ (.RESET_B(net110),
    .D(_0273_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3083_ (.RESET_B(net106),
    .D(net620),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[59] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3084_ (.RESET_B(net102),
    .D(net591),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[60] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3085_ (.RESET_B(net98),
    .D(_0276_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[61] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _3086_ (.RESET_B(net94),
    .D(_0277_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3087_ (.RESET_B(net90),
    .D(net651),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[63] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3088_ (.RESET_B(net86),
    .D(net348),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[64] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3089_ (.RESET_B(net82),
    .D(_0280_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3090_ (.RESET_B(net78),
    .D(_0281_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[66] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3091_ (.RESET_B(net74),
    .D(net575),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[67] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3092_ (.RESET_B(net70),
    .D(_0283_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[68] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _3093_ (.RESET_B(net66),
    .D(_0284_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3094_ (.RESET_B(net62),
    .D(net668),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[70] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3095_ (.RESET_B(net58),
    .D(net560),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[71] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3096_ (.RESET_B(net54),
    .D(_0287_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3097_ (.RESET_B(net51),
    .D(net631),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[73] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3098_ (.RESET_B(net47),
    .D(net608),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[74] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3099_ (.RESET_B(net43),
    .D(_0290_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[75] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3100_ (.RESET_B(net39),
    .D(_0291_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3101_ (.RESET_B(net35),
    .D(net653),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[77] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3102_ (.RESET_B(net31),
    .D(net365),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[78] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3103_ (.RESET_B(net191),
    .D(_0294_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[79] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3104_ (.RESET_B(net183),
    .D(_0295_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[80] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3105_ (.RESET_B(net176),
    .D(net701),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[81] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _3106_ (.RESET_B(net168),
    .D(net679),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[82] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _3107_ (.RESET_B(net160),
    .D(_0298_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[83] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _3108_ (.RESET_B(net151),
    .D(net359),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[84] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _3109_ (.RESET_B(net143),
    .D(_0300_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[85] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _3110_ (.RESET_B(net135),
    .D(net369),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3111_ (.RESET_B(net127),
    .D(net355),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[87] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3112_ (.RESET_B(net119),
    .D(_0303_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3113_ (.RESET_B(net112),
    .D(net615),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[89] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3114_ (.RESET_B(net104),
    .D(_0305_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3115_ (.RESET_B(net96),
    .D(net569),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[91] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3116_ (.RESET_B(net88),
    .D(_0307_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[92] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3117_ (.RESET_B(net80),
    .D(net641),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[93] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3118_ (.RESET_B(net72),
    .D(net598),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[94] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3119_ (.RESET_B(net64),
    .D(_0310_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[95] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3120_ (.RESET_B(net56),
    .D(_0311_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[96] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3121_ (.RESET_B(net49),
    .D(_0312_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3122_ (.RESET_B(net41),
    .D(net556),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[98] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3123_ (.RESET_B(net33),
    .D(net363),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[99] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3124_ (.RESET_B(net187),
    .D(_0315_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3125_ (.RESET_B(net172),
    .D(net626),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[101] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3126_ (.RESET_B(net156),
    .D(net595),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[102] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3127_ (.RESET_B(net139),
    .D(_0318_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[103] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3128_ (.RESET_B(net123),
    .D(_0319_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3129_ (.RESET_B(net108),
    .D(net750),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[105] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3130_ (.RESET_B(net92),
    .D(net613),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[106] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3131_ (.RESET_B(net76),
    .D(_0322_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3132_ (.RESET_B(net60),
    .D(_0323_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3133_ (.RESET_B(net45),
    .D(net605),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[109] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3134_ (.RESET_B(net29),
    .D(net583),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[110] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3135_ (.RESET_B(net164),
    .D(_0326_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3136_ (.RESET_B(net131),
    .D(_0327_),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3137_ (.RESET_B(net100),
    .D(net341),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3138_ (.RESET_B(net68),
    .D(net718),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3139_ (.RESET_B(net37),
    .D(net663),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _3140_ (.RESET_B(net147),
    .D(_0331_),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3141_ (.RESET_B(net84),
    .D(net332),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3142_ (.RESET_B(net193),
    .D(net696),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3143_ (.RESET_B(net194),
    .D(_0334_),
    .Q(\ppwm_i.u_ppwm.data_o ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3144_ (.RESET_B(net523),
    .D(_0074_),
    .Q(\sdr_i.mac1.products_ff[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3145_ (.RESET_B(net523),
    .D(_0075_),
    .Q(\sdr_i.mac1.products_ff[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3146_ (.RESET_B(net523),
    .D(_0054_),
    .Q(\sdr_i.mac1.products_ff[17] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3147_ (.RESET_B(net523),
    .D(_0055_),
    .Q(\sdr_i.mac1.products_ff[18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3148_ (.RESET_B(net526),
    .D(_0040_),
    .Q(\sdr_i.mac1.products_ff[34] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3149_ (.RESET_B(net526),
    .D(_0041_),
    .Q(\sdr_i.mac1.products_ff[35] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3150_ (.RESET_B(net536),
    .D(_0042_),
    .Q(\sdr_i.mac1.products_ff[51] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3151_ (.RESET_B(net535),
    .D(_0043_),
    .Q(\sdr_i.mac1.products_ff[52] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3152_ (.RESET_B(net529),
    .D(_0058_),
    .Q(\sdr_i.mac1.products_ff[68] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _3153_ (.RESET_B(net529),
    .D(_0059_),
    .Q(\sdr_i.mac1.products_ff[69] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _3154_ (.RESET_B(net531),
    .D(_0048_),
    .Q(\sdr_i.mac1.products_ff[85] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _3155_ (.RESET_B(net531),
    .D(_0049_),
    .Q(\sdr_i.mac1.products_ff[86] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _3156_ (.RESET_B(net528),
    .D(_0050_),
    .Q(\sdr_i.mac1.products_ff[102] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _3157_ (.RESET_B(net528),
    .D(_0051_),
    .Q(\sdr_i.mac1.products_ff[103] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _3158_ (.RESET_B(net530),
    .D(_0052_),
    .Q(\sdr_i.mac1.products_ff[119] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3159_ (.RESET_B(net530),
    .D(_0053_),
    .Q(\sdr_i.mac1.products_ff[120] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3160_ (.RESET_B(net522),
    .D(_0072_),
    .Q(\sdr_i.mac1.products_ff[136] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3161_ (.RESET_B(net522),
    .D(_0073_),
    .Q(\sdr_i.mac1.products_ff[137] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3162_ (.RESET_B(net533),
    .D(net218),
    .Q(\sdr_i.mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3163_ (.RESET_B(net526),
    .D(net735),
    .Q(\sdr_i.mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3164_ (.RESET_B(net526),
    .D(net314),
    .Q(\sdr_i.mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3165_ (.RESET_B(net526),
    .D(net779),
    .Q(\sdr_i.mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3166_ (.RESET_B(net531),
    .D(net308),
    .Q(\sdr_i.mac1.sum_lvl1_ff[16] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3167_ (.RESET_B(net531),
    .D(net742),
    .Q(\sdr_i.mac1.sum_lvl1_ff[17] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3168_ (.RESET_B(net529),
    .D(net231),
    .Q(\sdr_i.mac1.sum_lvl1_ff[24] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3169_ (.RESET_B(net530),
    .D(net763),
    .Q(\sdr_i.mac1.sum_lvl1_ff[25] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _3170_ (.RESET_B(net195),
    .D(_0003_),
    .Q(\ppwm_i.u_ppwm.u_mem.state_q[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _3171_ (.RESET_B(net196),
    .D(_0004_),
    .Q(\ppwm_i.u_ppwm.mem_write_done ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3172_ (.RESET_B(net197),
    .D(net325),
    .Q(\ppwm_i.u_ppwm.u_mem.state_q[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3173_ (.RESET_B(net522),
    .D(net201),
    .Q(\sdr_i.mac1.sum_lvl1_ff[32] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3174_ (.RESET_B(net522),
    .D(net207),
    .Q(\sdr_i.mac1.sum_lvl1_ff[33] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3175_ (.RESET_B(net533),
    .D(net216),
    .Q(\sdr_i.mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3176_ (.RESET_B(net533),
    .D(net738),
    .Q(\sdr_i.mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3177_ (.RESET_B(net531),
    .D(net268),
    .Q(\sdr_i.mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _3178_ (.RESET_B(net531),
    .D(net747),
    .Q(\sdr_i.mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3179_ (.RESET_B(net524),
    .D(net203),
    .Q(\sdr_i.mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3180_ (.RESET_B(net522),
    .D(net206),
    .Q(\sdr_i.mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3181_ (.RESET_B(net526),
    .D(net306),
    .Q(\sdr_i.mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3182_ (.RESET_B(net533),
    .D(net745),
    .Q(\sdr_i.mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _3183_ (.RESET_B(net526),
    .D(net210),
    .Q(\sdr_i.mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3184_ (.RESET_B(net524),
    .D(net205),
    .Q(\sdr_i.mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3185_ (.RESET_B(net525),
    .D(net262),
    .Q(\sdr_i.mac1.total_sum[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3186_ (.RESET_B(net525),
    .D(net775),
    .Q(\sdr_i.mac1.total_sum[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3187_ (.RESET_B(net525),
    .D(net554),
    .Q(\sdr_i.total_sum1[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3188_ (.RESET_B(net544),
    .D(_0056_),
    .Q(\sdr_i.mac2.products_ff[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3189_ (.RESET_B(net545),
    .D(_0057_),
    .Q(\sdr_i.mac2.products_ff[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3190_ (.RESET_B(net546),
    .D(_0060_),
    .Q(\sdr_i.mac2.products_ff[17] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3191_ (.RESET_B(net546),
    .D(_0061_),
    .Q(\sdr_i.mac2.products_ff[18] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3192_ (.RESET_B(net540),
    .D(_0062_),
    .Q(\sdr_i.mac2.products_ff[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3193_ (.RESET_B(net539),
    .D(_0063_),
    .Q(\sdr_i.mac2.products_ff[35] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3194_ (.RESET_B(net540),
    .D(_0064_),
    .Q(\sdr_i.mac2.products_ff[51] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3195_ (.RESET_B(net540),
    .D(_0065_),
    .Q(\sdr_i.mac2.products_ff[52] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3196_ (.RESET_B(net542),
    .D(_0046_),
    .Q(\sdr_i.mac2.products_ff[68] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3197_ (.RESET_B(net543),
    .D(_0047_),
    .Q(\sdr_i.mac2.products_ff[69] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3198_ (.RESET_B(net543),
    .D(_0066_),
    .Q(\sdr_i.mac2.products_ff[85] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3199_ (.RESET_B(net542),
    .D(_0067_),
    .Q(\sdr_i.mac2.products_ff[86] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3200_ (.RESET_B(net537),
    .D(_0044_),
    .Q(\sdr_i.mac2.products_ff[102] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3201_ (.RESET_B(net537),
    .D(_0045_),
    .Q(\sdr_i.mac2.products_ff[103] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3202_ (.RESET_B(net538),
    .D(_0068_),
    .Q(\sdr_i.mac2.products_ff[119] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3203_ (.RESET_B(net538),
    .D(_0069_),
    .Q(\sdr_i.mac2.products_ff[120] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3204_ (.RESET_B(net533),
    .D(_0070_),
    .Q(\sdr_i.mac2.products_ff[136] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3205_ (.RESET_B(net542),
    .D(_0071_),
    .Q(\sdr_i.mac2.products_ff[137] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3206_ (.RESET_B(net544),
    .D(net255),
    .Q(\sdr_i.mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3207_ (.RESET_B(net544),
    .D(net758),
    .Q(\sdr_i.mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3208_ (.RESET_B(net540),
    .D(net214),
    .Q(\sdr_i.mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3209_ (.RESET_B(net544),
    .D(net730),
    .Q(\sdr_i.mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3210_ (.RESET_B(net542),
    .D(net266),
    .Q(\sdr_i.mac2.sum_lvl1_ff[16] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3211_ (.RESET_B(net542),
    .D(net756),
    .Q(\sdr_i.mac2.sum_lvl1_ff[17] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3212_ (.RESET_B(net541),
    .D(net258),
    .Q(\sdr_i.mac2.sum_lvl1_ff[24] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3213_ (.RESET_B(net541),
    .D(net740),
    .Q(\sdr_i.mac2.sum_lvl1_ff[25] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3214_ (.RESET_B(net532),
    .D(net202),
    .Q(\sdr_i.mac2.sum_lvl1_ff[32] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3215_ (.RESET_B(net536),
    .D(net212),
    .Q(\sdr_i.mac2.sum_lvl1_ff[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3216_ (.RESET_B(net544),
    .D(net292),
    .Q(\sdr_i.mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3217_ (.RESET_B(net544),
    .D(net732),
    .Q(\sdr_i.mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3218_ (.RESET_B(net536),
    .D(net270),
    .Q(\sdr_i.mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3219_ (.RESET_B(net544),
    .D(net724),
    .Q(\sdr_i.mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3220_ (.RESET_B(net198),
    .D(net760),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3221_ (.RESET_B(net199),
    .D(net319),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3222_ (.RESET_B(net200),
    .D(_0002_),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3223_ (.RESET_B(net532),
    .D(net211),
    .Q(\sdr_i.mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3224_ (.RESET_B(net536),
    .D(net204),
    .Q(\sdr_i.mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3225_ (.RESET_B(net536),
    .D(net298),
    .Q(\sdr_i.mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _3226_ (.RESET_B(net537),
    .D(net765),
    .Q(\sdr_i.mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3227_ (.RESET_B(net532),
    .D(net208),
    .Q(\sdr_i.mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3228_ (.RESET_B(net526),
    .D(net209),
    .Q(\sdr_i.mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3229_ (.RESET_B(net525),
    .D(net260),
    .Q(\sdr_i.mac2.total_sum[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3230_ (.RESET_B(net525),
    .D(net783),
    .Q(\sdr_i.mac2.total_sum[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3231_ (.RESET_B(net525),
    .D(net603),
    .Q(\sdr_i.mac2.total_sum[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_tiehi _3134__29 (.L_HI(net29));
 sg13g2_tiehi _3060__30 (.L_HI(net30));
 sg13g2_tiehi _3102__31 (.L_HI(net31));
 sg13g2_tiehi _3059__32 (.L_HI(net32));
 sg13g2_tiehi _3123__33 (.L_HI(net33));
 sg13g2_tiehi _3058__34 (.L_HI(net34));
 sg13g2_tiehi _3101__35 (.L_HI(net35));
 sg13g2_tiehi _3057__36 (.L_HI(net36));
 sg13g2_tiehi _3139__37 (.L_HI(net37));
 sg13g2_tiehi _3056__38 (.L_HI(net38));
 sg13g2_tiehi _3100__39 (.L_HI(net39));
 sg13g2_tiehi _3055__40 (.L_HI(net40));
 sg13g2_tiehi _3122__41 (.L_HI(net41));
 sg13g2_tiehi _3054__42 (.L_HI(net42));
 sg13g2_tiehi _3099__43 (.L_HI(net43));
 sg13g2_tiehi _3053__44 (.L_HI(net44));
 sg13g2_tiehi _3133__45 (.L_HI(net45));
 sg13g2_tiehi _3052__46 (.L_HI(net46));
 sg13g2_tiehi _3098__47 (.L_HI(net47));
 sg13g2_tiehi _3051__48 (.L_HI(net48));
 sg13g2_tiehi _3121__49 (.L_HI(net49));
 sg13g2_tiehi _3050__50 (.L_HI(net50));
 sg13g2_tiehi _3097__51 (.L_HI(net51));
 sg13g2_tiehi _3049__52 (.L_HI(net52));
 sg13g2_tiehi _3048__53 (.L_HI(net53));
 sg13g2_tiehi _3096__54 (.L_HI(net54));
 sg13g2_tiehi _3047__55 (.L_HI(net55));
 sg13g2_tiehi _3120__56 (.L_HI(net56));
 sg13g2_tiehi _3046__57 (.L_HI(net57));
 sg13g2_tiehi _3095__58 (.L_HI(net58));
 sg13g2_tiehi _3045__59 (.L_HI(net59));
 sg13g2_tiehi _3132__60 (.L_HI(net60));
 sg13g2_tiehi _3044__61 (.L_HI(net61));
 sg13g2_tiehi _3094__62 (.L_HI(net62));
 sg13g2_tiehi _3043__63 (.L_HI(net63));
 sg13g2_tiehi _3119__64 (.L_HI(net64));
 sg13g2_tiehi _3042__65 (.L_HI(net65));
 sg13g2_tiehi _3093__66 (.L_HI(net66));
 sg13g2_tiehi _3041__67 (.L_HI(net67));
 sg13g2_tiehi _3138__68 (.L_HI(net68));
 sg13g2_tiehi _3040__69 (.L_HI(net69));
 sg13g2_tiehi _3092__70 (.L_HI(net70));
 sg13g2_tiehi _3039__71 (.L_HI(net71));
 sg13g2_tiehi _3118__72 (.L_HI(net72));
 sg13g2_tiehi _3038__73 (.L_HI(net73));
 sg13g2_tiehi _3091__74 (.L_HI(net74));
 sg13g2_tiehi _3037__75 (.L_HI(net75));
 sg13g2_tiehi _3131__76 (.L_HI(net76));
 sg13g2_tiehi _3036__77 (.L_HI(net77));
 sg13g2_tiehi _3090__78 (.L_HI(net78));
 sg13g2_tiehi _3035__79 (.L_HI(net79));
 sg13g2_tiehi _3117__80 (.L_HI(net80));
 sg13g2_tiehi _3034__81 (.L_HI(net81));
 sg13g2_tiehi _3089__82 (.L_HI(net82));
 sg13g2_tiehi _3033__83 (.L_HI(net83));
 sg13g2_tiehi _3141__84 (.L_HI(net84));
 sg13g2_tiehi _3032__85 (.L_HI(net85));
 sg13g2_tiehi _3088__86 (.L_HI(net86));
 sg13g2_tiehi _3031__87 (.L_HI(net87));
 sg13g2_tiehi _3116__88 (.L_HI(net88));
 sg13g2_tiehi _3030__89 (.L_HI(net89));
 sg13g2_tiehi _3087__90 (.L_HI(net90));
 sg13g2_tiehi _3029__91 (.L_HI(net91));
 sg13g2_tiehi _3130__92 (.L_HI(net92));
 sg13g2_tiehi _3028__93 (.L_HI(net93));
 sg13g2_tiehi _3086__94 (.L_HI(net94));
 sg13g2_tiehi _3027__95 (.L_HI(net95));
 sg13g2_tiehi _3115__96 (.L_HI(net96));
 sg13g2_tiehi _3026__97 (.L_HI(net97));
 sg13g2_tiehi _3085__98 (.L_HI(net98));
 sg13g2_tiehi _3025__99 (.L_HI(net99));
 sg13g2_tiehi _3137__100 (.L_HI(net100));
 sg13g2_tiehi _3024__101 (.L_HI(net101));
 sg13g2_tiehi _3084__102 (.L_HI(net102));
 sg13g2_tiehi _3023__103 (.L_HI(net103));
 sg13g2_tiehi _3114__104 (.L_HI(net104));
 sg13g2_tiehi _3022__105 (.L_HI(net105));
 sg13g2_tiehi _3083__106 (.L_HI(net106));
 sg13g2_tiehi _3021__107 (.L_HI(net107));
 sg13g2_tiehi _3129__108 (.L_HI(net108));
 sg13g2_tiehi _3020__109 (.L_HI(net109));
 sg13g2_tiehi _3082__110 (.L_HI(net110));
 sg13g2_tiehi _3019__111 (.L_HI(net111));
 sg13g2_tiehi _3113__112 (.L_HI(net112));
 sg13g2_tiehi _3018__113 (.L_HI(net113));
 sg13g2_tiehi _3081__114 (.L_HI(net114));
 sg13g2_tiehi _3017__115 (.L_HI(net115));
 sg13g2_tiehi _3016__116 (.L_HI(net116));
 sg13g2_tiehi _3080__117 (.L_HI(net117));
 sg13g2_tiehi _3015__118 (.L_HI(net118));
 sg13g2_tiehi _3112__119 (.L_HI(net119));
 sg13g2_tiehi _3014__120 (.L_HI(net120));
 sg13g2_tiehi _3079__121 (.L_HI(net121));
 sg13g2_tiehi _3013__122 (.L_HI(net122));
 sg13g2_tiehi _3128__123 (.L_HI(net123));
 sg13g2_tiehi _3012__124 (.L_HI(net124));
 sg13g2_tiehi _3078__125 (.L_HI(net125));
 sg13g2_tiehi _3011__126 (.L_HI(net126));
 sg13g2_tiehi _3111__127 (.L_HI(net127));
 sg13g2_tiehi _3010__128 (.L_HI(net128));
 sg13g2_tiehi _3077__129 (.L_HI(net129));
 sg13g2_tiehi _3009__130 (.L_HI(net130));
 sg13g2_tiehi _3136__131 (.L_HI(net131));
 sg13g2_tiehi _3008__132 (.L_HI(net132));
 sg13g2_tiehi _3076__133 (.L_HI(net133));
 sg13g2_tiehi _3007__134 (.L_HI(net134));
 sg13g2_tiehi _3110__135 (.L_HI(net135));
 sg13g2_tiehi _3006__136 (.L_HI(net136));
 sg13g2_tiehi _3075__137 (.L_HI(net137));
 sg13g2_tiehi _3005__138 (.L_HI(net138));
 sg13g2_tiehi _3127__139 (.L_HI(net139));
 sg13g2_tiehi _3004__140 (.L_HI(net140));
 sg13g2_tiehi _3074__141 (.L_HI(net141));
 sg13g2_tiehi _3003__142 (.L_HI(net142));
 sg13g2_tiehi _3109__143 (.L_HI(net143));
 sg13g2_tiehi _3002__144 (.L_HI(net144));
 sg13g2_tiehi _3073__145 (.L_HI(net145));
 sg13g2_tiehi _3001__146 (.L_HI(net146));
 sg13g2_tiehi _3140__147 (.L_HI(net147));
 sg13g2_tiehi _3000__148 (.L_HI(net148));
 sg13g2_tiehi _3072__149 (.L_HI(net149));
 sg13g2_tiehi _2999__150 (.L_HI(net150));
 sg13g2_tiehi _3108__151 (.L_HI(net151));
 sg13g2_tiehi _2998__152 (.L_HI(net152));
 sg13g2_tiehi _2997__153 (.L_HI(net153));
 sg13g2_tiehi _3071__154 (.L_HI(net154));
 sg13g2_tiehi _2996__155 (.L_HI(net155));
 sg13g2_tiehi _3126__156 (.L_HI(net156));
 sg13g2_tiehi _2995__157 (.L_HI(net157));
 sg13g2_tiehi _3070__158 (.L_HI(net158));
 sg13g2_tiehi _2994__159 (.L_HI(net159));
 sg13g2_tiehi _3107__160 (.L_HI(net160));
 sg13g2_tiehi _2993__161 (.L_HI(net161));
 sg13g2_tiehi _3069__162 (.L_HI(net162));
 sg13g2_tiehi _2992__163 (.L_HI(net163));
 sg13g2_tiehi _3135__164 (.L_HI(net164));
 sg13g2_tiehi _2991__165 (.L_HI(net165));
 sg13g2_tiehi _3068__166 (.L_HI(net166));
 sg13g2_tiehi _2990__167 (.L_HI(net167));
 sg13g2_tiehi _3106__168 (.L_HI(net168));
 sg13g2_tiehi _2989__169 (.L_HI(net169));
 sg13g2_tiehi _3067__170 (.L_HI(net170));
 sg13g2_tiehi _2988__171 (.L_HI(net171));
 sg13g2_tiehi _3125__172 (.L_HI(net172));
 sg13g2_tiehi _2987__173 (.L_HI(net173));
 sg13g2_tiehi _3066__174 (.L_HI(net174));
 sg13g2_tiehi _2986__175 (.L_HI(net175));
 sg13g2_tiehi _3105__176 (.L_HI(net176));
 sg13g2_tiehi _2985__177 (.L_HI(net177));
 sg13g2_tiehi _3065__178 (.L_HI(net178));
 sg13g2_tiehi _2984__179 (.L_HI(net179));
 sg13g2_tiehi _2983__180 (.L_HI(net180));
 sg13g2_tiehi _3064__181 (.L_HI(net181));
 sg13g2_tiehi _2982__182 (.L_HI(net182));
 sg13g2_tiehi _3104__183 (.L_HI(net183));
 sg13g2_tiehi _2981__184 (.L_HI(net184));
 sg13g2_tiehi _3063__185 (.L_HI(net185));
 sg13g2_tiehi _2980__186 (.L_HI(net186));
 sg13g2_tiehi _3124__187 (.L_HI(net187));
 sg13g2_tiehi _2979__188 (.L_HI(net188));
 sg13g2_tiehi _3062__189 (.L_HI(net189));
 sg13g2_tiehi _2978__190 (.L_HI(net190));
 sg13g2_tiehi _3103__191 (.L_HI(net191));
 sg13g2_tiehi _2977__192 (.L_HI(net192));
 sg13g2_tiehi _3142__193 (.L_HI(net193));
 sg13g2_tiehi _3143__194 (.L_HI(net194));
 sg13g2_tiehi _3170__195 (.L_HI(net195));
 sg13g2_tiehi _3171__196 (.L_HI(net196));
 sg13g2_tiehi _3172__197 (.L_HI(net197));
 sg13g2_tiehi _3220__198 (.L_HI(net198));
 sg13g2_tiehi _3221__199 (.L_HI(net199));
 sg13g2_tiehi _3222__200 (.L_HI(net200));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tiny_wrapper_17 (.L_LO(net17));
 sg13g2_tielo tiny_wrapper_18 (.L_LO(net18));
 sg13g2_tielo tiny_wrapper_19 (.L_LO(net19));
 sg13g2_tielo tiny_wrapper_20 (.L_LO(net20));
 sg13g2_tielo tiny_wrapper_21 (.L_LO(net21));
 sg13g2_tielo tiny_wrapper_22 (.L_LO(net22));
 sg13g2_tielo tiny_wrapper_23 (.L_LO(net23));
 sg13g2_tielo tiny_wrapper_24 (.L_LO(net24));
 sg13g2_tielo tiny_wrapper_25 (.L_LO(net25));
 sg13g2_tielo tiny_wrapper_26 (.L_LO(net26));
 sg13g2_tielo tiny_wrapper_27 (.L_LO(net27));
 sg13g2_tiehi _3061__28 (.L_HI(net28));
 sg13g2_buf_1 _3417_ (.A(net548),
    .X(net4));
 sg13g2_buf_1 _3418_ (.A(net549),
    .X(net5));
 sg13g2_buf_1 _3419_ (.A(net549),
    .X(net6));
 sg13g2_buf_1 _3420_ (.A(net549),
    .X(net7));
 sg13g2_buf_1 _3421_ (.A(net549),
    .X(net8));
 sg13g2_buf_1 _3422_ (.A(net548),
    .X(net9));
 sg13g2_buf_1 _3423_ (.A(net548),
    .X(net10));
 sg13g2_buf_1 _3424_ (.A(net549),
    .X(net11));
 sg13g2_buf_8 fanout370 (.A(_0861_),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(net373),
    .X(net371));
 sg13g2_buf_1 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(_0683_),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(_0860_),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(_0676_),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(_0673_),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(_0684_),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(_0684_),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(_0653_),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(_0671_),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net382),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(_0639_),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(_0639_),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(_0349_),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net388),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_1 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_0348_),
    .X(net389));
 sg13g2_buf_8 fanout390 (.A(_0336_),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(_0335_),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(_0335_),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(_1338_),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(_1325_),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(_1310_),
    .X(net396));
 sg13g2_buf_8 fanout397 (.A(_1310_),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net400),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(_1296_),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(_1295_),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_1295_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(_1352_),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_1346_),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net411),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(_0477_),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net415),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(net415),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net420),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net418),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(net420),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net424),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net422),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(\ppwm_i.rst_n ),
    .X(net424));
 sg13g2_buf_8 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net434),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net434),
    .X(net428));
 sg13g2_buf_1 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(net434),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net433),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net433),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(\ppwm_i.rst_n ),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(net437),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(\ppwm_i.rst_n ),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(_1283_),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(_1283_),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net441),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(_1283_),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(_1282_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_1282_),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net446),
    .X(net444));
 sg13g2_buf_1 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_1 fanout446 (.A(_1282_),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net449),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(_1280_),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net452),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(_1276_),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_1276_),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(net459),
    .X(net455));
 sg13g2_buf_1 fanout456 (.A(net459),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(net459),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(_1266_),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(_1233_),
    .X(net460));
 sg13g2_buf_1 fanout461 (.A(_1233_),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(net463),
    .X(net462));
 sg13g2_buf_8 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(net470),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(net467),
    .X(net465));
 sg13g2_buf_8 fanout466 (.A(net467),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net470),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(net470),
    .X(net468));
 sg13g2_buf_1 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net501),
    .X(net470));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_8 fanout472 (.A(net501),
    .X(net472));
 sg13g2_buf_8 fanout473 (.A(net476),
    .X(net473));
 sg13g2_buf_8 fanout474 (.A(net476),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_8 fanout476 (.A(net480),
    .X(net476));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_8 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net501),
    .X(net480));
 sg13g2_buf_8 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_8 fanout482 (.A(net486),
    .X(net482));
 sg13g2_buf_8 fanout483 (.A(net486),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net486),
    .X(net484));
 sg13g2_buf_8 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_8 fanout486 (.A(net501),
    .X(net486));
 sg13g2_buf_8 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net490),
    .X(net488));
 sg13g2_buf_8 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net500),
    .X(net490));
 sg13g2_buf_8 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_8 fanout492 (.A(net496),
    .X(net492));
 sg13g2_buf_8 fanout493 (.A(net496),
    .X(net493));
 sg13g2_buf_1 fanout494 (.A(net496),
    .X(net494));
 sg13g2_buf_8 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_8 fanout496 (.A(net500),
    .X(net496));
 sg13g2_buf_8 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_8 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_8 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_8 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_8 fanout501 (.A(net690),
    .X(net501));
 sg13g2_buf_8 fanout502 (.A(net836),
    .X(net502));
 sg13g2_buf_8 fanout503 (.A(net833),
    .X(net503));
 sg13g2_buf_8 fanout504 (.A(net830),
    .X(net504));
 sg13g2_buf_8 fanout505 (.A(net838),
    .X(net505));
 sg13g2_buf_8 fanout506 (.A(net770),
    .X(net506));
 sg13g2_buf_8 fanout507 (.A(net831),
    .X(net507));
 sg13g2_buf_8 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_8 fanout509 (.A(net835),
    .X(net509));
 sg13g2_buf_8 fanout510 (.A(net513),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net513),
    .X(net511));
 sg13g2_buf_8 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_8 fanout513 (.A(net827),
    .X(net513));
 sg13g2_buf_8 fanout514 (.A(net516),
    .X(net514));
 sg13g2_buf_8 fanout515 (.A(net825),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(\ppwm_i.u_ppwm.pc[1] ),
    .X(net516));
 sg13g2_buf_8 fanout517 (.A(net519),
    .X(net517));
 sg13g2_buf_8 fanout518 (.A(net788),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(\ppwm_i.u_ppwm.pc[0] ),
    .X(net519));
 sg13g2_buf_8 fanout520 (.A(net565),
    .X(net520));
 sg13g2_buf_8 fanout521 (.A(net524),
    .X(net521));
 sg13g2_buf_8 fanout522 (.A(net524),
    .X(net522));
 sg13g2_buf_8 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_8 fanout524 (.A(net547),
    .X(net524));
 sg13g2_buf_8 fanout525 (.A(net527),
    .X(net525));
 sg13g2_buf_8 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_8 fanout527 (.A(net547),
    .X(net527));
 sg13g2_buf_8 fanout528 (.A(net530),
    .X(net528));
 sg13g2_buf_8 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_8 fanout530 (.A(net534),
    .X(net530));
 sg13g2_buf_8 fanout531 (.A(net534),
    .X(net531));
 sg13g2_buf_8 fanout532 (.A(net534),
    .X(net532));
 sg13g2_buf_8 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_8 fanout534 (.A(net547),
    .X(net534));
 sg13g2_buf_8 fanout535 (.A(net537),
    .X(net535));
 sg13g2_buf_8 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_8 fanout537 (.A(net541),
    .X(net537));
 sg13g2_buf_8 fanout538 (.A(net540),
    .X(net538));
 sg13g2_buf_8 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_8 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_8 fanout541 (.A(net547),
    .X(net541));
 sg13g2_buf_8 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net547),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(net546),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_8 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(rst_n_sdr),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net1),
    .X(net548));
 sg13g2_buf_1 fanout549 (.A(net1),
    .X(net549));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[2]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[7]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[3]));
 sg13g2_tielo tiny_wrapper_16 (.L_LO(net16));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_46_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_19_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_22_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_29_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\sdr_i.mac1.products_ff[136] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold2 (.A(\sdr_i.mac2.products_ff[136] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold3 (.A(\sdr_i.mac1.sum_lvl1_ff[32] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold4 (.A(\sdr_i.mac2.sum_lvl1_ff[33] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold5 (.A(\sdr_i.mac1.sum_lvl2_ff[9] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sdr_i.mac1.sum_lvl1_ff[33] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold7 (.A(\sdr_i.mac1.products_ff[137] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold8 (.A(\sdr_i.mac2.sum_lvl2_ff[8] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold9 (.A(\sdr_i.mac2.sum_lvl2_ff[9] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold10 (.A(\sdr_i.mac1.sum_lvl2_ff[8] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold11 (.A(\sdr_i.mac2.sum_lvl1_ff[32] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold12 (.A(\sdr_i.mac2.products_ff[137] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold13 (.A(\sdr_i.mac2.products_ff[51] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0034_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold15 (.A(\sdr_i.mac1.sum_lvl1_ff[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0023_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold17 (.A(\sdr_i.mac1.products_ff[17] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0015_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold19 (.A(\sdr_i.DP_3.matrix[10] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold20 (.A(\sdr_i.DP_1.matrix[10] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold21 (.A(\sdr_i.DP_1.matrix[64] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold22 (.A(\sdr_i.DP_4.matrix[10] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold23 (.A(\sdr_i.DP_3.matrix[1] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold24 (.A(\sdr_i.DP_2.matrix[73] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold25 (.A(\sdr_i.DP_2.matrix[55] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold26 (.A(\sdr_i.DP_2.matrix[28] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold27 (.A(\sdr_i.DP_4.matrix[55] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold28 (.A(\sdr_i.DP_4.matrix[28] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold29 (.A(\sdr_i.DP_1.matrix[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold30 (.A(\sdr_i.mac1.products_ff[102] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0021_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold32 (.A(\sdr_i.DP_1.matrix[73] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold33 (.A(\sdr_i.DP_2.matrix[64] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold34 (.A(\sdr_i.DP_4.matrix[19] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold35 (.A(\sdr_i.DP_1.matrix[28] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold36 (.A(\sdr_i.DP_3.matrix[28] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold37 (.A(\sdr_i.DP_2.matrix[10] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold38 (.A(\sdr_i.DP_3.matrix[73] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold39 (.A(\sdr_i.DP_4.matrix[46] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold40 (.A(\sdr_i.DP_1.matrix[19] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold41 (.A(\sdr_i.DP_2.matrix[19] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold42 (.A(\sdr_i.DP_3.matrix[55] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold43 (.A(\sdr_i.DP_3.matrix[46] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold44 (.A(\sdr_i.DP_1.matrix[46] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold45 (.A(\sdr_i.DP_3.matrix[19] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold46 (.A(\sdr_i.DP_4.matrix[73] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold47 (.A(\sdr_i.DP_4.matrix[1] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold48 (.A(\sdr_i.DP_2.matrix[46] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold49 (.A(\sdr_i.DP_2.matrix[37] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold50 (.A(\sdr_i.DP_3.matrix[64] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold51 (.A(\sdr_i.DP_4.matrix[37] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold52 (.A(\sdr_i.DP_2.matrix[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold53 (.A(\sdr_i.DP_4.matrix[64] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold54 (.A(\sdr_i.mac2.products_ff[0] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0032_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold56 (.A(\sdr_i.DP_3.matrix[37] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold57 (.A(\sdr_i.mac2.products_ff[119] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0038_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold59 (.A(\sdr_i.mac2.sum_lvl3_ff[0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0007_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold61 (.A(\sdr_i.mac1.sum_lvl3_ff[0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0030_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold63 (.A(\sdr_i.DP_1.matrix[37] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold64 (.A(\sdr_i.DP_1.matrix[55] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold65 (.A(\sdr_i.mac2.products_ff[68] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0036_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold67 (.A(\sdr_i.mac1.sum_lvl1_ff[16] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0025_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold69 (.A(\sdr_i.mac2.sum_lvl1_ff[24] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0011_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold71 (.A(\sdr_i.DP_3.matrix[63] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold72 (.A(\sdr_i.DP_1.matrix[72] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold73 (.A(\sdr_i.DP_1.matrix[18] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold74 (.A(\sdr_i.DP_2.matrix[9] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold75 (.A(\sdr_i.DP_2.matrix[27] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold76 (.A(\sdr_i.DP_1.matrix[0] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold77 (.A(\sdr_i.DP_4.matrix[36] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold78 (.A(\sdr_i.DP_3.matrix[27] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold79 (.A(\sdr_i.DP_1.matrix[45] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold80 (.A(\sdr_i.DP_4.matrix[0] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold81 (.A(\sdr_i.DP_2.matrix[18] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold82 (.A(\sdr_i.DP_3.matrix[54] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold83 (.A(\sdr_i.DP_4.matrix[54] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold84 (.A(\sdr_i.DP_2.matrix[72] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold85 (.A(\sdr_i.DP_1.matrix[9] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold86 (.A(\sdr_i.DP_2.matrix[63] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold87 (.A(\sdr_i.DP_2.matrix[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold88 (.A(\sdr_i.DP_3.matrix[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold89 (.A(\sdr_i.DP_1.matrix[63] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold90 (.A(\sdr_i.DP_3.matrix[9] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold91 (.A(\sdr_i.mac2.sum_lvl1_ff[0] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0013_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold93 (.A(\sdr_i.DP_3.matrix[18] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold94 (.A(\sdr_i.DP_4.matrix[18] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold95 (.A(\sdr_i.DP_1.matrix[36] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold96 (.A(\sdr_i.DP_4.matrix[9] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold97 (.A(\sdr_i.mac2.sum_lvl2_ff[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0009_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold99 (.A(\sdr_i.DP_3.matrix[36] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold100 (.A(\sdr_i.DP_4.matrix[45] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold101 (.A(\sdr_i.DP_4.matrix[27] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold102 (.A(\sdr_i.DP_4.matrix[63] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold103 (.A(\sdr_i.DP_1.matrix[54] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold104 (.A(\sdr_i.DP_1.matrix[27] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold105 (.A(\sdr_i.mac1.sum_lvl2_ff[0] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0027_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold107 (.A(\sdr_i.mac1.products_ff[85] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0019_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold109 (.A(\sdr_i.DP_3.matrix[45] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold110 (.A(\sdr_i.DP_2.matrix[54] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold111 (.A(\sdr_i.DP_2.matrix[45] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold112 (.A(\sdr_i.DP_2.matrix[36] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold113 (.A(\sdr_i.mac1.products_ff[34] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0017_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold115 (.A(\sdr_i.DP_4.matrix[72] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold116 (.A(\sdr_i.DP_3.matrix[72] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ppwm_i.u_ppwm.u_ex.state_q[1] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0372_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0001_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ppwm_i.u_ppwm.global_counter[6] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0154_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0168_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ppwm_i.u_ppwm.u_mem.state_q[0] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0005_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ppwm_i.u_ppwm.period_start ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0148_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ppwm_i.u_ppwm.global_counter[19] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0167_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold131 (.A(_1076_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0332_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold133 (.A(\ppwm_i.u_ppwm.global_counter[5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0153_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ppwm_i.u_ppwm.global_counter[9] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0157_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0216_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold139 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold140 (.A(_1069_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0328_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold142 (.A(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ppwm_i.u_ppwm.u_mem.memory[1] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0215_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ppwm_i.u_ppwm.u_mem.memory[32] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0246_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0279_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ppwm_i.u_ppwm.u_ex.cmp_flag_q ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0550_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0193_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ppwm_i.u_ppwm.u_mem.memory[17] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0231_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0302_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0258_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ppwm_i.u_ppwm.u_mem.memory[85] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0299_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold160 (.A(\ppwm_i.u_ppwm.u_mem.memory[31] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0245_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0314_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ppwm_i.u_ppwm.u_mem.memory[79] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0293_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0265_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ppwm_i.u_ppwm.u_mem.memory[87] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0301_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold170 (.A(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0241_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold172 (.A(\sdr_i.mac1.sum_lvl3_ff[3] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0413_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0029_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold175 (.A(\ppwm_i.u_ppwm.u_mem.memory[99] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0313_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold177 (.A(\ppwm_i.u_ppwm.global_counter[10] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0158_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0286_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0223_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0272_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold185 (.A(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0506_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0188_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold188 (.A(\ppwm_i.u_ppwm.u_mem.memory[92] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0306_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0262_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ppwm_i.u_ppwm.global_counter[15] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0163_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold194 (.A(\ppwm_i.u_ppwm.u_mem.memory[68] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0282_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0244_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold198 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0169_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0175_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0325_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0250_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold206 (.A(\ppwm_i.u_ppwm.u_mem.memory[25] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0239_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ppwm_i.u_ppwm.u_mem.memory[15] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0229_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold210 (.A(\ppwm_i.u_ppwm.u_mem.memory[61] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0275_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold212 (.A(\ppwm_i.u_ppwm.u_mem.memory[46] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0260_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold214 (.A(\ppwm_i.u_ppwm.u_mem.memory[103] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0317_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ppwm_i.u_ppwm.u_mem.memory[28] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold217 (.A(\ppwm_i.u_ppwm.u_mem.memory[95] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0309_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold219 (.A(\ppwm_i.u_ppwm.u_mem.memory[24] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0238_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold221 (.A(\sdr_i.mac2.sum_lvl3_ff[3] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0417_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0006_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold224 (.A(\ppwm_i.u_ppwm.u_mem.memory[110] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0324_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold227 (.A(\ppwm_i.u_ppwm.u_mem.memory[75] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0289_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold229 (.A(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0227_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ppwm_i.u_ppwm.u_mem.memory[45] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold232 (.A(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0321_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold234 (.A(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0304_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold236 (.A(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0237_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold239 (.A(\ppwm_i.u_ppwm.u_mem.memory[60] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0274_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold241 (.A(\ppwm_i.u_ppwm.u_mem.memory[22] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0236_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold243 (.A(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0234_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold245 (.A(\ppwm_i.u_ppwm.u_mem.memory[102] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0316_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold247 (.A(\ppwm_i.u_ppwm.u_mem.memory[109] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold248 (.A(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0220_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold250 (.A(\ppwm_i.u_ppwm.u_mem.memory[74] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0288_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold252 (.A(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0271_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold254 (.A(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold255 (.A(\ppwm_i.u_ppwm.u_mem.memory[96] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold256 (.A(\ppwm_i.u_ppwm.u_mem.memory[29] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold257 (.A(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold258 (.A(\ppwm_i.u_ppwm.u_mem.memory[49] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold259 (.A(\ppwm_i.u_ppwm.u_mem.memory[50] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold260 (.A(\ppwm_i.u_ppwm.u_mem.memory[94] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0308_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold262 (.A(\ppwm_i.u_ppwm.u_mem.memory[10] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold263 (.A(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0252_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold265 (.A(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold266 (.A(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold267 (.A(\ppwm_i.u_ppwm.u_mem.memory[11] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0225_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold269 (.A(\ppwm_i.u_ppwm.u_mem.memory[101] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold270 (.A(\ppwm_i.u_ppwm.u_mem.memory[63] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0278_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold272 (.A(\ppwm_i.u_ppwm.u_mem.memory[77] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0292_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold274 (.A(\ppwm_i.u_ppwm.global_counter[7] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0155_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold276 (.A(\ppwm_i.u_ppwm.u_mem.memory[4] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold277 (.A(\ppwm_i.u_ppwm.u_mem.memory[52] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0267_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold279 (.A(\ppwm_i.u_ppwm.u_mem.memory[66] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold280 (.A(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold281 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold282 (.A(_1074_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0330_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold284 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0174_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold286 (.A(\ppwm_i.u_ppwm.u_mem.memory[14] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold287 (.A(\ppwm_i.u_ppwm.u_mem.memory[70] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0285_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold289 (.A(\ppwm_i.u_ppwm.u_mem.memory[54] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0269_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold291 (.A(\ppwm_i.u_ppwm.u_mem.memory[67] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold292 (.A(\ppwm_i.u_ppwm.u_mem.memory[93] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold293 (.A(\ppwm_i.u_ppwm.u_mem.memory[56] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0270_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold295 (.A(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0248_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold297 (.A(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold298 (.A(\ppwm_i.u_ppwm.u_mem.memory[83] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0297_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold300 (.A(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold301 (.A(\ppwm_i.u_ppwm.u_mem.memory[84] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold302 (.A(\ppwm_i.u_ppwm.u_mem.memory[42] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0257_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold304 (.A(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0219_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold306 (.A(\ppwm_i.u_ppwm.u_mem.memory[12] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold307 (.A(\ppwm_i.u_ppwm.u_mem.memory[89] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold308 (.A(\ppwm_i.u_ppwm.u_mem.memory[33] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0247_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold310 (.A(\ppwm_i.u_ppwm.u_mem.state_q[2] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold311 (.A(\ppwm_i.u_ppwm.u_mem.memory[26] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold312 (.A(\ppwm_i.u_ppwm.u_mem.memory[7] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0222_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold314 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[6] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1079_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0333_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold317 (.A(\ppwm_i.u_ppwm.u_mem.memory[18] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold318 (.A(\ppwm_i.u_ppwm.u_mem.memory[39] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold319 (.A(\ppwm_i.u_ppwm.u_mem.memory[40] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold320 (.A(\ppwm_i.u_ppwm.u_mem.memory[81] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0296_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold322 (.A(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold323 (.A(\ppwm_i.u_ppwm.u_mem.memory[47] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold324 (.A(\ppwm_i.u_ppwm.u_mem.memory[73] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold325 (.A(\ppwm_i.u_ppwm.u_mem.memory[19] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold326 (.A(\ppwm_i.u_ppwm.u_mem.memory[80] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold327 (.A(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0498_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0179_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold330 (.A(\ppwm_i.u_ppwm.global_counter[2] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0150_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold332 (.A(\ppwm_i.u_ppwm.polarity ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0194_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold334 (.A(\ppwm_i.u_ppwm.u_mem.memory[35] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold335 (.A(\ppwm_i.u_ppwm.mem_write_done ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold336 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[2] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold337 (.A(_1071_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0329_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold339 (.A(\ppwm_i.u_ppwm.global_counter[12] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0468_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0160_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold342 (.A(\sdr_i.mac2.sum_lvl1_ff[17] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0441_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0012_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold345 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[9] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold346 (.A(\ppwm_i.u_ppwm.u_mem.memory[53] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold347 (.A(\ppwm_i.u_ppwm.u_mem.memory[91] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold348 (.A(\ppwm_i.u_ppwm.u_mem.memory[59] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold349 (.A(\sdr_i.mac2.products_ff[34] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0035_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold351 (.A(\sdr_i.mac2.sum_lvl1_ff[8] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0014_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold353 (.A(\ppwm_i.u_ppwm.u_mem.memory[21] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold354 (.A(\sdr_i.mac1.products_ff[0] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0016_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold356 (.A(\sdr_i.mac1.sum_lvl1_ff[1] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0431_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0024_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold359 (.A(\sdr_i.mac2.products_ff[102] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0039_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold361 (.A(\sdr_i.mac1.products_ff[68] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0020_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold363 (.A(\sdr_i.mac1.sum_lvl2_ff[1] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0435_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0028_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold366 (.A(\sdr_i.mac1.sum_lvl1_ff[24] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0026_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold368 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold369 (.A(\ppwm_i.u_ppwm.u_mem.memory[105] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0320_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold371 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold372 (.A(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0514_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold374 (.A(\sdr_i.mac2.products_ff[69] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0409_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0037_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold377 (.A(\sdr_i.mac2.products_ff[17] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0033_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold379 (.A(\ppwm_i.u_ppwm.u_ex.state_q[0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0000_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold381 (.A(\sdr_i.mac1.products_ff[103] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0429_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0022_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold384 (.A(\sdr_i.mac2.sum_lvl2_ff[4] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0010_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold386 (.A(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0512_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold388 (.A(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold389 (.A(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold390 (.A(\ppwm_i.u_ppwm.pwm_value[3] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0483_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0171_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold393 (.A(\ppwm_i.u_ppwm.u_mem.memory[98] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold394 (.A(\sdr_i.mac1.sum_lvl3_ff[2] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0031_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold396 (.A(\ppwm_i.u_ppwm.global_counter[13] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0161_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold398 (.A(\sdr_i.mac1.products_ff[51] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0018_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold400 (.A(\ppwm_i.u_ppwm.global_counter[16] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0164_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold402 (.A(\sdr_i.mac2.sum_lvl3_ff[1] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0008_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold404 (.A(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold405 (.A(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold406 (.A(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold407 (.A(\ppwm_i.u_ppwm.global_counter[11] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold408 (.A(\ppwm_i.u_ppwm.pc[0] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold409 (.A(\ppwm_i.u_ppwm.global_counter[3] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0151_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold411 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0488_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold413 (.A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold414 (.A(\ppwm_i.u_ppwm.pwm_value[2] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0170_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold416 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0486_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold418 (.A(\ppwm_i.u_ppwm.global_counter[17] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0165_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold420 (.A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0195_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold422 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0494_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold424 (.A(\ppwm_i.u_ppwm.global_counter[18] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold425 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold426 (.A(\ppwm_i.u_ppwm.global_counter[4] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold427 (.A(\ppwm_i.u_ppwm.global_counter[8] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold428 (.A(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold429 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0213_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold431 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold432 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold433 (.A(\ppwm_i.u_ppwm.global_counter[14] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold434 (.A(\ppwm_i.u_ppwm.pwm_value[8] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0203_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold436 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold437 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold438 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold439 (.A(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold440 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold441 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold442 (.A(\ppwm_i.u_ppwm.global_counter[1] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0457_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0149_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold445 (.A(\ppwm_i.u_ppwm.pc[1] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold446 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold447 (.A(\ppwm_i.u_ppwm.pc[2] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold448 (.A(\ppwm_i.u_ppwm.pwm_value[5] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0200_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold450 (.A(\ppwm_i.u_ppwm.pwm_value[6] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold451 (.A(\ppwm_i.u_ppwm.pwm_value[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0196_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold453 (.A(\ppwm_i.u_ppwm.pwm_value[7] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0202_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold455 (.A(\ppwm_i.u_ppwm.pc[3] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold456 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0211_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold458 (.A(\ppwm_i.u_ppwm.pwm_value[4] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold459 (.A(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold460 (.A(_1094_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold461 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .X(net841));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_13 ();
 sg13g2_decap_8 FILLER_0_29 ();
 sg13g2_fill_2 FILLER_0_36 ();
 sg13g2_fill_2 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_61 ();
 sg13g2_decap_8 FILLER_0_68 ();
 sg13g2_decap_8 FILLER_0_75 ();
 sg13g2_decap_8 FILLER_0_82 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_137 ();
 sg13g2_decap_4 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_fill_2 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_4 FILLER_0_177 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_fill_2 FILLER_0_211 ();
 sg13g2_fill_1 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_fill_1 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_4 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_4 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_4 FILLER_0_321 ();
 sg13g2_fill_1 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_4 FILLER_0_365 ();
 sg13g2_fill_1 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_4 FILLER_0_423 ();
 sg13g2_fill_1 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_fill_2 FILLER_0_453 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_decap_8 FILLER_0_473 ();
 sg13g2_decap_8 FILLER_0_480 ();
 sg13g2_decap_4 FILLER_0_487 ();
 sg13g2_fill_1 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_496 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_fill_2 FILLER_0_527 ();
 sg13g2_fill_1 FILLER_0_529 ();
 sg13g2_decap_8 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_541 ();
 sg13g2_decap_8 FILLER_0_548 ();
 sg13g2_decap_8 FILLER_0_555 ();
 sg13g2_decap_8 FILLER_0_562 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_fill_1 FILLER_0_625 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_4 FILLER_0_658 ();
 sg13g2_fill_2 FILLER_0_662 ();
 sg13g2_decap_8 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_675 ();
 sg13g2_decap_8 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_64 ();
 sg13g2_fill_2 FILLER_1_106 ();
 sg13g2_decap_8 FILLER_1_135 ();
 sg13g2_fill_2 FILLER_1_142 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_2 FILLER_1_244 ();
 sg13g2_fill_1 FILLER_1_246 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_fill_2 FILLER_1_281 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_fill_2 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_348 ();
 sg13g2_decap_4 FILLER_1_355 ();
 sg13g2_fill_1 FILLER_1_364 ();
 sg13g2_fill_2 FILLER_1_393 ();
 sg13g2_fill_1 FILLER_1_422 ();
 sg13g2_decap_4 FILLER_1_477 ();
 sg13g2_fill_1 FILLER_1_481 ();
 sg13g2_fill_1 FILLER_1_524 ();
 sg13g2_decap_8 FILLER_1_552 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_601 ();
 sg13g2_decap_8 FILLER_1_608 ();
 sg13g2_decap_4 FILLER_1_615 ();
 sg13g2_fill_2 FILLER_1_619 ();
 sg13g2_decap_8 FILLER_1_648 ();
 sg13g2_fill_2 FILLER_1_655 ();
 sg13g2_fill_1 FILLER_1_657 ();
 sg13g2_fill_1 FILLER_1_688 ();
 sg13g2_decap_8 FILLER_1_716 ();
 sg13g2_decap_8 FILLER_1_723 ();
 sg13g2_decap_8 FILLER_1_730 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_decap_8 FILLER_1_751 ();
 sg13g2_decap_8 FILLER_1_758 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_decap_8 FILLER_1_772 ();
 sg13g2_decap_8 FILLER_1_779 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_821 ();
 sg13g2_decap_8 FILLER_1_828 ();
 sg13g2_decap_8 FILLER_1_835 ();
 sg13g2_decap_8 FILLER_1_842 ();
 sg13g2_decap_8 FILLER_1_849 ();
 sg13g2_decap_8 FILLER_1_856 ();
 sg13g2_decap_8 FILLER_1_863 ();
 sg13g2_decap_8 FILLER_1_870 ();
 sg13g2_decap_8 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_1_884 ();
 sg13g2_decap_8 FILLER_1_891 ();
 sg13g2_decap_8 FILLER_1_898 ();
 sg13g2_decap_8 FILLER_1_905 ();
 sg13g2_decap_8 FILLER_1_912 ();
 sg13g2_decap_8 FILLER_1_919 ();
 sg13g2_decap_8 FILLER_1_926 ();
 sg13g2_decap_8 FILLER_1_933 ();
 sg13g2_decap_8 FILLER_1_940 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_decap_8 FILLER_1_954 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_decap_8 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_989 ();
 sg13g2_decap_8 FILLER_1_996 ();
 sg13g2_decap_8 FILLER_1_1003 ();
 sg13g2_decap_8 FILLER_1_1010 ();
 sg13g2_decap_8 FILLER_1_1017 ();
 sg13g2_decap_4 FILLER_1_1024 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_fill_1 FILLER_2_8 ();
 sg13g2_decap_8 FILLER_2_13 ();
 sg13g2_fill_1 FILLER_2_20 ();
 sg13g2_decap_8 FILLER_2_30 ();
 sg13g2_decap_8 FILLER_2_37 ();
 sg13g2_decap_8 FILLER_2_44 ();
 sg13g2_decap_4 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_141 ();
 sg13g2_decap_8 FILLER_2_150 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_8 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_171 ();
 sg13g2_decap_4 FILLER_2_178 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_fill_2 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_fill_2 FILLER_2_362 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_fill_2 FILLER_2_387 ();
 sg13g2_decap_4 FILLER_2_394 ();
 sg13g2_fill_2 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_4 FILLER_2_418 ();
 sg13g2_fill_1 FILLER_2_454 ();
 sg13g2_fill_1 FILLER_2_470 ();
 sg13g2_fill_2 FILLER_2_485 ();
 sg13g2_decap_4 FILLER_2_500 ();
 sg13g2_decap_4 FILLER_2_509 ();
 sg13g2_decap_8 FILLER_2_538 ();
 sg13g2_decap_8 FILLER_2_545 ();
 sg13g2_decap_8 FILLER_2_552 ();
 sg13g2_fill_2 FILLER_2_559 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_603 ();
 sg13g2_decap_8 FILLER_2_610 ();
 sg13g2_decap_8 FILLER_2_617 ();
 sg13g2_decap_4 FILLER_2_624 ();
 sg13g2_fill_2 FILLER_2_628 ();
 sg13g2_fill_1 FILLER_2_639 ();
 sg13g2_decap_4 FILLER_2_670 ();
 sg13g2_fill_2 FILLER_2_674 ();
 sg13g2_fill_1 FILLER_2_685 ();
 sg13g2_fill_2 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_2 ();
 sg13g2_decap_8 FILLER_3_30 ();
 sg13g2_fill_2 FILLER_3_37 ();
 sg13g2_decap_8 FILLER_3_55 ();
 sg13g2_decap_8 FILLER_3_62 ();
 sg13g2_decap_8 FILLER_3_69 ();
 sg13g2_decap_8 FILLER_3_76 ();
 sg13g2_decap_4 FILLER_3_83 ();
 sg13g2_fill_1 FILLER_3_87 ();
 sg13g2_fill_1 FILLER_3_96 ();
 sg13g2_decap_8 FILLER_3_114 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_209 ();
 sg13g2_decap_4 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_223 ();
 sg13g2_decap_8 FILLER_3_251 ();
 sg13g2_decap_8 FILLER_3_258 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_4 FILLER_3_272 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_4 FILLER_3_314 ();
 sg13g2_fill_2 FILLER_3_318 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_4 FILLER_3_362 ();
 sg13g2_fill_2 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_fill_1 FILLER_3_392 ();
 sg13g2_fill_2 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_2 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_fill_1 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_fill_2 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_fill_1 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_fill_2 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_622 ();
 sg13g2_decap_8 FILLER_3_629 ();
 sg13g2_fill_2 FILLER_3_649 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_decap_4 FILLER_3_677 ();
 sg13g2_fill_2 FILLER_3_681 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_fill_2 FILLER_3_710 ();
 sg13g2_fill_1 FILLER_3_712 ();
 sg13g2_fill_1 FILLER_3_745 ();
 sg13g2_fill_2 FILLER_3_749 ();
 sg13g2_decap_4 FILLER_3_754 ();
 sg13g2_fill_1 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_fill_2 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_8 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_decap_8 FILLER_4_8 ();
 sg13g2_decap_8 FILLER_4_15 ();
 sg13g2_fill_2 FILLER_4_22 ();
 sg13g2_fill_1 FILLER_4_24 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_94 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_decap_8 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_decap_4 FILLER_4_151 ();
 sg13g2_fill_2 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_4 FILLER_4_191 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_2 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_208 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_4 FILLER_4_240 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_fill_2 FILLER_4_302 ();
 sg13g2_fill_1 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_339 ();
 sg13g2_decap_4 FILLER_4_346 ();
 sg13g2_fill_1 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_4 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_fill_2 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_8 FILLER_4_426 ();
 sg13g2_decap_4 FILLER_4_433 ();
 sg13g2_fill_1 FILLER_4_437 ();
 sg13g2_decap_8 FILLER_4_465 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_fill_2 FILLER_4_482 ();
 sg13g2_fill_1 FILLER_4_484 ();
 sg13g2_decap_8 FILLER_4_495 ();
 sg13g2_decap_8 FILLER_4_502 ();
 sg13g2_decap_8 FILLER_4_509 ();
 sg13g2_fill_2 FILLER_4_516 ();
 sg13g2_fill_1 FILLER_4_521 ();
 sg13g2_decap_8 FILLER_4_531 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_decap_8 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_552 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_8 FILLER_4_571 ();
 sg13g2_decap_4 FILLER_4_578 ();
 sg13g2_fill_1 FILLER_4_582 ();
 sg13g2_decap_4 FILLER_4_588 ();
 sg13g2_fill_2 FILLER_4_596 ();
 sg13g2_decap_8 FILLER_4_607 ();
 sg13g2_decap_4 FILLER_4_614 ();
 sg13g2_fill_2 FILLER_4_618 ();
 sg13g2_decap_8 FILLER_4_624 ();
 sg13g2_decap_4 FILLER_4_631 ();
 sg13g2_fill_2 FILLER_4_635 ();
 sg13g2_decap_4 FILLER_4_647 ();
 sg13g2_fill_1 FILLER_4_684 ();
 sg13g2_fill_1 FILLER_4_721 ();
 sg13g2_fill_1 FILLER_4_748 ();
 sg13g2_fill_2 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_decap_8 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_986 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_fill_2 FILLER_5_27 ();
 sg13g2_fill_1 FILLER_5_29 ();
 sg13g2_decap_8 FILLER_5_34 ();
 sg13g2_decap_8 FILLER_5_50 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_decap_8 FILLER_5_71 ();
 sg13g2_decap_4 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_111 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_4 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_4 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_296 ();
 sg13g2_fill_2 FILLER_5_329 ();
 sg13g2_fill_1 FILLER_5_331 ();
 sg13g2_fill_2 FILLER_5_343 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_decap_4 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_390 ();
 sg13g2_fill_1 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_405 ();
 sg13g2_fill_1 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_fill_2 FILLER_5_426 ();
 sg13g2_fill_1 FILLER_5_428 ();
 sg13g2_fill_1 FILLER_5_432 ();
 sg13g2_fill_1 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_4 FILLER_5_476 ();
 sg13g2_fill_1 FILLER_5_486 ();
 sg13g2_fill_2 FILLER_5_514 ();
 sg13g2_decap_4 FILLER_5_530 ();
 sg13g2_fill_1 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_4 FILLER_5_546 ();
 sg13g2_fill_1 FILLER_5_550 ();
 sg13g2_fill_2 FILLER_5_612 ();
 sg13g2_fill_1 FILLER_5_614 ();
 sg13g2_decap_4 FILLER_5_657 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_679 ();
 sg13g2_fill_1 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_4 FILLER_5_707 ();
 sg13g2_fill_2 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_743 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_decap_8 FILLER_5_757 ();
 sg13g2_decap_8 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_fill_1 FILLER_5_794 ();
 sg13g2_decap_8 FILLER_5_804 ();
 sg13g2_decap_8 FILLER_5_811 ();
 sg13g2_decap_8 FILLER_5_818 ();
 sg13g2_decap_8 FILLER_5_825 ();
 sg13g2_decap_8 FILLER_5_832 ();
 sg13g2_decap_8 FILLER_5_839 ();
 sg13g2_decap_8 FILLER_5_846 ();
 sg13g2_decap_8 FILLER_5_853 ();
 sg13g2_decap_8 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_4 FILLER_6_4 ();
 sg13g2_decap_4 FILLER_6_52 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_fill_2 FILLER_6_67 ();
 sg13g2_fill_1 FILLER_6_69 ();
 sg13g2_decap_8 FILLER_6_83 ();
 sg13g2_decap_8 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_97 ();
 sg13g2_decap_8 FILLER_6_104 ();
 sg13g2_decap_8 FILLER_6_111 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_decap_4 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_2 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_4 FILLER_6_364 ();
 sg13g2_decap_4 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_437 ();
 sg13g2_fill_2 FILLER_6_444 ();
 sg13g2_fill_1 FILLER_6_450 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_4 FILLER_6_462 ();
 sg13g2_fill_1 FILLER_6_466 ();
 sg13g2_decap_4 FILLER_6_472 ();
 sg13g2_fill_1 FILLER_6_476 ();
 sg13g2_fill_2 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_496 ();
 sg13g2_decap_8 FILLER_6_503 ();
 sg13g2_decap_8 FILLER_6_510 ();
 sg13g2_fill_1 FILLER_6_523 ();
 sg13g2_fill_1 FILLER_6_529 ();
 sg13g2_fill_1 FILLER_6_557 ();
 sg13g2_fill_2 FILLER_6_567 ();
 sg13g2_fill_1 FILLER_6_569 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_fill_2 FILLER_6_595 ();
 sg13g2_fill_1 FILLER_6_597 ();
 sg13g2_decap_4 FILLER_6_603 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_654 ();
 sg13g2_decap_8 FILLER_6_661 ();
 sg13g2_decap_8 FILLER_6_668 ();
 sg13g2_decap_8 FILLER_6_675 ();
 sg13g2_fill_2 FILLER_6_682 ();
 sg13g2_decap_8 FILLER_6_689 ();
 sg13g2_decap_8 FILLER_6_696 ();
 sg13g2_decap_8 FILLER_6_703 ();
 sg13g2_decap_8 FILLER_6_710 ();
 sg13g2_fill_2 FILLER_6_717 ();
 sg13g2_fill_1 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_4 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_fill_2 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_4 FILLER_6_795 ();
 sg13g2_fill_2 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_828 ();
 sg13g2_decap_8 FILLER_6_835 ();
 sg13g2_decap_8 FILLER_6_842 ();
 sg13g2_decap_8 FILLER_6_849 ();
 sg13g2_decap_8 FILLER_6_856 ();
 sg13g2_decap_8 FILLER_6_863 ();
 sg13g2_decap_8 FILLER_6_870 ();
 sg13g2_decap_8 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_6_884 ();
 sg13g2_decap_8 FILLER_6_891 ();
 sg13g2_decap_8 FILLER_6_898 ();
 sg13g2_decap_8 FILLER_6_905 ();
 sg13g2_decap_8 FILLER_6_912 ();
 sg13g2_decap_8 FILLER_6_919 ();
 sg13g2_decap_8 FILLER_6_926 ();
 sg13g2_decap_8 FILLER_6_933 ();
 sg13g2_decap_8 FILLER_6_940 ();
 sg13g2_decap_8 FILLER_6_947 ();
 sg13g2_decap_8 FILLER_6_954 ();
 sg13g2_decap_8 FILLER_6_961 ();
 sg13g2_decap_8 FILLER_6_968 ();
 sg13g2_decap_8 FILLER_6_975 ();
 sg13g2_decap_8 FILLER_6_982 ();
 sg13g2_decap_8 FILLER_6_989 ();
 sg13g2_decap_8 FILLER_6_996 ();
 sg13g2_decap_8 FILLER_6_1003 ();
 sg13g2_decap_8 FILLER_6_1010 ();
 sg13g2_decap_8 FILLER_6_1017 ();
 sg13g2_decap_4 FILLER_6_1024 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_4 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_8 ();
 sg13g2_decap_8 FILLER_7_13 ();
 sg13g2_fill_1 FILLER_7_20 ();
 sg13g2_decap_8 FILLER_7_30 ();
 sg13g2_decap_8 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_4 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_decap_8 FILLER_7_104 ();
 sg13g2_decap_4 FILLER_7_138 ();
 sg13g2_decap_4 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_296 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_315 ();
 sg13g2_fill_2 FILLER_7_326 ();
 sg13g2_decap_4 FILLER_7_337 ();
 sg13g2_fill_2 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_4 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_fill_2 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_425 ();
 sg13g2_fill_2 FILLER_7_437 ();
 sg13g2_fill_1 FILLER_7_439 ();
 sg13g2_fill_1 FILLER_7_445 ();
 sg13g2_decap_8 FILLER_7_478 ();
 sg13g2_fill_1 FILLER_7_485 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_fill_2 FILLER_7_509 ();
 sg13g2_fill_1 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_524 ();
 sg13g2_decap_8 FILLER_7_531 ();
 sg13g2_decap_8 FILLER_7_538 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_fill_2 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_583 ();
 sg13g2_decap_8 FILLER_7_590 ();
 sg13g2_decap_8 FILLER_7_597 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_fill_2 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_684 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_fill_2 FILLER_7_753 ();
 sg13g2_fill_1 FILLER_7_795 ();
 sg13g2_fill_1 FILLER_7_801 ();
 sg13g2_fill_2 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_decap_8 FILLER_7_829 ();
 sg13g2_decap_8 FILLER_7_836 ();
 sg13g2_decap_8 FILLER_7_843 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_decap_8 FILLER_7_857 ();
 sg13g2_decap_8 FILLER_7_864 ();
 sg13g2_decap_8 FILLER_7_871 ();
 sg13g2_decap_8 FILLER_7_878 ();
 sg13g2_decap_8 FILLER_7_885 ();
 sg13g2_decap_8 FILLER_7_892 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_906 ();
 sg13g2_decap_8 FILLER_7_913 ();
 sg13g2_decap_8 FILLER_7_920 ();
 sg13g2_decap_8 FILLER_7_927 ();
 sg13g2_decap_8 FILLER_7_934 ();
 sg13g2_decap_8 FILLER_7_941 ();
 sg13g2_decap_8 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_955 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_decap_8 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1004 ();
 sg13g2_decap_8 FILLER_7_1011 ();
 sg13g2_decap_8 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_decap_4 FILLER_8_30 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_85 ();
 sg13g2_decap_8 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_106 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_120 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_decap_4 FILLER_8_134 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_199 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_211 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_4 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_264 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_fill_2 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_383 ();
 sg13g2_fill_1 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_449 ();
 sg13g2_decap_8 FILLER_8_456 ();
 sg13g2_decap_4 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_467 ();
 sg13g2_decap_4 FILLER_8_489 ();
 sg13g2_fill_2 FILLER_8_493 ();
 sg13g2_decap_8 FILLER_8_499 ();
 sg13g2_fill_2 FILLER_8_506 ();
 sg13g2_fill_2 FILLER_8_524 ();
 sg13g2_fill_1 FILLER_8_526 ();
 sg13g2_fill_2 FILLER_8_537 ();
 sg13g2_fill_1 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_544 ();
 sg13g2_decap_8 FILLER_8_551 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_fill_2 FILLER_8_598 ();
 sg13g2_fill_2 FILLER_8_627 ();
 sg13g2_decap_4 FILLER_8_639 ();
 sg13g2_fill_2 FILLER_8_643 ();
 sg13g2_decap_8 FILLER_8_667 ();
 sg13g2_decap_8 FILLER_8_674 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_fill_2 FILLER_8_688 ();
 sg13g2_fill_2 FILLER_8_694 ();
 sg13g2_fill_1 FILLER_8_696 ();
 sg13g2_decap_8 FILLER_8_706 ();
 sg13g2_decap_8 FILLER_8_713 ();
 sg13g2_fill_1 FILLER_8_720 ();
 sg13g2_decap_8 FILLER_8_740 ();
 sg13g2_decap_8 FILLER_8_747 ();
 sg13g2_fill_1 FILLER_8_754 ();
 sg13g2_decap_8 FILLER_8_769 ();
 sg13g2_fill_2 FILLER_8_776 ();
 sg13g2_fill_1 FILLER_8_778 ();
 sg13g2_decap_4 FILLER_8_796 ();
 sg13g2_fill_1 FILLER_8_800 ();
 sg13g2_fill_1 FILLER_8_806 ();
 sg13g2_fill_1 FILLER_8_811 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_853 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_decap_8 FILLER_8_874 ();
 sg13g2_decap_8 FILLER_8_881 ();
 sg13g2_decap_8 FILLER_8_888 ();
 sg13g2_decap_8 FILLER_8_895 ();
 sg13g2_decap_8 FILLER_8_902 ();
 sg13g2_decap_8 FILLER_8_909 ();
 sg13g2_decap_8 FILLER_8_916 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_decap_8 FILLER_8_930 ();
 sg13g2_decap_8 FILLER_8_937 ();
 sg13g2_decap_8 FILLER_8_944 ();
 sg13g2_decap_8 FILLER_8_951 ();
 sg13g2_decap_8 FILLER_8_958 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_decap_8 FILLER_8_972 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_4 FILLER_9_18 ();
 sg13g2_fill_2 FILLER_9_22 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_36 ();
 sg13g2_decap_4 FILLER_9_43 ();
 sg13g2_fill_1 FILLER_9_69 ();
 sg13g2_fill_2 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_99 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_118 ();
 sg13g2_decap_4 FILLER_9_146 ();
 sg13g2_fill_1 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_decap_8 FILLER_9_183 ();
 sg13g2_decap_8 FILLER_9_190 ();
 sg13g2_decap_4 FILLER_9_197 ();
 sg13g2_fill_2 FILLER_9_201 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_fill_2 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_4 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_4 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_9_436 ();
 sg13g2_fill_2 FILLER_9_443 ();
 sg13g2_fill_1 FILLER_9_445 ();
 sg13g2_fill_2 FILLER_9_459 ();
 sg13g2_fill_1 FILLER_9_461 ();
 sg13g2_fill_2 FILLER_9_475 ();
 sg13g2_decap_8 FILLER_9_517 ();
 sg13g2_decap_8 FILLER_9_524 ();
 sg13g2_decap_4 FILLER_9_531 ();
 sg13g2_decap_8 FILLER_9_575 ();
 sg13g2_decap_8 FILLER_9_582 ();
 sg13g2_decap_8 FILLER_9_589 ();
 sg13g2_decap_8 FILLER_9_596 ();
 sg13g2_decap_8 FILLER_9_603 ();
 sg13g2_decap_8 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_617 ();
 sg13g2_fill_1 FILLER_9_635 ();
 sg13g2_decap_8 FILLER_9_663 ();
 sg13g2_fill_2 FILLER_9_670 ();
 sg13g2_fill_1 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_691 ();
 sg13g2_decap_8 FILLER_9_698 ();
 sg13g2_decap_8 FILLER_9_705 ();
 sg13g2_decap_4 FILLER_9_712 ();
 sg13g2_fill_1 FILLER_9_716 ();
 sg13g2_decap_4 FILLER_9_724 ();
 sg13g2_fill_2 FILLER_9_728 ();
 sg13g2_decap_4 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_771 ();
 sg13g2_fill_1 FILLER_9_778 ();
 sg13g2_fill_1 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_fill_1 FILLER_9_833 ();
 sg13g2_fill_2 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_decap_8 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_870 ();
 sg13g2_decap_8 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_9_884 ();
 sg13g2_decap_8 FILLER_9_891 ();
 sg13g2_decap_8 FILLER_9_898 ();
 sg13g2_decap_8 FILLER_9_905 ();
 sg13g2_decap_8 FILLER_9_912 ();
 sg13g2_decap_8 FILLER_9_919 ();
 sg13g2_decap_8 FILLER_9_926 ();
 sg13g2_decap_8 FILLER_9_933 ();
 sg13g2_decap_8 FILLER_9_940 ();
 sg13g2_decap_8 FILLER_9_947 ();
 sg13g2_decap_8 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_961 ();
 sg13g2_decap_8 FILLER_9_968 ();
 sg13g2_decap_8 FILLER_9_975 ();
 sg13g2_decap_8 FILLER_9_982 ();
 sg13g2_decap_8 FILLER_9_989 ();
 sg13g2_decap_8 FILLER_9_996 ();
 sg13g2_decap_8 FILLER_9_1003 ();
 sg13g2_decap_8 FILLER_9_1010 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_4 FILLER_9_1024 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_1 FILLER_10_8 ();
 sg13g2_decap_4 FILLER_10_13 ();
 sg13g2_fill_2 FILLER_10_17 ();
 sg13g2_decap_8 FILLER_10_40 ();
 sg13g2_fill_1 FILLER_10_47 ();
 sg13g2_decap_8 FILLER_10_75 ();
 sg13g2_decap_8 FILLER_10_82 ();
 sg13g2_fill_2 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_91 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_311 ();
 sg13g2_decap_4 FILLER_10_340 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_decap_4 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_fill_2 FILLER_10_414 ();
 sg13g2_fill_1 FILLER_10_416 ();
 sg13g2_fill_2 FILLER_10_453 ();
 sg13g2_fill_1 FILLER_10_469 ();
 sg13g2_fill_1 FILLER_10_481 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_fill_1 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_fill_1 FILLER_10_583 ();
 sg13g2_decap_4 FILLER_10_625 ();
 sg13g2_fill_2 FILLER_10_654 ();
 sg13g2_fill_1 FILLER_10_656 ();
 sg13g2_decap_4 FILLER_10_669 ();
 sg13g2_fill_1 FILLER_10_705 ();
 sg13g2_fill_2 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_757 ();
 sg13g2_decap_4 FILLER_10_764 ();
 sg13g2_fill_1 FILLER_10_768 ();
 sg13g2_decap_4 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_fill_1 FILLER_10_826 ();
 sg13g2_fill_1 FILLER_10_830 ();
 sg13g2_fill_2 FILLER_10_836 ();
 sg13g2_fill_1 FILLER_10_838 ();
 sg13g2_decap_8 FILLER_10_867 ();
 sg13g2_decap_8 FILLER_10_874 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_909 ();
 sg13g2_decap_8 FILLER_10_916 ();
 sg13g2_decap_8 FILLER_10_923 ();
 sg13g2_decap_8 FILLER_10_930 ();
 sg13g2_decap_8 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_951 ();
 sg13g2_decap_8 FILLER_10_958 ();
 sg13g2_decap_8 FILLER_10_965 ();
 sg13g2_decap_8 FILLER_10_972 ();
 sg13g2_decap_8 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_986 ();
 sg13g2_decap_8 FILLER_10_993 ();
 sg13g2_decap_8 FILLER_10_1000 ();
 sg13g2_decap_8 FILLER_10_1007 ();
 sg13g2_decap_8 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_fill_2 FILLER_11_75 ();
 sg13g2_decap_4 FILLER_11_85 ();
 sg13g2_fill_2 FILLER_11_89 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_decap_4 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_4 FILLER_11_180 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_4 FILLER_11_305 ();
 sg13g2_decap_4 FILLER_11_336 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_fill_1 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_4 FILLER_11_398 ();
 sg13g2_fill_1 FILLER_11_402 ();
 sg13g2_fill_1 FILLER_11_411 ();
 sg13g2_fill_2 FILLER_11_415 ();
 sg13g2_fill_1 FILLER_11_417 ();
 sg13g2_fill_2 FILLER_11_431 ();
 sg13g2_fill_1 FILLER_11_433 ();
 sg13g2_fill_2 FILLER_11_447 ();
 sg13g2_decap_4 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_468 ();
 sg13g2_fill_1 FILLER_11_475 ();
 sg13g2_decap_8 FILLER_11_499 ();
 sg13g2_decap_8 FILLER_11_506 ();
 sg13g2_decap_4 FILLER_11_513 ();
 sg13g2_fill_2 FILLER_11_517 ();
 sg13g2_fill_2 FILLER_11_524 ();
 sg13g2_fill_2 FILLER_11_584 ();
 sg13g2_decap_8 FILLER_11_594 ();
 sg13g2_fill_2 FILLER_11_601 ();
 sg13g2_fill_1 FILLER_11_603 ();
 sg13g2_decap_4 FILLER_11_613 ();
 sg13g2_fill_2 FILLER_11_617 ();
 sg13g2_fill_2 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_642 ();
 sg13g2_fill_2 FILLER_11_649 ();
 sg13g2_decap_8 FILLER_11_657 ();
 sg13g2_decap_8 FILLER_11_664 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_fill_1 FILLER_11_678 ();
 sg13g2_fill_1 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_fill_2 FILLER_11_707 ();
 sg13g2_decap_4 FILLER_11_717 ();
 sg13g2_fill_2 FILLER_11_721 ();
 sg13g2_fill_2 FILLER_11_726 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_decap_8 FILLER_11_761 ();
 sg13g2_decap_8 FILLER_11_768 ();
 sg13g2_decap_4 FILLER_11_775 ();
 sg13g2_decap_4 FILLER_11_785 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_decap_8 FILLER_11_800 ();
 sg13g2_fill_2 FILLER_11_807 ();
 sg13g2_fill_1 FILLER_11_809 ();
 sg13g2_fill_1 FILLER_11_823 ();
 sg13g2_fill_2 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_881 ();
 sg13g2_decap_8 FILLER_11_888 ();
 sg13g2_decap_8 FILLER_11_895 ();
 sg13g2_decap_8 FILLER_11_902 ();
 sg13g2_decap_8 FILLER_11_909 ();
 sg13g2_decap_8 FILLER_11_916 ();
 sg13g2_decap_8 FILLER_11_923 ();
 sg13g2_decap_8 FILLER_11_930 ();
 sg13g2_decap_8 FILLER_11_937 ();
 sg13g2_decap_8 FILLER_11_944 ();
 sg13g2_decap_8 FILLER_11_951 ();
 sg13g2_decap_8 FILLER_11_958 ();
 sg13g2_decap_8 FILLER_11_965 ();
 sg13g2_decap_8 FILLER_11_972 ();
 sg13g2_decap_8 FILLER_11_979 ();
 sg13g2_decap_8 FILLER_11_986 ();
 sg13g2_decap_8 FILLER_11_993 ();
 sg13g2_decap_8 FILLER_11_1000 ();
 sg13g2_decap_8 FILLER_11_1007 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_decap_8 FILLER_11_1021 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_fill_2 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_fill_1 FILLER_12_111 ();
 sg13g2_decap_8 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_decap_8 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_264 ();
 sg13g2_decap_4 FILLER_12_280 ();
 sg13g2_decap_4 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_300 ();
 sg13g2_decap_4 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_333 ();
 sg13g2_decap_4 FILLER_12_347 ();
 sg13g2_fill_2 FILLER_12_351 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_4 FILLER_12_386 ();
 sg13g2_fill_1 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_4 FILLER_12_448 ();
 sg13g2_fill_2 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_458 ();
 sg13g2_decap_4 FILLER_12_470 ();
 sg13g2_fill_2 FILLER_12_474 ();
 sg13g2_fill_1 FILLER_12_481 ();
 sg13g2_decap_8 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_fill_1 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_565 ();
 sg13g2_decap_8 FILLER_12_572 ();
 sg13g2_decap_4 FILLER_12_579 ();
 sg13g2_fill_2 FILLER_12_583 ();
 sg13g2_fill_1 FILLER_12_612 ();
 sg13g2_fill_2 FILLER_12_632 ();
 sg13g2_fill_1 FILLER_12_634 ();
 sg13g2_decap_4 FILLER_12_653 ();
 sg13g2_fill_1 FILLER_12_657 ();
 sg13g2_fill_1 FILLER_12_697 ();
 sg13g2_decap_4 FILLER_12_711 ();
 sg13g2_fill_2 FILLER_12_728 ();
 sg13g2_decap_4 FILLER_12_750 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_fill_2 FILLER_12_769 ();
 sg13g2_fill_1 FILLER_12_771 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_4 FILLER_12_840 ();
 sg13g2_fill_1 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_decap_8 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_12_884 ();
 sg13g2_decap_8 FILLER_12_891 ();
 sg13g2_decap_8 FILLER_12_898 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_decap_8 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_926 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_8 FILLER_12_940 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_decap_8 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_decap_8 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_975 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_decap_8 FILLER_12_989 ();
 sg13g2_decap_8 FILLER_12_996 ();
 sg13g2_decap_8 FILLER_12_1003 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_decap_8 FILLER_12_1017 ();
 sg13g2_decap_4 FILLER_12_1024 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_fill_1 FILLER_13_8 ();
 sg13g2_decap_8 FILLER_13_13 ();
 sg13g2_fill_1 FILLER_13_20 ();
 sg13g2_decap_4 FILLER_13_30 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_40 ();
 sg13g2_decap_8 FILLER_13_45 ();
 sg13g2_decap_4 FILLER_13_52 ();
 sg13g2_decap_8 FILLER_13_65 ();
 sg13g2_decap_8 FILLER_13_72 ();
 sg13g2_decap_8 FILLER_13_79 ();
 sg13g2_decap_8 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_decap_4 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_428 ();
 sg13g2_fill_2 FILLER_13_435 ();
 sg13g2_fill_1 FILLER_13_437 ();
 sg13g2_fill_2 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_decap_8 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_471 ();
 sg13g2_fill_1 FILLER_13_478 ();
 sg13g2_decap_8 FILLER_13_484 ();
 sg13g2_decap_8 FILLER_13_491 ();
 sg13g2_fill_2 FILLER_13_498 ();
 sg13g2_fill_1 FILLER_13_500 ();
 sg13g2_decap_8 FILLER_13_507 ();
 sg13g2_decap_8 FILLER_13_514 ();
 sg13g2_fill_1 FILLER_13_521 ();
 sg13g2_decap_4 FILLER_13_548 ();
 sg13g2_fill_2 FILLER_13_552 ();
 sg13g2_decap_8 FILLER_13_562 ();
 sg13g2_decap_8 FILLER_13_569 ();
 sg13g2_decap_8 FILLER_13_576 ();
 sg13g2_fill_2 FILLER_13_583 ();
 sg13g2_fill_1 FILLER_13_585 ();
 sg13g2_decap_8 FILLER_13_600 ();
 sg13g2_decap_8 FILLER_13_607 ();
 sg13g2_fill_2 FILLER_13_614 ();
 sg13g2_decap_4 FILLER_13_635 ();
 sg13g2_fill_1 FILLER_13_639 ();
 sg13g2_fill_2 FILLER_13_660 ();
 sg13g2_fill_1 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_667 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_fill_1 FILLER_13_681 ();
 sg13g2_fill_1 FILLER_13_687 ();
 sg13g2_decap_8 FILLER_13_696 ();
 sg13g2_fill_1 FILLER_13_703 ();
 sg13g2_fill_1 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_717 ();
 sg13g2_decap_8 FILLER_13_724 ();
 sg13g2_decap_4 FILLER_13_731 ();
 sg13g2_fill_1 FILLER_13_735 ();
 sg13g2_decap_4 FILLER_13_753 ();
 sg13g2_fill_1 FILLER_13_757 ();
 sg13g2_fill_2 FILLER_13_771 ();
 sg13g2_fill_1 FILLER_13_773 ();
 sg13g2_decap_8 FILLER_13_785 ();
 sg13g2_decap_8 FILLER_13_792 ();
 sg13g2_decap_4 FILLER_13_799 ();
 sg13g2_fill_1 FILLER_13_803 ();
 sg13g2_fill_1 FILLER_13_809 ();
 sg13g2_fill_1 FILLER_13_850 ();
 sg13g2_decap_8 FILLER_13_864 ();
 sg13g2_decap_8 FILLER_13_871 ();
 sg13g2_decap_8 FILLER_13_878 ();
 sg13g2_decap_8 FILLER_13_885 ();
 sg13g2_decap_8 FILLER_13_892 ();
 sg13g2_decap_8 FILLER_13_899 ();
 sg13g2_decap_8 FILLER_13_906 ();
 sg13g2_decap_8 FILLER_13_913 ();
 sg13g2_decap_8 FILLER_13_920 ();
 sg13g2_decap_8 FILLER_13_927 ();
 sg13g2_decap_8 FILLER_13_934 ();
 sg13g2_decap_8 FILLER_13_941 ();
 sg13g2_decap_8 FILLER_13_948 ();
 sg13g2_decap_8 FILLER_13_955 ();
 sg13g2_decap_8 FILLER_13_962 ();
 sg13g2_decap_8 FILLER_13_969 ();
 sg13g2_decap_8 FILLER_13_976 ();
 sg13g2_decap_8 FILLER_13_983 ();
 sg13g2_decap_8 FILLER_13_990 ();
 sg13g2_decap_8 FILLER_13_997 ();
 sg13g2_decap_8 FILLER_13_1004 ();
 sg13g2_decap_8 FILLER_13_1011 ();
 sg13g2_decap_8 FILLER_13_1018 ();
 sg13g2_decap_4 FILLER_13_1025 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_30 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_4 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_decap_4 FILLER_14_145 ();
 sg13g2_fill_2 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_fill_1 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_4 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_decap_4 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_4 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_14_417 ();
 sg13g2_fill_2 FILLER_14_421 ();
 sg13g2_decap_4 FILLER_14_464 ();
 sg13g2_fill_2 FILLER_14_468 ();
 sg13g2_decap_4 FILLER_14_486 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_decap_4 FILLER_14_521 ();
 sg13g2_fill_1 FILLER_14_525 ();
 sg13g2_decap_4 FILLER_14_539 ();
 sg13g2_fill_2 FILLER_14_543 ();
 sg13g2_fill_2 FILLER_14_561 ();
 sg13g2_decap_4 FILLER_14_603 ();
 sg13g2_fill_2 FILLER_14_607 ();
 sg13g2_decap_8 FILLER_14_629 ();
 sg13g2_decap_8 FILLER_14_636 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_fill_1 FILLER_14_650 ();
 sg13g2_fill_2 FILLER_14_660 ();
 sg13g2_fill_1 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_4 FILLER_14_700 ();
 sg13g2_fill_2 FILLER_14_708 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_4 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_4 FILLER_14_767 ();
 sg13g2_fill_2 FILLER_14_771 ();
 sg13g2_fill_2 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_fill_2 FILLER_14_812 ();
 sg13g2_fill_1 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_fill_1 FILLER_14_833 ();
 sg13g2_fill_1 FILLER_14_851 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_decap_8 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_decap_8 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_942 ();
 sg13g2_decap_8 FILLER_14_949 ();
 sg13g2_decap_8 FILLER_14_956 ();
 sg13g2_decap_8 FILLER_14_963 ();
 sg13g2_decap_8 FILLER_14_970 ();
 sg13g2_decap_8 FILLER_14_977 ();
 sg13g2_decap_8 FILLER_14_984 ();
 sg13g2_decap_8 FILLER_14_991 ();
 sg13g2_decap_8 FILLER_14_998 ();
 sg13g2_decap_8 FILLER_14_1005 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_fill_2 FILLER_14_1026 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_15_8 ();
 sg13g2_decap_8 FILLER_15_13 ();
 sg13g2_fill_2 FILLER_15_29 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_124 ();
 sg13g2_decap_8 FILLER_15_131 ();
 sg13g2_decap_8 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_4 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_4 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_fill_1 FILLER_15_376 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_1 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_4 FILLER_15_462 ();
 sg13g2_fill_2 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_fill_2 FILLER_15_512 ();
 sg13g2_decap_8 FILLER_15_523 ();
 sg13g2_decap_8 FILLER_15_530 ();
 sg13g2_decap_8 FILLER_15_548 ();
 sg13g2_fill_2 FILLER_15_555 ();
 sg13g2_fill_1 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_572 ();
 sg13g2_decap_8 FILLER_15_579 ();
 sg13g2_decap_8 FILLER_15_586 ();
 sg13g2_decap_8 FILLER_15_593 ();
 sg13g2_decap_8 FILLER_15_600 ();
 sg13g2_decap_4 FILLER_15_607 ();
 sg13g2_fill_1 FILLER_15_611 ();
 sg13g2_decap_8 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_decap_8 FILLER_15_639 ();
 sg13g2_fill_1 FILLER_15_646 ();
 sg13g2_fill_2 FILLER_15_655 ();
 sg13g2_fill_1 FILLER_15_657 ();
 sg13g2_decap_8 FILLER_15_698 ();
 sg13g2_decap_4 FILLER_15_705 ();
 sg13g2_fill_1 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_716 ();
 sg13g2_decap_4 FILLER_15_723 ();
 sg13g2_fill_2 FILLER_15_727 ();
 sg13g2_decap_8 FILLER_15_750 ();
 sg13g2_decap_8 FILLER_15_757 ();
 sg13g2_fill_1 FILLER_15_764 ();
 sg13g2_fill_2 FILLER_15_808 ();
 sg13g2_fill_1 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_fill_1 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_871 ();
 sg13g2_decap_8 FILLER_15_878 ();
 sg13g2_decap_8 FILLER_15_885 ();
 sg13g2_decap_8 FILLER_15_892 ();
 sg13g2_decap_8 FILLER_15_899 ();
 sg13g2_decap_8 FILLER_15_906 ();
 sg13g2_decap_8 FILLER_15_913 ();
 sg13g2_decap_8 FILLER_15_920 ();
 sg13g2_decap_8 FILLER_15_927 ();
 sg13g2_decap_8 FILLER_15_934 ();
 sg13g2_decap_8 FILLER_15_941 ();
 sg13g2_decap_8 FILLER_15_948 ();
 sg13g2_decap_8 FILLER_15_955 ();
 sg13g2_decap_8 FILLER_15_962 ();
 sg13g2_decap_8 FILLER_15_969 ();
 sg13g2_decap_8 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_983 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_decap_8 FILLER_15_997 ();
 sg13g2_decap_8 FILLER_15_1004 ();
 sg13g2_decap_8 FILLER_15_1011 ();
 sg13g2_decap_8 FILLER_15_1018 ();
 sg13g2_decap_4 FILLER_15_1025 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_29 ();
 sg13g2_decap_8 FILLER_16_58 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_94 ();
 sg13g2_decap_8 FILLER_16_101 ();
 sg13g2_decap_8 FILLER_16_108 ();
 sg13g2_decap_4 FILLER_16_128 ();
 sg13g2_decap_4 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_4 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_424 ();
 sg13g2_decap_4 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_16_433 ();
 sg13g2_decap_8 FILLER_16_439 ();
 sg13g2_decap_8 FILLER_16_446 ();
 sg13g2_fill_2 FILLER_16_453 ();
 sg13g2_fill_1 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_461 ();
 sg13g2_fill_2 FILLER_16_468 ();
 sg13g2_decap_4 FILLER_16_478 ();
 sg13g2_fill_1 FILLER_16_482 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_decap_8 FILLER_16_494 ();
 sg13g2_fill_2 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_4 FILLER_16_583 ();
 sg13g2_fill_2 FILLER_16_587 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_4 FILLER_16_609 ();
 sg13g2_fill_2 FILLER_16_613 ();
 sg13g2_fill_1 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_633 ();
 sg13g2_decap_8 FILLER_16_640 ();
 sg13g2_fill_1 FILLER_16_647 ();
 sg13g2_fill_1 FILLER_16_653 ();
 sg13g2_fill_1 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_fill_2 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_731 ();
 sg13g2_fill_1 FILLER_16_738 ();
 sg13g2_decap_8 FILLER_16_766 ();
 sg13g2_fill_1 FILLER_16_773 ();
 sg13g2_fill_2 FILLER_16_786 ();
 sg13g2_fill_1 FILLER_16_788 ();
 sg13g2_decap_4 FILLER_16_821 ();
 sg13g2_fill_2 FILLER_16_825 ();
 sg13g2_decap_4 FILLER_16_831 ();
 sg13g2_fill_1 FILLER_16_835 ();
 sg13g2_decap_4 FILLER_16_851 ();
 sg13g2_fill_2 FILLER_16_855 ();
 sg13g2_decap_8 FILLER_16_885 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_8 FILLER_16_899 ();
 sg13g2_decap_8 FILLER_16_906 ();
 sg13g2_decap_8 FILLER_16_913 ();
 sg13g2_decap_8 FILLER_16_920 ();
 sg13g2_decap_8 FILLER_16_927 ();
 sg13g2_decap_8 FILLER_16_934 ();
 sg13g2_decap_8 FILLER_16_941 ();
 sg13g2_decap_8 FILLER_16_948 ();
 sg13g2_decap_8 FILLER_16_955 ();
 sg13g2_decap_8 FILLER_16_962 ();
 sg13g2_decap_8 FILLER_16_969 ();
 sg13g2_decap_8 FILLER_16_976 ();
 sg13g2_decap_8 FILLER_16_983 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_decap_8 FILLER_16_997 ();
 sg13g2_decap_8 FILLER_16_1004 ();
 sg13g2_decap_8 FILLER_16_1011 ();
 sg13g2_decap_8 FILLER_16_1018 ();
 sg13g2_decap_4 FILLER_16_1025 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_30 ();
 sg13g2_decap_8 FILLER_17_37 ();
 sg13g2_decap_8 FILLER_17_44 ();
 sg13g2_decap_8 FILLER_17_51 ();
 sg13g2_decap_4 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_decap_4 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_4 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_465 ();
 sg13g2_decap_4 FILLER_17_472 ();
 sg13g2_decap_8 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_487 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_fill_2 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_fill_2 FILLER_17_542 ();
 sg13g2_fill_1 FILLER_17_544 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_fill_2 FILLER_17_612 ();
 sg13g2_decap_8 FILLER_17_663 ();
 sg13g2_decap_8 FILLER_17_670 ();
 sg13g2_decap_8 FILLER_17_677 ();
 sg13g2_decap_8 FILLER_17_684 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_decap_8 FILLER_17_715 ();
 sg13g2_decap_4 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_726 ();
 sg13g2_fill_1 FILLER_17_733 ();
 sg13g2_fill_1 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_748 ();
 sg13g2_decap_4 FILLER_17_755 ();
 sg13g2_decap_4 FILLER_17_764 ();
 sg13g2_fill_1 FILLER_17_768 ();
 sg13g2_fill_2 FILLER_17_781 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_803 ();
 sg13g2_fill_1 FILLER_17_816 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_18_8 ();
 sg13g2_decap_4 FILLER_18_13 ();
 sg13g2_fill_2 FILLER_18_17 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_decap_8 FILLER_18_90 ();
 sg13g2_decap_4 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_4 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_208 ();
 sg13g2_decap_8 FILLER_18_215 ();
 sg13g2_decap_8 FILLER_18_222 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_decap_8 FILLER_18_243 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_4 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_fill_1 FILLER_18_410 ();
 sg13g2_decap_4 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_429 ();
 sg13g2_decap_4 FILLER_18_436 ();
 sg13g2_fill_2 FILLER_18_440 ();
 sg13g2_fill_2 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_461 ();
 sg13g2_fill_2 FILLER_18_499 ();
 sg13g2_decap_8 FILLER_18_505 ();
 sg13g2_decap_8 FILLER_18_512 ();
 sg13g2_decap_4 FILLER_18_519 ();
 sg13g2_fill_1 FILLER_18_523 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_554 ();
 sg13g2_decap_4 FILLER_18_561 ();
 sg13g2_fill_2 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_621 ();
 sg13g2_decap_4 FILLER_18_628 ();
 sg13g2_decap_8 FILLER_18_636 ();
 sg13g2_decap_8 FILLER_18_643 ();
 sg13g2_decap_8 FILLER_18_650 ();
 sg13g2_decap_8 FILLER_18_657 ();
 sg13g2_decap_8 FILLER_18_664 ();
 sg13g2_fill_1 FILLER_18_671 ();
 sg13g2_fill_2 FILLER_18_698 ();
 sg13g2_decap_4 FILLER_18_725 ();
 sg13g2_fill_1 FILLER_18_734 ();
 sg13g2_decap_4 FILLER_18_770 ();
 sg13g2_fill_2 FILLER_18_774 ();
 sg13g2_decap_4 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_856 ();
 sg13g2_fill_2 FILLER_18_863 ();
 sg13g2_decap_8 FILLER_18_869 ();
 sg13g2_decap_8 FILLER_18_876 ();
 sg13g2_decap_8 FILLER_18_883 ();
 sg13g2_decap_8 FILLER_18_890 ();
 sg13g2_decap_8 FILLER_18_897 ();
 sg13g2_decap_8 FILLER_18_904 ();
 sg13g2_decap_8 FILLER_18_911 ();
 sg13g2_decap_8 FILLER_18_918 ();
 sg13g2_decap_8 FILLER_18_925 ();
 sg13g2_decap_8 FILLER_18_932 ();
 sg13g2_decap_8 FILLER_18_939 ();
 sg13g2_decap_8 FILLER_18_946 ();
 sg13g2_decap_8 FILLER_18_953 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_decap_8 FILLER_18_967 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_decap_8 FILLER_18_981 ();
 sg13g2_decap_8 FILLER_18_988 ();
 sg13g2_decap_8 FILLER_18_995 ();
 sg13g2_decap_8 FILLER_18_1002 ();
 sg13g2_decap_8 FILLER_18_1009 ();
 sg13g2_decap_8 FILLER_18_1016 ();
 sg13g2_decap_4 FILLER_18_1023 ();
 sg13g2_fill_2 FILLER_18_1027 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_55 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_decap_8 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_decap_8 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_142 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_1 FILLER_19_407 ();
 sg13g2_fill_1 FILLER_19_439 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_4 FILLER_19_525 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_fill_2 FILLER_19_541 ();
 sg13g2_fill_1 FILLER_19_543 ();
 sg13g2_fill_1 FILLER_19_549 ();
 sg13g2_decap_8 FILLER_19_563 ();
 sg13g2_decap_8 FILLER_19_570 ();
 sg13g2_decap_4 FILLER_19_577 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_fill_2 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_617 ();
 sg13g2_fill_1 FILLER_19_624 ();
 sg13g2_decap_4 FILLER_19_638 ();
 sg13g2_decap_8 FILLER_19_646 ();
 sg13g2_decap_4 FILLER_19_662 ();
 sg13g2_decap_4 FILLER_19_685 ();
 sg13g2_fill_2 FILLER_19_689 ();
 sg13g2_fill_1 FILLER_19_695 ();
 sg13g2_fill_1 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_decap_4 FILLER_19_727 ();
 sg13g2_fill_2 FILLER_19_731 ();
 sg13g2_fill_2 FILLER_19_738 ();
 sg13g2_decap_8 FILLER_19_744 ();
 sg13g2_decap_4 FILLER_19_751 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_4 FILLER_19_774 ();
 sg13g2_fill_2 FILLER_19_778 ();
 sg13g2_fill_2 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_790 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_fill_2 FILLER_19_819 ();
 sg13g2_fill_1 FILLER_19_821 ();
 sg13g2_fill_2 FILLER_19_848 ();
 sg13g2_fill_1 FILLER_19_850 ();
 sg13g2_decap_8 FILLER_19_888 ();
 sg13g2_decap_8 FILLER_19_895 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_8 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_930 ();
 sg13g2_decap_8 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_944 ();
 sg13g2_decap_8 FILLER_19_951 ();
 sg13g2_decap_8 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_decap_8 FILLER_19_1000 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1021 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_4 FILLER_20_18 ();
 sg13g2_fill_2 FILLER_20_22 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_decap_4 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_4 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_decap_4 FILLER_20_438 ();
 sg13g2_fill_2 FILLER_20_442 ();
 sg13g2_decap_4 FILLER_20_478 ();
 sg13g2_decap_8 FILLER_20_492 ();
 sg13g2_fill_2 FILLER_20_499 ();
 sg13g2_fill_2 FILLER_20_506 ();
 sg13g2_decap_8 FILLER_20_513 ();
 sg13g2_fill_2 FILLER_20_520 ();
 sg13g2_decap_8 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_542 ();
 sg13g2_fill_1 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_549 ();
 sg13g2_fill_2 FILLER_20_556 ();
 sg13g2_fill_1 FILLER_20_558 ();
 sg13g2_decap_4 FILLER_20_572 ();
 sg13g2_fill_2 FILLER_20_576 ();
 sg13g2_decap_4 FILLER_20_591 ();
 sg13g2_fill_1 FILLER_20_595 ();
 sg13g2_fill_2 FILLER_20_600 ();
 sg13g2_fill_1 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_fill_1 FILLER_20_664 ();
 sg13g2_decap_4 FILLER_20_682 ();
 sg13g2_fill_1 FILLER_20_704 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_4 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_4 FILLER_20_770 ();
 sg13g2_fill_2 FILLER_20_774 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_4 FILLER_20_818 ();
 sg13g2_fill_1 FILLER_20_822 ();
 sg13g2_decap_4 FILLER_20_845 ();
 sg13g2_fill_1 FILLER_20_849 ();
 sg13g2_decap_8 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_20_884 ();
 sg13g2_decap_8 FILLER_20_891 ();
 sg13g2_decap_8 FILLER_20_898 ();
 sg13g2_decap_8 FILLER_20_905 ();
 sg13g2_decap_8 FILLER_20_912 ();
 sg13g2_decap_8 FILLER_20_919 ();
 sg13g2_decap_8 FILLER_20_926 ();
 sg13g2_decap_8 FILLER_20_933 ();
 sg13g2_decap_8 FILLER_20_940 ();
 sg13g2_decap_8 FILLER_20_947 ();
 sg13g2_decap_8 FILLER_20_954 ();
 sg13g2_decap_8 FILLER_20_961 ();
 sg13g2_decap_8 FILLER_20_968 ();
 sg13g2_decap_8 FILLER_20_975 ();
 sg13g2_decap_8 FILLER_20_982 ();
 sg13g2_decap_8 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_996 ();
 sg13g2_decap_8 FILLER_20_1003 ();
 sg13g2_decap_8 FILLER_20_1010 ();
 sg13g2_decap_8 FILLER_20_1017 ();
 sg13g2_decap_4 FILLER_20_1024 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_1 FILLER_21_8 ();
 sg13g2_decap_4 FILLER_21_13 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_decap_8 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_66 ();
 sg13g2_decap_8 FILLER_21_73 ();
 sg13g2_decap_4 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_99 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_148 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_400 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_21_435 ();
 sg13g2_decap_8 FILLER_21_442 ();
 sg13g2_decap_4 FILLER_21_449 ();
 sg13g2_fill_2 FILLER_21_453 ();
 sg13g2_decap_8 FILLER_21_468 ();
 sg13g2_decap_8 FILLER_21_496 ();
 sg13g2_fill_1 FILLER_21_508 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_8 FILLER_21_540 ();
 sg13g2_decap_8 FILLER_21_547 ();
 sg13g2_fill_1 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_597 ();
 sg13g2_decap_4 FILLER_21_604 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_decap_8 FILLER_21_619 ();
 sg13g2_fill_2 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_fill_2 FILLER_21_665 ();
 sg13g2_fill_1 FILLER_21_670 ();
 sg13g2_fill_2 FILLER_21_676 ();
 sg13g2_fill_1 FILLER_21_678 ();
 sg13g2_decap_4 FILLER_21_706 ();
 sg13g2_fill_1 FILLER_21_710 ();
 sg13g2_decap_4 FILLER_21_721 ();
 sg13g2_fill_2 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_737 ();
 sg13g2_decap_4 FILLER_21_744 ();
 sg13g2_fill_1 FILLER_21_775 ();
 sg13g2_fill_2 FILLER_21_788 ();
 sg13g2_fill_1 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_4 FILLER_21_826 ();
 sg13g2_fill_2 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_863 ();
 sg13g2_decap_8 FILLER_21_870 ();
 sg13g2_decap_8 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_21_884 ();
 sg13g2_decap_8 FILLER_21_891 ();
 sg13g2_decap_8 FILLER_21_898 ();
 sg13g2_decap_8 FILLER_21_905 ();
 sg13g2_decap_8 FILLER_21_912 ();
 sg13g2_decap_8 FILLER_21_919 ();
 sg13g2_decap_8 FILLER_21_926 ();
 sg13g2_decap_8 FILLER_21_933 ();
 sg13g2_decap_8 FILLER_21_940 ();
 sg13g2_decap_8 FILLER_21_947 ();
 sg13g2_decap_8 FILLER_21_954 ();
 sg13g2_decap_8 FILLER_21_961 ();
 sg13g2_decap_8 FILLER_21_968 ();
 sg13g2_decap_8 FILLER_21_975 ();
 sg13g2_decap_8 FILLER_21_982 ();
 sg13g2_decap_8 FILLER_21_989 ();
 sg13g2_decap_8 FILLER_21_996 ();
 sg13g2_decap_8 FILLER_21_1003 ();
 sg13g2_decap_8 FILLER_21_1010 ();
 sg13g2_decap_8 FILLER_21_1017 ();
 sg13g2_decap_4 FILLER_21_1024 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_22_27 ();
 sg13g2_decap_8 FILLER_22_34 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_decap_8 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_decap_4 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_4 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_22_458 ();
 sg13g2_decap_8 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_479 ();
 sg13g2_decap_8 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_493 ();
 sg13g2_decap_8 FILLER_22_500 ();
 sg13g2_decap_8 FILLER_22_507 ();
 sg13g2_decap_4 FILLER_22_514 ();
 sg13g2_decap_8 FILLER_22_535 ();
 sg13g2_decap_8 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_549 ();
 sg13g2_decap_8 FILLER_22_556 ();
 sg13g2_fill_2 FILLER_22_563 ();
 sg13g2_decap_4 FILLER_22_570 ();
 sg13g2_fill_2 FILLER_22_578 ();
 sg13g2_fill_1 FILLER_22_580 ();
 sg13g2_decap_4 FILLER_22_604 ();
 sg13g2_fill_1 FILLER_22_608 ();
 sg13g2_decap_8 FILLER_22_614 ();
 sg13g2_decap_8 FILLER_22_621 ();
 sg13g2_decap_8 FILLER_22_628 ();
 sg13g2_fill_1 FILLER_22_635 ();
 sg13g2_fill_2 FILLER_22_663 ();
 sg13g2_fill_1 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_689 ();
 sg13g2_fill_1 FILLER_22_696 ();
 sg13g2_decap_4 FILLER_22_702 ();
 sg13g2_fill_2 FILLER_22_706 ();
 sg13g2_fill_2 FILLER_22_716 ();
 sg13g2_fill_1 FILLER_22_718 ();
 sg13g2_decap_4 FILLER_22_747 ();
 sg13g2_fill_2 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_decap_8 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_780 ();
 sg13g2_fill_1 FILLER_22_794 ();
 sg13g2_decap_4 FILLER_22_798 ();
 sg13g2_fill_2 FILLER_22_807 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_fill_1 FILLER_22_823 ();
 sg13g2_decap_4 FILLER_22_827 ();
 sg13g2_fill_1 FILLER_22_831 ();
 sg13g2_fill_2 FILLER_22_845 ();
 sg13g2_fill_1 FILLER_22_856 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_decap_8 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_891 ();
 sg13g2_decap_8 FILLER_22_898 ();
 sg13g2_decap_8 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_912 ();
 sg13g2_decap_8 FILLER_22_919 ();
 sg13g2_decap_8 FILLER_22_926 ();
 sg13g2_decap_8 FILLER_22_933 ();
 sg13g2_decap_8 FILLER_22_940 ();
 sg13g2_decap_8 FILLER_22_947 ();
 sg13g2_decap_8 FILLER_22_954 ();
 sg13g2_decap_8 FILLER_22_961 ();
 sg13g2_decap_8 FILLER_22_968 ();
 sg13g2_decap_8 FILLER_22_975 ();
 sg13g2_decap_8 FILLER_22_982 ();
 sg13g2_decap_8 FILLER_22_989 ();
 sg13g2_decap_8 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1010 ();
 sg13g2_decap_8 FILLER_22_1017 ();
 sg13g2_decap_4 FILLER_22_1024 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_78 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_2 FILLER_23_202 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_decap_4 FILLER_23_253 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_4 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_413 ();
 sg13g2_fill_1 FILLER_23_415 ();
 sg13g2_fill_2 FILLER_23_421 ();
 sg13g2_fill_1 FILLER_23_423 ();
 sg13g2_decap_4 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_23_433 ();
 sg13g2_decap_8 FILLER_23_439 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_decap_8 FILLER_23_457 ();
 sg13g2_fill_1 FILLER_23_464 ();
 sg13g2_decap_4 FILLER_23_492 ();
 sg13g2_decap_8 FILLER_23_524 ();
 sg13g2_decap_8 FILLER_23_531 ();
 sg13g2_fill_2 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_540 ();
 sg13g2_decap_8 FILLER_23_554 ();
 sg13g2_decap_8 FILLER_23_561 ();
 sg13g2_decap_8 FILLER_23_568 ();
 sg13g2_fill_2 FILLER_23_575 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_597 ();
 sg13g2_decap_8 FILLER_23_622 ();
 sg13g2_decap_8 FILLER_23_629 ();
 sg13g2_decap_4 FILLER_23_636 ();
 sg13g2_fill_2 FILLER_23_640 ();
 sg13g2_decap_8 FILLER_23_646 ();
 sg13g2_decap_8 FILLER_23_653 ();
 sg13g2_decap_8 FILLER_23_660 ();
 sg13g2_decap_4 FILLER_23_667 ();
 sg13g2_fill_1 FILLER_23_671 ();
 sg13g2_decap_8 FILLER_23_689 ();
 sg13g2_decap_8 FILLER_23_696 ();
 sg13g2_fill_2 FILLER_23_708 ();
 sg13g2_fill_1 FILLER_23_719 ();
 sg13g2_fill_2 FILLER_23_733 ();
 sg13g2_decap_4 FILLER_23_748 ();
 sg13g2_fill_1 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_fill_2 FILLER_23_772 ();
 sg13g2_fill_1 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_4 FILLER_23_829 ();
 sg13g2_fill_2 FILLER_23_833 ();
 sg13g2_decap_4 FILLER_23_840 ();
 sg13g2_fill_2 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_873 ();
 sg13g2_decap_8 FILLER_23_880 ();
 sg13g2_decap_8 FILLER_23_887 ();
 sg13g2_decap_8 FILLER_23_894 ();
 sg13g2_decap_8 FILLER_23_901 ();
 sg13g2_decap_8 FILLER_23_908 ();
 sg13g2_decap_8 FILLER_23_915 ();
 sg13g2_decap_8 FILLER_23_922 ();
 sg13g2_decap_8 FILLER_23_929 ();
 sg13g2_decap_8 FILLER_23_936 ();
 sg13g2_decap_8 FILLER_23_943 ();
 sg13g2_decap_8 FILLER_23_950 ();
 sg13g2_decap_8 FILLER_23_957 ();
 sg13g2_decap_8 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_971 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_8 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_999 ();
 sg13g2_decap_8 FILLER_23_1006 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_decap_8 FILLER_23_1020 ();
 sg13g2_fill_2 FILLER_23_1027 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_34 ();
 sg13g2_decap_4 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_390 ();
 sg13g2_decap_4 FILLER_24_430 ();
 sg13g2_fill_1 FILLER_24_446 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_4 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_517 ();
 sg13g2_decap_4 FILLER_24_524 ();
 sg13g2_fill_2 FILLER_24_528 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_fill_1 FILLER_24_546 ();
 sg13g2_decap_4 FILLER_24_575 ();
 sg13g2_fill_2 FILLER_24_579 ();
 sg13g2_decap_4 FILLER_24_586 ();
 sg13g2_fill_2 FILLER_24_590 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_4 FILLER_24_606 ();
 sg13g2_fill_2 FILLER_24_610 ();
 sg13g2_decap_4 FILLER_24_625 ();
 sg13g2_fill_1 FILLER_24_629 ();
 sg13g2_decap_4 FILLER_24_643 ();
 sg13g2_fill_2 FILLER_24_647 ();
 sg13g2_fill_2 FILLER_24_676 ();
 sg13g2_decap_4 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_fill_2 FILLER_24_796 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_fill_1 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_fill_2 FILLER_24_834 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_decap_8 FILLER_24_875 ();
 sg13g2_decap_8 FILLER_24_882 ();
 sg13g2_decap_8 FILLER_24_889 ();
 sg13g2_decap_8 FILLER_24_896 ();
 sg13g2_decap_8 FILLER_24_903 ();
 sg13g2_decap_8 FILLER_24_910 ();
 sg13g2_decap_8 FILLER_24_917 ();
 sg13g2_decap_8 FILLER_24_924 ();
 sg13g2_decap_8 FILLER_24_931 ();
 sg13g2_decap_8 FILLER_24_938 ();
 sg13g2_decap_8 FILLER_24_945 ();
 sg13g2_decap_8 FILLER_24_952 ();
 sg13g2_decap_8 FILLER_24_959 ();
 sg13g2_decap_8 FILLER_24_966 ();
 sg13g2_decap_8 FILLER_24_973 ();
 sg13g2_decap_8 FILLER_24_980 ();
 sg13g2_decap_8 FILLER_24_987 ();
 sg13g2_decap_8 FILLER_24_994 ();
 sg13g2_decap_8 FILLER_24_1001 ();
 sg13g2_decap_8 FILLER_24_1008 ();
 sg13g2_decap_8 FILLER_24_1015 ();
 sg13g2_decap_8 FILLER_24_1022 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_29 ();
 sg13g2_decap_4 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_8 FILLER_25_134 ();
 sg13g2_decap_8 FILLER_25_141 ();
 sg13g2_decap_8 FILLER_25_148 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_436 ();
 sg13g2_decap_4 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_447 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_fill_1 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_484 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_8 FILLER_25_512 ();
 sg13g2_fill_2 FILLER_25_519 ();
 sg13g2_decap_8 FILLER_25_533 ();
 sg13g2_decap_8 FILLER_25_540 ();
 sg13g2_decap_4 FILLER_25_547 ();
 sg13g2_fill_1 FILLER_25_551 ();
 sg13g2_decap_4 FILLER_25_556 ();
 sg13g2_fill_2 FILLER_25_564 ();
 sg13g2_fill_1 FILLER_25_566 ();
 sg13g2_decap_8 FILLER_25_576 ();
 sg13g2_decap_8 FILLER_25_583 ();
 sg13g2_decap_8 FILLER_25_590 ();
 sg13g2_fill_2 FILLER_25_597 ();
 sg13g2_fill_2 FILLER_25_612 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_fill_1 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_fill_2 FILLER_25_693 ();
 sg13g2_fill_1 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_4 FILLER_25_749 ();
 sg13g2_fill_1 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_766 ();
 sg13g2_decap_8 FILLER_25_773 ();
 sg13g2_fill_2 FILLER_25_780 ();
 sg13g2_fill_2 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_822 ();
 sg13g2_fill_2 FILLER_25_829 ();
 sg13g2_decap_8 FILLER_25_859 ();
 sg13g2_decap_8 FILLER_25_866 ();
 sg13g2_decap_8 FILLER_25_873 ();
 sg13g2_decap_8 FILLER_25_880 ();
 sg13g2_decap_8 FILLER_25_887 ();
 sg13g2_decap_8 FILLER_25_894 ();
 sg13g2_decap_8 FILLER_25_901 ();
 sg13g2_decap_8 FILLER_25_908 ();
 sg13g2_decap_8 FILLER_25_915 ();
 sg13g2_decap_8 FILLER_25_922 ();
 sg13g2_decap_8 FILLER_25_929 ();
 sg13g2_decap_8 FILLER_25_936 ();
 sg13g2_decap_8 FILLER_25_943 ();
 sg13g2_decap_8 FILLER_25_950 ();
 sg13g2_decap_8 FILLER_25_957 ();
 sg13g2_decap_8 FILLER_25_964 ();
 sg13g2_decap_8 FILLER_25_971 ();
 sg13g2_decap_8 FILLER_25_978 ();
 sg13g2_decap_8 FILLER_25_985 ();
 sg13g2_decap_8 FILLER_25_992 ();
 sg13g2_decap_8 FILLER_25_999 ();
 sg13g2_decap_8 FILLER_25_1006 ();
 sg13g2_decap_8 FILLER_25_1013 ();
 sg13g2_decap_8 FILLER_25_1020 ();
 sg13g2_fill_2 FILLER_25_1027 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_4 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_439 ();
 sg13g2_decap_8 FILLER_26_446 ();
 sg13g2_decap_8 FILLER_26_453 ();
 sg13g2_fill_2 FILLER_26_460 ();
 sg13g2_fill_1 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_473 ();
 sg13g2_fill_1 FILLER_26_492 ();
 sg13g2_decap_8 FILLER_26_537 ();
 sg13g2_decap_4 FILLER_26_544 ();
 sg13g2_fill_1 FILLER_26_548 ();
 sg13g2_decap_8 FILLER_26_557 ();
 sg13g2_decap_8 FILLER_26_564 ();
 sg13g2_fill_2 FILLER_26_571 ();
 sg13g2_fill_1 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_fill_2 FILLER_26_586 ();
 sg13g2_decap_4 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_604 ();
 sg13g2_fill_2 FILLER_26_611 ();
 sg13g2_fill_1 FILLER_26_613 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_4 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_fill_1 FILLER_26_684 ();
 sg13g2_fill_2 FILLER_26_703 ();
 sg13g2_fill_2 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_4 FILLER_26_742 ();
 sg13g2_fill_2 FILLER_26_749 ();
 sg13g2_fill_1 FILLER_26_751 ();
 sg13g2_fill_2 FILLER_26_775 ();
 sg13g2_fill_2 FILLER_26_790 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_fill_2 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_836 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_8 FILLER_26_850 ();
 sg13g2_decap_8 FILLER_26_857 ();
 sg13g2_decap_8 FILLER_26_864 ();
 sg13g2_decap_8 FILLER_26_871 ();
 sg13g2_decap_8 FILLER_26_878 ();
 sg13g2_decap_8 FILLER_26_885 ();
 sg13g2_decap_8 FILLER_26_892 ();
 sg13g2_decap_8 FILLER_26_899 ();
 sg13g2_decap_8 FILLER_26_906 ();
 sg13g2_decap_8 FILLER_26_913 ();
 sg13g2_decap_8 FILLER_26_920 ();
 sg13g2_decap_8 FILLER_26_927 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_941 ();
 sg13g2_decap_8 FILLER_26_948 ();
 sg13g2_decap_8 FILLER_26_955 ();
 sg13g2_decap_8 FILLER_26_962 ();
 sg13g2_decap_8 FILLER_26_969 ();
 sg13g2_decap_8 FILLER_26_976 ();
 sg13g2_decap_8 FILLER_26_983 ();
 sg13g2_decap_8 FILLER_26_990 ();
 sg13g2_decap_8 FILLER_26_997 ();
 sg13g2_decap_8 FILLER_26_1004 ();
 sg13g2_decap_8 FILLER_26_1011 ();
 sg13g2_decap_8 FILLER_26_1018 ();
 sg13g2_decap_4 FILLER_26_1025 ();
 sg13g2_decap_4 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_8 ();
 sg13g2_decap_8 FILLER_27_13 ();
 sg13g2_fill_1 FILLER_27_33 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_80 ();
 sg13g2_decap_4 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_decap_8 FILLER_27_424 ();
 sg13g2_decap_8 FILLER_27_431 ();
 sg13g2_decap_4 FILLER_27_438 ();
 sg13g2_fill_2 FILLER_27_442 ();
 sg13g2_decap_8 FILLER_27_472 ();
 sg13g2_decap_4 FILLER_27_479 ();
 sg13g2_fill_1 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_4 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_533 ();
 sg13g2_fill_2 FILLER_27_540 ();
 sg13g2_fill_1 FILLER_27_562 ();
 sg13g2_decap_4 FILLER_27_576 ();
 sg13g2_fill_2 FILLER_27_580 ();
 sg13g2_fill_2 FILLER_27_607 ();
 sg13g2_fill_2 FILLER_27_621 ();
 sg13g2_decap_8 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_638 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_4 FILLER_27_651 ();
 sg13g2_fill_2 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_670 ();
 sg13g2_decap_4 FILLER_27_677 ();
 sg13g2_fill_1 FILLER_27_681 ();
 sg13g2_decap_4 FILLER_27_749 ();
 sg13g2_fill_1 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_781 ();
 sg13g2_decap_4 FILLER_27_788 ();
 sg13g2_fill_1 FILLER_27_792 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_68 ();
 sg13g2_decap_8 FILLER_28_75 ();
 sg13g2_decap_8 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_89 ();
 sg13g2_decap_8 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_460 ();
 sg13g2_decap_8 FILLER_28_467 ();
 sg13g2_decap_8 FILLER_28_474 ();
 sg13g2_decap_8 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_488 ();
 sg13g2_decap_4 FILLER_28_495 ();
 sg13g2_decap_8 FILLER_28_507 ();
 sg13g2_decap_8 FILLER_28_514 ();
 sg13g2_decap_8 FILLER_28_521 ();
 sg13g2_decap_8 FILLER_28_528 ();
 sg13g2_decap_8 FILLER_28_556 ();
 sg13g2_decap_8 FILLER_28_563 ();
 sg13g2_decap_8 FILLER_28_570 ();
 sg13g2_decap_8 FILLER_28_577 ();
 sg13g2_fill_2 FILLER_28_584 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_4 FILLER_28_609 ();
 sg13g2_fill_2 FILLER_28_613 ();
 sg13g2_decap_4 FILLER_28_628 ();
 sg13g2_fill_2 FILLER_28_632 ();
 sg13g2_decap_8 FILLER_28_640 ();
 sg13g2_decap_8 FILLER_28_647 ();
 sg13g2_fill_1 FILLER_28_654 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_fill_2 FILLER_28_704 ();
 sg13g2_fill_1 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_fill_1 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_4 FILLER_28_753 ();
 sg13g2_fill_1 FILLER_28_757 ();
 sg13g2_decap_8 FILLER_28_775 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_decap_4 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_decap_8 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_decap_8 FILLER_28_876 ();
 sg13g2_decap_8 FILLER_28_883 ();
 sg13g2_decap_8 FILLER_28_890 ();
 sg13g2_decap_8 FILLER_28_897 ();
 sg13g2_decap_8 FILLER_28_904 ();
 sg13g2_decap_8 FILLER_28_911 ();
 sg13g2_decap_8 FILLER_28_918 ();
 sg13g2_decap_8 FILLER_28_925 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_8 FILLER_28_939 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_decap_8 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_28_1002 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_decap_4 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_8 ();
 sg13g2_decap_8 FILLER_29_13 ();
 sg13g2_fill_2 FILLER_29_20 ();
 sg13g2_decap_4 FILLER_29_39 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_4 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_4 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_fill_2 FILLER_29_405 ();
 sg13g2_fill_1 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_29_436 ();
 sg13g2_fill_2 FILLER_29_466 ();
 sg13g2_fill_1 FILLER_29_468 ();
 sg13g2_decap_4 FILLER_29_482 ();
 sg13g2_fill_1 FILLER_29_486 ();
 sg13g2_fill_2 FILLER_29_493 ();
 sg13g2_fill_1 FILLER_29_495 ();
 sg13g2_decap_8 FILLER_29_530 ();
 sg13g2_decap_8 FILLER_29_537 ();
 sg13g2_fill_2 FILLER_29_544 ();
 sg13g2_decap_4 FILLER_29_560 ();
 sg13g2_fill_2 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_fill_2 FILLER_29_595 ();
 sg13g2_fill_1 FILLER_29_597 ();
 sg13g2_decap_8 FILLER_29_608 ();
 sg13g2_fill_2 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_617 ();
 sg13g2_decap_4 FILLER_29_627 ();
 sg13g2_fill_1 FILLER_29_631 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_fill_2 FILLER_29_651 ();
 sg13g2_fill_1 FILLER_29_653 ();
 sg13g2_fill_1 FILLER_29_659 ();
 sg13g2_decap_8 FILLER_29_664 ();
 sg13g2_decap_8 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_717 ();
 sg13g2_decap_4 FILLER_29_738 ();
 sg13g2_fill_2 FILLER_29_742 ();
 sg13g2_fill_1 FILLER_29_752 ();
 sg13g2_fill_2 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_773 ();
 sg13g2_decap_8 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_787 ();
 sg13g2_decap_8 FILLER_29_794 ();
 sg13g2_decap_8 FILLER_29_801 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_8 FILLER_29_857 ();
 sg13g2_decap_8 FILLER_29_864 ();
 sg13g2_decap_8 FILLER_29_871 ();
 sg13g2_decap_8 FILLER_29_878 ();
 sg13g2_decap_8 FILLER_29_885 ();
 sg13g2_decap_8 FILLER_29_892 ();
 sg13g2_decap_8 FILLER_29_899 ();
 sg13g2_decap_8 FILLER_29_906 ();
 sg13g2_decap_8 FILLER_29_913 ();
 sg13g2_decap_8 FILLER_29_920 ();
 sg13g2_decap_8 FILLER_29_927 ();
 sg13g2_decap_8 FILLER_29_934 ();
 sg13g2_decap_8 FILLER_29_941 ();
 sg13g2_decap_8 FILLER_29_948 ();
 sg13g2_decap_8 FILLER_29_955 ();
 sg13g2_decap_8 FILLER_29_962 ();
 sg13g2_decap_8 FILLER_29_969 ();
 sg13g2_decap_8 FILLER_29_976 ();
 sg13g2_decap_8 FILLER_29_983 ();
 sg13g2_decap_8 FILLER_29_990 ();
 sg13g2_decap_8 FILLER_29_997 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_decap_8 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1018 ();
 sg13g2_decap_4 FILLER_29_1025 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_76 ();
 sg13g2_decap_8 FILLER_30_83 ();
 sg13g2_decap_8 FILLER_30_90 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_decap_4 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_decap_4 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_397 ();
 sg13g2_fill_2 FILLER_30_418 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_438 ();
 sg13g2_fill_2 FILLER_30_445 ();
 sg13g2_decap_8 FILLER_30_463 ();
 sg13g2_decap_8 FILLER_30_470 ();
 sg13g2_decap_8 FILLER_30_477 ();
 sg13g2_decap_4 FILLER_30_492 ();
 sg13g2_fill_1 FILLER_30_496 ();
 sg13g2_fill_1 FILLER_30_510 ();
 sg13g2_decap_8 FILLER_30_533 ();
 sg13g2_fill_1 FILLER_30_540 ();
 sg13g2_decap_8 FILLER_30_554 ();
 sg13g2_decap_8 FILLER_30_561 ();
 sg13g2_decap_8 FILLER_30_568 ();
 sg13g2_decap_8 FILLER_30_575 ();
 sg13g2_decap_8 FILLER_30_582 ();
 sg13g2_decap_4 FILLER_30_589 ();
 sg13g2_fill_2 FILLER_30_593 ();
 sg13g2_decap_8 FILLER_30_617 ();
 sg13g2_fill_1 FILLER_30_624 ();
 sg13g2_fill_1 FILLER_30_654 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_fill_1 FILLER_30_681 ();
 sg13g2_fill_2 FILLER_30_710 ();
 sg13g2_fill_1 FILLER_30_712 ();
 sg13g2_fill_1 FILLER_30_741 ();
 sg13g2_decap_8 FILLER_30_783 ();
 sg13g2_decap_8 FILLER_30_790 ();
 sg13g2_decap_8 FILLER_30_797 ();
 sg13g2_decap_8 FILLER_30_804 ();
 sg13g2_decap_8 FILLER_30_811 ();
 sg13g2_decap_8 FILLER_30_818 ();
 sg13g2_decap_8 FILLER_30_825 ();
 sg13g2_decap_8 FILLER_30_832 ();
 sg13g2_decap_8 FILLER_30_839 ();
 sg13g2_decap_8 FILLER_30_846 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_decap_8 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_867 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_decap_8 FILLER_30_881 ();
 sg13g2_decap_8 FILLER_30_888 ();
 sg13g2_decap_8 FILLER_30_895 ();
 sg13g2_decap_8 FILLER_30_902 ();
 sg13g2_decap_8 FILLER_30_909 ();
 sg13g2_decap_8 FILLER_30_916 ();
 sg13g2_decap_8 FILLER_30_923 ();
 sg13g2_decap_8 FILLER_30_930 ();
 sg13g2_decap_8 FILLER_30_937 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_decap_8 FILLER_30_951 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_decap_8 FILLER_30_965 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_986 ();
 sg13g2_decap_8 FILLER_30_993 ();
 sg13g2_decap_8 FILLER_30_1000 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_8 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1021 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_248 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_4 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_360 ();
 sg13g2_decap_4 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_387 ();
 sg13g2_decap_4 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_443 ();
 sg13g2_decap_8 FILLER_31_459 ();
 sg13g2_decap_8 FILLER_31_472 ();
 sg13g2_decap_4 FILLER_31_479 ();
 sg13g2_fill_1 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_496 ();
 sg13g2_decap_4 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_507 ();
 sg13g2_decap_8 FILLER_31_517 ();
 sg13g2_decap_8 FILLER_31_524 ();
 sg13g2_decap_8 FILLER_31_531 ();
 sg13g2_fill_2 FILLER_31_542 ();
 sg13g2_fill_1 FILLER_31_544 ();
 sg13g2_fill_1 FILLER_31_548 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_4 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_585 ();
 sg13g2_decap_4 FILLER_31_592 ();
 sg13g2_fill_1 FILLER_31_596 ();
 sg13g2_decap_8 FILLER_31_618 ();
 sg13g2_decap_8 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_632 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_fill_1 FILLER_31_640 ();
 sg13g2_fill_1 FILLER_31_663 ();
 sg13g2_decap_4 FILLER_31_672 ();
 sg13g2_fill_1 FILLER_31_686 ();
 sg13g2_fill_1 FILLER_31_691 ();
 sg13g2_decap_8 FILLER_31_698 ();
 sg13g2_decap_8 FILLER_31_705 ();
 sg13g2_decap_8 FILLER_31_712 ();
 sg13g2_decap_8 FILLER_31_719 ();
 sg13g2_fill_1 FILLER_31_726 ();
 sg13g2_decap_4 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_8 FILLER_31_856 ();
 sg13g2_decap_8 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_870 ();
 sg13g2_decap_8 FILLER_31_877 ();
 sg13g2_decap_8 FILLER_31_884 ();
 sg13g2_decap_8 FILLER_31_891 ();
 sg13g2_decap_8 FILLER_31_898 ();
 sg13g2_decap_8 FILLER_31_905 ();
 sg13g2_decap_8 FILLER_31_912 ();
 sg13g2_decap_8 FILLER_31_919 ();
 sg13g2_decap_8 FILLER_31_926 ();
 sg13g2_decap_8 FILLER_31_933 ();
 sg13g2_decap_8 FILLER_31_940 ();
 sg13g2_decap_8 FILLER_31_947 ();
 sg13g2_decap_8 FILLER_31_954 ();
 sg13g2_decap_8 FILLER_31_961 ();
 sg13g2_decap_8 FILLER_31_968 ();
 sg13g2_decap_8 FILLER_31_975 ();
 sg13g2_decap_8 FILLER_31_982 ();
 sg13g2_decap_8 FILLER_31_989 ();
 sg13g2_decap_8 FILLER_31_996 ();
 sg13g2_decap_8 FILLER_31_1003 ();
 sg13g2_decap_8 FILLER_31_1010 ();
 sg13g2_decap_8 FILLER_31_1017 ();
 sg13g2_decap_4 FILLER_31_1024 ();
 sg13g2_fill_1 FILLER_31_1028 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_decap_8 FILLER_32_36 ();
 sg13g2_fill_2 FILLER_32_43 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_decap_4 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_405 ();
 sg13g2_decap_4 FILLER_32_411 ();
 sg13g2_decap_8 FILLER_32_439 ();
 sg13g2_decap_8 FILLER_32_446 ();
 sg13g2_fill_2 FILLER_32_453 ();
 sg13g2_decap_4 FILLER_32_459 ();
 sg13g2_decap_8 FILLER_32_474 ();
 sg13g2_decap_8 FILLER_32_481 ();
 sg13g2_fill_1 FILLER_32_488 ();
 sg13g2_decap_4 FILLER_32_501 ();
 sg13g2_fill_2 FILLER_32_505 ();
 sg13g2_fill_1 FILLER_32_528 ();
 sg13g2_decap_8 FILLER_32_555 ();
 sg13g2_fill_2 FILLER_32_562 ();
 sg13g2_fill_1 FILLER_32_564 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_4 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_fill_2 FILLER_32_630 ();
 sg13g2_decap_4 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_677 ();
 sg13g2_decap_8 FILLER_32_684 ();
 sg13g2_decap_8 FILLER_32_691 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_decap_4 FILLER_32_705 ();
 sg13g2_fill_1 FILLER_32_709 ();
 sg13g2_decap_8 FILLER_32_727 ();
 sg13g2_decap_4 FILLER_32_734 ();
 sg13g2_fill_2 FILLER_32_738 ();
 sg13g2_fill_2 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_828 ();
 sg13g2_decap_8 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_842 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_8 FILLER_32_856 ();
 sg13g2_decap_8 FILLER_32_863 ();
 sg13g2_decap_8 FILLER_32_870 ();
 sg13g2_decap_8 FILLER_32_877 ();
 sg13g2_decap_8 FILLER_32_884 ();
 sg13g2_decap_8 FILLER_32_891 ();
 sg13g2_decap_8 FILLER_32_898 ();
 sg13g2_decap_8 FILLER_32_905 ();
 sg13g2_decap_8 FILLER_32_912 ();
 sg13g2_decap_8 FILLER_32_919 ();
 sg13g2_decap_8 FILLER_32_926 ();
 sg13g2_decap_8 FILLER_32_933 ();
 sg13g2_decap_8 FILLER_32_940 ();
 sg13g2_decap_8 FILLER_32_947 ();
 sg13g2_decap_8 FILLER_32_954 ();
 sg13g2_decap_8 FILLER_32_961 ();
 sg13g2_decap_8 FILLER_32_968 ();
 sg13g2_decap_8 FILLER_32_975 ();
 sg13g2_decap_8 FILLER_32_982 ();
 sg13g2_decap_8 FILLER_32_989 ();
 sg13g2_decap_8 FILLER_32_996 ();
 sg13g2_decap_8 FILLER_32_1003 ();
 sg13g2_decap_8 FILLER_32_1010 ();
 sg13g2_decap_8 FILLER_32_1017 ();
 sg13g2_decap_4 FILLER_32_1024 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_13 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_decap_4 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_8 FILLER_33_404 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_decap_4 FILLER_33_421 ();
 sg13g2_decap_4 FILLER_33_430 ();
 sg13g2_decap_4 FILLER_33_447 ();
 sg13g2_decap_8 FILLER_33_474 ();
 sg13g2_decap_8 FILLER_33_481 ();
 sg13g2_fill_2 FILLER_33_488 ();
 sg13g2_decap_8 FILLER_33_503 ();
 sg13g2_decap_8 FILLER_33_510 ();
 sg13g2_decap_8 FILLER_33_517 ();
 sg13g2_fill_2 FILLER_33_534 ();
 sg13g2_fill_1 FILLER_33_536 ();
 sg13g2_fill_2 FILLER_33_541 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_fill_2 FILLER_33_555 ();
 sg13g2_decap_8 FILLER_33_563 ();
 sg13g2_decap_8 FILLER_33_570 ();
 sg13g2_decap_8 FILLER_33_582 ();
 sg13g2_decap_8 FILLER_33_589 ();
 sg13g2_decap_4 FILLER_33_596 ();
 sg13g2_fill_2 FILLER_33_600 ();
 sg13g2_decap_8 FILLER_33_614 ();
 sg13g2_decap_8 FILLER_33_621 ();
 sg13g2_decap_4 FILLER_33_628 ();
 sg13g2_fill_1 FILLER_33_640 ();
 sg13g2_decap_8 FILLER_33_649 ();
 sg13g2_decap_8 FILLER_33_656 ();
 sg13g2_decap_8 FILLER_33_663 ();
 sg13g2_fill_2 FILLER_33_670 ();
 sg13g2_fill_1 FILLER_33_682 ();
 sg13g2_decap_8 FILLER_33_711 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_4 FILLER_33_753 ();
 sg13g2_fill_1 FILLER_33_757 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_8 FILLER_33_783 ();
 sg13g2_decap_8 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_797 ();
 sg13g2_decap_8 FILLER_33_804 ();
 sg13g2_decap_8 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_853 ();
 sg13g2_decap_8 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_33_867 ();
 sg13g2_decap_8 FILLER_33_874 ();
 sg13g2_decap_8 FILLER_33_881 ();
 sg13g2_decap_8 FILLER_33_888 ();
 sg13g2_decap_8 FILLER_33_895 ();
 sg13g2_decap_8 FILLER_33_902 ();
 sg13g2_decap_8 FILLER_33_909 ();
 sg13g2_decap_8 FILLER_33_916 ();
 sg13g2_decap_8 FILLER_33_923 ();
 sg13g2_decap_8 FILLER_33_930 ();
 sg13g2_decap_8 FILLER_33_937 ();
 sg13g2_decap_8 FILLER_33_944 ();
 sg13g2_decap_8 FILLER_33_951 ();
 sg13g2_decap_8 FILLER_33_958 ();
 sg13g2_decap_8 FILLER_33_965 ();
 sg13g2_decap_8 FILLER_33_972 ();
 sg13g2_decap_8 FILLER_33_979 ();
 sg13g2_decap_8 FILLER_33_986 ();
 sg13g2_decap_8 FILLER_33_993 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_decap_8 FILLER_33_1007 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_decap_8 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_decap_4 FILLER_34_234 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_decap_8 FILLER_34_323 ();
 sg13g2_decap_8 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_4 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_8 FILLER_34_426 ();
 sg13g2_decap_8 FILLER_34_433 ();
 sg13g2_decap_8 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_447 ();
 sg13g2_decap_4 FILLER_34_454 ();
 sg13g2_fill_2 FILLER_34_458 ();
 sg13g2_fill_1 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_478 ();
 sg13g2_decap_4 FILLER_34_485 ();
 sg13g2_fill_2 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_508 ();
 sg13g2_decap_8 FILLER_34_515 ();
 sg13g2_decap_4 FILLER_34_522 ();
 sg13g2_fill_1 FILLER_34_526 ();
 sg13g2_fill_1 FILLER_34_537 ();
 sg13g2_decap_4 FILLER_34_542 ();
 sg13g2_fill_2 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_fill_2 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_599 ();
 sg13g2_decap_8 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_613 ();
 sg13g2_decap_4 FILLER_34_620 ();
 sg13g2_fill_2 FILLER_34_624 ();
 sg13g2_fill_2 FILLER_34_634 ();
 sg13g2_fill_1 FILLER_34_636 ();
 sg13g2_decap_8 FILLER_34_645 ();
 sg13g2_decap_8 FILLER_34_652 ();
 sg13g2_decap_8 FILLER_34_659 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_fill_2 FILLER_34_686 ();
 sg13g2_fill_1 FILLER_34_688 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_fill_2 FILLER_34_707 ();
 sg13g2_fill_1 FILLER_34_709 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_fill_2 FILLER_34_737 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_8 FILLER_34_896 ();
 sg13g2_decap_8 FILLER_34_903 ();
 sg13g2_decap_8 FILLER_34_910 ();
 sg13g2_decap_8 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_13 ();
 sg13g2_fill_2 FILLER_35_17 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_34 ();
 sg13g2_decap_4 FILLER_35_41 ();
 sg13g2_decap_4 FILLER_35_54 ();
 sg13g2_fill_2 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_fill_2 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_129 ();
 sg13g2_fill_2 FILLER_35_136 ();
 sg13g2_fill_1 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_4 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_2 FILLER_35_387 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_447 ();
 sg13g2_decap_4 FILLER_35_454 ();
 sg13g2_decap_8 FILLER_35_474 ();
 sg13g2_decap_4 FILLER_35_481 ();
 sg13g2_fill_1 FILLER_35_485 ();
 sg13g2_decap_4 FILLER_35_513 ();
 sg13g2_fill_1 FILLER_35_517 ();
 sg13g2_fill_2 FILLER_35_523 ();
 sg13g2_fill_1 FILLER_35_525 ();
 sg13g2_fill_2 FILLER_35_538 ();
 sg13g2_fill_2 FILLER_35_549 ();
 sg13g2_fill_1 FILLER_35_551 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_decap_8 FILLER_35_572 ();
 sg13g2_decap_8 FILLER_35_579 ();
 sg13g2_decap_8 FILLER_35_586 ();
 sg13g2_fill_2 FILLER_35_593 ();
 sg13g2_decap_8 FILLER_35_599 ();
 sg13g2_decap_8 FILLER_35_606 ();
 sg13g2_decap_8 FILLER_35_613 ();
 sg13g2_decap_4 FILLER_35_620 ();
 sg13g2_fill_1 FILLER_35_639 ();
 sg13g2_decap_4 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_648 ();
 sg13g2_decap_4 FILLER_35_653 ();
 sg13g2_fill_1 FILLER_35_657 ();
 sg13g2_decap_4 FILLER_35_667 ();
 sg13g2_fill_2 FILLER_35_671 ();
 sg13g2_decap_4 FILLER_35_686 ();
 sg13g2_fill_1 FILLER_35_690 ();
 sg13g2_decap_4 FILLER_35_700 ();
 sg13g2_fill_2 FILLER_35_704 ();
 sg13g2_decap_4 FILLER_35_724 ();
 sg13g2_fill_1 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_fill_2 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_8 FILLER_35_857 ();
 sg13g2_decap_8 FILLER_35_864 ();
 sg13g2_decap_8 FILLER_35_871 ();
 sg13g2_decap_8 FILLER_35_878 ();
 sg13g2_decap_8 FILLER_35_885 ();
 sg13g2_decap_8 FILLER_35_892 ();
 sg13g2_decap_8 FILLER_35_899 ();
 sg13g2_decap_8 FILLER_35_906 ();
 sg13g2_decap_8 FILLER_35_913 ();
 sg13g2_decap_8 FILLER_35_920 ();
 sg13g2_decap_8 FILLER_35_927 ();
 sg13g2_decap_8 FILLER_35_934 ();
 sg13g2_decap_8 FILLER_35_941 ();
 sg13g2_decap_8 FILLER_35_948 ();
 sg13g2_decap_8 FILLER_35_955 ();
 sg13g2_decap_8 FILLER_35_962 ();
 sg13g2_decap_8 FILLER_35_969 ();
 sg13g2_decap_8 FILLER_35_976 ();
 sg13g2_decap_8 FILLER_35_983 ();
 sg13g2_decap_8 FILLER_35_990 ();
 sg13g2_decap_8 FILLER_35_997 ();
 sg13g2_decap_8 FILLER_35_1004 ();
 sg13g2_decap_8 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1018 ();
 sg13g2_decap_4 FILLER_35_1025 ();
 sg13g2_fill_2 FILLER_36_27 ();
 sg13g2_fill_1 FILLER_36_29 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_78 ();
 sg13g2_decap_4 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_97 ();
 sg13g2_fill_2 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_decap_4 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_decap_4 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_fill_1 FILLER_36_411 ();
 sg13g2_decap_8 FILLER_36_416 ();
 sg13g2_decap_4 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_fill_2 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_483 ();
 sg13g2_decap_4 FILLER_36_496 ();
 sg13g2_decap_8 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_520 ();
 sg13g2_fill_2 FILLER_36_527 ();
 sg13g2_decap_8 FILLER_36_534 ();
 sg13g2_decap_8 FILLER_36_541 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_decap_8 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_decap_4 FILLER_36_576 ();
 sg13g2_decap_4 FILLER_36_584 ();
 sg13g2_fill_2 FILLER_36_588 ();
 sg13g2_fill_2 FILLER_36_618 ();
 sg13g2_fill_1 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_627 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_fill_2 FILLER_36_652 ();
 sg13g2_fill_2 FILLER_36_659 ();
 sg13g2_fill_1 FILLER_36_661 ();
 sg13g2_fill_2 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_683 ();
 sg13g2_decap_4 FILLER_36_690 ();
 sg13g2_decap_8 FILLER_36_734 ();
 sg13g2_decap_8 FILLER_36_741 ();
 sg13g2_decap_8 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_8 FILLER_36_835 ();
 sg13g2_decap_8 FILLER_36_842 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_8 FILLER_36_856 ();
 sg13g2_decap_8 FILLER_36_863 ();
 sg13g2_decap_8 FILLER_36_870 ();
 sg13g2_decap_8 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_36_884 ();
 sg13g2_decap_8 FILLER_36_891 ();
 sg13g2_decap_8 FILLER_36_898 ();
 sg13g2_decap_8 FILLER_36_905 ();
 sg13g2_decap_8 FILLER_36_912 ();
 sg13g2_decap_8 FILLER_36_919 ();
 sg13g2_decap_8 FILLER_36_926 ();
 sg13g2_decap_8 FILLER_36_933 ();
 sg13g2_decap_8 FILLER_36_940 ();
 sg13g2_decap_8 FILLER_36_947 ();
 sg13g2_decap_8 FILLER_36_954 ();
 sg13g2_decap_8 FILLER_36_961 ();
 sg13g2_decap_8 FILLER_36_968 ();
 sg13g2_decap_8 FILLER_36_975 ();
 sg13g2_decap_8 FILLER_36_982 ();
 sg13g2_decap_8 FILLER_36_989 ();
 sg13g2_decap_8 FILLER_36_996 ();
 sg13g2_decap_8 FILLER_36_1003 ();
 sg13g2_decap_8 FILLER_36_1010 ();
 sg13g2_decap_8 FILLER_36_1017 ();
 sg13g2_decap_4 FILLER_36_1024 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_13 ();
 sg13g2_fill_1 FILLER_37_20 ();
 sg13g2_fill_2 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_decap_4 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_265 ();
 sg13g2_decap_8 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_279 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_decap_4 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_decap_4 FILLER_37_353 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_fill_2 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_444 ();
 sg13g2_decap_8 FILLER_37_451 ();
 sg13g2_decap_8 FILLER_37_458 ();
 sg13g2_decap_8 FILLER_37_478 ();
 sg13g2_decap_8 FILLER_37_485 ();
 sg13g2_decap_8 FILLER_37_492 ();
 sg13g2_decap_4 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_503 ();
 sg13g2_decap_8 FILLER_37_519 ();
 sg13g2_decap_8 FILLER_37_526 ();
 sg13g2_decap_8 FILLER_37_533 ();
 sg13g2_decap_8 FILLER_37_540 ();
 sg13g2_decap_8 FILLER_37_547 ();
 sg13g2_decap_8 FILLER_37_554 ();
 sg13g2_fill_2 FILLER_37_561 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_fill_2 FILLER_37_595 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_fill_2 FILLER_37_612 ();
 sg13g2_fill_1 FILLER_37_614 ();
 sg13g2_decap_8 FILLER_37_628 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_2 FILLER_37_639 ();
 sg13g2_decap_8 FILLER_37_652 ();
 sg13g2_decap_8 FILLER_37_659 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_decap_8 FILLER_37_684 ();
 sg13g2_decap_4 FILLER_37_691 ();
 sg13g2_fill_1 FILLER_37_695 ();
 sg13g2_decap_8 FILLER_37_705 ();
 sg13g2_decap_8 FILLER_37_712 ();
 sg13g2_decap_8 FILLER_37_719 ();
 sg13g2_fill_1 FILLER_37_726 ();
 sg13g2_fill_2 FILLER_37_744 ();
 sg13g2_decap_8 FILLER_37_774 ();
 sg13g2_decap_8 FILLER_37_781 ();
 sg13g2_decap_8 FILLER_37_788 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_816 ();
 sg13g2_decap_8 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_858 ();
 sg13g2_decap_8 FILLER_37_865 ();
 sg13g2_decap_8 FILLER_37_872 ();
 sg13g2_decap_8 FILLER_37_879 ();
 sg13g2_decap_8 FILLER_37_886 ();
 sg13g2_decap_8 FILLER_37_893 ();
 sg13g2_decap_8 FILLER_37_900 ();
 sg13g2_decap_8 FILLER_37_907 ();
 sg13g2_decap_8 FILLER_37_914 ();
 sg13g2_decap_8 FILLER_37_921 ();
 sg13g2_decap_8 FILLER_37_928 ();
 sg13g2_decap_8 FILLER_37_935 ();
 sg13g2_decap_8 FILLER_37_942 ();
 sg13g2_decap_8 FILLER_37_949 ();
 sg13g2_decap_8 FILLER_37_956 ();
 sg13g2_decap_8 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_970 ();
 sg13g2_decap_8 FILLER_37_977 ();
 sg13g2_decap_8 FILLER_37_984 ();
 sg13g2_decap_8 FILLER_37_991 ();
 sg13g2_decap_8 FILLER_37_998 ();
 sg13g2_decap_8 FILLER_37_1005 ();
 sg13g2_decap_8 FILLER_37_1012 ();
 sg13g2_decap_8 FILLER_37_1019 ();
 sg13g2_fill_2 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_34 ();
 sg13g2_fill_1 FILLER_38_36 ();
 sg13g2_decap_4 FILLER_38_69 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_107 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_4 FILLER_38_379 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_425 ();
 sg13g2_decap_8 FILLER_38_437 ();
 sg13g2_decap_8 FILLER_38_444 ();
 sg13g2_decap_8 FILLER_38_451 ();
 sg13g2_fill_2 FILLER_38_458 ();
 sg13g2_fill_1 FILLER_38_460 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_fill_2 FILLER_38_490 ();
 sg13g2_fill_1 FILLER_38_497 ();
 sg13g2_fill_2 FILLER_38_508 ();
 sg13g2_fill_1 FILLER_38_510 ();
 sg13g2_decap_8 FILLER_38_526 ();
 sg13g2_fill_1 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_559 ();
 sg13g2_decap_8 FILLER_38_566 ();
 sg13g2_fill_2 FILLER_38_573 ();
 sg13g2_decap_8 FILLER_38_593 ();
 sg13g2_fill_2 FILLER_38_600 ();
 sg13g2_fill_1 FILLER_38_602 ();
 sg13g2_fill_2 FILLER_38_615 ();
 sg13g2_fill_1 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_626 ();
 sg13g2_decap_8 FILLER_38_633 ();
 sg13g2_decap_8 FILLER_38_640 ();
 sg13g2_fill_2 FILLER_38_647 ();
 sg13g2_fill_2 FILLER_38_655 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_decap_4 FILLER_38_662 ();
 sg13g2_fill_2 FILLER_38_666 ();
 sg13g2_fill_2 FILLER_38_671 ();
 sg13g2_fill_1 FILLER_38_673 ();
 sg13g2_decap_8 FILLER_38_678 ();
 sg13g2_fill_2 FILLER_38_685 ();
 sg13g2_fill_1 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_716 ();
 sg13g2_decap_8 FILLER_38_723 ();
 sg13g2_decap_8 FILLER_38_730 ();
 sg13g2_decap_8 FILLER_38_737 ();
 sg13g2_decap_8 FILLER_38_744 ();
 sg13g2_fill_2 FILLER_38_751 ();
 sg13g2_fill_1 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_37 ();
 sg13g2_decap_4 FILLER_39_44 ();
 sg13g2_fill_1 FILLER_39_48 ();
 sg13g2_decap_4 FILLER_39_58 ();
 sg13g2_fill_1 FILLER_39_62 ();
 sg13g2_decap_8 FILLER_39_76 ();
 sg13g2_decap_8 FILLER_39_83 ();
 sg13g2_decap_8 FILLER_39_90 ();
 sg13g2_decap_8 FILLER_39_97 ();
 sg13g2_decap_4 FILLER_39_104 ();
 sg13g2_fill_2 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_123 ();
 sg13g2_fill_1 FILLER_39_125 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_4 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_262 ();
 sg13g2_decap_8 FILLER_39_269 ();
 sg13g2_fill_2 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_300 ();
 sg13g2_decap_8 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_fill_2 FILLER_39_387 ();
 sg13g2_fill_1 FILLER_39_394 ();
 sg13g2_decap_4 FILLER_39_399 ();
 sg13g2_fill_2 FILLER_39_403 ();
 sg13g2_decap_8 FILLER_39_414 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_39_450 ();
 sg13g2_decap_8 FILLER_39_457 ();
 sg13g2_fill_2 FILLER_39_464 ();
 sg13g2_decap_4 FILLER_39_485 ();
 sg13g2_fill_2 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_510 ();
 sg13g2_decap_8 FILLER_39_517 ();
 sg13g2_decap_8 FILLER_39_524 ();
 sg13g2_decap_8 FILLER_39_531 ();
 sg13g2_fill_2 FILLER_39_538 ();
 sg13g2_decap_4 FILLER_39_546 ();
 sg13g2_fill_1 FILLER_39_550 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_fill_2 FILLER_39_570 ();
 sg13g2_fill_1 FILLER_39_572 ();
 sg13g2_fill_2 FILLER_39_582 ();
 sg13g2_fill_1 FILLER_39_584 ();
 sg13g2_decap_8 FILLER_39_594 ();
 sg13g2_decap_4 FILLER_39_601 ();
 sg13g2_decap_8 FILLER_39_613 ();
 sg13g2_decap_4 FILLER_39_620 ();
 sg13g2_fill_2 FILLER_39_644 ();
 sg13g2_fill_1 FILLER_39_646 ();
 sg13g2_decap_8 FILLER_39_666 ();
 sg13g2_decap_8 FILLER_39_673 ();
 sg13g2_fill_1 FILLER_39_680 ();
 sg13g2_decap_8 FILLER_39_698 ();
 sg13g2_decap_4 FILLER_39_705 ();
 sg13g2_fill_1 FILLER_39_709 ();
 sg13g2_fill_2 FILLER_39_713 ();
 sg13g2_fill_1 FILLER_39_715 ();
 sg13g2_decap_8 FILLER_39_720 ();
 sg13g2_fill_2 FILLER_39_736 ();
 sg13g2_fill_1 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_747 ();
 sg13g2_fill_1 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_778 ();
 sg13g2_decap_8 FILLER_39_785 ();
 sg13g2_decap_8 FILLER_39_792 ();
 sg13g2_decap_8 FILLER_39_799 ();
 sg13g2_decap_8 FILLER_39_806 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_decap_8 FILLER_39_841 ();
 sg13g2_decap_8 FILLER_39_848 ();
 sg13g2_decap_8 FILLER_39_855 ();
 sg13g2_decap_8 FILLER_39_862 ();
 sg13g2_decap_8 FILLER_39_869 ();
 sg13g2_decap_8 FILLER_39_876 ();
 sg13g2_decap_8 FILLER_39_883 ();
 sg13g2_decap_8 FILLER_39_890 ();
 sg13g2_decap_8 FILLER_39_897 ();
 sg13g2_decap_8 FILLER_39_904 ();
 sg13g2_decap_8 FILLER_39_911 ();
 sg13g2_decap_8 FILLER_39_918 ();
 sg13g2_decap_8 FILLER_39_925 ();
 sg13g2_decap_8 FILLER_39_932 ();
 sg13g2_decap_8 FILLER_39_939 ();
 sg13g2_decap_8 FILLER_39_946 ();
 sg13g2_decap_8 FILLER_39_953 ();
 sg13g2_decap_8 FILLER_39_960 ();
 sg13g2_decap_8 FILLER_39_967 ();
 sg13g2_decap_8 FILLER_39_974 ();
 sg13g2_decap_8 FILLER_39_981 ();
 sg13g2_decap_8 FILLER_39_988 ();
 sg13g2_decap_8 FILLER_39_995 ();
 sg13g2_decap_8 FILLER_39_1002 ();
 sg13g2_decap_8 FILLER_39_1009 ();
 sg13g2_decap_8 FILLER_39_1016 ();
 sg13g2_decap_4 FILLER_39_1023 ();
 sg13g2_fill_2 FILLER_39_1027 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_13 ();
 sg13g2_fill_1 FILLER_40_20 ();
 sg13g2_decap_8 FILLER_40_30 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_decap_8 FILLER_40_65 ();
 sg13g2_fill_2 FILLER_40_72 ();
 sg13g2_decap_8 FILLER_40_87 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_8 FILLER_40_108 ();
 sg13g2_decap_8 FILLER_40_115 ();
 sg13g2_decap_8 FILLER_40_122 ();
 sg13g2_decap_4 FILLER_40_129 ();
 sg13g2_decap_8 FILLER_40_150 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_205 ();
 sg13g2_decap_8 FILLER_40_212 ();
 sg13g2_decap_4 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_229 ();
 sg13g2_decap_8 FILLER_40_236 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_265 ();
 sg13g2_decap_8 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_decap_4 FILLER_40_297 ();
 sg13g2_decap_8 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_337 ();
 sg13g2_decap_4 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_4 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_421 ();
 sg13g2_decap_4 FILLER_40_428 ();
 sg13g2_decap_8 FILLER_40_442 ();
 sg13g2_decap_4 FILLER_40_449 ();
 sg13g2_fill_2 FILLER_40_453 ();
 sg13g2_fill_1 FILLER_40_460 ();
 sg13g2_decap_4 FILLER_40_466 ();
 sg13g2_decap_8 FILLER_40_481 ();
 sg13g2_decap_4 FILLER_40_488 ();
 sg13g2_decap_8 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_decap_4 FILLER_40_519 ();
 sg13g2_decap_8 FILLER_40_536 ();
 sg13g2_decap_8 FILLER_40_543 ();
 sg13g2_decap_8 FILLER_40_550 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_fill_2 FILLER_40_577 ();
 sg13g2_fill_1 FILLER_40_579 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_594 ();
 sg13g2_decap_4 FILLER_40_601 ();
 sg13g2_decap_8 FILLER_40_610 ();
 sg13g2_decap_8 FILLER_40_617 ();
 sg13g2_decap_8 FILLER_40_624 ();
 sg13g2_decap_8 FILLER_40_631 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_fill_2 FILLER_40_645 ();
 sg13g2_fill_1 FILLER_40_647 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_decap_8 FILLER_40_675 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_4 FILLER_40_693 ();
 sg13g2_fill_2 FILLER_40_697 ();
 sg13g2_decap_4 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_decap_8 FILLER_40_794 ();
 sg13g2_decap_8 FILLER_40_801 ();
 sg13g2_decap_8 FILLER_40_808 ();
 sg13g2_decap_8 FILLER_40_815 ();
 sg13g2_decap_8 FILLER_40_822 ();
 sg13g2_decap_8 FILLER_40_829 ();
 sg13g2_decap_8 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_40_843 ();
 sg13g2_decap_8 FILLER_40_850 ();
 sg13g2_decap_8 FILLER_40_857 ();
 sg13g2_decap_8 FILLER_40_864 ();
 sg13g2_decap_8 FILLER_40_871 ();
 sg13g2_decap_8 FILLER_40_878 ();
 sg13g2_decap_8 FILLER_40_885 ();
 sg13g2_decap_8 FILLER_40_892 ();
 sg13g2_decap_8 FILLER_40_899 ();
 sg13g2_decap_8 FILLER_40_906 ();
 sg13g2_decap_8 FILLER_40_913 ();
 sg13g2_decap_8 FILLER_40_920 ();
 sg13g2_decap_8 FILLER_40_927 ();
 sg13g2_decap_8 FILLER_40_934 ();
 sg13g2_decap_8 FILLER_40_941 ();
 sg13g2_decap_8 FILLER_40_948 ();
 sg13g2_decap_8 FILLER_40_955 ();
 sg13g2_decap_8 FILLER_40_962 ();
 sg13g2_decap_8 FILLER_40_969 ();
 sg13g2_decap_8 FILLER_40_976 ();
 sg13g2_decap_8 FILLER_40_983 ();
 sg13g2_decap_8 FILLER_40_990 ();
 sg13g2_decap_8 FILLER_40_997 ();
 sg13g2_decap_8 FILLER_40_1004 ();
 sg13g2_decap_8 FILLER_40_1011 ();
 sg13g2_decap_8 FILLER_40_1018 ();
 sg13g2_decap_4 FILLER_40_1025 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_decap_8 FILLER_41_30 ();
 sg13g2_fill_1 FILLER_41_37 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_4 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_62 ();
 sg13g2_decap_8 FILLER_41_131 ();
 sg13g2_decap_8 FILLER_41_138 ();
 sg13g2_fill_2 FILLER_41_145 ();
 sg13g2_fill_2 FILLER_41_151 ();
 sg13g2_fill_2 FILLER_41_161 ();
 sg13g2_decap_4 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_decap_8 FILLER_41_213 ();
 sg13g2_decap_4 FILLER_41_220 ();
 sg13g2_fill_2 FILLER_41_224 ();
 sg13g2_fill_2 FILLER_41_267 ();
 sg13g2_decap_4 FILLER_41_325 ();
 sg13g2_fill_1 FILLER_41_337 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_4 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_415 ();
 sg13g2_decap_8 FILLER_41_422 ();
 sg13g2_decap_4 FILLER_41_437 ();
 sg13g2_decap_4 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_452 ();
 sg13g2_decap_8 FILLER_41_457 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_fill_2 FILLER_41_478 ();
 sg13g2_fill_1 FILLER_41_480 ();
 sg13g2_decap_4 FILLER_41_495 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_decap_8 FILLER_41_505 ();
 sg13g2_fill_2 FILLER_41_512 ();
 sg13g2_fill_1 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_533 ();
 sg13g2_fill_2 FILLER_41_540 ();
 sg13g2_fill_1 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_563 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_576 ();
 sg13g2_decap_8 FILLER_41_583 ();
 sg13g2_decap_8 FILLER_41_590 ();
 sg13g2_fill_2 FILLER_41_597 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_decap_4 FILLER_41_650 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_688 ();
 sg13g2_decap_8 FILLER_41_695 ();
 sg13g2_decap_8 FILLER_41_702 ();
 sg13g2_decap_4 FILLER_41_709 ();
 sg13g2_fill_2 FILLER_41_713 ();
 sg13g2_decap_8 FILLER_41_719 ();
 sg13g2_decap_8 FILLER_41_726 ();
 sg13g2_fill_2 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_4 FILLER_41_752 ();
 sg13g2_fill_1 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_8 FILLER_41_857 ();
 sg13g2_decap_8 FILLER_41_864 ();
 sg13g2_decap_8 FILLER_41_871 ();
 sg13g2_decap_8 FILLER_41_878 ();
 sg13g2_decap_8 FILLER_41_885 ();
 sg13g2_decap_8 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_899 ();
 sg13g2_decap_8 FILLER_41_906 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_8 FILLER_41_948 ();
 sg13g2_decap_8 FILLER_41_955 ();
 sg13g2_decap_8 FILLER_41_962 ();
 sg13g2_decap_8 FILLER_41_969 ();
 sg13g2_decap_8 FILLER_41_976 ();
 sg13g2_decap_8 FILLER_41_983 ();
 sg13g2_decap_8 FILLER_41_990 ();
 sg13g2_decap_8 FILLER_41_997 ();
 sg13g2_decap_8 FILLER_41_1004 ();
 sg13g2_decap_8 FILLER_41_1011 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_13 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_decap_8 FILLER_42_43 ();
 sg13g2_decap_8 FILLER_42_50 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_4 FILLER_42_113 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_decap_8 FILLER_42_163 ();
 sg13g2_decap_4 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_202 ();
 sg13g2_decap_8 FILLER_42_209 ();
 sg13g2_decap_8 FILLER_42_216 ();
 sg13g2_decap_8 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_230 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_249 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_decap_4 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_274 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_295 ();
 sg13g2_decap_8 FILLER_42_302 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_fill_2 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_fill_1 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_431 ();
 sg13g2_fill_2 FILLER_42_442 ();
 sg13g2_decap_4 FILLER_42_449 ();
 sg13g2_fill_1 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_470 ();
 sg13g2_fill_1 FILLER_42_484 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_536 ();
 sg13g2_fill_2 FILLER_42_565 ();
 sg13g2_fill_2 FILLER_42_580 ();
 sg13g2_decap_8 FILLER_42_593 ();
 sg13g2_decap_8 FILLER_42_600 ();
 sg13g2_fill_1 FILLER_42_607 ();
 sg13g2_decap_8 FILLER_42_612 ();
 sg13g2_decap_4 FILLER_42_619 ();
 sg13g2_fill_1 FILLER_42_623 ();
 sg13g2_fill_1 FILLER_42_629 ();
 sg13g2_decap_4 FILLER_42_663 ();
 sg13g2_fill_1 FILLER_42_667 ();
 sg13g2_decap_8 FILLER_42_677 ();
 sg13g2_decap_8 FILLER_42_684 ();
 sg13g2_fill_1 FILLER_42_691 ();
 sg13g2_decap_4 FILLER_42_696 ();
 sg13g2_fill_2 FILLER_42_700 ();
 sg13g2_fill_2 FILLER_42_715 ();
 sg13g2_fill_1 FILLER_42_717 ();
 sg13g2_fill_1 FILLER_42_722 ();
 sg13g2_decap_4 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_decap_8 FILLER_42_874 ();
 sg13g2_decap_8 FILLER_42_881 ();
 sg13g2_decap_8 FILLER_42_888 ();
 sg13g2_decap_8 FILLER_42_895 ();
 sg13g2_decap_8 FILLER_42_902 ();
 sg13g2_decap_8 FILLER_42_909 ();
 sg13g2_decap_8 FILLER_42_916 ();
 sg13g2_decap_8 FILLER_42_923 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_8 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_8 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_83 ();
 sg13g2_decap_8 FILLER_43_90 ();
 sg13g2_fill_2 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_decap_4 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_113 ();
 sg13g2_decap_8 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_decap_8 FILLER_43_145 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_4 FILLER_43_166 ();
 sg13g2_decap_8 FILLER_43_232 ();
 sg13g2_decap_8 FILLER_43_239 ();
 sg13g2_fill_1 FILLER_43_246 ();
 sg13g2_decap_8 FILLER_43_251 ();
 sg13g2_decap_4 FILLER_43_258 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_279 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_decap_8 FILLER_43_311 ();
 sg13g2_fill_2 FILLER_43_318 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_4 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_361 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_decap_4 FILLER_43_430 ();
 sg13g2_fill_1 FILLER_43_434 ();
 sg13g2_fill_1 FILLER_43_445 ();
 sg13g2_decap_8 FILLER_43_461 ();
 sg13g2_decap_8 FILLER_43_468 ();
 sg13g2_decap_8 FILLER_43_475 ();
 sg13g2_decap_8 FILLER_43_482 ();
 sg13g2_decap_8 FILLER_43_494 ();
 sg13g2_decap_8 FILLER_43_501 ();
 sg13g2_decap_8 FILLER_43_508 ();
 sg13g2_fill_1 FILLER_43_515 ();
 sg13g2_decap_8 FILLER_43_526 ();
 sg13g2_decap_8 FILLER_43_533 ();
 sg13g2_fill_2 FILLER_43_540 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_8 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_decap_4 FILLER_43_593 ();
 sg13g2_fill_1 FILLER_43_597 ();
 sg13g2_decap_8 FILLER_43_608 ();
 sg13g2_decap_8 FILLER_43_615 ();
 sg13g2_decap_8 FILLER_43_622 ();
 sg13g2_decap_8 FILLER_43_629 ();
 sg13g2_decap_8 FILLER_43_636 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_fill_2 FILLER_43_654 ();
 sg13g2_fill_1 FILLER_43_656 ();
 sg13g2_decap_4 FILLER_43_666 ();
 sg13g2_fill_2 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_680 ();
 sg13g2_decap_8 FILLER_43_724 ();
 sg13g2_decap_8 FILLER_43_731 ();
 sg13g2_fill_1 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_decap_8 FILLER_43_915 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_decap_8 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_8 FILLER_43_985 ();
 sg13g2_decap_8 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_fill_2 FILLER_43_1027 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_fill_1 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_65 ();
 sg13g2_fill_2 FILLER_44_72 ();
 sg13g2_fill_2 FILLER_44_101 ();
 sg13g2_decap_8 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_fill_1 FILLER_44_191 ();
 sg13g2_fill_2 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_4 FILLER_44_224 ();
 sg13g2_decap_4 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_241 ();
 sg13g2_fill_2 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_314 ();
 sg13g2_decap_4 FILLER_44_321 ();
 sg13g2_decap_8 FILLER_44_341 ();
 sg13g2_decap_8 FILLER_44_348 ();
 sg13g2_decap_8 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_decap_8 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_44_415 ();
 sg13g2_decap_4 FILLER_44_435 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_fill_1 FILLER_44_452 ();
 sg13g2_decap_8 FILLER_44_456 ();
 sg13g2_decap_8 FILLER_44_463 ();
 sg13g2_fill_2 FILLER_44_470 ();
 sg13g2_fill_1 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_486 ();
 sg13g2_decap_4 FILLER_44_493 ();
 sg13g2_fill_2 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_fill_1 FILLER_44_522 ();
 sg13g2_decap_4 FILLER_44_527 ();
 sg13g2_fill_2 FILLER_44_531 ();
 sg13g2_decap_4 FILLER_44_552 ();
 sg13g2_fill_1 FILLER_44_556 ();
 sg13g2_decap_4 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_4 FILLER_44_602 ();
 sg13g2_fill_2 FILLER_44_610 ();
 sg13g2_fill_1 FILLER_44_612 ();
 sg13g2_fill_2 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_decap_4 FILLER_44_641 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_decap_8 FILLER_44_657 ();
 sg13g2_decap_4 FILLER_44_664 ();
 sg13g2_fill_1 FILLER_44_668 ();
 sg13g2_decap_8 FILLER_44_678 ();
 sg13g2_decap_8 FILLER_44_685 ();
 sg13g2_decap_8 FILLER_44_692 ();
 sg13g2_fill_1 FILLER_44_699 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_fill_2 FILLER_44_737 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_decap_8 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_44_928 ();
 sg13g2_decap_8 FILLER_44_935 ();
 sg13g2_decap_8 FILLER_44_942 ();
 sg13g2_decap_8 FILLER_44_949 ();
 sg13g2_decap_8 FILLER_44_956 ();
 sg13g2_decap_8 FILLER_44_963 ();
 sg13g2_decap_8 FILLER_44_970 ();
 sg13g2_decap_8 FILLER_44_977 ();
 sg13g2_decap_8 FILLER_44_984 ();
 sg13g2_decap_8 FILLER_44_991 ();
 sg13g2_decap_8 FILLER_44_998 ();
 sg13g2_decap_8 FILLER_44_1005 ();
 sg13g2_decap_8 FILLER_44_1012 ();
 sg13g2_decap_8 FILLER_44_1019 ();
 sg13g2_fill_2 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_4 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_46 ();
 sg13g2_decap_8 FILLER_45_60 ();
 sg13g2_decap_8 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_74 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_decap_8 FILLER_45_88 ();
 sg13g2_decap_4 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_99 ();
 sg13g2_decap_4 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_117 ();
 sg13g2_fill_2 FILLER_45_124 ();
 sg13g2_decap_4 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_144 ();
 sg13g2_decap_8 FILLER_45_151 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_decap_4 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_256 ();
 sg13g2_fill_2 FILLER_45_263 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_decap_4 FILLER_45_284 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_4 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_319 ();
 sg13g2_fill_2 FILLER_45_326 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_4 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_decap_4 FILLER_45_377 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_4 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_decap_4 FILLER_45_427 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_fill_1 FILLER_45_487 ();
 sg13g2_fill_2 FILLER_45_503 ();
 sg13g2_fill_2 FILLER_45_518 ();
 sg13g2_fill_1 FILLER_45_525 ();
 sg13g2_decap_4 FILLER_45_530 ();
 sg13g2_fill_2 FILLER_45_534 ();
 sg13g2_fill_2 FILLER_45_548 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_fill_2 FILLER_45_584 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_fill_2 FILLER_45_592 ();
 sg13g2_fill_1 FILLER_45_594 ();
 sg13g2_decap_4 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_614 ();
 sg13g2_decap_4 FILLER_45_621 ();
 sg13g2_fill_1 FILLER_45_625 ();
 sg13g2_fill_2 FILLER_45_642 ();
 sg13g2_decap_4 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_666 ();
 sg13g2_decap_8 FILLER_45_685 ();
 sg13g2_fill_1 FILLER_45_692 ();
 sg13g2_decap_8 FILLER_45_710 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_decap_8 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_8 FILLER_45_856 ();
 sg13g2_decap_8 FILLER_45_863 ();
 sg13g2_decap_8 FILLER_45_870 ();
 sg13g2_decap_8 FILLER_45_877 ();
 sg13g2_decap_8 FILLER_45_884 ();
 sg13g2_decap_8 FILLER_45_891 ();
 sg13g2_decap_8 FILLER_45_898 ();
 sg13g2_decap_8 FILLER_45_905 ();
 sg13g2_decap_8 FILLER_45_912 ();
 sg13g2_decap_8 FILLER_45_919 ();
 sg13g2_decap_8 FILLER_45_926 ();
 sg13g2_decap_8 FILLER_45_933 ();
 sg13g2_decap_8 FILLER_45_940 ();
 sg13g2_decap_8 FILLER_45_947 ();
 sg13g2_decap_8 FILLER_45_954 ();
 sg13g2_decap_8 FILLER_45_961 ();
 sg13g2_decap_8 FILLER_45_968 ();
 sg13g2_decap_8 FILLER_45_975 ();
 sg13g2_decap_8 FILLER_45_982 ();
 sg13g2_decap_8 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_996 ();
 sg13g2_decap_8 FILLER_45_1003 ();
 sg13g2_decap_8 FILLER_45_1010 ();
 sg13g2_decap_8 FILLER_45_1017 ();
 sg13g2_decap_4 FILLER_45_1024 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_decap_8 FILLER_46_5 ();
 sg13g2_fill_1 FILLER_46_12 ();
 sg13g2_decap_4 FILLER_46_17 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_32 ();
 sg13g2_fill_1 FILLER_46_34 ();
 sg13g2_decap_8 FILLER_46_39 ();
 sg13g2_decap_4 FILLER_46_46 ();
 sg13g2_fill_2 FILLER_46_50 ();
 sg13g2_fill_1 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_decap_8 FILLER_46_102 ();
 sg13g2_fill_2 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_decap_4 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_decap_4 FILLER_46_209 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_fill_2 FILLER_46_232 ();
 sg13g2_decap_8 FILLER_46_243 ();
 sg13g2_decap_4 FILLER_46_250 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_fill_2 FILLER_46_302 ();
 sg13g2_fill_1 FILLER_46_304 ();
 sg13g2_decap_8 FILLER_46_318 ();
 sg13g2_fill_1 FILLER_46_353 ();
 sg13g2_fill_1 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_372 ();
 sg13g2_decap_4 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_fill_1 FILLER_46_435 ();
 sg13g2_decap_8 FILLER_46_446 ();
 sg13g2_decap_8 FILLER_46_453 ();
 sg13g2_decap_8 FILLER_46_460 ();
 sg13g2_decap_4 FILLER_46_467 ();
 sg13g2_fill_1 FILLER_46_471 ();
 sg13g2_decap_8 FILLER_46_478 ();
 sg13g2_decap_8 FILLER_46_485 ();
 sg13g2_decap_4 FILLER_46_505 ();
 sg13g2_fill_2 FILLER_46_509 ();
 sg13g2_decap_4 FILLER_46_519 ();
 sg13g2_fill_1 FILLER_46_536 ();
 sg13g2_decap_8 FILLER_46_550 ();
 sg13g2_decap_8 FILLER_46_557 ();
 sg13g2_decap_4 FILLER_46_564 ();
 sg13g2_fill_1 FILLER_46_568 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_fill_1 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_593 ();
 sg13g2_decap_4 FILLER_46_600 ();
 sg13g2_fill_2 FILLER_46_609 ();
 sg13g2_fill_1 FILLER_46_611 ();
 sg13g2_decap_4 FILLER_46_624 ();
 sg13g2_fill_1 FILLER_46_628 ();
 sg13g2_decap_8 FILLER_46_639 ();
 sg13g2_fill_2 FILLER_46_646 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_fill_2 FILLER_46_672 ();
 sg13g2_fill_1 FILLER_46_674 ();
 sg13g2_decap_8 FILLER_46_682 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_4 FILLER_46_696 ();
 sg13g2_fill_2 FILLER_46_728 ();
 sg13g2_fill_1 FILLER_46_730 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_8 FILLER_46_857 ();
 sg13g2_decap_8 FILLER_46_864 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_decap_8 FILLER_46_878 ();
 sg13g2_decap_8 FILLER_46_885 ();
 sg13g2_decap_8 FILLER_46_892 ();
 sg13g2_decap_8 FILLER_46_899 ();
 sg13g2_decap_8 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_913 ();
 sg13g2_decap_8 FILLER_46_920 ();
 sg13g2_decap_8 FILLER_46_927 ();
 sg13g2_decap_8 FILLER_46_934 ();
 sg13g2_decap_8 FILLER_46_941 ();
 sg13g2_decap_8 FILLER_46_948 ();
 sg13g2_decap_8 FILLER_46_955 ();
 sg13g2_decap_8 FILLER_46_962 ();
 sg13g2_decap_8 FILLER_46_969 ();
 sg13g2_decap_8 FILLER_46_976 ();
 sg13g2_decap_8 FILLER_46_983 ();
 sg13g2_decap_8 FILLER_46_990 ();
 sg13g2_decap_8 FILLER_46_997 ();
 sg13g2_decap_8 FILLER_46_1004 ();
 sg13g2_decap_8 FILLER_46_1011 ();
 sg13g2_decap_8 FILLER_46_1018 ();
 sg13g2_decap_4 FILLER_46_1025 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_decap_8 FILLER_47_79 ();
 sg13g2_decap_8 FILLER_47_86 ();
 sg13g2_decap_8 FILLER_47_93 ();
 sg13g2_decap_8 FILLER_47_100 ();
 sg13g2_decap_8 FILLER_47_107 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_decap_8 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_128 ();
 sg13g2_fill_2 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_fill_2 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_191 ();
 sg13g2_fill_1 FILLER_47_193 ();
 sg13g2_fill_2 FILLER_47_215 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_260 ();
 sg13g2_decap_8 FILLER_47_265 ();
 sg13g2_decap_8 FILLER_47_272 ();
 sg13g2_fill_2 FILLER_47_279 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_decap_8 FILLER_47_299 ();
 sg13g2_decap_4 FILLER_47_306 ();
 sg13g2_decap_8 FILLER_47_319 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_decap_4 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_fill_2 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_4 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_400 ();
 sg13g2_decap_8 FILLER_47_415 ();
 sg13g2_fill_1 FILLER_47_431 ();
 sg13g2_decap_8 FILLER_47_437 ();
 sg13g2_decap_4 FILLER_47_444 ();
 sg13g2_fill_2 FILLER_47_448 ();
 sg13g2_fill_1 FILLER_47_455 ();
 sg13g2_fill_1 FILLER_47_460 ();
 sg13g2_decap_8 FILLER_47_470 ();
 sg13g2_decap_8 FILLER_47_477 ();
 sg13g2_decap_8 FILLER_47_484 ();
 sg13g2_fill_2 FILLER_47_491 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_decap_8 FILLER_47_514 ();
 sg13g2_fill_2 FILLER_47_521 ();
 sg13g2_decap_4 FILLER_47_528 ();
 sg13g2_fill_2 FILLER_47_532 ();
 sg13g2_fill_2 FILLER_47_556 ();
 sg13g2_fill_1 FILLER_47_558 ();
 sg13g2_decap_4 FILLER_47_568 ();
 sg13g2_fill_1 FILLER_47_572 ();
 sg13g2_decap_8 FILLER_47_582 ();
 sg13g2_decap_4 FILLER_47_607 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_fill_2 FILLER_47_647 ();
 sg13g2_decap_8 FILLER_47_660 ();
 sg13g2_fill_2 FILLER_47_667 ();
 sg13g2_fill_1 FILLER_47_669 ();
 sg13g2_fill_2 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_698 ();
 sg13g2_decap_8 FILLER_47_705 ();
 sg13g2_decap_4 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_101 ();
 sg13g2_fill_2 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_decap_4 FILLER_48_169 ();
 sg13g2_fill_2 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_decap_8 FILLER_48_237 ();
 sg13g2_decap_8 FILLER_48_244 ();
 sg13g2_decap_8 FILLER_48_251 ();
 sg13g2_decap_8 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_265 ();
 sg13g2_decap_8 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_279 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_decap_4 FILLER_48_348 ();
 sg13g2_decap_8 FILLER_48_384 ();
 sg13g2_fill_2 FILLER_48_391 ();
 sg13g2_fill_1 FILLER_48_393 ();
 sg13g2_fill_2 FILLER_48_431 ();
 sg13g2_fill_1 FILLER_48_433 ();
 sg13g2_fill_2 FILLER_48_462 ();
 sg13g2_decap_4 FILLER_48_504 ();
 sg13g2_fill_1 FILLER_48_508 ();
 sg13g2_fill_2 FILLER_48_541 ();
 sg13g2_fill_1 FILLER_48_543 ();
 sg13g2_fill_2 FILLER_48_640 ();
 sg13g2_fill_1 FILLER_48_645 ();
 sg13g2_fill_2 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_716 ();
 sg13g2_decap_8 FILLER_48_723 ();
 sg13g2_decap_8 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_8 FILLER_48_744 ();
 sg13g2_decap_8 FILLER_48_751 ();
 sg13g2_decap_8 FILLER_48_758 ();
 sg13g2_decap_8 FILLER_48_765 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_decap_8 FILLER_48_877 ();
 sg13g2_decap_8 FILLER_48_884 ();
 sg13g2_decap_8 FILLER_48_891 ();
 sg13g2_decap_8 FILLER_48_898 ();
 sg13g2_decap_8 FILLER_48_905 ();
 sg13g2_decap_8 FILLER_48_912 ();
 sg13g2_decap_8 FILLER_48_919 ();
 sg13g2_decap_8 FILLER_48_926 ();
 sg13g2_decap_8 FILLER_48_933 ();
 sg13g2_decap_8 FILLER_48_940 ();
 sg13g2_decap_8 FILLER_48_947 ();
 sg13g2_decap_8 FILLER_48_954 ();
 sg13g2_decap_8 FILLER_48_961 ();
 sg13g2_decap_8 FILLER_48_968 ();
 sg13g2_decap_8 FILLER_48_975 ();
 sg13g2_decap_8 FILLER_48_982 ();
 sg13g2_decap_8 FILLER_48_989 ();
 sg13g2_decap_8 FILLER_48_996 ();
 sg13g2_decap_8 FILLER_48_1003 ();
 sg13g2_decap_8 FILLER_48_1010 ();
 sg13g2_decap_8 FILLER_48_1017 ();
 sg13g2_decap_4 FILLER_48_1024 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_5 ();
 sg13g2_decap_8 FILLER_49_12 ();
 sg13g2_decap_8 FILLER_49_19 ();
 sg13g2_decap_8 FILLER_49_26 ();
 sg13g2_decap_8 FILLER_49_33 ();
 sg13g2_decap_8 FILLER_49_40 ();
 sg13g2_decap_8 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_58 ();
 sg13g2_decap_4 FILLER_49_69 ();
 sg13g2_decap_8 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_89 ();
 sg13g2_decap_8 FILLER_49_96 ();
 sg13g2_decap_8 FILLER_49_103 ();
 sg13g2_decap_8 FILLER_49_110 ();
 sg13g2_decap_8 FILLER_49_117 ();
 sg13g2_decap_8 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_138 ();
 sg13g2_decap_8 FILLER_49_145 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_177 ();
 sg13g2_decap_8 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_decap_8 FILLER_49_198 ();
 sg13g2_decap_8 FILLER_49_205 ();
 sg13g2_decap_8 FILLER_49_212 ();
 sg13g2_decap_8 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_8 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_247 ();
 sg13g2_decap_8 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_275 ();
 sg13g2_decap_8 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_decap_4 FILLER_49_302 ();
 sg13g2_fill_1 FILLER_49_306 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_4 FILLER_49_357 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_decap_4 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_decap_8 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_421 ();
 sg13g2_decap_8 FILLER_49_428 ();
 sg13g2_decap_4 FILLER_49_435 ();
 sg13g2_decap_8 FILLER_49_443 ();
 sg13g2_decap_8 FILLER_49_450 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_decap_4 FILLER_49_464 ();
 sg13g2_fill_1 FILLER_49_468 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_4 FILLER_49_487 ();
 sg13g2_fill_1 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_4 FILLER_49_508 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_fill_2 FILLER_49_546 ();
 sg13g2_fill_1 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_fill_2 FILLER_49_574 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_621 ();
 sg13g2_decap_8 FILLER_49_628 ();
 sg13g2_decap_8 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_8 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_decap_8 FILLER_49_663 ();
 sg13g2_decap_8 FILLER_49_670 ();
 sg13g2_decap_8 FILLER_49_677 ();
 sg13g2_decap_8 FILLER_49_684 ();
 sg13g2_decap_4 FILLER_49_691 ();
 sg13g2_fill_2 FILLER_49_695 ();
 sg13g2_decap_8 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_713 ();
 sg13g2_decap_8 FILLER_49_720 ();
 sg13g2_decap_8 FILLER_49_727 ();
 sg13g2_decap_8 FILLER_49_734 ();
 sg13g2_decap_8 FILLER_49_741 ();
 sg13g2_decap_8 FILLER_49_748 ();
 sg13g2_decap_8 FILLER_49_755 ();
 sg13g2_decap_8 FILLER_49_762 ();
 sg13g2_decap_8 FILLER_49_769 ();
 sg13g2_decap_8 FILLER_49_776 ();
 sg13g2_decap_8 FILLER_49_783 ();
 sg13g2_decap_8 FILLER_49_790 ();
 sg13g2_decap_8 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_804 ();
 sg13g2_decap_8 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_decap_8 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_49_867 ();
 sg13g2_decap_8 FILLER_49_874 ();
 sg13g2_decap_8 FILLER_49_881 ();
 sg13g2_decap_8 FILLER_49_888 ();
 sg13g2_decap_8 FILLER_49_895 ();
 sg13g2_decap_8 FILLER_49_902 ();
 sg13g2_decap_8 FILLER_49_909 ();
 sg13g2_decap_8 FILLER_49_916 ();
 sg13g2_decap_8 FILLER_49_923 ();
 sg13g2_decap_8 FILLER_49_930 ();
 sg13g2_decap_8 FILLER_49_937 ();
 sg13g2_decap_8 FILLER_49_944 ();
 sg13g2_decap_8 FILLER_49_951 ();
 sg13g2_decap_8 FILLER_49_958 ();
 sg13g2_decap_8 FILLER_49_965 ();
 sg13g2_decap_8 FILLER_49_972 ();
 sg13g2_decap_8 FILLER_49_979 ();
 sg13g2_decap_8 FILLER_49_986 ();
 sg13g2_decap_8 FILLER_49_993 ();
 sg13g2_decap_8 FILLER_49_1000 ();
 sg13g2_decap_8 FILLER_49_1007 ();
 sg13g2_decap_8 FILLER_49_1014 ();
 sg13g2_decap_8 FILLER_49_1021 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule
