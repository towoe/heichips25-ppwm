* NGSPICE file created from heichips25_ppwm.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

.subckt heichips25_ppwm VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_28_918 VPWR VGND sg13g2_decap_8
XFILLER_36_19 VPWR VGND sg13g2_fill_1
XFILLER_23_601 VPWR VGND sg13g2_decap_8
XFILLER_36_984 VPWR VGND sg13g2_decap_8
XFILLER_22_111 VPWR VGND sg13g2_decap_8
XFILLER_23_678 VPWR VGND sg13g2_decap_8
XFILLER_2_527 VPWR VGND sg13g2_decap_8
XFILLER_18_417 VPWR VGND sg13g2_fill_2
XFILLER_19_918 VPWR VGND sg13g2_decap_8
XFILLER_46_748 VPWR VGND sg13g2_decap_8
XFILLER_33_409 VPWR VGND sg13g2_fill_2
XFILLER_14_601 VPWR VGND sg13g2_decap_8
XFILLER_27_984 VPWR VGND sg13g2_decap_8
XFILLER_42_943 VPWR VGND sg13g2_decap_8
XFILLER_41_453 VPWR VGND sg13g2_decap_8
XFILLER_14_678 VPWR VGND sg13g2_decap_8
XFILLER_6_800 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__182_ net547 u_ppwm_u_pwm__182_/B hold180/A VPWR VGND sg13g2_nor2_1
XFILLER_6_877 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_37_759 VPWR VGND sg13g2_decap_8
XFILLER_18_995 VPWR VGND sg13g2_decap_8
XFILLER_33_932 VPWR VGND sg13g2_decap_8
XFILLER_20_648 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0995_ net358 u_ppwm_u_ex__0995_/B u_ppwm_u_ex__1000_/B VPWR VGND sg13g2_nor2_1
XFILLER_41_1013 VPWR VGND sg13g2_decap_8
XFILLER_28_715 VPWR VGND sg13g2_decap_8
XFILLER_36_781 VPWR VGND sg13g2_decap_8
XFILLER_23_442 VPWR VGND sg13g2_decap_8
XFILLER_23_453 VPWR VGND sg13g2_fill_1
XFILLER_24_976 VPWR VGND sg13g2_decap_8
XFILLER_11_637 VPWR VGND sg13g2_decap_8
XFILLER_7_619 VPWR VGND sg13g2_decap_8
XFILLER_3_814 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_2_335 VPWR VGND sg13g2_decap_4
Xhold170 hold170/A VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold181 hold181/A VPWR VGND net549 sg13g2_dlygate4sd3_1
Xhold192 hold192/A VPWR VGND net560 sg13g2_dlygate4sd3_1
XFILLER_19_715 VPWR VGND sg13g2_decap_8
XFILLER_46_545 VPWR VGND sg13g2_decap_8
XFILLER_18_236 VPWR VGND sg13g2_fill_2
XFILLER_27_781 VPWR VGND sg13g2_decap_8
XFILLER_42_740 VPWR VGND sg13g2_decap_8
XFILLER_15_943 VPWR VGND sg13g2_decap_8
XFILLER_41_250 VPWR VGND sg13g2_fill_2
XFILLER_30_924 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0992_ net497 VPWR u_ppwm_u_mem__0992_/Y VGND net413 net228 sg13g2_o21ai_1
Xu_ppwm_u_ex__0780_ u_ppwm_u_ex__0781_/A u_ppwm_u_ex__0819_/C u_ppwm_u_ex__0780_/X
+ VPWR VGND sg13g2_and2_1
Xu_ppwm_u_pwm__234_ net177 VGND VPWR net210 hold11/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__165_ VGND VPWR net549 u_ppwm_u_pwm__163_/A hold182/A u_ppwm_u_pwm__164_/Y
+ sg13g2_a21oi_1
XFILLER_6_674 VPWR VGND sg13g2_decap_8
XFILLER_2_891 VPWR VGND sg13g2_decap_8
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_556 VPWR VGND sg13g2_decap_8
XFILLER_25_729 VPWR VGND sg13g2_decap_8
XFILLER_18_792 VPWR VGND sg13g2_decap_8
XFILLER_21_946 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0978_ VGND VPWR u_ppwm_u_ex__0970_/Y u_ppwm_u_ex__0976_/Y u_ppwm_u_ex__1114_/D
+ u_ppwm_u_ex__0977_/Y sg13g2_a21oi_1
XFILLER_20_445 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
XFILLER_0_817 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_11 VPWR VGND uio_out[0] sg13g2_tielo
Xheichips25_ppwm_22 VPWR VGND uo_out[4] sg13g2_tielo
XFILLER_28_589 VPWR VGND sg13g2_decap_8
XFILLER_43_559 VPWR VGND sg13g2_decap_8
XFILLER_15_239 VPWR VGND sg13g2_decap_8
XFILLER_12_902 VPWR VGND sg13g2_decap_8
XFILLER_24_773 VPWR VGND sg13g2_decap_8
XFILLER_12_979 VPWR VGND sg13g2_decap_8
XFILLER_3_611 VPWR VGND sg13g2_decap_8
XFILLER_3_688 VPWR VGND sg13g2_decap_8
Xfanout491 net492 net491 VPWR VGND sg13g2_buf_1
XFILLER_19_512 VPWR VGND sg13g2_decap_8
Xfanout480 net487 net480 VPWR VGND sg13g2_buf_8
XFILLER_47_865 VPWR VGND sg13g2_decap_8
XFILLER_46_342 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1146__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_0_35 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1191_ net170 VGND VPWR net539 hold203/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_589 VPWR VGND sg13g2_decap_8
XFILLER_34_548 VPWR VGND sg13g2_decap_8
XFILLER_15_740 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0901_ u_ppwm_u_ex__0880_/Y VPWR u_ppwm_u_ex__0901_/Y VGND u_ppwm_u_ex__0881_/Y
+ u_ppwm_u_ex__0884_/Y sg13g2_o21ai_1
XFILLER_30_721 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0832_ u_ppwm_u_ex__0831_/Y VPWR u_ppwm_u_ex__0833_/C VGND net360 u_ppwm_u_ex__0830_/Y
+ sg13g2_o21ai_1
XFILLER_30_798 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0975_ VGND VPWR net415 u_ppwm_u_mem__0667_/Y hold118/A u_ppwm_u_mem__0974_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__217_ VPWR VGND u_ppwm_u_pwm__203_/Y u_ppwm_u_pwm__216_/Y u_ppwm_u_pwm__215_/Y
+ u_ppwm_u_pwm__206_/Y u_ppwm_u_pwm__222_/A u_ppwm_u_pwm__209_/D sg13g2_a221oi_1
Xu_ppwm_u_ex__0763_ u_ppwm_u_ex__0763_/A u_ppwm_u_ex__0762_/Y u_ppwm_u_ex__0763_/Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
XFILLER_6_471 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0694_ hold310/A u_ppwm_u_ex__0998_/B2 u_ppwm_u_ex__0694_/Y VPWR VGND
+ sg13g2_nor2b_1
Xu_ppwm_u_pwm__148_ VGND VPWR u_ppwm_u_pwm__132_/Y net390 hold166/A u_ppwm_u_pwm__147_/Y
+ sg13g2_a21oi_1
XFILLER_9_1013 VPWR VGND sg13g2_decap_8
XFILLER_38_865 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__097_ VGND VPWR u_ppwm_u_global_counter__056_/Y u_ppwm_u_global_counter__093_/Y
+ hold255/A u_ppwm_u_global_counter__099_/B sg13g2_a21oi_1
XFILLER_25_526 VPWR VGND sg13g2_decap_8
XFILLER_37_386 VPWR VGND sg13g2_fill_2
XFILLER_21_743 VPWR VGND sg13g2_decap_8
XFILLER_0_614 VPWR VGND sg13g2_decap_8
XFILLER_48_607 VPWR VGND sg13g2_decap_8
XFILLER_47_106 VPWR VGND sg13g2_fill_2
XFILLER_29_854 VPWR VGND sg13g2_decap_8
XFILLER_44_813 VPWR VGND sg13g2_decap_8
XFILLER_16_559 VPWR VGND sg13g2_decap_8
XFILLER_24_570 VPWR VGND sg13g2_decap_8
XFILLER_12_776 VPWR VGND sg13g2_decap_8
XFILLER_8_758 VPWR VGND sg13g2_decap_8
XFILLER_7_257 VPWR VGND sg13g2_decap_8
XFILLER_11_297 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0760_ u_ppwm_u_mem__0760_/Y net395 u_ppwm_u_mem__0760_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_4_953 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0691_ VPWR u_ppwm_u_mem__0691_/Y net314 VGND sg13g2_inv_1
XFILLER_3_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1100_ net51 VGND VPWR u_ppwm_u_ex__1100_/D hold321/A clknet_5_25__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1031_ u_ppwm_u_ex__1030_/Y VPWR u_ppwm_u_ex__1035_/C VGND u_ppwm_u_ex__1054_/A
+ u_ppwm_u_ex__1029_/Y sg13g2_o21ai_1
XFILLER_47_662 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1174_ net119 VGND VPWR u_ppwm_u_mem__1174_/D hold94/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_46_183 VPWR VGND sg13g2_fill_1
XFILLER_35_857 VPWR VGND sg13g2_decap_8
XFILLER_22_507 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0815_ net466 hold292/A net386 u_ppwm_u_ex__0816_/B VPWR VGND sg13g2_mux2_1
XFILLER_30_595 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0746_ u_ppwm_u_ex__0746_/Y net466 net445 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0958_ net510 VPWR u_ppwm_u_mem__0958_/Y VGND net429 net309 sg13g2_o21ai_1
XFILLER_7_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0677_ u_ppwm_u_ex__0676_/Y VPWR u_ppwm_u_ex__0678_/C VGND u_ppwm_u_ex__0732_/B
+ hold240/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0889_ VGND VPWR net423 u_ppwm_u_mem__0710_/Y u_ppwm_u_mem__1121_/D
+ u_ppwm_u_mem__0888_/Y sg13g2_a21oi_1
XFILLER_29_139 VPWR VGND sg13g2_fill_1
XFILLER_26_813 VPWR VGND sg13g2_decap_8
XFILLER_37_150 VPWR VGND sg13g2_fill_2
XFILLER_38_662 VPWR VGND sg13g2_decap_8
XFILLER_13_507 VPWR VGND sg13g2_decap_8
XFILLER_25_356 VPWR VGND sg13g2_decap_8
XFILLER_25_367 VPWR VGND sg13g2_fill_2
XFILLER_41_838 VPWR VGND sg13g2_decap_8
XFILLER_21_540 VPWR VGND sg13g2_decap_8
XFILLER_5_717 VPWR VGND sg13g2_decap_8
XFILLER_4_216 VPWR VGND sg13g2_decap_8
XFILLER_0_411 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
XFILLER_49_949 VPWR VGND sg13g2_decap_8
Xhold30 hold30/A VPWR VGND net228 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1173__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_48_404 VPWR VGND sg13g2_decap_8
Xhold41 hold41/A VPWR VGND net239 sg13g2_dlygate4sd3_1
XFILLER_0_488 VPWR VGND sg13g2_decap_8
Xhold74 hold74/A VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold52 hold52/A VPWR VGND net250 sg13g2_dlygate4sd3_1
Xhold63 hold63/A VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold85 hold85/A VPWR VGND net283 sg13g2_dlygate4sd3_1
XFILLER_29_651 VPWR VGND sg13g2_decap_8
Xhold96 hold96/A VPWR VGND net294 sg13g2_dlygate4sd3_1
XFILLER_44_610 VPWR VGND sg13g2_decap_8
XFILLER_17_824 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_decap_8
XFILLER_25_890 VPWR VGND sg13g2_decap_8
XFILLER_12_573 VPWR VGND sg13g2_decap_8
XFILLER_8_555 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0600_ u_ppwm_u_ex__0600_/Y net446 u_ppwm_u_ex__0601_/C VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0812_ hold107/A hold141/A net480 u_ppwm_u_mem__0812_/X VPWR VGND sg13g2_mux2_1
XFILLER_6_67 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0743_ u_ppwm_u_mem__0743_/Y net396 u_ppwm_u_mem__0743_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_4_750 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0674_ VPWR u_ppwm_u_mem__0674_/Y net245 VGND sg13g2_inv_1
XFILLER_48_971 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1014_ u_ppwm_u_ex__1014_/A u_ppwm_u_ex__1012_/Y u_ppwm_u_ex__1117_/D
+ VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__1226_ net176 VGND VPWR net334 hold135/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1157_ net167 VGND VPWR net246 hold173/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_654 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1088_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1088_/B u_ppwm_u_mem__1090_/B
+ u_ppwm_u_mem__1219_/D VPWR VGND sg13g2_nor3_1
XFILLER_34_186 VPWR VGND sg13g2_fill_1
XFILLER_2_709 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0729_ net460 net449 u_ppwm_u_ex__0730_/D VPWR VGND sg13g2_xor2_1
XFILLER_45_429 VPWR VGND sg13g2_decap_8
XFILLER_26_610 VPWR VGND sg13g2_decap_8
XFILLER_26_687 VPWR VGND sg13g2_decap_8
XFILLER_41_635 VPWR VGND sg13g2_decap_8
XFILLER_25_186 VPWR VGND sg13g2_fill_2
XFILLER_22_871 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_21_381 VPWR VGND sg13g2_fill_1
XFILLER_5_514 VPWR VGND sg13g2_decap_8
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_48_201 VPWR VGND sg13g2_decap_8
XFILLER_0_241 VPWR VGND sg13g2_decap_8
XFILLER_49_746 VPWR VGND sg13g2_decap_8
XFILLER_48_278 VPWR VGND sg13g2_decap_8
XFILLER_17_621 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1011_ VGND VPWR net410 u_ppwm_u_mem__0649_/Y hold148/A u_ppwm_u_mem__1010_/Y
+ sg13g2_a21oi_1
XFILLER_45_996 VPWR VGND sg13g2_decap_8
XFILLER_44_484 VPWR VGND sg13g2_decap_8
XFILLER_16_164 VPWR VGND sg13g2_decap_8
XFILLER_16_175 VPWR VGND sg13g2_fill_2
XFILLER_17_698 VPWR VGND sg13g2_decap_8
XFILLER_13_871 VPWR VGND sg13g2_decap_8
XFILLER_32_668 VPWR VGND sg13g2_decap_8
XFILLER_9_831 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_8_341 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0726_ VPWR u_ppwm_u_mem__0726_/Y net333 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0657_ VPWR u_ppwm_u_mem__0657_/Y net297 VGND sg13g2_inv_1
XFILLER_27_407 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1209_ net168 VGND VPWR u_ppwm_u_mem__1209_/D hold120/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_963 VPWR VGND sg13g2_decap_8
XFILLER_23_657 VPWR VGND sg13g2_decap_8
XFILLER_11_819 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1163__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_2_506 VPWR VGND sg13g2_decap_8
XFILLER_46_727 VPWR VGND sg13g2_decap_8
XFILLER_45_226 VPWR VGND sg13g2_decap_8
XFILLER_27_963 VPWR VGND sg13g2_decap_8
XFILLER_42_922 VPWR VGND sg13g2_decap_8
XFILLER_41_432 VPWR VGND sg13g2_decap_8
XFILLER_13_101 VPWR VGND sg13g2_decap_8
XFILLER_14_657 VPWR VGND sg13g2_decap_8
XFILLER_42_999 VPWR VGND sg13g2_decap_8
XFILLER_13_167 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__181_ u_ppwm_u_pwm__182_/B net489 hold269/A VPWR VGND sg13g2_nand2_1
XFILLER_10_885 VPWR VGND sg13g2_decap_8
XFILLER_6_856 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_37_738 VPWR VGND sg13g2_decap_8
XFILLER_18_974 VPWR VGND sg13g2_decap_8
XFILLER_33_911 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
XFILLER_17_495 VPWR VGND sg13g2_decap_8
XFILLER_33_988 VPWR VGND sg13g2_decap_8
XFILLER_20_627 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0994_ u_ppwm_u_ex__0995_/B u_ppwm_u_ex__0994_/A u_ppwm_u_ex__0994_/B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_34_1010 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0709_ VPWR u_ppwm_u_mem__0709_/Y net551 VGND sg13g2_inv_1
XFILLER_36_760 VPWR VGND sg13g2_decap_8
XFILLER_24_955 VPWR VGND sg13g2_decap_8
XFILLER_11_616 VPWR VGND sg13g2_decap_8
Xhold160 hold160/A VPWR VGND net528 sg13g2_dlygate4sd3_1
Xhold171 hold171/A VPWR VGND net539 sg13g2_dlygate4sd3_1
Xhold182 hold182/A VPWR VGND net550 sg13g2_dlygate4sd3_1
Xhold193 hold193/A VPWR VGND net561 sg13g2_dlygate4sd3_1
XFILLER_46_524 VPWR VGND sg13g2_decap_8
XFILLER_18_204 VPWR VGND sg13g2_fill_1
XFILLER_15_922 VPWR VGND sg13g2_decap_8
XFILLER_27_760 VPWR VGND sg13g2_decap_8
XFILLER_18_1016 VPWR VGND sg13g2_decap_8
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_30_903 VPWR VGND sg13g2_decap_8
XFILLER_42_796 VPWR VGND sg13g2_decap_8
XFILLER_41_262 VPWR VGND sg13g2_fill_1
XFILLER_15_999 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0991_ VGND VPWR net413 u_ppwm_u_mem__0659_/Y hold31/A u_ppwm_u_mem__0990_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__233_ net179 VGND VPWR net261 hold62/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_6_653 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_10_682 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__164_ net489 VPWR u_ppwm_u_pwm__164_/Y VGND net549 u_ppwm_u_pwm__163_/A
+ sg13g2_o21ai_1
XFILLER_5_152 VPWR VGND sg13g2_decap_8
XFILLER_2_870 VPWR VGND sg13g2_decap_8
XFILLER_25_1009 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_25_708 VPWR VGND sg13g2_decap_8
XFILLER_37_535 VPWR VGND sg13g2_decap_8
XFILLER_18_771 VPWR VGND sg13g2_decap_8
XFILLER_45_590 VPWR VGND sg13g2_decap_8
XFILLER_17_292 VPWR VGND sg13g2_decap_8
XFILLER_21_925 VPWR VGND sg13g2_decap_8
XFILLER_32_262 VPWR VGND sg13g2_fill_2
XFILLER_33_785 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0977_ net492 VPWR u_ppwm_u_ex__0977_/Y VGND net454 net353 sg13g2_o21ai_1
Xheichips25_ppwm_23 VPWR VGND uo_out[5] sg13g2_tielo
Xheichips25_ppwm_12 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_28_568 VPWR VGND sg13g2_decap_8
XFILLER_43_538 VPWR VGND sg13g2_decap_8
XFILLER_24_752 VPWR VGND sg13g2_decap_8
XFILLER_12_958 VPWR VGND sg13g2_decap_8
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_3_667 VPWR VGND sg13g2_decap_8
XFILLER_2_155 VPWR VGND sg13g2_fill_2
Xfanout492 net493 net492 VPWR VGND sg13g2_buf_8
Xfanout470 hold305/A net470 VPWR VGND sg13g2_buf_8
Xfanout481 net487 net481 VPWR VGND sg13g2_buf_8
XFILLER_47_844 VPWR VGND sg13g2_decap_8
XFILLER_46_321 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1190_ net55 VGND VPWR u_ppwm_u_mem__1190_/D hold128/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_19_568 VPWR VGND sg13g2_decap_8
XFILLER_46_398 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0900_ u_ppwm_u_ex__0900_/A u_ppwm_u_ex__0898_/Y u_ppwm_u_ex__1109_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_14_262 VPWR VGND sg13g2_decap_4
XFILLER_15_796 VPWR VGND sg13g2_decap_8
XFILLER_30_700 VPWR VGND sg13g2_decap_8
XFILLER_42_593 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0831_ u_ppwm_u_ex__0831_/Y net678 u_ppwm_u_ex__0831_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0974_ net498 VPWR u_ppwm_u_mem__0974_/Y VGND net415 hold163/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0762_ VPWR VGND u_ppwm_u_ex__0757_/A u_ppwm_u_ex__0761_/Y hold262/A
+ u_ppwm_u_ex__0954_/A u_ppwm_u_ex__0762_/Y net442 sg13g2_a221oi_1
XFILLER_30_777 VPWR VGND sg13g2_decap_8
XFILLER_31_1024 VPWR VGND sg13g2_decap_4
XFILLER_7_962 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__216_ u_ppwm_u_pwm__216_/A u_ppwm_u_pwm__216_/B u_ppwm_u_pwm__216_/C
+ u_ppwm_u_pwm__216_/Y VPWR VGND sg13g2_nor3_1
XFILLER_11_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0693_ u_ppwm_u_ex__0693_/Y hold314/A u_ppwm_u_ex__0693_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_pwm__147_ net490 VPWR u_ppwm_u_pwm__147_/Y VGND hold324/A net390 sg13g2_o21ai_1
XFILLER_38_844 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__096_ net392 u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__099_/B
+ VPWR VGND sg13g2_and2_1
XFILLER_25_505 VPWR VGND sg13g2_decap_8
XFILLER_21_722 VPWR VGND sg13g2_decap_8
XFILLER_33_582 VPWR VGND sg13g2_decap_8
XFILLER_21_799 VPWR VGND sg13g2_decap_8
XFILLER_18_10 VPWR VGND sg13g2_fill_1
XFILLER_47_129 VPWR VGND sg13g2_decap_8
XFILLER_29_833 VPWR VGND sg13g2_decap_8
XFILLER_16_538 VPWR VGND sg13g2_decap_8
XFILLER_28_376 VPWR VGND sg13g2_decap_4
XFILLER_44_869 VPWR VGND sg13g2_decap_8
XFILLER_34_20 VPWR VGND sg13g2_fill_2
XFILLER_12_755 VPWR VGND sg13g2_decap_8
XFILLER_8_737 VPWR VGND sg13g2_decap_8
XFILLER_7_225 VPWR VGND sg13g2_fill_2
XFILLER_4_932 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0690_ VPWR u_ppwm_u_mem__0690_/Y net545 VGND sg13g2_inv_1
XFILLER_3_464 VPWR VGND sg13g2_decap_8
XFILLER_39_619 VPWR VGND sg13g2_decap_8
XFILLER_47_641 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1030_ VGND VPWR u_ppwm_u_ex__1054_/A u_ppwm_u_ex__1029_/Y u_ppwm_u_ex__1030_/Y
+ net357 sg13g2_a21oi_1
Xu_ppwm_u_mem__1173_ net123 VGND VPWR u_ppwm_u_mem__1173_/D hold30/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_35_836 VPWR VGND sg13g2_decap_8
XFILLER_34_368 VPWR VGND sg13g2_decap_8
XFILLER_34_379 VPWR VGND sg13g2_fill_2
XFILLER_15_593 VPWR VGND sg13g2_decap_8
XFILLER_30_574 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0814_ VPWR u_ppwm_u_ex__0814_/Y u_ppwm_u_ex__0814_/A VGND sg13g2_inv_1
Xu_ppwm_u_ex__0745_ net464 net444 u_ppwm_u_ex__0745_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0957_ VGND VPWR net419 u_ppwm_u_mem__0676_/Y u_ppwm_u_mem__1155_/D
+ u_ppwm_u_mem__0956_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0676_ u_ppwm_u_ex__0676_/Y net458 hold254/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0888_ net513 VPWR u_ppwm_u_mem__0888_/Y VGND net423 net275 sg13g2_o21ai_1
XFILLER_41_0 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1204__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_38_641 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__079_ net441 u_ppwm_u_global_counter__082_/D net442 u_ppwm_u_global_counter__083_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_26_869 VPWR VGND sg13g2_decap_8
XFILLER_38_1019 VPWR VGND sg13g2_decap_8
XFILLER_41_817 VPWR VGND sg13g2_decap_8
XFILLER_34_891 VPWR VGND sg13g2_decap_8
XFILLER_21_596 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_49_928 VPWR VGND sg13g2_decap_8
Xhold31 hold31/A VPWR VGND net229 sg13g2_dlygate4sd3_1
XFILLER_0_467 VPWR VGND sg13g2_decap_8
Xhold20 hold20/A VPWR VGND net218 sg13g2_dlygate4sd3_1
Xhold53 hold53/A VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold42 hold42/A VPWR VGND net240 sg13g2_dlygate4sd3_1
XFILLER_29_630 VPWR VGND sg13g2_decap_8
Xhold64 hold64/A VPWR VGND net262 sg13g2_dlygate4sd3_1
XFILLER_17_803 VPWR VGND sg13g2_decap_8
XFILLER_21_1023 VPWR VGND sg13g2_decap_4
Xhold86 hold86/A VPWR VGND net284 sg13g2_dlygate4sd3_1
Xhold97 hold97/A VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold75 hold75/A VPWR VGND net273 sg13g2_dlygate4sd3_1
XFILLER_44_666 VPWR VGND sg13g2_decap_8
XFILLER_28_195 VPWR VGND sg13g2_fill_2
XFILLER_24_390 VPWR VGND sg13g2_fill_1
XFILLER_12_552 VPWR VGND sg13g2_decap_8
XFILLER_40_894 VPWR VGND sg13g2_decap_8
XFILLER_8_534 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0811_ net476 u_ppwm_u_mem__0616_/Y u_ppwm_u_mem__0810_/Y u_ppwm_u_mem__0811_/X
+ VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_mem__0742_ hold88/A hold69/A net481 u_ppwm_u_mem__0743_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0673_ VPWR u_ppwm_u_mem__0673_/Y net536 VGND sg13g2_inv_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1017 VPWR VGND sg13g2_decap_8
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_48_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1225_ net175 VGND VPWR net567 hold197/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1013_ net508 VPWR u_ppwm_u_ex__1014_/A VGND net451 net350 sg13g2_o21ai_1
XFILLER_35_633 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1156_ net169 VGND VPWR u_ppwm_u_mem__1156_/D hold111/A clknet_5_30__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_mem__1087_ net617 net400 u_ppwm_u_mem__1090_/B VPWR VGND sg13g2_and2_1
XFILLER_23_839 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1102__47 VPWR VGND net47 sg13g2_tiehi
Xu_ppwm_u_ex__0728_ net462 hold313/A u_ppwm_u_ex__0730_/C VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_ex__0659_ u_ppwm_u_ex__0660_/B u_ppwm_u_ex__0659_/B u_ppwm_u_ex__0656_/Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
XFILLER_46_909 VPWR VGND sg13g2_decap_8
XFILLER_45_408 VPWR VGND sg13g2_decap_8
XFILLER_39_983 VPWR VGND sg13g2_decap_8
XFILLER_26_666 VPWR VGND sg13g2_decap_8
XFILLER_41_614 VPWR VGND sg13g2_decap_8
XFILLER_14_839 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_15_22 VPWR VGND sg13g2_fill_2
XFILLER_9_309 VPWR VGND sg13g2_decap_8
XFILLER_22_850 VPWR VGND sg13g2_decap_8
XFILLER_31_32 VPWR VGND sg13g2_fill_2
XFILLER_0_220 VPWR VGND sg13g2_decap_8
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_49_725 VPWR VGND sg13g2_decap_8
XFILLER_0_264 VPWR VGND sg13g2_fill_1
XFILLER_0_297 VPWR VGND sg13g2_decap_4
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_48_257 VPWR VGND sg13g2_decap_8
XFILLER_17_600 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1010_ net495 VPWR u_ppwm_u_mem__1010_/Y VGND net410 hold172/A sg13g2_o21ai_1
XFILLER_45_975 VPWR VGND sg13g2_decap_8
XFILLER_44_463 VPWR VGND sg13g2_decap_8
XFILLER_17_677 VPWR VGND sg13g2_decap_8
XFILLER_32_647 VPWR VGND sg13g2_decap_8
XFILLER_9_810 VPWR VGND sg13g2_decap_8
XFILLER_13_850 VPWR VGND sg13g2_decap_8
XFILLER_20_809 VPWR VGND sg13g2_decap_8
XFILLER_31_146 VPWR VGND sg13g2_fill_1
XFILLER_31_168 VPWR VGND sg13g2_fill_2
XFILLER_40_691 VPWR VGND sg13g2_decap_8
XFILLER_9_887 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0725_ u_ppwm_u_mem__1094_/A net488 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0656_ VPWR u_ppwm_u_mem__0656_/Y net579 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1208_ net57 VGND VPWR u_ppwm_u_mem__1208_/D hold55/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_942 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_3 VPWR VGND uio_oe[0] sg13g2_tielo
Xu_ppwm_u_mem__1139_ net84 VGND VPWR net227 hold191/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_636 VPWR VGND sg13g2_decap_8
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
Xhold320 hold320/A VPWR VGND net688 sg13g2_dlygate4sd3_1
XFILLER_46_706 VPWR VGND sg13g2_decap_8
XFILLER_39_780 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_942 VPWR VGND sg13g2_decap_8
XFILLER_42_901 VPWR VGND sg13g2_decap_8
XFILLER_26_463 VPWR VGND sg13g2_fill_2
XFILLER_14_636 VPWR VGND sg13g2_decap_8
XFILLER_42_978 VPWR VGND sg13g2_decap_8
XFILLER_41_488 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__180_ net636 u_ppwm_u_pwm__180_/C net546 hold269/A VPWR VGND sg13g2_nand3_1
XFILLER_6_835 VPWR VGND sg13g2_decap_8
XFILLER_10_864 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_fill_1
XFILLER_3_47 VPWR VGND sg13g2_fill_2
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_49_599 VPWR VGND sg13g2_decap_8
XFILLER_37_717 VPWR VGND sg13g2_decap_8
XFILLER_18_953 VPWR VGND sg13g2_decap_8
XFILLER_29_290 VPWR VGND sg13g2_fill_2
XFILLER_36_227 VPWR VGND sg13g2_decap_8
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_20_606 VPWR VGND sg13g2_decap_8
XFILLER_33_967 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0993_ net380 net453 u_ppwm_u_ex__0994_/B VPWR VGND sg13g2_xor2_1
XFILLER_9_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0708_ VPWR u_ppwm_u_mem__0708_/Y net543 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0639_ VPWR u_ppwm_u_mem__0639_/Y net568 VGND sg13g2_inv_1
XFILLER_27_227 VPWR VGND sg13g2_fill_1
XFILLER_24_934 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__234__177 VPWR VGND net177 sg13g2_tiehi
Xhold150 hold150/A VPWR VGND net348 sg13g2_dlygate4sd3_1
XFILLER_3_849 VPWR VGND sg13g2_decap_8
Xhold161 hold161/A VPWR VGND net529 sg13g2_dlygate4sd3_1
Xhold194 hold194/A VPWR VGND net562 sg13g2_dlygate4sd3_1
Xhold183 hold183/A VPWR VGND net551 sg13g2_dlygate4sd3_1
Xhold172 hold172/A VPWR VGND net540 sg13g2_dlygate4sd3_1
XFILLER_46_503 VPWR VGND sg13g2_decap_8
XFILLER_15_901 VPWR VGND sg13g2_decap_8
XFILLER_34_709 VPWR VGND sg13g2_decap_8
XFILLER_26_282 VPWR VGND sg13g2_decap_8
XFILLER_33_219 VPWR VGND sg13g2_fill_2
XFILLER_15_978 VPWR VGND sg13g2_decap_8
XFILLER_42_775 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0990_ net497 VPWR u_ppwm_u_mem__0990_/Y VGND net413 hold105/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__232_ net181 VGND VPWR net208 hold9/A clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_10_661 VPWR VGND sg13g2_decap_8
XFILLER_6_632 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__163_ u_ppwm_u_pwm__163_/A u_ppwm_u_pwm__163_/B u_ppwm_u_pwm__238_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_197 VPWR VGND sg13g2_decap_4
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_514 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_18_750 VPWR VGND sg13g2_decap_8
XFILLER_21_904 VPWR VGND sg13g2_decap_8
XFILLER_33_764 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0976_ VGND VPWR u_ppwm_u_ex__0820_/C u_ppwm_u_ex__0972_/Y u_ppwm_u_ex__0976_/Y
+ u_ppwm_u_ex__0975_/Y sg13g2_a21oi_1
Xheichips25_ppwm_24 VPWR VGND uo_out[6] sg13g2_tielo
Xheichips25_ppwm_13 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_28_547 VPWR VGND sg13g2_decap_8
XFILLER_43_517 VPWR VGND sg13g2_decap_8
XFILLER_24_731 VPWR VGND sg13g2_decap_8
XFILLER_12_937 VPWR VGND sg13g2_decap_8
XFILLER_8_919 VPWR VGND sg13g2_decap_8
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_3_646 VPWR VGND sg13g2_decap_8
XFILLER_2_134 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1176__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_2_189 VPWR VGND sg13g2_decap_4
XFILLER_47_823 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_fill_2
XFILLER_46_300 VPWR VGND sg13g2_decap_8
Xfanout471 net472 net471 VPWR VGND sg13g2_buf_8
Xfanout460 net676 net460 VPWR VGND sg13g2_buf_8
Xfanout493 rst_n net493 VPWR VGND sg13g2_buf_8
Xfanout482 net483 net482 VPWR VGND sg13g2_buf_8
XFILLER_19_547 VPWR VGND sg13g2_decap_8
XFILLER_46_377 VPWR VGND sg13g2_decap_8
XFILLER_42_572 VPWR VGND sg13g2_decap_8
XFILLER_15_775 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0830_ u_ppwm_u_ex__0830_/Y net365 u_ppwm_u_ex__0998_/B2 net366 net444
+ VPWR VGND sg13g2_a22oi_1
XFILLER_30_756 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0973_ VGND VPWR net420 u_ppwm_u_mem__0668_/Y u_ppwm_u_mem__1163_/D
+ u_ppwm_u_mem__0972_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0761_ net457 u_ppwm_u_ex__0761_/B u_ppwm_u_ex__0761_/C u_ppwm_u_ex__0761_/Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_31_1003 VPWR VGND sg13g2_decap_8
XFILLER_7_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__215_ u_ppwm_u_pwm__216_/A u_ppwm_u_pwm__215_/B u_ppwm_u_pwm__215_/C
+ u_ppwm_u_pwm__216_/C u_ppwm_u_pwm__215_/Y VPWR VGND sg13g2_nor4_1
Xu_ppwm_u_ex__0692_ VPWR VGND u_ppwm_u_ex__0682_/Y u_ppwm_u_ex__0691_/Y u_ppwm_u_ex__0688_/Y
+ u_ppwm_u_ex__0688_/A u_ppwm_u_ex__0769_/B u_ppwm_u_ex__0686_/Y sg13g2_a221oi_1
Xu_ppwm_u_pwm__146_ VGND VPWR u_ppwm_u_pwm__133_/Y net391 hold6/A u_ppwm_u_pwm__145_/Y
+ sg13g2_a21oi_1
XFILLER_43_4 VPWR VGND sg13g2_fill_2
XFILLER_38_823 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__095_ u_ppwm_u_global_counter__103_/C net608 net622 u_ppwm_u_global_counter__095_/C
+ VPWR VGND sg13g2_and3_2
XFILLER_37_399 VPWR VGND sg13g2_decap_4
XFILLER_40_509 VPWR VGND sg13g2_decap_8
XFILLER_21_701 VPWR VGND sg13g2_decap_8
XFILLER_33_561 VPWR VGND sg13g2_decap_8
XFILLER_20_266 VPWR VGND sg13g2_decap_8
XFILLER_21_778 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0959_ u_ppwm_u_ex__0958_/Y VPWR u_ppwm_u_ex__0959_/Y VGND u_ppwm_u_ex__0839_/Y
+ u_ppwm_u_ex__0847_/Y sg13g2_o21ai_1
XFILLER_20_288 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1207__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_0_649 VPWR VGND sg13g2_decap_8
XFILLER_47_108 VPWR VGND sg13g2_fill_1
XFILLER_29_812 VPWR VGND sg13g2_decap_8
XFILLER_28_355 VPWR VGND sg13g2_fill_1
XFILLER_29_889 VPWR VGND sg13g2_decap_8
XFILLER_44_848 VPWR VGND sg13g2_decap_8
XFILLER_16_517 VPWR VGND sg13g2_decap_8
XFILLER_12_734 VPWR VGND sg13g2_decap_8
XFILLER_8_716 VPWR VGND sg13g2_decap_8
XFILLER_7_204 VPWR VGND sg13g2_decap_8
XFILLER_11_233 VPWR VGND sg13g2_fill_2
XFILLER_4_911 VPWR VGND sg13g2_decap_8
XFILLER_3_443 VPWR VGND sg13g2_decap_8
XFILLER_4_988 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_47_620 VPWR VGND sg13g2_decap_8
XFILLER_19_300 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1172_ net127 VGND VPWR net229 hold105/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_815 VPWR VGND sg13g2_decap_8
XFILLER_47_697 VPWR VGND sg13g2_decap_8
XFILLER_43_881 VPWR VGND sg13g2_decap_8
XFILLER_15_572 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0813_ u_ppwm_u_ex__0799_/A u_ppwm_u_ex__0925_/B net377 u_ppwm_u_ex__0814_/A
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_553 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0744_ u_ppwm_u_ex__0718_/X VPWR u_ppwm_u_ex__0769_/D VGND u_ppwm_u_ex__0740_/Y
+ u_ppwm_u_ex__0743_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__0956_ net502 VPWR u_ppwm_u_mem__0956_/Y VGND net419 net240 sg13g2_o21ai_1
Xu_ppwm_u_ex__0675_ u_ppwm_u_ex__0674_/Y VPWR u_ppwm_u_ex__0678_/B VGND net460 u_ppwm_u_ex__0693_/B
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0887_ VGND VPWR net432 u_ppwm_u_mem__0711_/Y hold78/A u_ppwm_u_mem__0886_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__129_ VPWR u_ppwm_u_pwm__129_/Y net209 VGND sg13g2_inv_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_38_620 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_26_848 VPWR VGND sg13g2_decap_8
XFILLER_38_697 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__078_ u_ppwm_u_global_counter__082_/D net201 hold4/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__1089_ u_ppwm_u_ex__1079_/Y VPWR u_ppwm_u_ex__1089_/Y VGND u_ppwm_u_ex__1078_/Y
+ u_ppwm_u_ex__1080_/Y sg13g2_o21ai_1
XFILLER_25_336 VPWR VGND sg13g2_fill_1
XFILLER_34_870 VPWR VGND sg13g2_decap_8
XFILLER_21_575 VPWR VGND sg13g2_decap_8
XFILLER_4_229 VPWR VGND sg13g2_fill_2
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_49_907 VPWR VGND sg13g2_decap_8
XFILLER_0_446 VPWR VGND sg13g2_decap_8
Xhold10 hold10/A VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold21 hold21/A VPWR VGND net219 sg13g2_dlygate4sd3_1
Xhold32 hold32/A VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_48_439 VPWR VGND sg13g2_decap_8
Xhold54 hold54/A VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold43 hold43/A VPWR VGND net241 sg13g2_dlygate4sd3_1
XFILLER_21_1002 VPWR VGND sg13g2_decap_8
Xhold65 hold65/A VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold76 hold76/A VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold87 hold87/A VPWR VGND net285 sg13g2_dlygate4sd3_1
XFILLER_28_130 VPWR VGND sg13g2_fill_2
Xhold98 hold98/A VPWR VGND net296 sg13g2_dlygate4sd3_1
XFILLER_29_686 VPWR VGND sg13g2_decap_8
XFILLER_44_645 VPWR VGND sg13g2_decap_8
XFILLER_17_859 VPWR VGND sg13g2_decap_8
XFILLER_32_829 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1110__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_40_873 VPWR VGND sg13g2_decap_8
XFILLER_8_513 VPWR VGND sg13g2_decap_8
XFILLER_12_531 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0810_ net471 VPWR u_ppwm_u_mem__0810_/Y VGND hold120/A net476 sg13g2_o21ai_1
Xu_ppwm_u_mem__0741_ hold150/A hold215/A net478 u_ppwm_u_mem__0741_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0672_ VPWR u_ppwm_u_mem__0672_/Y net553 VGND sg13g2_inv_1
XFILLER_4_785 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1224_ net69 VGND VPWR net589 hold219/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1012_ u_ppwm_u_ex__1012_/B net350 u_ppwm_u_ex__1012_/A u_ppwm_u_ex__1012_/Y
+ VPWR VGND u_ppwm_u_ex__1012_/D sg13g2_nand4_1
XFILLER_35_612 VPWR VGND sg13g2_decap_8
XFILLER_47_494 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1155_ net171 VGND VPWR u_ppwm_u_mem__1155_/D hold42/A clknet_5_27__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_34_122 VPWR VGND sg13g2_fill_1
XFILLER_23_818 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1086_ net617 net400 u_ppwm_u_mem__1088_/B VPWR VGND sg13g2_nor2_1
XFILLER_35_689 VPWR VGND sg13g2_decap_8
XFILLER_16_881 VPWR VGND sg13g2_decap_8
XFILLER_31_884 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0727_ net459 hold299/A u_ppwm_u_ex__0732_/C VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0939_ VGND VPWR net421 u_ppwm_u_mem__0685_/Y hold76/A u_ppwm_u_mem__0938_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0658_ u_ppwm_u_ex__0659_/B u_ppwm_u_ex__0660_/A u_ppwm_u_ex__0658_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0589_ VPWR u_ppwm_u_ex__0755_/B hold222/A VGND sg13g2_inv_1
XFILLER_39_962 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_26_645 VPWR VGND sg13g2_decap_8
XFILLER_38_494 VPWR VGND sg13g2_decap_8
XFILLER_14_818 VPWR VGND sg13g2_decap_8
XFILLER_13_317 VPWR VGND sg13g2_decap_4
XFILLER_25_188 VPWR VGND sg13g2_fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_5_549 VPWR VGND sg13g2_decap_8
XFILLER_1_700 VPWR VGND sg13g2_decap_8
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_0_276 VPWR VGND sg13g2_decap_8
XFILLER_48_236 VPWR VGND sg13g2_decap_8
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_17_656 VPWR VGND sg13g2_decap_8
XFILLER_29_483 VPWR VGND sg13g2_fill_2
XFILLER_44_442 VPWR VGND sg13g2_decap_8
XFILLER_32_626 VPWR VGND sg13g2_decap_8
XFILLER_40_670 VPWR VGND sg13g2_decap_8
XFILLER_9_866 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0724_ VPWR u_ppwm_u_mem__0724_/Y u_ppwm_u_mem__1108_/Q VGND sg13g2_inv_1
Xu_ppwm_u_mem__0655_ VPWR u_ppwm_u_mem__0655_/Y net348 VGND sg13g2_inv_1
XFILLER_4_582 VPWR VGND sg13g2_decap_8
XFILLER_36_921 VPWR VGND sg13g2_decap_8
XFILLER_47_291 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1207_ net65 VGND VPWR net254 hold60/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
Xheichips25_ppwm_4 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_23_615 VPWR VGND sg13g2_decap_8
XFILLER_36_998 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1138_ net86 VGND VPWR u_ppwm_u_mem__1138_/D hold126/A clknet_5_30__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1069_ VGND VPWR net401 u_ppwm_u_mem__0620_/Y hold146/A u_ppwm_u_mem__1068_/Y
+ sg13g2_a21oi_1
XFILLER_31_681 VPWR VGND sg13g2_decap_8
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
Xhold310 hold310/A VPWR VGND net678 sg13g2_dlygate4sd3_1
Xhold321 hold321/A VPWR VGND net689 sg13g2_dlygate4sd3_1
XFILLER_27_921 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_38_291 VPWR VGND sg13g2_decap_4
XFILLER_26_55 VPWR VGND sg13g2_fill_1
XFILLER_27_998 VPWR VGND sg13g2_decap_8
XFILLER_42_957 VPWR VGND sg13g2_decap_8
XFILLER_14_615 VPWR VGND sg13g2_decap_8
XFILLER_26_99 VPWR VGND sg13g2_fill_2
XFILLER_41_467 VPWR VGND sg13g2_decap_8
XFILLER_10_843 VPWR VGND sg13g2_decap_8
XFILLER_6_814 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_49_578 VPWR VGND sg13g2_decap_8
XFILLER_18_932 VPWR VGND sg13g2_decap_8
XFILLER_45_751 VPWR VGND sg13g2_decap_8
XFILLER_32_412 VPWR VGND sg13g2_fill_1
XFILLER_33_946 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0992_ net453 net380 u_ppwm_u_ex__0992_/X VPWR VGND sg13g2_and2_1
XFILLER_32_456 VPWR VGND sg13g2_fill_1
XFILLER_9_663 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0707_ VPWR u_ppwm_u_mem__0707_/Y net558 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0638_ VPWR u_ppwm_u_mem__0638_/Y net230 VGND sg13g2_inv_1
XFILLER_41_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_729 VPWR VGND sg13g2_decap_8
XFILLER_24_913 VPWR VGND sg13g2_decap_8
XFILLER_36_795 VPWR VGND sg13g2_decap_8
XFILLER_23_489 VPWR VGND sg13g2_decap_8
XFILLER_32_990 VPWR VGND sg13g2_decap_8
XFILLER_3_828 VPWR VGND sg13g2_decap_8
Xhold151 hold151/A VPWR VGND net519 sg13g2_dlygate4sd3_1
Xhold140 hold140/A VPWR VGND net338 sg13g2_dlygate4sd3_1
Xhold162 hold162/A VPWR VGND net530 sg13g2_dlygate4sd3_1
Xhold173 hold173/A VPWR VGND net541 sg13g2_dlygate4sd3_1
Xhold184 hold184/A VPWR VGND net552 sg13g2_dlygate4sd3_1
Xhold195 hold195/A VPWR VGND net563 sg13g2_dlygate4sd3_1
XFILLER_19_729 VPWR VGND sg13g2_decap_8
XFILLER_46_559 VPWR VGND sg13g2_decap_8
XFILLER_2_1010 VPWR VGND sg13g2_decap_8
XFILLER_37_43 VPWR VGND sg13g2_fill_1
XFILLER_27_795 VPWR VGND sg13g2_decap_8
XFILLER_42_754 VPWR VGND sg13g2_decap_8
XFILLER_15_957 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_41_286 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_pwm__231_ net183 VGND VPWR net534 hold165/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_6_611 VPWR VGND sg13g2_decap_8
XFILLER_10_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__162_ net489 VPWR u_ppwm_u_pwm__163_/B VGND net625 net647 sg13g2_o21ai_1
XFILLER_6_688 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_33_743 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_32_264 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0975_ net353 VPWR u_ppwm_u_ex__0975_/Y VGND net361 u_ppwm_u_ex__0974_/Y
+ sg13g2_o21ai_1
XFILLER_20_459 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1201__113 VPWR VGND net113 sg13g2_tiehi
Xheichips25_ppwm_25 VPWR VGND uo_out[7] sg13g2_tielo
Xheichips25_ppwm_14 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_24_710 VPWR VGND sg13g2_decap_8
XFILLER_23_220 VPWR VGND sg13g2_decap_4
XFILLER_36_592 VPWR VGND sg13g2_decap_8
XFILLER_12_916 VPWR VGND sg13g2_decap_8
XFILLER_24_787 VPWR VGND sg13g2_decap_8
XFILLER_23_275 VPWR VGND sg13g2_decap_4
XFILLER_23_297 VPWR VGND sg13g2_fill_2
XFILLER_3_625 VPWR VGND sg13g2_decap_8
XFILLER_2_113 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_157 VPWR VGND sg13g2_fill_1
XFILLER_48_42 VPWR VGND sg13g2_decap_8
Xfanout450 net681 net450 VPWR VGND sg13g2_buf_8
XFILLER_24_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_802 VPWR VGND sg13g2_decap_8
Xfanout461 hold308/A net461 VPWR VGND sg13g2_buf_1
Xfanout472 hold321/A net472 VPWR VGND sg13g2_buf_8
Xfanout483 net486 net483 VPWR VGND sg13g2_buf_8
XFILLER_19_526 VPWR VGND sg13g2_decap_8
Xfanout494 net495 net494 VPWR VGND sg13g2_buf_8
XFILLER_47_879 VPWR VGND sg13g2_decap_8
XFILLER_46_356 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_15_754 VPWR VGND sg13g2_decap_8
XFILLER_27_592 VPWR VGND sg13g2_decap_8
XFILLER_42_551 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1126__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_30_735 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0972_ net503 VPWR u_ppwm_u_mem__0972_/Y VGND net420 net286 sg13g2_o21ai_1
Xu_ppwm_u_ex__0760_ u_ppwm_u_ex__0760_/A u_ppwm_u_ex__0761_/C u_ppwm_u_ex__0760_/C
+ u_ppwm_u_ex__0760_/D u_ppwm_u_ex__0763_/A VPWR VGND sg13g2_nor4_1
XFILLER_7_920 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__214_ hold233/A u_ppwm_u_pwm__214_/B u_ppwm_u_pwm__216_/C VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_ex__0691_ VPWR u_ppwm_u_ex__0691_/Y net366 VGND sg13g2_inv_1
Xu_ppwm_u_pwm__145_ net493 VPWR u_ppwm_u_pwm__145_/Y VGND net463 net390 sg13g2_o21ai_1
Xu_ppwm_u_mem__1216__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_7_997 VPWR VGND sg13g2_decap_8
XFILLER_6_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1120__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_802 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_37_323 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__094_ net609 u_ppwm_u_global_counter__093_/Y hold242/A VPWR
+ VGND sg13g2_nor2b_1
XFILLER_38_879 VPWR VGND sg13g2_decap_8
XFILLER_33_540 VPWR VGND sg13g2_decap_8
XFILLER_20_223 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0958_ u_ppwm_u_ex__0958_/Y u_ppwm_u_ex__0870_/Y net368 u_ppwm_u_ex__0838_/B
+ u_ppwm_u_ex__0799_/A VPWR VGND sg13g2_a22oi_1
XFILLER_21_757 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0889_ u_ppwm_u_ex__0888_/Y VPWR u_ppwm_u_ex__0890_/B VGND u_ppwm_u_ex__0795_/Y
+ u_ppwm_u_ex__0839_/Y sg13g2_o21ai_1
XFILLER_0_628 VPWR VGND sg13g2_decap_8
XFILLER_18_45 VPWR VGND sg13g2_fill_1
XFILLER_29_868 VPWR VGND sg13g2_decap_8
XFILLER_44_827 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1143__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_12_713 VPWR VGND sg13g2_decap_8
XFILLER_24_584 VPWR VGND sg13g2_decap_8
XFILLER_7_227 VPWR VGND sg13g2_fill_1
XFILLER_4_967 VPWR VGND sg13g2_decap_8
XFILLER_3_422 VPWR VGND sg13g2_decap_8
XFILLER_3_499 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1171_ net131 VGND VPWR net304 hold53/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_676 VPWR VGND sg13g2_decap_8
XFILLER_34_304 VPWR VGND sg13g2_fill_1
XFILLER_46_197 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_34_359 VPWR VGND sg13g2_fill_2
XFILLER_43_860 VPWR VGND sg13g2_decap_8
XFILLER_15_551 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0812_ u_ppwm_u_ex__0651_/A u_ppwm_u_ex__0758_/A u_ppwm_u_ex__0979_/A
+ u_ppwm_u_ex__0812_/X VPWR VGND sg13g2_mux2_1
XFILLER_30_532 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1114__46 VPWR VGND net46 sg13g2_tiehi
Xu_ppwm_u_mem__0955_ VGND VPWR net419 u_ppwm_u_mem__0677_/Y hold43/A u_ppwm_u_mem__0954_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0743_ net356 VPWR u_ppwm_u_ex__0743_/Y VGND u_ppwm_u_ex__0739_/A u_ppwm_u_ex__0737_/Y
+ sg13g2_o21ai_1
XFILLER_7_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0674_ u_ppwm_u_ex__0674_/Y hold254/A net458 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0886_ net513 VPWR u_ppwm_u_mem__0886_/Y VGND net432 hold95/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__128_ VPWR u_ppwm_u_pwm__128_/Y net211 VGND sg13g2_inv_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_37_142 VPWR VGND sg13g2_fill_2
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_26_827 VPWR VGND sg13g2_decap_8
XFILLER_38_676 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1088_ u_ppwm_u_ex__1088_/A u_ppwm_u_ex__1086_/Y u_ppwm_u_ex__1123_/D
+ VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_global_counter__077_ u_ppwm_u_global_counter__082_/D net631 hold264/A VPWR
+ VGND sg13g2_nor2_1
XFILLER_19_890 VPWR VGND sg13g2_decap_8
XFILLER_21_554 VPWR VGND sg13g2_decap_8
XFILLER_14_1021 VPWR VGND sg13g2_decap_8
XFILLER_0_425 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
XFILLER_48_418 VPWR VGND sg13g2_decap_8
Xhold11 hold11/A VPWR VGND net209 sg13g2_dlygate4sd3_1
Xhold22 hold22/A VPWR VGND net220 sg13g2_dlygate4sd3_1
Xhold55 hold55/A VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold44 hold44/A VPWR VGND net242 sg13g2_dlygate4sd3_1
Xhold33 hold33/A VPWR VGND net231 sg13g2_dlygate4sd3_1
Xhold66 hold66/A VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold88 hold88/A VPWR VGND net286 sg13g2_dlygate4sd3_1
Xhold99 hold99/A VPWR VGND net297 sg13g2_dlygate4sd3_1
Xhold77 hold77/A VPWR VGND net275 sg13g2_dlygate4sd3_1
XFILLER_29_665 VPWR VGND sg13g2_decap_8
XFILLER_44_624 VPWR VGND sg13g2_decap_8
XFILLER_17_838 VPWR VGND sg13g2_decap_8
XFILLER_16_326 VPWR VGND sg13g2_fill_1
XFILLER_32_808 VPWR VGND sg13g2_decap_8
XFILLER_12_510 VPWR VGND sg13g2_decap_8
XFILLER_40_852 VPWR VGND sg13g2_decap_8
XFILLER_12_587 VPWR VGND sg13g2_decap_8
XFILLER_8_569 VPWR VGND sg13g2_decap_8
XFILLER_6_15 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0740_ u_ppwm_u_mem__0739_/Y VPWR u_ppwm_u_mem__1228_/D VGND net619
+ u_ppwm_u_mem__0737_/D sg13g2_o21ai_1
Xu_ppwm_u_mem__0671_ VPWR u_ppwm_u_mem__0671_/Y net271 VGND sg13g2_inv_1
XFILLER_4_764 VPWR VGND sg13g2_decap_8
XFILLER_0_992 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1223_ net133 VGND VPWR u_ppwm_u_mem__1223_/D hold250/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1011_ u_ppwm_u_ex__1012_/D u_ppwm_u_ex__1010_/Y u_ppwm_u_ex__0784_/A
+ u_ppwm_u_ex__1007_/Y u_ppwm_u_ex__1017_/B VPWR VGND sg13g2_a22oi_1
XFILLER_48_985 VPWR VGND sg13g2_decap_8
XFILLER_47_473 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1154_ net173 VGND VPWR net241 hold71/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_860 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1085_ u_ppwm_u_mem__1103_/A net488 u_ppwm_u_mem__1085_/B VPWR VGND
+ sg13g2_nand2_2
XFILLER_35_668 VPWR VGND sg13g2_decap_8
XFILLER_31_863 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0938_ net502 VPWR u_ppwm_u_mem__0938_/Y VGND net421 hold137/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0726_ hold299/A net459 u_ppwm_u_ex__0730_/A VPWR VGND sg13g2_nor2b_1
XFILLER_7_591 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0657_ net441 hold289/A u_ppwm_u_ex__0660_/A VPWR VGND sg13g2_xor2_1
Xu_ppwm_u_mem__0869_ VGND VPWR net433 u_ppwm_u_mem__0720_/Y u_ppwm_u_mem__1111_/D
+ u_ppwm_u_mem__0868_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0588_ VPWR u_ppwm_u_ex__0761_/B hold236/A VGND sg13g2_inv_1
XFILLER_39_941 VPWR VGND sg13g2_decap_8
XFILLER_26_624 VPWR VGND sg13g2_decap_8
XFILLER_41_649 VPWR VGND sg13g2_decap_8
XFILLER_22_885 VPWR VGND sg13g2_decap_8
XFILLER_5_528 VPWR VGND sg13g2_decap_8
XFILLER_0_255 VPWR VGND sg13g2_decap_8
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_48_215 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_44_421 VPWR VGND sg13g2_decap_8
XFILLER_17_635 VPWR VGND sg13g2_decap_8
XFILLER_32_605 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_9_845 VPWR VGND sg13g2_decap_8
XFILLER_13_885 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0723_ VPWR u_ppwm_u_mem__0723_/Y net577 VGND sg13g2_inv_1
XFILLER_4_561 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0654_ VPWR u_ppwm_u_mem__0654_/Y net265 VGND sg13g2_inv_1
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
XFILLER_48_782 VPWR VGND sg13g2_decap_8
XFILLER_36_900 VPWR VGND sg13g2_decap_8
XFILLER_47_270 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1206_ net73 VGND VPWR net259 hold103/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
Xheichips25_ppwm_5 VPWR VGND uio_oe[2] sg13g2_tielo
Xu_ppwm_u_mem__1137_ net88 VGND VPWR net325 hold186/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_977 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1068_ net488 VPWR u_ppwm_u_mem__1068_/Y VGND net401 hold169/A sg13g2_o21ai_1
XFILLER_31_660 VPWR VGND sg13g2_decap_8
Xhold300 hold300/A VPWR VGND net668 sg13g2_dlygate4sd3_1
Xhold311 hold311/A VPWR VGND net679 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0709_ u_ppwm_u_ex__0709_/Y u_ppwm_u_ex__0973_/A hold217/A VPWR VGND
+ sg13g2_nand2_1
Xhold322 hold324/A VPWR VGND net690 sg13g2_dlygate4sd3_1
XFILLER_27_900 VPWR VGND sg13g2_decap_8
XFILLER_38_270 VPWR VGND sg13g2_fill_1
XFILLER_27_977 VPWR VGND sg13g2_decap_8
XFILLER_42_936 VPWR VGND sg13g2_decap_8
XFILLER_26_78 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_decap_4
XFILLER_41_446 VPWR VGND sg13g2_decap_8
XFILLER_10_822 VPWR VGND sg13g2_decap_8
XFILLER_22_682 VPWR VGND sg13g2_decap_8
XFILLER_10_899 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_18_911 VPWR VGND sg13g2_decap_8
XFILLER_45_730 VPWR VGND sg13g2_decap_8
XFILLER_18_988 VPWR VGND sg13g2_decap_8
XFILLER_29_292 VPWR VGND sg13g2_fill_1
XFILLER_33_925 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0991_ u_ppwm_u_ex__0991_/A u_ppwm_u_ex__0991_/B u_ppwm_u_ex__1115_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_1024 VPWR VGND sg13g2_decap_4
XFILLER_9_642 VPWR VGND sg13g2_decap_8
XFILLER_13_682 VPWR VGND sg13g2_decap_8
XFILLER_5_892 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0706_ VPWR u_ppwm_u_mem__0706_/Y net529 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0637_ VPWR u_ppwm_u_mem__0637_/Y net305 VGND sg13g2_inv_1
XFILLER_41_1006 VPWR VGND sg13g2_decap_8
XFILLER_28_708 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1130__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_36_774 VPWR VGND sg13g2_decap_8
XFILLER_24_969 VPWR VGND sg13g2_decap_8
XFILLER_10_107 VPWR VGND sg13g2_decap_4
XFILLER_3_807 VPWR VGND sg13g2_decap_8
XFILLER_2_339 VPWR VGND sg13g2_fill_1
Xhold130 hold130/A VPWR VGND net328 sg13g2_dlygate4sd3_1
Xhold141 hold141/A VPWR VGND net339 sg13g2_dlygate4sd3_1
Xhold152 hold152/A VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold185 hold185/A VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold163 hold163/A VPWR VGND net531 sg13g2_dlygate4sd3_1
Xhold174 hold174/A VPWR VGND net542 sg13g2_dlygate4sd3_1
Xhold196 hold196/A VPWR VGND net564 sg13g2_dlygate4sd3_1
XFILLER_19_708 VPWR VGND sg13g2_decap_8
XFILLER_46_538 VPWR VGND sg13g2_decap_8
XFILLER_18_229 VPWR VGND sg13g2_decap_8
XFILLER_15_936 VPWR VGND sg13g2_decap_8
XFILLER_27_774 VPWR VGND sg13g2_decap_8
XFILLER_42_733 VPWR VGND sg13g2_decap_8
XFILLER_41_232 VPWR VGND sg13g2_fill_1
XFILLER_30_917 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__230_ net185 VGND VPWR net204 hold5/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__161_ net625 net647 u_ppwm_u_pwm__163_/A VPWR VGND sg13g2_and2_1
XFILLER_10_696 VPWR VGND sg13g2_decap_8
XFILLER_6_667 VPWR VGND sg13g2_decap_8
XFILLER_2_884 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_37_549 VPWR VGND sg13g2_decap_8
XFILLER_17_273 VPWR VGND sg13g2_fill_2
XFILLER_18_785 VPWR VGND sg13g2_decap_8
XFILLER_33_722 VPWR VGND sg13g2_decap_8
XFILLER_21_939 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0974_ VPWR VGND hold217/A u_ppwm_u_ex__0973_/Y net364 net441 u_ppwm_u_ex__0974_/Y
+ net366 sg13g2_a221oi_1
XFILLER_20_438 VPWR VGND sg13g2_decap_8
XFILLER_33_799 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_15 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_36_571 VPWR VGND sg13g2_decap_8
XFILLER_23_232 VPWR VGND sg13g2_decap_8
XFILLER_23_243 VPWR VGND sg13g2_fill_2
XFILLER_23_254 VPWR VGND sg13g2_fill_1
XFILLER_24_766 VPWR VGND sg13g2_decap_8
XFILLER_23_57 VPWR VGND sg13g2_fill_1
XFILLER_3_604 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 net633 net440 VPWR VGND sg13g2_buf_8
XFILLER_48_65 VPWR VGND sg13g2_fill_1
Xfanout462 net690 net462 VPWR VGND sg13g2_buf_8
XFILLER_19_505 VPWR VGND sg13g2_decap_8
Xfanout451 net668 net451 VPWR VGND sg13g2_buf_8
Xfanout473 net475 net473 VPWR VGND sg13g2_buf_8
Xfanout484 net486 net484 VPWR VGND sg13g2_buf_8
Xfanout495 net500 net495 VPWR VGND sg13g2_buf_8
XFILLER_47_858 VPWR VGND sg13g2_decap_8
XFILLER_46_335 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_27_571 VPWR VGND sg13g2_decap_8
XFILLER_42_530 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_15_733 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0971_ VGND VPWR net419 u_ppwm_u_mem__0669_/Y hold89/A u_ppwm_u_mem__0970_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__213_ hold284/A u_ppwm_u_pwm__213_/B u_ppwm_u_pwm__215_/C VPWR VGND
+ sg13g2_nor2_1
XFILLER_11_994 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0690_ net379 u_ppwm_u_ex__0983_/B fanout367/A VPWR VGND sg13g2_and2_1
XFILLER_7_976 VPWR VGND sg13g2_decap_8
XFILLER_6_442 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__144_ VGND VPWR u_ppwm_u_pwm__134_/Y net390 hold18/A u_ppwm_u_pwm__143_/Y
+ sg13g2_a21oi_1
XFILLER_6_464 VPWR VGND sg13g2_decap_8
XFILLER_9_1006 VPWR VGND sg13g2_decap_8
XFILLER_2_681 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_49_151 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__093_ fanout392/A u_ppwm_u_global_counter__095_/C net608
+ u_ppwm_u_global_counter__093_/Y VPWR VGND sg13g2_nand3_1
XFILLER_38_858 VPWR VGND sg13g2_decap_8
XFILLER_25_519 VPWR VGND sg13g2_decap_8
XFILLER_18_582 VPWR VGND sg13g2_decap_8
XFILLER_20_202 VPWR VGND sg13g2_fill_1
XFILLER_21_736 VPWR VGND sg13g2_decap_8
XFILLER_33_596 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0957_ u_ppwm_u_ex__0956_/Y VPWR u_ppwm_u_ex__0964_/B VGND u_ppwm_u_ex__0953_/Y
+ u_ppwm_u_ex__0955_/X sg13g2_o21ai_1
Xu_ppwm_u_ex__0888_ u_ppwm_u_ex__0888_/Y net368 u_ppwm_u_ex__0800_/X VPWR VGND sg13g2_nand2b_1
XFILLER_47_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_607 VPWR VGND sg13g2_decap_8
XFILLER_29_847 VPWR VGND sg13g2_decap_8
XFILLER_44_806 VPWR VGND sg13g2_decap_8
XFILLER_36_390 VPWR VGND sg13g2_fill_2
XFILLER_24_563 VPWR VGND sg13g2_decap_8
XFILLER_12_769 VPWR VGND sg13g2_decap_8
Xclkload0 VPWR clkload0/Y clknet_5_1__leaf_clk VGND sg13g2_inv_1
XFILLER_11_268 VPWR VGND sg13g2_decap_4
XFILLER_4_946 VPWR VGND sg13g2_decap_8
XFILLER_3_478 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_655 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1170_ net135 VGND VPWR net252 hold69/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_335 VPWR VGND sg13g2_fill_2
XFILLER_15_530 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0811_ net459 hold299/A net386 u_ppwm_u_ex__0925_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0954_ net502 VPWR u_ppwm_u_mem__0954_/Y VGND net419 hold71/A sg13g2_o21ai_1
XFILLER_30_588 VPWR VGND sg13g2_decap_8
XFILLER_11_791 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0742_ net387 net363 fanout356/A VPWR VGND sg13g2_nor2_2
XFILLER_7_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0673_ net463 u_ppwm_u_ex__0673_/B u_ppwm_u_ex__0673_/C u_ppwm_u_ex__0678_/A
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__0885_ VGND VPWR net432 u_ppwm_u_mem__0712_/Y hold96/A u_ppwm_u_mem__0884_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__127_ VPWR u_ppwm_u_pwm__218_/B net238 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1159__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_26_806 VPWR VGND sg13g2_decap_8
XFILLER_37_132 VPWR VGND sg13g2_fill_2
XFILLER_38_655 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__076_ VGND VPWR net604 u_ppwm_u_global_counter__073_/B hold263/A
+ net630 sg13g2_a21oi_1
Xu_ppwm_u_ex__1087_ net491 VPWR u_ppwm_u_ex__1088_/A VGND net663 net349 sg13g2_o21ai_1
XFILLER_25_349 VPWR VGND sg13g2_decap_8
XFILLER_21_533 VPWR VGND sg13g2_decap_8
XFILLER_14_1000 VPWR VGND sg13g2_decap_8
XFILLER_0_404 VPWR VGND sg13g2_decap_8
XFILLER_1_938 VPWR VGND sg13g2_decap_8
Xhold12 hold12/A VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold23 hold23/A VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold56 hold56/A VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold34 hold34/A VPWR VGND net232 sg13g2_dlygate4sd3_1
Xhold45 hold45/A VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold89 hold89/A VPWR VGND net287 sg13g2_dlygate4sd3_1
Xhold67 hold67/A VPWR VGND net265 sg13g2_dlygate4sd3_1
XFILLER_28_132 VPWR VGND sg13g2_fill_1
XFILLER_29_644 VPWR VGND sg13g2_decap_8
Xhold78 hold78/A VPWR VGND net276 sg13g2_dlygate4sd3_1
XFILLER_44_603 VPWR VGND sg13g2_decap_8
XFILLER_17_817 VPWR VGND sg13g2_decap_8
XFILLER_28_143 VPWR VGND sg13g2_fill_2
XFILLER_25_883 VPWR VGND sg13g2_decap_8
XFILLER_40_831 VPWR VGND sg13g2_decap_8
XFILLER_12_566 VPWR VGND sg13g2_decap_8
XFILLER_8_548 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0670_ VPWR u_ppwm_u_mem__0670_/Y net317 VGND sg13g2_inv_1
XFILLER_4_743 VPWR VGND sg13g2_decap_8
XFILLER_10_91 VPWR VGND sg13g2_fill_2
XFILLER_0_971 VPWR VGND sg13g2_decap_8
XFILLER_48_964 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1010_ u_ppwm_u_ex__1010_/Y u_ppwm_u_ex__1010_/A u_ppwm_u_ex__1010_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1222_ net172 VGND VPWR u_ppwm_u_mem__1222_/D hold238/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_47_452 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1153_ net56 VGND VPWR net270 hold174/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_647 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1084_ u_ppwm_u_mem__1085_/B net333 VPWR VGND net400 sg13g2_nand2b_2
XFILLER_22_308 VPWR VGND sg13g2_fill_2
XFILLER_37_1011 VPWR VGND sg13g2_decap_8
XFILLER_31_842 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0725_ u_ppwm_u_ex__0724_/Y VPWR u_ppwm_u_ex__0725_/Y VGND net452 u_ppwm_u_ex__0850_/A
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0937_ VGND VPWR net417 u_ppwm_u_mem__0686_/Y u_ppwm_u_mem__1145_/D
+ u_ppwm_u_mem__0936_/Y sg13g2_a21oi_1
XFILLER_7_570 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0868_ net515 VPWR u_ppwm_u_mem__0868_/Y VGND net433 net242 sg13g2_o21ai_1
Xu_ppwm_u_ex__0656_ u_ppwm_u_ex__0655_/Y VPWR u_ppwm_u_ex__0656_/Y VGND u_ppwm_u_ex__0735_/A
+ hold262/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0799_ u_ppwm_u_mem__0799_/Y net472 u_ppwm_u_mem__0799_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_ex__0587_ VPWR u_ppwm_u_ex__0673_/B net440 VGND sg13g2_inv_1
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_920 VPWR VGND sg13g2_decap_8
XFILLER_39_997 VPWR VGND sg13g2_decap_8
XFILLER_26_603 VPWR VGND sg13g2_decap_8
XFILLER_38_441 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__059_ VPWR u_ppwm_u_global_counter__075_/A net398 VGND sg13g2_inv_1
XFILLER_41_628 VPWR VGND sg13g2_decap_8
XFILLER_33_190 VPWR VGND sg13g2_fill_1
XFILLER_22_864 VPWR VGND sg13g2_decap_8
XFILLER_5_507 VPWR VGND sg13g2_decap_8
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_0_234 VPWR VGND sg13g2_fill_2
XFILLER_49_739 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_44_400 VPWR VGND sg13g2_decap_8
XFILLER_17_614 VPWR VGND sg13g2_decap_8
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_44_477 VPWR VGND sg13g2_decap_8
XFILLER_25_680 VPWR VGND sg13g2_decap_8
XFILLER_9_824 VPWR VGND sg13g2_decap_8
XFILLER_13_864 VPWR VGND sg13g2_decap_8
XFILLER_8_356 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0722_ VPWR u_ppwm_u_mem__0722_/Y net341 VGND sg13g2_inv_1
XFILLER_4_540 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0653_ VPWR u_ppwm_u_mem__0653_/Y net255 VGND sg13g2_inv_1
XFILLER_48_761 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1205_ net81 VGND VPWR net302 hold114/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1117__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_36_956 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_6 VPWR VGND uio_oe[3] sg13g2_tielo
Xu_ppwm_u_mem__1136_ net90 VGND VPWR net555 hold131/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1067_ VGND VPWR net401 u_ppwm_u_mem__0621_/Y u_ppwm_u_mem__1210_/D
+ u_ppwm_u_mem__1066_/Y sg13g2_a21oi_1
Xhold301 hold301/A VPWR VGND net669 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0708_ u_ppwm_u_ex__0707_/Y VPWR u_ppwm_u_ex__0708_/Y VGND u_ppwm_u_ex__0704_/Y
+ u_ppwm_u_ex__0706_/Y sg13g2_o21ai_1
Xhold312 hold312/A VPWR VGND net680 sg13g2_dlygate4sd3_1
Xhold323 hold323/A VPWR VGND net691 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0639_ net501 VPWR hold316/A VGND net468 net447 sg13g2_o21ai_1
XFILLER_39_794 VPWR VGND sg13g2_decap_8
XFILLER_27_956 VPWR VGND sg13g2_decap_8
XFILLER_42_915 VPWR VGND sg13g2_decap_8
XFILLER_41_425 VPWR VGND sg13g2_decap_8
XFILLER_10_801 VPWR VGND sg13g2_decap_8
XFILLER_22_661 VPWR VGND sg13g2_decap_8
XFILLER_10_878 VPWR VGND sg13g2_decap_8
XFILLER_6_849 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_4
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_17_400 VPWR VGND sg13g2_decap_4
XFILLER_29_260 VPWR VGND sg13g2_fill_2
XFILLER_17_433 VPWR VGND sg13g2_fill_2
XFILLER_18_967 VPWR VGND sg13g2_decap_8
XFILLER_33_904 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_8
XFILLER_17_488 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0990_ u_ppwm_u_ex__0989_/Y VPWR u_ppwm_u_ex__0991_/B VGND net660 net350
+ sg13g2_o21ai_1
XFILLER_13_661 VPWR VGND sg13g2_decap_8
XFILLER_34_1003 VPWR VGND sg13g2_decap_8
XFILLER_41_992 VPWR VGND sg13g2_decap_8
XFILLER_9_621 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1227__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_9_698 VPWR VGND sg13g2_decap_8
XFILLER_5_871 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0705_ VPWR u_ppwm_u_mem__0705_/Y net331 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0636_ VPWR u_ppwm_u_mem__0636_/Y net232 VGND sg13g2_inv_1
XFILLER_36_753 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1119_ net124 VGND VPWR net294 hold164/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_24_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1210__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_11_609 VPWR VGND sg13g2_decap_8
XFILLER_2_307 VPWR VGND sg13g2_fill_2
Xhold131 hold131/A VPWR VGND net329 sg13g2_dlygate4sd3_1
Xhold120 hold120/A VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold142 hold142/A VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold153 hold153/A VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold164 hold164/A VPWR VGND net532 sg13g2_dlygate4sd3_1
Xhold186 hold186/A VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold175 hold175/A VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold197 hold197/A VPWR VGND net565 sg13g2_dlygate4sd3_1
XFILLER_46_517 VPWR VGND sg13g2_decap_8
XFILLER_27_753 VPWR VGND sg13g2_decap_8
XFILLER_39_591 VPWR VGND sg13g2_decap_8
XFILLER_42_712 VPWR VGND sg13g2_decap_8
XFILLER_15_915 VPWR VGND sg13g2_decap_8
XFILLER_26_252 VPWR VGND sg13g2_fill_2
XFILLER_18_1009 VPWR VGND sg13g2_decap_8
XFILLER_26_296 VPWR VGND sg13g2_decap_8
XFILLER_42_789 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__160_ VGND VPWR u_ppwm_u_pwm__223_/B net390 hold102/A u_ppwm_u_pwm__159_/Y
+ sg13g2_a21oi_1
XFILLER_5_112 VPWR VGND sg13g2_fill_1
XFILLER_10_675 VPWR VGND sg13g2_decap_8
XFILLER_6_646 VPWR VGND sg13g2_decap_8
XFILLER_2_863 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_37_528 VPWR VGND sg13g2_decap_8
XFILLER_18_764 VPWR VGND sg13g2_decap_8
XFILLER_33_701 VPWR VGND sg13g2_decap_8
XFILLER_45_583 VPWR VGND sg13g2_decap_8
XFILLER_21_918 VPWR VGND sg13g2_decap_8
XFILLER_32_255 VPWR VGND sg13g2_decap_8
XFILLER_33_778 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0973_ u_ppwm_u_ex__0973_/A net366 net364 u_ppwm_u_ex__0973_/Y VPWR VGND
+ sg13g2_nor3_1
XFILLER_9_495 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0619_ VPWR u_ppwm_u_mem__0619_/Y net307 VGND sg13g2_inv_1
Xheichips25_ppwm_16 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_36_550 VPWR VGND sg13g2_decap_8
XFILLER_24_745 VPWR VGND sg13g2_decap_8
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
XFILLER_20_984 VPWR VGND sg13g2_decap_8
XFILLER_2_148 VPWR VGND sg13g2_decap_8
Xfanout430 net431 net430 VPWR VGND sg13g2_buf_1
Xfanout441 net639 net441 VPWR VGND sg13g2_buf_8
Xfanout463 net680 net463 VPWR VGND sg13g2_buf_8
Xfanout452 hold300/A net452 VPWR VGND sg13g2_buf_1
Xfanout474 net475 net474 VPWR VGND sg13g2_buf_1
XFILLER_47_837 VPWR VGND sg13g2_decap_8
XFILLER_46_314 VPWR VGND sg13g2_decap_8
Xfanout496 net499 net496 VPWR VGND sg13g2_buf_8
Xfanout485 net486 net485 VPWR VGND sg13g2_buf_8
XFILLER_15_712 VPWR VGND sg13g2_decap_8
XFILLER_27_550 VPWR VGND sg13g2_decap_8
XFILLER_14_255 VPWR VGND sg13g2_decap_8
XFILLER_42_586 VPWR VGND sg13g2_decap_8
XFILLER_14_266 VPWR VGND sg13g2_fill_1
XFILLER_15_789 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0970_ net503 VPWR u_ppwm_u_mem__0970_/Y VGND net419 hold119/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__212_ u_ppwm_u_pwm__213_/B hold284/A u_ppwm_u_pwm__210_/Y u_ppwm_u_pwm__215_/B
+ VPWR VGND sg13g2_a21o_1
XFILLER_14_299 VPWR VGND sg13g2_decap_8
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_31_1017 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_955 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__143_ net492 VPWR u_ppwm_u_pwm__143_/Y VGND net465 net390 sg13g2_o21ai_1
XFILLER_2_660 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_38_837 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__092_ VGND VPWR net392 u_ppwm_u_global_counter__095_/C hold241/A
+ net608 sg13g2_a21oi_1
XFILLER_18_561 VPWR VGND sg13g2_decap_8
XFILLER_46_881 VPWR VGND sg13g2_decap_8
XFILLER_45_380 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1117__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_21_715 VPWR VGND sg13g2_decap_8
XFILLER_33_575 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0956_ VGND VPWR u_ppwm_u_ex__0953_/Y u_ppwm_u_ex__0955_/X u_ppwm_u_ex__0956_/Y
+ net357 sg13g2_a21oi_1
Xu_ppwm_u_ex__0887_ u_ppwm_u_ex__0820_/C VPWR u_ppwm_u_ex__0890_/A VGND u_ppwm_u_ex__0816_/B
+ u_ppwm_u_ex__0842_/B sg13g2_o21ai_1
XFILLER_29_826 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_fill_2
XFILLER_28_369 VPWR VGND sg13g2_decap_8
XFILLER_37_892 VPWR VGND sg13g2_decap_8
XFILLER_24_542 VPWR VGND sg13g2_decap_8
XFILLER_11_203 VPWR VGND sg13g2_fill_2
XFILLER_11_214 VPWR VGND sg13g2_decap_4
XFILLER_12_748 VPWR VGND sg13g2_decap_8
XFILLER_7_218 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_5_3__leaf_clk clkload1/X VPWR VGND sg13g2_buf_1
XFILLER_20_781 VPWR VGND sg13g2_decap_8
XFILLER_4_925 VPWR VGND sg13g2_decap_8
XFILLER_3_457 VPWR VGND sg13g2_decap_8
XFILLER_47_634 VPWR VGND sg13g2_decap_8
XFILLER_46_111 VPWR VGND sg13g2_fill_2
XFILLER_46_155 VPWR VGND sg13g2_fill_1
XFILLER_35_829 VPWR VGND sg13g2_decap_8
XFILLER_43_895 VPWR VGND sg13g2_decap_8
XFILLER_15_586 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0810_ VGND VPWR u_ppwm_u_ex__0787_/Y u_ppwm_u_ex__0808_/X hold293/A
+ u_ppwm_u_ex__0809_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0953_ VGND VPWR net428 u_ppwm_u_mem__0678_/Y hold72/A u_ppwm_u_mem__0952_/Y
+ sg13g2_a21oi_1
XFILLER_11_770 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0741_ fanout363/A net382 net370 VPWR VGND sg13g2_nand2_1
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_7_752 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__126_ VPWR u_ppwm_u_pwm__223_/B net299 VGND sg13g2_inv_1
XFILLER_6_262 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0672_ u_ppwm_u_ex__0671_/Y VPWR u_ppwm_u_ex__0672_/Y VGND u_ppwm_u_ex__0668_/Y
+ u_ppwm_u_ex__0670_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__0884_ net515 VPWR u_ppwm_u_mem__0884_/Y VGND net432 hold164/A sg13g2_o21ai_1
XFILLER_41_4 VPWR VGND sg13g2_fill_1
XFILLER_37_111 VPWR VGND sg13g2_decap_4
XFILLER_38_634 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__075_ u_ppwm_u_global_counter__075_/A u_ppwm_u_global_counter__085_/A
+ net666 u_ppwm_u_global_counter__082_/D VPWR VGND sg13g2_nor3_2
Xu_ppwm_u_ex__1086_ net349 u_ppwm_u_ex__1086_/C u_ppwm_u_ex__1086_/A u_ppwm_u_ex__1086_/Y
+ VPWR VGND u_ppwm_u_ex__1086_/D sg13g2_nand4_1
XFILLER_21_512 VPWR VGND sg13g2_decap_8
XFILLER_34_884 VPWR VGND sg13g2_decap_8
XFILLER_21_589 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1127__108 VPWR VGND net108 sg13g2_tiehi
Xu_ppwm_u_ex__0939_ VGND VPWR u_ppwm_u_ex__0937_/Y u_ppwm_u_ex__0950_/D u_ppwm_u_ex__0939_/Y
+ net357 sg13g2_a21oi_1
XFILLER_1_917 VPWR VGND sg13g2_decap_8
Xhold13 hold13/A VPWR VGND net211 sg13g2_dlygate4sd3_1
XFILLER_29_35 VPWR VGND sg13g2_fill_1
Xhold46 hold46/A VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold35 hold35/A VPWR VGND net233 sg13g2_dlygate4sd3_1
Xhold24 hold24/A VPWR VGND net222 sg13g2_dlygate4sd3_1
Xhold57 hold57/A VPWR VGND net255 sg13g2_dlygate4sd3_1
Xhold68 hold68/A VPWR VGND net266 sg13g2_dlygate4sd3_1
XFILLER_21_1016 VPWR VGND sg13g2_decap_8
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_29_79 VPWR VGND sg13g2_decap_4
XFILLER_29_623 VPWR VGND sg13g2_decap_8
Xhold79 hold79/A VPWR VGND net277 sg13g2_dlygate4sd3_1
XFILLER_16_317 VPWR VGND sg13g2_decap_4
XFILLER_16_339 VPWR VGND sg13g2_decap_4
XFILLER_44_659 VPWR VGND sg13g2_decap_8
XFILLER_43_158 VPWR VGND sg13g2_fill_2
XFILLER_25_862 VPWR VGND sg13g2_decap_8
XFILLER_40_810 VPWR VGND sg13g2_decap_8
XFILLER_12_545 VPWR VGND sg13g2_decap_8
XFILLER_40_887 VPWR VGND sg13g2_decap_8
XFILLER_8_527 VPWR VGND sg13g2_decap_8
XFILLER_6_28 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1111__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_4_722 VPWR VGND sg13g2_decap_8
XFILLER_4_799 VPWR VGND sg13g2_decap_8
XFILLER_0_950 VPWR VGND sg13g2_decap_8
XFILLER_48_943 VPWR VGND sg13g2_decap_8
XFILLER_47_431 VPWR VGND sg13g2_decap_8
XFILLER_19_122 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1221_ net85 VGND VPWR net613 hold243/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1152_ net58 VGND VPWR u_ppwm_u_mem__1152_/D hold80/A clknet_5_27__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_626 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1083_ VGND VPWR u_ppwm_u_mem__0730_/A net400 u_ppwm_u_mem__1218_/D
+ u_ppwm_u_mem__1082_/Y sg13g2_a21oi_1
XFILLER_34_158 VPWR VGND sg13g2_fill_2
XFILLER_16_895 VPWR VGND sg13g2_decap_8
XFILLER_31_821 VPWR VGND sg13g2_decap_8
XFILLER_43_692 VPWR VGND sg13g2_decap_8
XFILLER_31_898 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0724_ u_ppwm_u_ex__0724_/Y net462 hold313/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0936_ net502 VPWR u_ppwm_u_mem__0936_/Y VGND net426 net320 sg13g2_o21ai_1
Xu_ppwm_u_ex__0655_ u_ppwm_u_ex__0655_/Y hold295/A net442 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0867_ VGND VPWR net437 u_ppwm_u_mem__0721_/Y hold45/A u_ppwm_u_mem__0866_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1189__59 VPWR VGND net59 sg13g2_tiehi
Xu_ppwm_u_mem__0798_ hold36/A hold38/A net478 u_ppwm_u_mem__0799_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0586_ VPWR u_ppwm_u_ex__0693_/B hold240/A VGND sg13g2_inv_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_4
XFILLER_39_976 VPWR VGND sg13g2_decap_8
XFILLER_41_607 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1069_ u_ppwm_u_ex__1069_/Y net356 net630 net363 hold296/A VPWR VGND
+ sg13g2_a22oi_1
Xu_ppwm_u_global_counter__058_ VPWR u_ppwm_u_global_counter__058_/Y net620 VGND sg13g2_inv_1
XFILLER_26_659 VPWR VGND sg13g2_decap_8
XFILLER_22_843 VPWR VGND sg13g2_decap_8
XFILLER_34_681 VPWR VGND sg13g2_decap_8
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_0_213 VPWR VGND sg13g2_decap_8
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_16_114 VPWR VGND sg13g2_fill_2
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_44_456 VPWR VGND sg13g2_decap_8
XFILLER_13_843 VPWR VGND sg13g2_decap_8
XFILLER_9_803 VPWR VGND sg13g2_decap_8
XFILLER_40_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0721_ VPWR u_ppwm_u_mem__0721_/Y net242 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0652_ VPWR u_ppwm_u_mem__0652_/Y net234 VGND sg13g2_inv_1
XFILLER_4_596 VPWR VGND sg13g2_decap_8
XFILLER_48_740 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1204_ net89 VGND VPWR net313 hold130/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_935 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1135_ net92 VGND VPWR net330 hold90/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_629 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_7 VPWR VGND uio_oe[4] sg13g2_tielo
Xu_ppwm_u_mem__1066_ net494 VPWR u_ppwm_u_mem__1066_/Y VGND net401 net528 sg13g2_o21ai_1
XFILLER_16_692 VPWR VGND sg13g2_decap_8
XFILLER_15_191 VPWR VGND sg13g2_fill_2
XFILLER_31_695 VPWR VGND sg13g2_decap_8
XFILLER_8_891 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0707_ u_ppwm_u_ex__0707_/Y net439 u_ppwm_u_ex__1049_/A hold277/A u_ppwm_u_ex__0735_/A
+ VPWR VGND sg13g2_a22oi_1
Xhold302 hold302/A VPWR VGND net670 sg13g2_dlygate4sd3_1
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0919_ VGND VPWR net438 u_ppwm_u_mem__0695_/Y hold187/A u_ppwm_u_mem__0918_/Y
+ sg13g2_a21oi_1
Xhold324 hold324/A VPWR VGND net692 sg13g2_dlygate4sd3_1
Xhold313 hold313/A VPWR VGND net681 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0638_ VGND VPWR u_ppwm_u_ex__0623_/B u_ppwm_u_ex__0634_/Y u_ppwm_u_ex__0640_/A
+ u_ppwm_u_ex__0637_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0569_ u_ppwm_u_ex__1025_/A net449 VPWR VGND sg13g2_inv_2
XFILLER_26_412 VPWR VGND sg13g2_fill_2
XFILLER_27_935 VPWR VGND sg13g2_decap_8
XFILLER_39_773 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_26_47 VPWR VGND sg13g2_decap_4
XFILLER_14_629 VPWR VGND sg13g2_decap_8
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_22_640 VPWR VGND sg13g2_decap_8
XFILLER_6_828 VPWR VGND sg13g2_decap_8
XFILLER_10_857 VPWR VGND sg13g2_decap_8
XFILLER_5_338 VPWR VGND sg13g2_decap_4
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_18_946 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
XFILLER_41_971 VPWR VGND sg13g2_decap_8
XFILLER_9_600 VPWR VGND sg13g2_decap_8
XFILLER_13_640 VPWR VGND sg13g2_decap_8
XFILLER_40_481 VPWR VGND sg13g2_decap_8
XFILLER_8_121 VPWR VGND sg13g2_decap_8
XFILLER_9_677 VPWR VGND sg13g2_decap_8
XFILLER_5_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0704_ VPWR u_ppwm_u_mem__0704_/Y net347 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0635_ VPWR u_ppwm_u_mem__0635_/Y net257 VGND sg13g2_inv_1
XFILLER_36_732 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1182__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_24_927 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1118_ net126 VGND VPWR u_ppwm_u_mem__1118_/D hold82/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1049_ VGND VPWR net417 u_ppwm_u_mem__0630_/Y hold142/A u_ppwm_u_mem__1048_/Y
+ sg13g2_a21oi_1
Xhold110 hold110/A VPWR VGND net308 sg13g2_dlygate4sd3_1
Xhold121 hold121/A VPWR VGND net319 sg13g2_dlygate4sd3_1
Xhold132 hold132/A VPWR VGND net330 sg13g2_dlygate4sd3_1
Xhold143 hold143/A VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold154 hold154/A VPWR VGND net522 sg13g2_dlygate4sd3_1
Xhold165 hold165/A VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold176 hold176/A VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold198 hold198/A VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold187 hold187/A VPWR VGND net555 sg13g2_dlygate4sd3_1
XFILLER_39_570 VPWR VGND sg13g2_decap_8
XFILLER_2_1024 VPWR VGND sg13g2_decap_4
XFILLER_27_732 VPWR VGND sg13g2_decap_8
XFILLER_42_768 VPWR VGND sg13g2_decap_8
XFILLER_23_993 VPWR VGND sg13g2_decap_8
XFILLER_10_654 VPWR VGND sg13g2_decap_8
XFILLER_6_625 VPWR VGND sg13g2_decap_8
XFILLER_2_842 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_37_507 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_18_743 VPWR VGND sg13g2_decap_8
XFILLER_45_562 VPWR VGND sg13g2_decap_8
XFILLER_17_275 VPWR VGND sg13g2_fill_1
XFILLER_17_286 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0972_ u_ppwm_u_ex__0971_/Y VPWR u_ppwm_u_ex__0972_/Y VGND u_ppwm_u_ex__0812_/X
+ u_ppwm_u_ex__0842_/B sg13g2_o21ai_1
XFILLER_33_757 VPWR VGND sg13g2_decap_8
XFILLER_14_993 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0618_ VPWR u_ppwm_u_mem__0618_/Y net290 VGND sg13g2_inv_1
Xheichips25_ppwm_17 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_23_201 VPWR VGND sg13g2_decap_8
XFILLER_24_724 VPWR VGND sg13g2_decap_8
XFILLER_23_15 VPWR VGND sg13g2_decap_8
XFILLER_20_963 VPWR VGND sg13g2_decap_8
XFILLER_3_639 VPWR VGND sg13g2_decap_8
XFILLER_2_127 VPWR VGND sg13g2_decap_8
Xfanout420 net421 net420 VPWR VGND sg13g2_buf_8
Xfanout431 net438 net431 VPWR VGND sg13g2_buf_2
XFILLER_48_56 VPWR VGND sg13g2_decap_8
Xfanout442 net201 net442 VPWR VGND sg13g2_buf_8
Xfanout464 net465 net464 VPWR VGND sg13g2_buf_8
Xfanout453 net678 net453 VPWR VGND sg13g2_buf_8
XFILLER_24_1025 VPWR VGND sg13g2_decap_4
Xfanout475 net689 net475 VPWR VGND sg13g2_buf_8
XFILLER_47_816 VPWR VGND sg13g2_decap_8
Xfanout497 net499 net497 VPWR VGND sg13g2_buf_1
Xfanout486 net487 net486 VPWR VGND sg13g2_buf_8
XFILLER_14_212 VPWR VGND sg13g2_fill_1
XFILLER_42_565 VPWR VGND sg13g2_decap_8
XFILLER_15_768 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__211_ VGND VPWR hold284/A u_ppwm_u_pwm__213_/B u_ppwm_u_pwm__216_/B
+ u_ppwm_u_pwm__210_/Y sg13g2_a21oi_1
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_23_790 VPWR VGND sg13g2_decap_8
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_7_934 VPWR VGND sg13g2_decap_8
XFILLER_6_422 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__142_ VGND VPWR u_ppwm_u_pwm__135_/Y net390 hold2/A u_ppwm_u_pwm__141_/Y
+ sg13g2_a21oi_1
XFILLER_6_499 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_4
XFILLER_38_816 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__091_ hold267/A u_ppwm_u_global_counter__095_/C net392 net634
+ u_ppwm_u_global_counter__055_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_46_860 VPWR VGND sg13g2_decap_8
XFILLER_18_540 VPWR VGND sg13g2_decap_8
XFILLER_33_554 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0955_ net372 net455 u_ppwm_u_ex__0955_/X VPWR VGND sg13g2_xor2_1
XFILLER_14_790 VPWR VGND sg13g2_decap_8
XFILLER_20_215 VPWR VGND sg13g2_fill_2
XFILLER_20_237 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0886_ u_ppwm_u_ex__0884_/Y u_ppwm_u_ex__0881_/Y u_ppwm_u_ex__0885_/Y
+ u_ppwm_u_ex__0898_/B VPWR VGND sg13g2_a21o_1
XFILLER_9_293 VPWR VGND sg13g2_decap_8
XFILLER_9_271 VPWR VGND sg13g2_decap_4
XFILLER_29_805 VPWR VGND sg13g2_decap_8
XFILLER_18_15 VPWR VGND sg13g2_fill_2
XFILLER_43_307 VPWR VGND sg13g2_decap_8
XFILLER_37_871 VPWR VGND sg13g2_decap_8
XFILLER_24_521 VPWR VGND sg13g2_decap_8
XFILLER_34_14 VPWR VGND sg13g2_fill_2
XFILLER_12_727 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1108__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_8_709 VPWR VGND sg13g2_decap_8
XFILLER_24_598 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_5_6__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_20_760 VPWR VGND sg13g2_decap_8
XFILLER_4_904 VPWR VGND sg13g2_decap_8
XFILLER_3_436 VPWR VGND sg13g2_decap_8
XFILLER_47_613 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_4
XFILLER_19_337 VPWR VGND sg13g2_fill_1
XFILLER_35_808 VPWR VGND sg13g2_decap_8
XFILLER_43_874 VPWR VGND sg13g2_decap_8
XFILLER_15_565 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0952_ net510 VPWR u_ppwm_u_mem__0952_/Y VGND net427 hold174/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0740_ VGND VPWR u_ppwm_u_ex__0734_/X u_ppwm_u_ex__0735_/Y u_ppwm_u_ex__0740_/Y
+ u_ppwm_u_ex__0739_/Y sg13g2_a21oi_1
XFILLER_7_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__125_ VPWR u_ppwm_u_pwm__183_/A net593 VGND sg13g2_inv_1
XFILLER_6_230 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0671_ u_ppwm_u_ex__0671_/Y net440 u_ppwm_u_ex__0850_/A u_ppwm_u_ex__1020_/B2
+ u_ppwm_u_ex__0576_/Y VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__0883_ VGND VPWR net433 u_ppwm_u_mem__0713_/Y u_ppwm_u_mem__1118_/D
+ u_ppwm_u_mem__0882_/Y sg13g2_a21oi_1
XFILLER_6_285 VPWR VGND sg13g2_fill_2
XFILLER_38_613 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__074_ hold297/A net604 net653 hold298/A VPWR VGND net630
+ sg13g2_nand4_1
Xu_ppwm_u_ex__1085_ u_ppwm_u_ex__1084_/Y u_ppwm_u_ex__1083_/Y net361 u_ppwm_u_ex__1086_/D
+ VPWR VGND sg13g2_a21o_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_25_329 VPWR VGND sg13g2_decap_8
XFILLER_34_863 VPWR VGND sg13g2_decap_8
XFILLER_21_568 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0938_ u_ppwm_u_ex__0950_/D net664 net371 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__0869_ hold296/A net385 u_ppwm_u_ex__0869_/Y VPWR VGND sg13g2_nor2_1
Xhold14 hold14/A VPWR VGND net212 sg13g2_dlygate4sd3_1
XFILLER_0_439 VPWR VGND sg13g2_decap_8
Xhold36 hold36/A VPWR VGND net234 sg13g2_dlygate4sd3_1
Xhold47 hold47/A VPWR VGND net245 sg13g2_dlygate4sd3_1
Xu_ppwm_u_pwm__246__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_29_602 VPWR VGND sg13g2_decap_8
Xhold25 hold25/A VPWR VGND net223 sg13g2_dlygate4sd3_1
Xhold69 hold69/A VPWR VGND net267 sg13g2_dlygate4sd3_1
Xhold58 hold58/A VPWR VGND net256 sg13g2_dlygate4sd3_1
XFILLER_29_679 VPWR VGND sg13g2_decap_8
XFILLER_44_638 VPWR VGND sg13g2_decap_8
XFILLER_25_841 VPWR VGND sg13g2_decap_8
XFILLER_12_524 VPWR VGND sg13g2_decap_8
XFILLER_40_866 VPWR VGND sg13g2_decap_8
XFILLER_8_506 VPWR VGND sg13g2_decap_8
XFILLER_4_701 VPWR VGND sg13g2_decap_8
XFILLER_4_778 VPWR VGND sg13g2_decap_8
XFILLER_10_93 VPWR VGND sg13g2_fill_1
XFILLER_48_922 VPWR VGND sg13g2_decap_8
XFILLER_47_410 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1220_ net117 VGND VPWR u_ppwm_u_mem__1220_/D hold323/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1151_ net60 VGND VPWR net279 hold112/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_605 VPWR VGND sg13g2_decap_8
XFILLER_48_999 VPWR VGND sg13g2_decap_8
XFILLER_47_487 VPWR VGND sg13g2_decap_8
XFILLER_19_167 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1082_ net488 VPWR u_ppwm_u_mem__1082_/Y VGND net535 net401 sg13g2_o21ai_1
XFILLER_43_671 VPWR VGND sg13g2_decap_8
XFILLER_16_874 VPWR VGND sg13g2_decap_8
XFILLER_31_800 VPWR VGND sg13g2_decap_8
XFILLER_15_373 VPWR VGND sg13g2_decap_4
XFILLER_31_877 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0723_ VPWR VGND u_ppwm_u_ex__0721_/Y u_ppwm_u_ex__0722_/Y u_ppwm_u_ex__0720_/Y
+ net452 u_ppwm_u_ex__0723_/Y u_ppwm_u_ex__0850_/A sg13g2_a221oi_1
Xu_ppwm_u_mem__0935_ VGND VPWR net426 u_ppwm_u_mem__0687_/Y hold123/A u_ppwm_u_mem__0934_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0654_ u_ppwm_u_ex__0653_/Y VPWR u_ppwm_u_ex__0654_/Y VGND hold303/A
+ u_ppwm_u_ex__0761_/B sg13g2_o21ai_1
Xu_ppwm_u_mem__0866_ net516 VPWR u_ppwm_u_mem__0866_/Y VGND net437 hold143/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0585_ VPWR u_ppwm_u_ex__0585_/Y hold252/A VGND sg13g2_inv_1
Xu_ppwm_u_mem__0797_ VGND VPWR net395 u_ppwm_u_mem__0796_/X u_ppwm_u_mem__0797_/Y
+ net394 sg13g2_a21oi_1
XFILLER_39_955 VPWR VGND sg13g2_decap_8
XFILLER_38_410 VPWR VGND sg13g2_fill_2
XFILLER_26_638 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__057_ VPWR u_ppwm_u_global_counter__057_/Y net645 VGND sg13g2_inv_1
Xu_ppwm_u_ex__1068_ u_ppwm_u_ex__1068_/Y net645 net355 VPWR VGND sg13g2_nand2_1
XFILLER_34_660 VPWR VGND sg13g2_decap_8
XFILLER_40_129 VPWR VGND sg13g2_fill_2
XFILLER_22_822 VPWR VGND sg13g2_decap_8
XFILLER_22_899 VPWR VGND sg13g2_decap_8
XFILLER_31_48 VPWR VGND sg13g2_fill_2
XFILLER_0_236 VPWR VGND sg13g2_fill_1
XFILLER_0_269 VPWR VGND sg13g2_fill_2
XFILLER_48_229 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_decap_8
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_44_435 VPWR VGND sg13g2_decap_8
XFILLER_17_649 VPWR VGND sg13g2_decap_8
XFILLER_32_619 VPWR VGND sg13g2_decap_8
XFILLER_13_822 VPWR VGND sg13g2_decap_8
XFILLER_40_663 VPWR VGND sg13g2_decap_8
XFILLER_9_859 VPWR VGND sg13g2_decap_8
XFILLER_13_899 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0720_ VPWR u_ppwm_u_mem__0720_/Y net277 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0651_ VPWR u_ppwm_u_mem__0651_/Y net244 VGND sg13g2_inv_1
XFILLER_4_575 VPWR VGND sg13g2_decap_8
XFILLER_11_6 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1203_ net97 VGND VPWR u_ppwm_u_mem__1203_/D hold15/A clknet_5_25__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_48_796 VPWR VGND sg13g2_decap_8
XFILLER_36_914 VPWR VGND sg13g2_decap_8
XFILLER_47_284 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1134_ net94 VGND VPWR net289 hold202/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_435 VPWR VGND sg13g2_decap_4
XFILLER_23_608 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_8 VPWR VGND uio_oe[5] sg13g2_tielo
Xu_ppwm_u_mem__1065_ VGND VPWR net403 u_ppwm_u_mem__0622_/Y u_ppwm_u_mem__1209_/D
+ u_ppwm_u_mem__1064_/Y sg13g2_a21oi_1
XFILLER_16_671 VPWR VGND sg13g2_decap_8
XFILLER_22_118 VPWR VGND sg13g2_fill_1
XFILLER_31_674 VPWR VGND sg13g2_decap_8
XFILLER_8_870 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0706_ u_ppwm_u_ex__0705_/Y VPWR u_ppwm_u_ex__0706_/Y VGND u_ppwm_u_ex__0651_/A
+ hold254/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0918_ net512 VPWR u_ppwm_u_mem__0918_/Y VGND net426 net329 sg13g2_o21ai_1
Xhold303 hold303/A VPWR VGND net671 sg13g2_dlygate4sd3_1
Xhold314 hold314/A VPWR VGND net682 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0637_ net447 VPWR u_ppwm_u_ex__0637_/Y VGND u_ppwm_u_ex__0635_/Y u_ppwm_u_ex__0636_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0849_ hold169/A hold167/A net476 u_ppwm_u_mem__0850_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0568_ hold299/A u_ppwm_u_ex__0651_/A VPWR VGND sg13g2_inv_4
XFILLER_39_752 VPWR VGND sg13g2_decap_8
XFILLER_27_914 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__109_ net508 VGND VPWR net600 hold231/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_38_284 VPWR VGND sg13g2_decap_8
XFILLER_38_295 VPWR VGND sg13g2_fill_1
XFILLER_14_608 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_4
XFILLER_10_836 VPWR VGND sg13g2_decap_8
XFILLER_22_696 VPWR VGND sg13g2_decap_8
XFILLER_6_807 VPWR VGND sg13g2_decap_8
XFILLER_27_1012 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_fill_2
XFILLER_18_925 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1116__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_45_744 VPWR VGND sg13g2_decap_8
XFILLER_17_435 VPWR VGND sg13g2_fill_1
XFILLER_33_939 VPWR VGND sg13g2_decap_8
XFILLER_41_950 VPWR VGND sg13g2_decap_8
XFILLER_40_460 VPWR VGND sg13g2_decap_8
XFILLER_8_111 VPWR VGND sg13g2_fill_1
XFILLER_12_151 VPWR VGND sg13g2_fill_2
XFILLER_13_696 VPWR VGND sg13g2_decap_8
XFILLER_9_656 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0703_ VPWR u_ppwm_u_mem__0703_/Y net282 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0634_ VPWR u_ppwm_u_mem__0634_/Y net205 VGND sg13g2_inv_1
XFILLER_36_711 VPWR VGND sg13g2_decap_8
XFILLER_48_593 VPWR VGND sg13g2_decap_8
XFILLER_24_906 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1117_ net128 VGND VPWR net281 hold195/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_788 VPWR VGND sg13g2_decap_8
XFILLER_35_276 VPWR VGND sg13g2_decap_8
XFILLER_35_298 VPWR VGND sg13g2_decap_4
XFILLER_23_449 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1048_ net501 VPWR u_ppwm_u_mem__1048_/Y VGND net418 hold152/A sg13g2_o21ai_1
XFILLER_32_983 VPWR VGND sg13g2_decap_8
Xhold100 hold100/A VPWR VGND net298 sg13g2_dlygate4sd3_1
Xhold133 hold133/A VPWR VGND net331 sg13g2_dlygate4sd3_1
Xhold144 hold144/A VPWR VGND net342 sg13g2_dlygate4sd3_1
Xhold122 hold122/A VPWR VGND net320 sg13g2_dlygate4sd3_1
Xhold111 hold111/A VPWR VGND net309 sg13g2_dlygate4sd3_1
Xhold166 hold166/A VPWR VGND net534 sg13g2_dlygate4sd3_1
Xhold177 hold177/A VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold155 hold155/A VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold199 hold199/A VPWR VGND net567 sg13g2_dlygate4sd3_1
Xhold188 hold188/A VPWR VGND net556 sg13g2_dlygate4sd3_1
XFILLER_2_1003 VPWR VGND sg13g2_decap_8
XFILLER_27_711 VPWR VGND sg13g2_decap_8
XFILLER_27_788 VPWR VGND sg13g2_decap_8
XFILLER_42_747 VPWR VGND sg13g2_decap_8
XFILLER_41_213 VPWR VGND sg13g2_decap_4
XFILLER_23_972 VPWR VGND sg13g2_decap_8
XFILLER_10_633 VPWR VGND sg13g2_decap_8
XFILLER_22_493 VPWR VGND sg13g2_decap_8
XFILLER_6_604 VPWR VGND sg13g2_decap_8
XFILLER_2_821 VPWR VGND sg13g2_decap_8
XFILLER_2_898 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_40_1020 VPWR VGND sg13g2_decap_8
XFILLER_18_722 VPWR VGND sg13g2_decap_8
XFILLER_45_541 VPWR VGND sg13g2_decap_8
XFILLER_17_243 VPWR VGND sg13g2_fill_2
XFILLER_18_799 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_fill_2
XFILLER_33_736 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0971_ u_ppwm_u_ex__0971_/Y u_ppwm_u_ex__0892_/Y net368 u_ppwm_u_ex__0871_/X
+ u_ppwm_u_ex__0838_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_14_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0617_ VPWR u_ppwm_u_mem__0617_/Y net222 VGND sg13g2_inv_1
Xheichips25_ppwm_18 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_48_390 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__240__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_24_703 VPWR VGND sg13g2_decap_8
XFILLER_36_585 VPWR VGND sg13g2_decap_8
XFILLER_12_909 VPWR VGND sg13g2_decap_8
XFILLER_23_224 VPWR VGND sg13g2_fill_2
XFILLER_23_268 VPWR VGND sg13g2_decap_8
XFILLER_23_279 VPWR VGND sg13g2_fill_1
XFILLER_20_942 VPWR VGND sg13g2_decap_8
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_32_780 VPWR VGND sg13g2_decap_8
XFILLER_3_618 VPWR VGND sg13g2_decap_8
XFILLER_2_106 VPWR VGND sg13g2_decap_8
Xfanout421 net422 net421 VPWR VGND sg13g2_buf_2
Xfanout432 net435 net432 VPWR VGND sg13g2_buf_8
Xfanout410 net411 net410 VPWR VGND sg13g2_buf_2
XFILLER_48_35 VPWR VGND sg13g2_decap_8
Xfanout454 net675 net454 VPWR VGND sg13g2_buf_8
Xfanout443 net655 net443 VPWR VGND sg13g2_buf_8
Xfanout465 net687 net465 VPWR VGND sg13g2_buf_8
XFILLER_24_1004 VPWR VGND sg13g2_decap_8
Xfanout498 net499 net498 VPWR VGND sg13g2_buf_8
XFILLER_19_519 VPWR VGND sg13g2_decap_8
Xfanout487 fanout487/A net487 VPWR VGND sg13g2_buf_8
Xfanout476 net479 net476 VPWR VGND sg13g2_buf_8
XFILLER_46_349 VPWR VGND sg13g2_decap_8
XFILLER_27_585 VPWR VGND sg13g2_decap_8
XFILLER_42_544 VPWR VGND sg13g2_decap_8
XFILLER_14_235 VPWR VGND sg13g2_fill_2
XFILLER_15_747 VPWR VGND sg13g2_decap_8
XFILLER_30_728 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__210_ hold62/A hold233/A u_ppwm_u_pwm__210_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_7_913 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__141_ net492 VPWR u_ppwm_u_pwm__141_/Y VGND net466 net390 sg13g2_o21ai_1
XFILLER_6_478 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_fill_2
XFILLER_2_695 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__090_ u_ppwm_u_global_counter__095_/C net633 u_ppwm_u_ex__1020_/B2
+ net398 VPWR VGND sg13g2_and3_2
Xu_ppwm_u_mem__1137__88 VPWR VGND net88 sg13g2_tiehi
Xu_ppwm_u_mem__1152__58 VPWR VGND net58 sg13g2_tiehi
XFILLER_18_596 VPWR VGND sg13g2_decap_8
XFILLER_33_533 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0954_ u_ppwm_u_ex__0954_/A u_ppwm_u_ex__1049_/B u_ppwm_u_ex__0954_/Y
+ VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0885_ u_ppwm_u_ex__0780_/X VPWR u_ppwm_u_ex__0885_/Y VGND u_ppwm_u_ex__0881_/Y
+ u_ppwm_u_ex__0884_/Y sg13g2_o21ai_1
XFILLER_47_1026 VPWR VGND sg13g2_fill_2
XFILLER_37_850 VPWR VGND sg13g2_decap_8
XFILLER_24_500 VPWR VGND sg13g2_decap_8
XFILLER_36_382 VPWR VGND sg13g2_decap_4
XFILLER_12_706 VPWR VGND sg13g2_decap_8
XFILLER_24_577 VPWR VGND sg13g2_decap_8
Xclkload3 clknet_5_14__leaf_clk clkload3/X VPWR VGND sg13g2_buf_1
XFILLER_3_415 VPWR VGND sg13g2_decap_8
XFILLER_47_669 VPWR VGND sg13g2_decap_8
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_43_853 VPWR VGND sg13g2_decap_8
XFILLER_15_544 VPWR VGND sg13g2_decap_8
XFILLER_42_341 VPWR VGND sg13g2_fill_1
XFILLER_30_525 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0951_ VGND VPWR net427 u_ppwm_u_mem__0679_/Y u_ppwm_u_mem__1152_/D
+ u_ppwm_u_mem__0950_/Y sg13g2_a21oi_1
XFILLER_24_70 VPWR VGND sg13g2_decap_4
XFILLER_10_271 VPWR VGND sg13g2_decap_4
XFILLER_10_260 VPWR VGND sg13g2_fill_1
XFILLER_7_710 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0882_ net515 VPWR u_ppwm_u_mem__0882_/Y VGND net433 net280 sg13g2_o21ai_1
XFILLER_10_293 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0670_ VGND VPWR u_ppwm_u_ex__0666_/Y u_ppwm_u_ex__0669_/Y u_ppwm_u_ex__0670_/Y
+ u_ppwm_u_ex__0665_/Y sg13g2_a21oi_1
XFILLER_7_787 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__230__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_3_982 VPWR VGND sg13g2_decap_8
XFILLER_2_492 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1084_ u_ppwm_u_ex__1084_/Y net356 net442 net363 hold304/A VPWR VGND
+ sg13g2_a22oi_1
Xu_ppwm_u_global_counter__073_ u_ppwm_u_global_counter__073_/B net604 hold237/A VPWR
+ VGND sg13g2_xor2_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_38_669 VPWR VGND sg13g2_decap_8
XFILLER_19_883 VPWR VGND sg13g2_decap_8
XFILLER_34_842 VPWR VGND sg13g2_decap_8
XFILLER_21_547 VPWR VGND sg13g2_decap_8
XFILLER_33_385 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0937_ VGND VPWR u_ppwm_u_ex__0924_/A u_ppwm_u_ex__0924_/B u_ppwm_u_ex__0937_/Y
+ u_ppwm_u_ex__0950_/B sg13g2_a21oi_1
XFILLER_14_1014 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1113__50 VPWR VGND net50 sg13g2_tiehi
Xu_ppwm_u_ex__0868_ u_ppwm_u_ex__0867_/Y VPWR u_ppwm_u_ex__0868_/Y VGND u_ppwm_u_ex__0820_/B
+ u_ppwm_u_ex__0839_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__0799_ VPWR u_ppwm_u_ex__0799_/Y u_ppwm_u_ex__0799_/A VGND sg13g2_inv_1
XFILLER_0_418 VPWR VGND sg13g2_decap_8
Xhold26 hold26/A VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold37 hold37/A VPWR VGND net235 sg13g2_dlygate4sd3_1
XFILLER_29_59 VPWR VGND sg13g2_fill_2
Xhold15 hold15/A VPWR VGND net213 sg13g2_dlygate4sd3_1
Xhold48 hold48/A VPWR VGND net246 sg13g2_dlygate4sd3_1
Xhold59 hold59/A VPWR VGND net257 sg13g2_dlygate4sd3_1
XFILLER_29_658 VPWR VGND sg13g2_decap_8
XFILLER_45_25 VPWR VGND sg13g2_fill_2
XFILLER_44_617 VPWR VGND sg13g2_decap_8
XFILLER_25_820 VPWR VGND sg13g2_decap_8
XFILLER_43_138 VPWR VGND sg13g2_fill_2
XFILLER_36_190 VPWR VGND sg13g2_fill_1
XFILLER_40_845 VPWR VGND sg13g2_decap_8
XFILLER_25_897 VPWR VGND sg13g2_decap_8
XFILLER_4_757 VPWR VGND sg13g2_decap_8
XFILLER_3_234 VPWR VGND sg13g2_decap_4
XFILLER_48_901 VPWR VGND sg13g2_decap_8
XFILLER_0_985 VPWR VGND sg13g2_decap_8
XFILLER_48_978 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1150_ net62 VGND VPWR net311 hold154/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_466 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1081_ VGND VPWR u_ppwm_u_mem__0613_/Y net400 u_ppwm_u_mem__1217_/D
+ u_ppwm_u_mem__1080_/Y sg13g2_a21oi_1
XFILLER_16_853 VPWR VGND sg13g2_decap_8
XFILLER_28_680 VPWR VGND sg13g2_decap_8
XFILLER_43_650 VPWR VGND sg13g2_decap_8
XFILLER_15_341 VPWR VGND sg13g2_decap_8
XFILLER_37_1025 VPWR VGND sg13g2_decap_4
XFILLER_42_171 VPWR VGND sg13g2_fill_2
XFILLER_31_856 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1126__110 VPWR VGND net110 sg13g2_tiehi
Xu_ppwm_u_ex__0722_ net465 net453 u_ppwm_u_ex__0722_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0934_ net510 VPWR u_ppwm_u_mem__0934_/Y VGND net426 hold139/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0653_ u_ppwm_u_ex__0653_/Y u_ppwm_u_ex__0735_/A hold262/A VPWR VGND
+ sg13g2_nand2_1
XFILLER_7_584 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0865_ VGND VPWR net435 u_ppwm_u_mem__0722_/Y hold144/A u_ppwm_u_mem__0864_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__1110__31 VPWR VGND net31 sg13g2_tiehi
Xu_ppwm_u_mem__0796_ hold32/A hold152/A net480 u_ppwm_u_mem__0796_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0584_ VPWR u_ppwm_u_ex__0605_/A net399 VGND sg13g2_inv_1
XFILLER_39_934 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__125_ net505 VGND VPWR net586 hold217/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_617 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__056_ VPWR u_ppwm_u_global_counter__056_/Y net622 VGND sg13g2_inv_1
Xu_ppwm_u_ex__1067_ u_ppwm_u_ex__1066_/Y VPWR u_ppwm_u_ex__1067_/Y VGND u_ppwm_u_ex__1064_/Y
+ u_ppwm_u_ex__1075_/C sg13g2_o21ai_1
XFILLER_19_680 VPWR VGND sg13g2_decap_8
XFILLER_22_801 VPWR VGND sg13g2_decap_8
XFILLER_22_878 VPWR VGND sg13g2_decap_8
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_48_208 VPWR VGND sg13g2_decap_8
XFILLER_0_248 VPWR VGND sg13g2_decap_8
XFILLER_29_444 VPWR VGND sg13g2_fill_1
XFILLER_45_926 VPWR VGND sg13g2_decap_8
XFILLER_44_414 VPWR VGND sg13g2_decap_8
XFILLER_17_628 VPWR VGND sg13g2_decap_8
XFILLER_16_116 VPWR VGND sg13g2_fill_1
XFILLER_16_127 VPWR VGND sg13g2_fill_1
XFILLER_13_801 VPWR VGND sg13g2_decap_8
XFILLER_25_694 VPWR VGND sg13g2_decap_8
XFILLER_40_642 VPWR VGND sg13g2_decap_8
XFILLER_13_878 VPWR VGND sg13g2_decap_8
XFILLER_9_838 VPWR VGND sg13g2_decap_8
XFILLER_8_348 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0650_ VPWR u_ppwm_u_mem__0650_/Y net540 VGND sg13g2_inv_1
XFILLER_4_554 VPWR VGND sg13g2_decap_8
XFILLER_0_782 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1202_ net105 VGND VPWR net214 hold141/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1156__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_48_775 VPWR VGND sg13g2_decap_8
XFILLER_47_263 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1133_ net96 VGND VPWR u_ppwm_u_mem__1133_/D hold138/A clknet_5_31__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_16_650 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_9 VPWR VGND uio_oe[6] sg13g2_tielo
Xu_ppwm_u_mem__1064_ net494 VPWR u_ppwm_u_mem__1064_/Y VGND net403 net318 sg13g2_o21ai_1
XFILLER_44_981 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
XFILLER_31_653 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0705_ u_ppwm_u_ex__0705_/Y net448 net439 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0917_ VGND VPWR net425 u_ppwm_u_mem__0696_/Y hold132/A u_ppwm_u_mem__0916_/Y
+ sg13g2_a21oi_1
Xhold304 hold304/A VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold315 hold315/A VPWR VGND net683 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0636_ u_ppwm_u_ex__0636_/Y u_ppwm_u_ex__0636_/A u_ppwm_u_ex__0636_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0848_ hold59/A hold130/A net476 u_ppwm_u_mem__0848_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0779_ hold57/A hold51/A net478 u_ppwm_u_mem__0780_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0567_ u_ppwm_u_ex__1049_/A net448 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__1185__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_39_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1119_ net26 VGND VPWR u_ppwm_u_ex__1119_/D hold314/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_global_counter__108_ net508 VGND VPWR net656 hold291/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_26_414 VPWR VGND sg13g2_fill_1
XFILLER_42_929 VPWR VGND sg13g2_decap_8
XFILLER_41_439 VPWR VGND sg13g2_decap_8
XFILLER_13_108 VPWR VGND sg13g2_fill_2
XFILLER_21_130 VPWR VGND sg13g2_decap_8
XFILLER_10_815 VPWR VGND sg13g2_decap_8
XFILLER_22_675 VPWR VGND sg13g2_decap_8
XFILLER_5_307 VPWR VGND sg13g2_fill_1
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_18_904 VPWR VGND sg13g2_decap_8
XFILLER_45_723 VPWR VGND sg13g2_decap_8
XFILLER_33_918 VPWR VGND sg13g2_decap_8
XFILLER_26_981 VPWR VGND sg13g2_decap_8
XFILLER_25_491 VPWR VGND sg13g2_decap_8
XFILLER_9_635 VPWR VGND sg13g2_decap_8
XFILLER_13_675 VPWR VGND sg13g2_decap_8
XFILLER_34_1017 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0702_ VPWR u_ppwm_u_mem__0702_/Y net524 VGND sg13g2_inv_1
XFILLER_5_885 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0633_ VPWR u_ppwm_u_mem__0633_/Y net526 VGND sg13g2_inv_1
XFILLER_48_572 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1116_ net130 VGND VPWR u_ppwm_u_mem__1116_/D hold193/A clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_767 VPWR VGND sg13g2_decap_8
XFILLER_17_992 VPWR VGND sg13g2_decap_8
XFILLER_35_288 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1047_ VGND VPWR net418 u_ppwm_u_mem__0631_/Y hold153/A u_ppwm_u_mem__1046_/Y
+ sg13g2_a21oi_1
XFILLER_32_962 VPWR VGND sg13g2_decap_8
XFILLER_31_472 VPWR VGND sg13g2_fill_2
Xhold101 hold101/A VPWR VGND net299 sg13g2_dlygate4sd3_1
Xhold112 hold112/A VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold123 hold123/A VPWR VGND net321 sg13g2_dlygate4sd3_1
Xhold134 hold134/A VPWR VGND net332 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0619_ u_ppwm_u_ex__0636_/B u_ppwm_u_ex__0619_/B u_ppwm_u_ex__0619_/C
+ u_ppwm_u_ex__0619_/X VPWR VGND sg13g2_or3_1
Xhold167 hold167/A VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold145 hold145/A VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold156 hold156/A VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold189 hold189/A VPWR VGND net557 sg13g2_dlygate4sd3_1
Xhold178 hold178/A VPWR VGND net546 sg13g2_dlygate4sd3_1
XFILLER_27_767 VPWR VGND sg13g2_decap_8
XFILLER_42_726 VPWR VGND sg13g2_decap_8
XFILLER_15_929 VPWR VGND sg13g2_decap_8
XFILLER_23_951 VPWR VGND sg13g2_decap_8
XFILLER_10_612 VPWR VGND sg13g2_decap_8
XFILLER_22_472 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_fill_2
XFILLER_10_689 VPWR VGND sg13g2_decap_8
XFILLER_2_800 VPWR VGND sg13g2_decap_8
XFILLER_2_877 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1149__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_18_701 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1192__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_45_520 VPWR VGND sg13g2_decap_8
XFILLER_18_778 VPWR VGND sg13g2_decap_8
XFILLER_45_597 VPWR VGND sg13g2_decap_8
XFILLER_33_715 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0970_ u_ppwm_u_ex__0969_/Y VPWR u_ppwm_u_ex__0970_/Y VGND u_ppwm_u_ex__0967_/Y
+ u_ppwm_u_ex__0968_/Y sg13g2_o21ai_1
XFILLER_14_951 VPWR VGND sg13g2_decap_8
XFILLER_17_299 VPWR VGND sg13g2_decap_8
XFILLER_43_80 VPWR VGND sg13g2_decap_8
XFILLER_13_472 VPWR VGND sg13g2_fill_1
XFILLER_5_682 VPWR VGND sg13g2_decap_8
XFILLER_4_192 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0616_ VPWR u_ppwm_u_mem__0616_/Y net527 VGND sg13g2_inv_1
Xheichips25_ppwm_19 VPWR VGND uo_out[1] sg13g2_tielo
XFILLER_36_564 VPWR VGND sg13g2_decap_8
XFILLER_24_759 VPWR VGND sg13g2_decap_8
XFILLER_20_921 VPWR VGND sg13g2_decap_8
XFILLER_20_998 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout400 net402 net400 VPWR VGND sg13g2_buf_8
Xfanout422 fanout438/A net422 VPWR VGND sg13g2_buf_8
Xfanout411 net422 net411 VPWR VGND sg13g2_buf_8
Xfanout455 net672 net455 VPWR VGND sg13g2_buf_8
Xfanout444 net665 net444 VPWR VGND sg13g2_buf_8
Xfanout466 fanout466/A net466 VPWR VGND sg13g2_buf_8
Xfanout433 net435 net433 VPWR VGND sg13g2_buf_8
XFILLER_48_69 VPWR VGND sg13g2_fill_2
Xfanout488 net489 net488 VPWR VGND sg13g2_buf_8
Xfanout477 net479 net477 VPWR VGND sg13g2_buf_8
Xfanout499 net500 net499 VPWR VGND sg13g2_buf_8
XFILLER_46_328 VPWR VGND sg13g2_decap_8
XFILLER_15_726 VPWR VGND sg13g2_decap_8
XFILLER_27_564 VPWR VGND sg13g2_decap_8
XFILLER_42_523 VPWR VGND sg13g2_decap_8
XFILLER_11_910 VPWR VGND sg13g2_decap_8
XFILLER_30_707 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__140_ u_ppwm_u_pwm__140_/B u_ppwm_u_pwm__140_/C u_ppwm_u_pwm__140_/A
+ fanout391/A VPWR VGND sg13g2_nand3_1
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_13_72 VPWR VGND sg13g2_fill_1
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_2_674 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_144 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_895 VPWR VGND sg13g2_decap_8
XFILLER_18_575 VPWR VGND sg13g2_decap_8
XFILLER_45_394 VPWR VGND sg13g2_decap_8
XFILLER_21_729 VPWR VGND sg13g2_decap_8
XFILLER_33_589 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0953_ u_ppwm_u_ex__0952_/X VPWR u_ppwm_u_ex__0953_/Y VGND u_ppwm_u_ex__0884_/Y
+ u_ppwm_u_ex__0950_/X sg13g2_o21ai_1
Xu_ppwm_u_ex__0884_ VGND VPWR u_ppwm_u_ex__0883_/Y u_ppwm_u_ex__0884_/Y u_ppwm_u_ex__0882_/Y
+ u_ppwm_u_ex__0849_/Y sg13g2_a21oi_2
XFILLER_47_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1215__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_18_17 VPWR VGND sg13g2_fill_1
XFILLER_24_556 VPWR VGND sg13g2_decap_8
XFILLER_34_38 VPWR VGND sg13g2_fill_1
Xclkload4 clknet_5_16__leaf_clk clkload4/X VPWR VGND sg13g2_buf_1
XFILLER_20_795 VPWR VGND sg13g2_decap_8
XFILLER_4_939 VPWR VGND sg13g2_decap_8
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1221__85 VPWR VGND net85 sg13g2_tiehi
XFILLER_47_648 VPWR VGND sg13g2_decap_8
XFILLER_28_862 VPWR VGND sg13g2_decap_8
XFILLER_34_309 VPWR VGND sg13g2_fill_2
XFILLER_43_832 VPWR VGND sg13g2_decap_8
XFILLER_42_320 VPWR VGND sg13g2_fill_2
XFILLER_15_523 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0950_ net510 VPWR u_ppwm_u_mem__0950_/Y VGND net427 net278 sg13g2_o21ai_1
XFILLER_11_784 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0881_ VGND VPWR net433 u_ppwm_u_mem__0714_/Y hold83/A u_ppwm_u_mem__0880_/Y
+ sg13g2_a21oi_1
XFILLER_7_766 VPWR VGND sg13g2_decap_8
XFILLER_6_232 VPWR VGND sg13g2_fill_1
XFILLER_3_961 VPWR VGND sg13g2_decap_8
XFILLER_2_471 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__072_ u_ppwm_u_global_counter__073_/B net628 hold261/A VPWR
+ VGND sg13g2_nor2_1
Xu_ppwm_u_ex__1083_ u_ppwm_u_ex__1083_/Y hold252/A net355 VPWR VGND sg13g2_nand2_1
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_125 VPWR VGND sg13g2_decap_8
XFILLER_38_648 VPWR VGND sg13g2_decap_8
XFILLER_19_862 VPWR VGND sg13g2_decap_8
XFILLER_46_692 VPWR VGND sg13g2_decap_8
XFILLER_18_372 VPWR VGND sg13g2_decap_8
XFILLER_18_383 VPWR VGND sg13g2_fill_1
XFILLER_34_821 VPWR VGND sg13g2_decap_8
XFILLER_21_526 VPWR VGND sg13g2_decap_8
XFILLER_34_898 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1166__149 VPWR VGND net149 sg13g2_tiehi
Xu_ppwm_u_ex__0936_ u_ppwm_u_ex__0936_/A u_ppwm_u_ex__0936_/B u_ppwm_u_ex__1111_/D
+ VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0867_ u_ppwm_u_ex__0867_/A u_ppwm_u_ex__0867_/B u_ppwm_u_ex__0867_/Y
+ VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0798_ net461 net449 net386 u_ppwm_u_ex__0799_/A VPWR VGND sg13g2_mux2_1
Xhold27 hold27/A VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold38 hold38/A VPWR VGND net236 sg13g2_dlygate4sd3_1
Xhold16 hold16/A VPWR VGND net214 sg13g2_dlygate4sd3_1
Xhold49 hold49/A VPWR VGND net247 sg13g2_dlygate4sd3_1
XFILLER_29_637 VPWR VGND sg13g2_decap_8
XFILLER_24_320 VPWR VGND sg13g2_decap_8
XFILLER_25_876 VPWR VGND sg13g2_decap_8
XFILLER_40_824 VPWR VGND sg13g2_decap_8
XFILLER_12_559 VPWR VGND sg13g2_decap_8
XFILLER_20_592 VPWR VGND sg13g2_decap_8
XFILLER_3_202 VPWR VGND sg13g2_fill_2
XFILLER_4_736 VPWR VGND sg13g2_decap_8
XFILLER_0_964 VPWR VGND sg13g2_decap_8
XFILLER_19_103 VPWR VGND sg13g2_decap_4
XFILLER_48_957 VPWR VGND sg13g2_decap_8
XFILLER_47_445 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1080_ net494 VPWR u_ppwm_u_mem__1080_/Y VGND net400 net295 sg13g2_o21ai_1
XFILLER_16_832 VPWR VGND sg13g2_decap_8
XFILLER_37_1004 VPWR VGND sg13g2_decap_8
XFILLER_31_835 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0721_ net466 hold292/A u_ppwm_u_ex__0721_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0933_ VGND VPWR net426 u_ppwm_u_mem__0688_/Y hold140/A u_ppwm_u_mem__0932_/Y
+ sg13g2_a21oi_1
XFILLER_11_581 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0652_ VPWR VGND u_ppwm_u_ex__0650_/Y u_ppwm_u_ex__0651_/Y u_ppwm_u_ex__0642_/Y
+ net448 u_ppwm_u_ex__0652_/Y u_ppwm_u_ex__0761_/B sg13g2_a221oi_1
XFILLER_7_563 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0864_ net516 VPWR u_ppwm_u_mem__0864_/Y VGND net433 hold209/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0583_ VPWR fanout370/A net377 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0795_ u_ppwm_u_mem__0795_/Y net471 u_ppwm_u_mem__0795_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_39_913 VPWR VGND sg13g2_decap_8
XFILLER_38_412 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_global_counter__124_ net505 VGND VPWR net621 hold252/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__055_ VPWR u_ppwm_u_global_counter__055_/Y u_ppwm_u_ex__1020_/B2
+ VGND sg13g2_inv_1
Xu_ppwm_u_ex__1066_ VGND VPWR u_ppwm_u_ex__1064_/Y u_ppwm_u_ex__1075_/C u_ppwm_u_ex__1066_/Y
+ net358 sg13g2_a21oi_1
XFILLER_15_18 VPWR VGND sg13g2_decap_4
XFILLER_33_150 VPWR VGND sg13g2_fill_2
XFILLER_34_695 VPWR VGND sg13g2_decap_8
XFILLER_22_857 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0919_ net456 net371 u_ppwm_u_ex__0950_/B VPWR VGND sg13g2_and2_1
XFILLER_0_227 VPWR VGND sg13g2_decap_8
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_17_607 VPWR VGND sg13g2_decap_8
XFILLER_40_621 VPWR VGND sg13g2_decap_8
XFILLER_25_673 VPWR VGND sg13g2_decap_8
XFILLER_9_817 VPWR VGND sg13g2_decap_8
XFILLER_12_345 VPWR VGND sg13g2_fill_1
XFILLER_13_857 VPWR VGND sg13g2_decap_8
XFILLER_8_327 VPWR VGND sg13g2_fill_2
XFILLER_40_698 VPWR VGND sg13g2_decap_8
XFILLER_21_890 VPWR VGND sg13g2_decap_8
XFILLER_4_533 VPWR VGND sg13g2_decap_8
XFILLER_0_761 VPWR VGND sg13g2_decap_8
XFILLER_48_754 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1201_ net113 VGND VPWR net340 hold152/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_242 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1132_ net98 VGND VPWR u_ppwm_u_mem__1132_/D hold64/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_949 VPWR VGND sg13g2_decap_8
XFILLER_44_960 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1063_ VGND VPWR net403 u_ppwm_u_mem__0623_/Y u_ppwm_u_mem__1208_/D
+ u_ppwm_u_mem__1062_/Y sg13g2_a21oi_1
XFILLER_31_632 VPWR VGND sg13g2_decap_8
XFILLER_7_30 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0704_ u_ppwm_u_ex__0704_/Y u_ppwm_u_ex__0693_/Y u_ppwm_u_ex__0703_/Y
+ hold254/A u_ppwm_u_ex__0651_/A VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__0916_ net512 VPWR u_ppwm_u_mem__0916_/Y VGND net425 net288 sg13g2_o21ai_1
Xu_ppwm_u_ex__0635_ VGND VPWR net469 u_ppwm_u_ex__0622_/B u_ppwm_u_ex__0635_/Y net468
+ sg13g2_a21oi_1
Xhold316 hold316/A VPWR VGND net684 sg13g2_dlygate4sd3_1
Xhold305 hold305/A VPWR VGND net673 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0847_ VGND VPWR net395 u_ppwm_u_mem__0846_/X u_ppwm_u_mem__0847_/Y
+ net470 sg13g2_a21oi_1
Xu_ppwm_u_ex__0566_ hold294/A u_ppwm_u_ex__0735_/A VPWR VGND sg13g2_inv_4
Xu_ppwm_u_mem__0778_ VGND VPWR net395 u_ppwm_u_mem__0777_/X u_ppwm_u_mem__0778_/Y
+ net394 sg13g2_a21oi_1
XFILLER_30_0 VPWR VGND sg13g2_decap_4
XFILLER_39_710 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__243__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_39_787 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__107_ net508 VGND VPWR u_ppwm_u_global_counter__107_/D hold297/A
+ clknet_5_20__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1118_ net30 VGND VPWR u_ppwm_u_ex__1118_/D hold313/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_27_949 VPWR VGND sg13g2_decap_8
XFILLER_42_908 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1049_ u_ppwm_u_ex__1049_/A u_ppwm_u_ex__1049_/B u_ppwm_u_ex__1049_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_41_418 VPWR VGND sg13g2_decap_8
XFILLER_22_654 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_45_702 VPWR VGND sg13g2_decap_8
XFILLER_17_404 VPWR VGND sg13g2_fill_1
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_44_256 VPWR VGND sg13g2_fill_2
XFILLER_26_960 VPWR VGND sg13g2_decap_8
XFILLER_41_985 VPWR VGND sg13g2_decap_8
XFILLER_9_614 VPWR VGND sg13g2_decap_8
XFILLER_13_654 VPWR VGND sg13g2_decap_8
XFILLER_40_495 VPWR VGND sg13g2_decap_8
XFILLER_12_175 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0701_ VPWR u_ppwm_u_mem__0701_/Y net581 VGND sg13g2_inv_1
XFILLER_5_864 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0632_ VPWR u_ppwm_u_mem__0632_/Y net582 VGND sg13g2_inv_1
XFILLER_48_551 VPWR VGND sg13g2_decap_8
XFILLER_36_746 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1115_ net132 VGND VPWR net562 hold100/A clknet_5_23__leaf_clk sg13g2_dfrbpq_2
XFILLER_17_971 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1046_ net503 VPWR u_ppwm_u_mem__1046_/Y VGND net418 hold214/A sg13g2_o21ai_1
XFILLER_32_941 VPWR VGND sg13g2_decap_8
Xhold124 hold124/A VPWR VGND net322 sg13g2_dlygate4sd3_1
Xhold102 hold102/A VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold135 hold135/A VPWR VGND net333 sg13g2_dlygate4sd3_1
Xhold113 hold113/A VPWR VGND net311 sg13g2_dlygate4sd3_1
Xhold168 hold168/A VPWR VGND net536 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0618_ u_ppwm_u_ex__0619_/C net483 net385 u_ppwm_u_ex__0618_/C VPWR VGND
+ sg13g2_and3_1
Xhold157 hold157/A VPWR VGND net525 sg13g2_dlygate4sd3_1
Xhold146 hold146/A VPWR VGND net344 sg13g2_dlygate4sd3_1
Xhold179 hold179/A VPWR VGND net547 sg13g2_dlygate4sd3_1
XFILLER_26_212 VPWR VGND sg13g2_decap_4
XFILLER_39_584 VPWR VGND sg13g2_decap_8
XFILLER_42_705 VPWR VGND sg13g2_decap_8
XFILLER_15_908 VPWR VGND sg13g2_decap_8
XFILLER_27_746 VPWR VGND sg13g2_decap_8
XFILLER_26_289 VPWR VGND sg13g2_decap_8
XFILLER_23_930 VPWR VGND sg13g2_decap_8
XFILLER_22_451 VPWR VGND sg13g2_decap_8
XFILLER_10_668 VPWR VGND sg13g2_decap_8
XFILLER_6_639 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_decap_8
XFILLER_2_856 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_18_757 VPWR VGND sg13g2_decap_8
XFILLER_45_576 VPWR VGND sg13g2_decap_8
XFILLER_14_930 VPWR VGND sg13g2_decap_8
XFILLER_41_782 VPWR VGND sg13g2_decap_8
XFILLER_40_292 VPWR VGND sg13g2_decap_8
XFILLER_9_488 VPWR VGND sg13g2_decap_8
XFILLER_5_661 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0615_ VPWR u_ppwm_u_mem__0615_/Y net295 VGND sg13g2_inv_1
XFILLER_49_893 VPWR VGND sg13g2_decap_8
XFILLER_36_510 VPWR VGND sg13g2_fill_2
XFILLER_36_543 VPWR VGND sg13g2_decap_8
XFILLER_24_738 VPWR VGND sg13g2_decap_8
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_20_900 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1029_ VGND VPWR net405 u_ppwm_u_mem__0640_/Y hold171/A u_ppwm_u_mem__1028_/Y
+ sg13g2_a21oi_1
XFILLER_20_977 VPWR VGND sg13g2_decap_8
Xfanout412 net416 net412 VPWR VGND sg13g2_buf_8
Xfanout423 net424 net423 VPWR VGND sg13g2_buf_8
Xfanout401 net402 net401 VPWR VGND sg13g2_buf_1
Xfanout456 net677 net456 VPWR VGND sg13g2_buf_8
Xfanout445 net653 net445 VPWR VGND sg13g2_buf_8
Xfanout434 net435 net434 VPWR VGND sg13g2_buf_8
XFILLER_46_307 VPWR VGND sg13g2_decap_8
Xfanout489 net493 net489 VPWR VGND sg13g2_buf_8
Xfanout467 hold315/A net467 VPWR VGND sg13g2_buf_8
Xfanout478 net479 net478 VPWR VGND sg13g2_buf_8
XFILLER_27_510 VPWR VGND sg13g2_fill_1
XFILLER_27_543 VPWR VGND sg13g2_decap_8
XFILLER_42_502 VPWR VGND sg13g2_decap_8
XFILLER_15_705 VPWR VGND sg13g2_decap_8
XFILLER_14_237 VPWR VGND sg13g2_fill_1
XFILLER_42_579 VPWR VGND sg13g2_decap_8
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_2_653 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_1_185 VPWR VGND sg13g2_fill_2
XFILLER_46_874 VPWR VGND sg13g2_decap_8
XFILLER_18_554 VPWR VGND sg13g2_decap_8
XFILLER_45_373 VPWR VGND sg13g2_decap_8
XFILLER_21_708 VPWR VGND sg13g2_decap_8
XFILLER_33_568 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0952_ u_ppwm_u_ex__0952_/A u_ppwm_u_ex__0952_/B u_ppwm_u_ex__0952_/X
+ VPWR VGND sg13g2_and2_1
XFILLER_13_292 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0883_ VGND VPWR u_ppwm_u_ex__0576_/Y u_ppwm_u_ex__0850_/A u_ppwm_u_ex__0883_/Y
+ u_ppwm_u_ex__1049_/B sg13g2_a21oi_1
Xu_ppwm_u_mem__1199__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_47_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__199_ u_ppwm_u_pwm__199_/Y hold17/A hold181/A VPWR VGND sg13g2_nand2b_1
XFILLER_29_819 VPWR VGND sg13g2_decap_8
XFILLER_49_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1136__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_37_885 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1151__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_24_535 VPWR VGND sg13g2_decap_8
XFILLER_11_218 VPWR VGND sg13g2_fill_1
Xclkload5 clknet_5_18__leaf_clk clkload5/X VPWR VGND sg13g2_buf_1
XFILLER_20_774 VPWR VGND sg13g2_decap_8
XFILLER_4_918 VPWR VGND sg13g2_decap_8
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_627 VPWR VGND sg13g2_decap_8
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_43_811 VPWR VGND sg13g2_decap_8
XFILLER_15_502 VPWR VGND sg13g2_decap_8
XFILLER_27_362 VPWR VGND sg13g2_fill_1
XFILLER_43_888 VPWR VGND sg13g2_decap_8
XFILLER_15_579 VPWR VGND sg13g2_decap_8
XFILLER_24_94 VPWR VGND sg13g2_fill_2
XFILLER_6_200 VPWR VGND sg13g2_fill_1
XFILLER_11_763 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0880_ net516 VPWR u_ppwm_u_mem__0880_/Y VGND net433 hold195/A sg13g2_o21ai_1
XFILLER_7_745 VPWR VGND sg13g2_decap_8
XFILLER_6_266 VPWR VGND sg13g2_fill_1
XFILLER_6_255 VPWR VGND sg13g2_decap_8
XFILLER_40_93 VPWR VGND sg13g2_fill_1
XFILLER_3_940 VPWR VGND sg13g2_decap_8
XFILLER_2_450 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_37_115 VPWR VGND sg13g2_fill_1
XFILLER_38_627 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__071_ VGND VPWR net590 u_ppwm_u_global_counter__068_/B hold260/A
+ net627 sg13g2_a21oi_1
Xu_ppwm_u_ex__1082_ u_ppwm_u_ex__1081_/Y VPWR u_ppwm_u_ex__1086_/C VGND u_ppwm_u_ex__1078_/Y
+ u_ppwm_u_ex__1080_/Y sg13g2_o21ai_1
XFILLER_19_841 VPWR VGND sg13g2_decap_8
XFILLER_46_671 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_34_800 VPWR VGND sg13g2_decap_8
XFILLER_34_877 VPWR VGND sg13g2_decap_8
XFILLER_21_505 VPWR VGND sg13g2_decap_8
XFILLER_33_365 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0935_ net491 VPWR u_ppwm_u_ex__0936_/B VGND net456 net352 sg13g2_o21ai_1
Xu_ppwm_u_ex__0866_ net375 net378 u_ppwm_u_ex__0866_/C u_ppwm_u_ex__0867_/B VPWR VGND
+ sg13g2_nor3_1
Xu_ppwm_u_ex__0797_ u_ppwm_u_ex__0843_/A u_ppwm_u_ex__0796_/Y u_ppwm_u_ex__0797_/Y
+ VPWR VGND sg13g2_nor2b_2
Xu_ppwm_u_mem__1203__97 VPWR VGND net97 sg13g2_tiehi
Xhold17 hold17/A VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold28 hold28/A VPWR VGND net226 sg13g2_dlygate4sd3_1
Xhold39 hold39/A VPWR VGND net237 sg13g2_dlygate4sd3_1
XFILLER_21_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_616 VPWR VGND sg13g2_decap_8
XFILLER_37_682 VPWR VGND sg13g2_decap_8
XFILLER_40_803 VPWR VGND sg13g2_decap_8
XFILLER_25_855 VPWR VGND sg13g2_decap_8
XFILLER_12_538 VPWR VGND sg13g2_decap_8
XFILLER_20_571 VPWR VGND sg13g2_decap_8
XFILLER_4_715 VPWR VGND sg13g2_decap_8
XFILLER_0_943 VPWR VGND sg13g2_decap_8
XFILLER_48_936 VPWR VGND sg13g2_decap_8
XFILLER_47_424 VPWR VGND sg13g2_decap_8
XFILLER_35_619 VPWR VGND sg13g2_decap_8
XFILLER_16_811 VPWR VGND sg13g2_decap_8
XFILLER_34_118 VPWR VGND sg13g2_decap_4
XFILLER_43_685 VPWR VGND sg13g2_decap_8
XFILLER_42_173 VPWR VGND sg13g2_fill_1
XFILLER_16_888 VPWR VGND sg13g2_decap_8
XFILLER_31_814 VPWR VGND sg13g2_decap_8
XFILLER_30_335 VPWR VGND sg13g2_fill_2
XFILLER_11_560 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0720_ u_ppwm_u_ex__0720_/Y net465 net453 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0932_ net512 VPWR u_ppwm_u_mem__0932_/Y VGND net425 net220 sg13g2_o21ai_1
XFILLER_7_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0651_ u_ppwm_u_ex__0651_/A hold259/A u_ppwm_u_ex__0651_/Y VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_mem__0863_ VGND VPWR net434 u_ppwm_u_mem__0723_/Y hold210/A u_ppwm_u_mem__0862_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0582_ net373 u_ppwm_u_ex__1049_/B VPWR VGND sg13g2_inv_4
Xu_ppwm_u_mem__0794_ hold55/A hold24/A net476 u_ppwm_u_mem__0795_/B VPWR VGND sg13g2_mux2_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
XFILLER_39_969 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__123_ net505 VGND VPWR net646 hold277/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1065_ u_ppwm_u_ex__1075_/C net662 net373 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_global_counter__054_ VPWR u_ppwm_u_global_counter__054_/Y u_ppwm_u_ex__0998_/B2
+ VGND sg13g2_inv_1
XFILLER_47_991 VPWR VGND sg13g2_decap_8
XFILLER_22_836 VPWR VGND sg13g2_decap_8
XFILLER_34_674 VPWR VGND sg13g2_decap_8
XFILLER_21_335 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0918_ net456 net371 u_ppwm_u_ex__0950_/A VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0849_ u_ppwm_u_ex__0825_/Y VPWR u_ppwm_u_ex__0849_/Y VGND u_ppwm_u_ex__0782_/Y
+ u_ppwm_u_ex__0826_/Y sg13g2_o21ai_1
XFILLER_1_707 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1188__63 VPWR VGND net63 sg13g2_tiehi
XFILLER_0_206 VPWR VGND sg13g2_decap_8
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
XFILLER_38_991 VPWR VGND sg13g2_decap_8
XFILLER_44_449 VPWR VGND sg13g2_decap_8
XFILLER_25_652 VPWR VGND sg13g2_decap_8
XFILLER_40_600 VPWR VGND sg13g2_decap_8
XFILLER_13_836 VPWR VGND sg13g2_decap_8
XFILLER_40_677 VPWR VGND sg13g2_decap_8
XFILLER_8_317 VPWR VGND sg13g2_fill_2
XFILLER_4_512 VPWR VGND sg13g2_decap_8
XFILLER_4_589 VPWR VGND sg13g2_decap_8
XFILLER_0_740 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1195__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_48_733 VPWR VGND sg13g2_decap_8
XFILLER_47_221 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1200_ net121 VGND VPWR net521 hold214/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_928 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1131_ net100 VGND VPWR net263 hold213/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_298 VPWR VGND sg13g2_decap_8
XFILLER_29_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1062_ net494 VPWR u_ppwm_u_mem__1062_/Y VGND net403 net253 sg13g2_o21ai_1
XFILLER_16_685 VPWR VGND sg13g2_decap_8
XFILLER_31_611 VPWR VGND sg13g2_decap_8
XFILLER_43_482 VPWR VGND sg13g2_decap_8
XFILLER_31_688 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0703_ u_ppwm_u_ex__0702_/Y VPWR u_ppwm_u_ex__0703_/Y VGND u_ppwm_u_ex__0697_/Y
+ u_ppwm_u_ex__0699_/Y sg13g2_o21ai_1
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
XFILLER_30_198 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0915_ VGND VPWR net425 u_ppwm_u_mem__0697_/Y hold91/A u_ppwm_u_mem__0914_/Y
+ sg13g2_a21oi_1
XFILLER_8_884 VPWR VGND sg13g2_decap_8
XFILLER_7_383 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0634_ u_ppwm_u_ex__0634_/Y u_ppwm_u_ex__0634_/A u_ppwm_u_ex__0634_/B
+ VPWR VGND sg13g2_xnor2_1
Xhold317 hold317/A VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold306 hold306/A VPWR VGND net674 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0846_ hold224/A hold211/A net479 u_ppwm_u_mem__0846_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0565_ u_ppwm_u_ex__0711_/A hold295/A VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0777_ hold200/A hold214/A net480 u_ppwm_u_mem__0777_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_global_counter__106_ net508 VGND VPWR u_ppwm_u_global_counter__106_/D hold285/A
+ clknet_5_21__leaf_clk sg13g2_dfrbpq_2
XFILLER_27_928 VPWR VGND sg13g2_decap_8
XFILLER_39_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1117_ net34 VGND VPWR u_ppwm_u_ex__1117_/D hold300/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_26_18 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1048_ u_ppwm_u_ex__1048_/A u_ppwm_u_ex__1046_/Y u_ppwm_u_ex__1120_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_22_633 VPWR VGND sg13g2_decap_8
XFILLER_21_154 VPWR VGND sg13g2_decap_4
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_508 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1155__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_18_939 VPWR VGND sg13g2_decap_8
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_17_449 VPWR VGND sg13g2_decap_4
XFILLER_25_460 VPWR VGND sg13g2_decap_4
XFILLER_13_633 VPWR VGND sg13g2_decap_8
XFILLER_41_964 VPWR VGND sg13g2_decap_8
XFILLER_40_441 VPWR VGND sg13g2_fill_2
XFILLER_40_474 VPWR VGND sg13g2_decap_8
XFILLER_32_61 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0700_ VPWR u_ppwm_u_mem__0700_/Y net262 VGND sg13g2_inv_1
XFILLER_5_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0631_ VPWR u_ppwm_u_mem__0631_/Y net520 VGND sg13g2_inv_1
XFILLER_48_530 VPWR VGND sg13g2_decap_8
XFILLER_36_725 VPWR VGND sg13g2_decap_8
XFILLER_17_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1114_ net134 VGND VPWR u_ppwm_u_mem__1114_/D hold86/A clknet_5_22__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1045_ VGND VPWR net407 u_ppwm_u_mem__0632_/Y u_ppwm_u_mem__1199_/D
+ u_ppwm_u_mem__1044_/Y sg13g2_a21oi_1
XFILLER_32_920 VPWR VGND sg13g2_decap_8
XFILLER_31_474 VPWR VGND sg13g2_fill_1
XFILLER_32_997 VPWR VGND sg13g2_decap_8
XFILLER_8_681 VPWR VGND sg13g2_decap_8
Xhold114 hold114/A VPWR VGND net312 sg13g2_dlygate4sd3_1
Xhold103 hold103/A VPWR VGND net301 sg13g2_dlygate4sd3_1
Xhold125 hold125/A VPWR VGND net323 sg13g2_dlygate4sd3_1
Xhold136 hold136/A VPWR VGND net334 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0617_ VGND VPWR net483 net385 u_ppwm_u_ex__0619_/B u_ppwm_u_ex__0618_/C
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0829_ net471 VPWR u_ppwm_u_mem__0829_/Y VGND hold160/A net476 sg13g2_o21ai_1
Xhold158 hold158/A VPWR VGND net526 sg13g2_dlygate4sd3_1
Xhold147 hold147/A VPWR VGND net345 sg13g2_dlygate4sd3_1
Xhold169 hold169/A VPWR VGND net537 sg13g2_dlygate4sd3_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_725 VPWR VGND sg13g2_decap_8
XFILLER_39_563 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1181__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_35_780 VPWR VGND sg13g2_decap_8
XFILLER_22_430 VPWR VGND sg13g2_decap_8
XFILLER_23_986 VPWR VGND sg13g2_decap_8
XFILLER_6_618 VPWR VGND sg13g2_decap_8
XFILLER_10_647 VPWR VGND sg13g2_decap_8
XFILLER_2_835 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_18_736 VPWR VGND sg13g2_decap_8
XFILLER_45_555 VPWR VGND sg13g2_decap_8
XFILLER_41_761 VPWR VGND sg13g2_decap_8
XFILLER_32_249 VPWR VGND sg13g2_fill_1
XFILLER_40_271 VPWR VGND sg13g2_decap_8
XFILLER_14_986 VPWR VGND sg13g2_decap_8
XFILLER_5_640 VPWR VGND sg13g2_decap_8
XFILLER_4_194 VPWR VGND sg13g2_fill_1
XFILLER_4_32 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0614_ VPWR u_ppwm_u_mem__0730_/A net1 VGND sg13g2_inv_1
XFILLER_4_65 VPWR VGND sg13g2_fill_1
XFILLER_49_872 VPWR VGND sg13g2_decap_8
XFILLER_36_522 VPWR VGND sg13g2_decap_8
XFILLER_24_717 VPWR VGND sg13g2_decap_8
XFILLER_36_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1028_ net495 VPWR u_ppwm_u_mem__1028_/Y VGND net405 hold203/A sg13g2_o21ai_1
XFILLER_31_271 VPWR VGND sg13g2_fill_2
XFILLER_32_794 VPWR VGND sg13g2_decap_8
XFILLER_20_956 VPWR VGND sg13g2_decap_8
Xfanout413 net416 net413 VPWR VGND sg13g2_buf_2
Xfanout402 net406 net402 VPWR VGND sg13g2_buf_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
Xfanout457 hold309/A net457 VPWR VGND sg13g2_buf_2
Xfanout446 net686 net446 VPWR VGND sg13g2_buf_8
XFILLER_24_1018 VPWR VGND sg13g2_decap_8
Xfanout424 net425 net424 VPWR VGND sg13g2_buf_8
Xfanout435 net437 net435 VPWR VGND sg13g2_buf_8
XFILLER_47_809 VPWR VGND sg13g2_decap_8
Xfanout468 net683 net468 VPWR VGND sg13g2_buf_1
Xfanout479 net487 net479 VPWR VGND sg13g2_buf_8
XFILLER_27_522 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1113__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_27_599 VPWR VGND sg13g2_decap_8
XFILLER_42_558 VPWR VGND sg13g2_decap_8
XFILLER_23_783 VPWR VGND sg13g2_decap_8
XFILLER_11_945 VPWR VGND sg13g2_decap_8
XFILLER_7_927 VPWR VGND sg13g2_decap_8
XFILLER_2_632 VPWR VGND sg13g2_decap_8
XFILLER_38_809 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_46_853 VPWR VGND sg13g2_decap_8
XFILLER_45_330 VPWR VGND sg13g2_decap_4
XFILLER_18_533 VPWR VGND sg13g2_decap_8
XFILLER_45_352 VPWR VGND sg13g2_decap_8
XFILLER_33_514 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0951_ net371 VPWR u_ppwm_u_ex__0952_/B VGND hold296/A net456 sg13g2_o21ai_1
XFILLER_33_547 VPWR VGND sg13g2_decap_8
XFILLER_14_783 VPWR VGND sg13g2_decap_8
XFILLER_13_271 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0882_ u_ppwm_u_ex__0882_/A u_ppwm_u_ex__0882_/B u_ppwm_u_ex__0882_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_286 VPWR VGND sg13g2_decap_8
XFILLER_6_982 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__198_ u_ppwm_u_pwm__198_/Y hold1/A hold279/A VPWR VGND sg13g2_nand2b_1
XFILLER_37_864 VPWR VGND sg13g2_decap_8
XFILLER_24_514 VPWR VGND sg13g2_decap_8
XFILLER_32_591 VPWR VGND sg13g2_decap_8
Xclkload6 clknet_5_20__leaf_clk clkload6/X VPWR VGND sg13g2_buf_1
XFILLER_20_753 VPWR VGND sg13g2_decap_8
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1206__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_3_429 VPWR VGND sg13g2_decap_8
XFILLER_47_606 VPWR VGND sg13g2_decap_8
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_fill_2
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_43_867 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_fill_1
XFILLER_15_558 VPWR VGND sg13g2_decap_8
XFILLER_24_40 VPWR VGND sg13g2_fill_2
XFILLER_11_742 VPWR VGND sg13g2_decap_8
XFILLER_23_580 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_7_724 VPWR VGND sg13g2_decap_8
XFILLER_3_996 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_4
XFILLER_49_92 VPWR VGND sg13g2_fill_1
XFILLER_38_606 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1081_ VGND VPWR u_ppwm_u_ex__1078_/Y u_ppwm_u_ex__1080_/Y u_ppwm_u_ex__1081_/Y
+ net357 sg13g2_a21oi_1
Xu_ppwm_u_global_counter__070_ u_ppwm_u_global_counter__070_/A u_ppwm_u_global_counter__085_/A
+ u_ppwm_u_global_counter__073_/B VPWR VGND sg13g2_nor2_1
XFILLER_19_820 VPWR VGND sg13g2_decap_8
XFILLER_37_138 VPWR VGND sg13g2_decap_4
XFILLER_46_650 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_19_897 VPWR VGND sg13g2_decap_8
XFILLER_34_856 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0934_ VGND VPWR u_ppwm_u_ex__0780_/X u_ppwm_u_ex__0924_/X u_ppwm_u_ex__0936_/A
+ u_ppwm_u_ex__0933_/Y sg13g2_a21oi_1
XFILLER_14_580 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0865_ u_ppwm_u_ex__0864_/Y VPWR u_ppwm_u_ex__0877_/B VGND u_ppwm_u_ex__0882_/B
+ u_ppwm_u_ex__0863_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__0796_ net382 u_ppwm_u_ex__1049_/B u_ppwm_u_ex__0796_/Y VPWR VGND sg13g2_nor2_1
Xhold29 hold29/A VPWR VGND net227 sg13g2_dlygate4sd3_1
Xhold18 hold18/A VPWR VGND net216 sg13g2_dlygate4sd3_1
XFILLER_37_661 VPWR VGND sg13g2_decap_8
XFILLER_25_834 VPWR VGND sg13g2_decap_8
XFILLER_12_517 VPWR VGND sg13g2_decap_8
XFILLER_40_859 VPWR VGND sg13g2_decap_8
XFILLER_20_550 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_fill_1
XFILLER_0_922 VPWR VGND sg13g2_decap_8
XFILLER_48_915 VPWR VGND sg13g2_decap_8
XFILLER_47_403 VPWR VGND sg13g2_decap_8
XFILLER_0_999 VPWR VGND sg13g2_decap_8
XFILLER_19_127 VPWR VGND sg13g2_fill_2
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_16_867 VPWR VGND sg13g2_decap_8
XFILLER_27_193 VPWR VGND sg13g2_fill_2
XFILLER_43_664 VPWR VGND sg13g2_decap_8
XFILLER_15_366 VPWR VGND sg13g2_decap_8
XFILLER_15_377 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1165__151 VPWR VGND net151 sg13g2_tiehi
Xu_ppwm_u_mem__0931_ VGND VPWR net425 u_ppwm_u_mem__0689_/Y hold23/A u_ppwm_u_mem__0930_/Y
+ sg13g2_a21oi_1
XFILLER_7_521 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0650_ u_ppwm_u_ex__0649_/Y VPWR u_ppwm_u_ex__0650_/Y VGND u_ppwm_u_ex__0646_/Y
+ u_ppwm_u_ex__0648_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__0862_ net514 VPWR u_ppwm_u_mem__0862_/Y VGND net434 u_ppwm_u_mem__1108_/Q
+ sg13g2_o21ai_1
XFILLER_7_598 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0581_ u_ppwm_u_ex__0979_/A net386 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0793_ u_ppwm_u_mem__0792_/X u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0783_/Y
+ fanout388/A VPWR VGND sg13g2_a21o_2
XFILLER_3_793 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_39_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__122_ net505 VGND VPWR u_ppwm_u_global_counter__122_/D hold286/A
+ clknet_5_17__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1064_ VGND VPWR u_ppwm_u_ex__1051_/A u_ppwm_u_ex__1055_/X u_ppwm_u_ex__1064_/Y
+ u_ppwm_u_ex__1049_/Y sg13g2_a21oi_1
Xu_ppwm_u_global_counter__053_ VPWR u_ppwm_u_global_counter__066_/A net599 VGND sg13g2_inv_1
XFILLER_47_970 VPWR VGND sg13g2_decap_8
XFILLER_18_160 VPWR VGND sg13g2_fill_2
XFILLER_19_694 VPWR VGND sg13g2_decap_8
XFILLER_34_653 VPWR VGND sg13g2_decap_8
XFILLER_22_815 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0917_ u_ppwm_u_ex__0917_/A u_ppwm_u_ex__0915_/Y hold302/A VPWR VGND
+ sg13g2_nor2b_1
Xu_ppwm_u_ex__0848_ VPWR VGND u_ppwm_u_ex__0797_/Y u_ppwm_u_ex__0843_/Y u_ppwm_u_ex__0847_/A
+ u_ppwm_u_ex__0790_/Y u_ppwm_u_ex__1012_/A u_ppwm_u_ex__0801_/X sg13g2_a221oi_1
Xu_ppwm_u_ex__0779_ net388 u_ppwm/instr\[1\] u_ppwm_u_ex__0819_/C VPWR VGND sg13g2_nor2b_2
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
XFILLER_44_428 VPWR VGND sg13g2_decap_8
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_25_631 VPWR VGND sg13g2_decap_8
XFILLER_13_815 VPWR VGND sg13g2_decap_8
XFILLER_40_656 VPWR VGND sg13g2_decap_8
XFILLER_4_568 VPWR VGND sg13g2_decap_8
XFILLER_48_712 VPWR VGND sg13g2_decap_8
XFILLER_43_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_200 VPWR VGND sg13g2_decap_8
XFILLER_0_796 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1130_ net102 VGND VPWR u_ppwm_u_mem__1130_/D hold156/A clknet_5_23__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_907 VPWR VGND sg13g2_decap_8
XFILLER_48_789 VPWR VGND sg13g2_decap_8
XFILLER_47_277 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1061_ VGND VPWR net403 u_ppwm_u_mem__0624_/Y hold56/A u_ppwm_u_mem__1060_/Y
+ sg13g2_a21oi_1
XFILLER_35_439 VPWR VGND sg13g2_fill_1
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_43_461 VPWR VGND sg13g2_decap_8
XFILLER_15_152 VPWR VGND sg13g2_decap_8
XFILLER_16_664 VPWR VGND sg13g2_decap_8
XFILLER_31_667 VPWR VGND sg13g2_decap_8
XFILLER_12_881 VPWR VGND sg13g2_decap_8
XFILLER_8_863 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0702_ VPWR VGND u_ppwm_u_ex__0700_/Y u_ppwm_u_ex__0701_/Y u_ppwm_u_ex__0696_/Y
+ u_ppwm_u_ex__1025_/A u_ppwm_u_ex__0702_/Y hold240/A sg13g2_a221oi_1
Xu_ppwm_u_mem__0914_ net512 VPWR u_ppwm_u_mem__0914_/Y VGND net426 hold202/A sg13g2_o21ai_1
XFILLER_7_76 VPWR VGND sg13g2_fill_2
Xhold307 hold307/A VPWR VGND net675 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0633_ u_ppwm_u_ex__0634_/B net468 net375 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__0845_ u_ppwm_u_mem__0845_/Y net471 u_ppwm_u_mem__0845_/B VPWR VGND
+ sg13g2_nand2_1
Xhold318 hold318/A VPWR VGND net686 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0564_ u_ppwm_u_ex__0973_/A hold289/A VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0776_ u_ppwm_u_mem__0776_/Y net471 u_ppwm_u_mem__0776_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_3_590 VPWR VGND sg13g2_decap_8
XFILLER_39_745 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__105_ u_ppwm_u_global_counter__105_/B net585 hold218/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__1116_ net38 VGND VPWR net679 hold310/A clknet_5_18__leaf_clk sg13g2_dfrbpq_2
XFILLER_27_907 VPWR VGND sg13g2_decap_8
XFILLER_38_255 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1047_ net506 VPWR u_ppwm_u_ex__1048_/A VGND net667 net351 sg13g2_o21ai_1
XFILLER_19_491 VPWR VGND sg13g2_decap_8
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_22_612 VPWR VGND sg13g2_decap_8
XFILLER_34_483 VPWR VGND sg13g2_fill_2
XFILLER_10_829 VPWR VGND sg13g2_decap_8
XFILLER_22_689 VPWR VGND sg13g2_decap_8
XFILLER_27_1005 VPWR VGND sg13g2_decap_8
XFILLER_18_918 VPWR VGND sg13g2_decap_8
XFILLER_45_737 VPWR VGND sg13g2_decap_8
XFILLER_44_258 VPWR VGND sg13g2_fill_1
XFILLER_41_943 VPWR VGND sg13g2_decap_8
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_13_612 VPWR VGND sg13g2_decap_8
XFILLER_26_995 VPWR VGND sg13g2_decap_8
XFILLER_40_453 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_9_649 VPWR VGND sg13g2_decap_8
XFILLER_12_177 VPWR VGND sg13g2_fill_1
XFILLER_13_689 VPWR VGND sg13g2_decap_8
XFILLER_32_40 VPWR VGND sg13g2_fill_1
XFILLER_5_822 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1123__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_4_310 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0630_ VPWR u_ppwm_u_mem__0630_/Y net339 VGND sg13g2_inv_1
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_4_365 VPWR VGND sg13g2_fill_2
XFILLER_0_593 VPWR VGND sg13g2_decap_8
XFILLER_48_586 VPWR VGND sg13g2_decap_8
XFILLER_36_704 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1113_ net136 VGND VPWR net285 hold192/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_247 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1044_ net495 VPWR u_ppwm_u_mem__1044_/Y VGND net405 net526 sg13g2_o21ai_1
XFILLER_35_269 VPWR VGND sg13g2_decap_8
XFILLER_44_792 VPWR VGND sg13g2_decap_8
XFILLER_32_976 VPWR VGND sg13g2_decap_8
XFILLER_8_660 VPWR VGND sg13g2_decap_8
Xhold104 hold104/A VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold115 hold115/A VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold126 hold126/A VPWR VGND net324 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0616_ net383 net473 u_ppwm_u_ex__0618_/C VPWR VGND sg13g2_xor2_1
Xu_ppwm_u_mem__0828_ hold97/A net476 u_ppwm_u_mem__0828_/Y VPWR VGND sg13g2_nor2b_1
Xhold159 hold159/A VPWR VGND net527 sg13g2_dlygate4sd3_1
Xhold137 hold137/A VPWR VGND net335 sg13g2_dlygate4sd3_1
Xhold148 hold148/A VPWR VGND net346 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0759_ hold170/A hold158/A net477 u_ppwm_u_mem__0760_/B VPWR VGND sg13g2_mux2_1
XFILLER_39_542 VPWR VGND sg13g2_decap_8
XFILLER_27_704 VPWR VGND sg13g2_decap_8
XFILLER_14_409 VPWR VGND sg13g2_fill_2
XFILLER_41_217 VPWR VGND sg13g2_fill_2
XFILLER_23_965 VPWR VGND sg13g2_decap_8
XFILLER_10_626 VPWR VGND sg13g2_decap_8
XFILLER_22_486 VPWR VGND sg13g2_decap_8
XFILLER_2_814 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_40_1013 VPWR VGND sg13g2_decap_8
XFILLER_18_715 VPWR VGND sg13g2_decap_8
XFILLER_45_534 VPWR VGND sg13g2_decap_8
XFILLER_17_236 VPWR VGND sg13g2_decap_8
XFILLER_17_258 VPWR VGND sg13g2_fill_2
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_33_729 VPWR VGND sg13g2_decap_8
XFILLER_26_792 VPWR VGND sg13g2_decap_8
XFILLER_41_740 VPWR VGND sg13g2_decap_8
XFILLER_14_965 VPWR VGND sg13g2_decap_8
XFILLER_13_486 VPWR VGND sg13g2_fill_1
XFILLER_9_457 VPWR VGND sg13g2_fill_2
XFILLER_5_696 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0613_ VPWR u_ppwm_u_mem__0613_/Y net535 VGND sg13g2_inv_1
XFILLER_49_851 VPWR VGND sg13g2_decap_8
XFILLER_0_390 VPWR VGND sg13g2_decap_8
XFILLER_36_512 VPWR VGND sg13g2_fill_1
XFILLER_48_383 VPWR VGND sg13g2_decap_8
XFILLER_36_578 VPWR VGND sg13g2_decap_8
XFILLER_23_239 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1027_ VGND VPWR net404 u_ppwm_u_mem__0641_/Y u_ppwm_u_mem__1190_/D
+ u_ppwm_u_mem__1026_/Y sg13g2_a21oi_1
XFILLER_20_935 VPWR VGND sg13g2_decap_8
XFILLER_32_773 VPWR VGND sg13g2_decap_8
Xfanout414 net415 net414 VPWR VGND sg13g2_buf_8
Xfanout403 net404 net403 VPWR VGND sg13g2_buf_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
Xfanout447 net686 net447 VPWR VGND sg13g2_buf_1
Xfanout425 fanout438/A net425 VPWR VGND sg13g2_buf_8
Xfanout436 net437 net436 VPWR VGND sg13g2_buf_8
Xfanout458 net669 net458 VPWR VGND sg13g2_buf_8
Xfanout469 net673 net469 VPWR VGND sg13g2_buf_8
XFILLER_39_372 VPWR VGND sg13g2_fill_1
XFILLER_27_578 VPWR VGND sg13g2_decap_8
XFILLER_42_537 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_decap_8
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_23_762 VPWR VGND sg13g2_decap_8
XFILLER_7_906 VPWR VGND sg13g2_decap_8
XFILLER_22_283 VPWR VGND sg13g2_fill_1
XFILLER_6_449 VPWR VGND sg13g2_fill_2
XFILLER_2_611 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1200__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_2_688 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_46_832 VPWR VGND sg13g2_decap_8
XFILLER_18_512 VPWR VGND sg13g2_decap_8
XFILLER_18_589 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0950_ u_ppwm_u_ex__0950_/A u_ppwm_u_ex__0950_/B u_ppwm_u_ex__0950_/C
+ u_ppwm_u_ex__0950_/D u_ppwm_u_ex__0950_/X VPWR VGND sg13g2_or4_1
XFILLER_14_762 VPWR VGND sg13g2_decap_8
XFILLER_9_221 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0881_ u_ppwm_u_ex__0881_/Y net460 net372 VPWR VGND sg13g2_xnor2_1
XFILLER_10_990 VPWR VGND sg13g2_decap_8
XFILLER_6_961 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__197_ hold17/A hold181/A u_ppwm_u_pwm__197_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_47_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_493 VPWR VGND sg13g2_decap_8
XFILLER_48_180 VPWR VGND sg13g2_decap_8
XFILLER_37_843 VPWR VGND sg13g2_decap_8
XFILLER_20_732 VPWR VGND sg13g2_decap_8
XFILLER_32_570 VPWR VGND sg13g2_decap_8
Xclkload7 clknet_5_22__leaf_clk clkload7/X VPWR VGND sg13g2_buf_1
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
XFILLER_3_408 VPWR VGND sg13g2_decap_8
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_43_846 VPWR VGND sg13g2_decap_8
XFILLER_15_537 VPWR VGND sg13g2_decap_8
XFILLER_30_507 VPWR VGND sg13g2_fill_1
XFILLER_11_721 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_fill_1
XFILLER_7_703 VPWR VGND sg13g2_decap_8
XFILLER_24_96 VPWR VGND sg13g2_fill_1
XFILLER_10_275 VPWR VGND sg13g2_fill_1
XFILLER_10_264 VPWR VGND sg13g2_fill_2
XFILLER_11_798 VPWR VGND sg13g2_decap_8
XFILLER_40_62 VPWR VGND sg13g2_fill_1
XFILLER_3_975 VPWR VGND sg13g2_decap_8
XFILLER_2_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1080_ u_ppwm_u_ex__1080_/Y hold295/A net371 VPWR VGND sg13g2_xnor2_1
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_876 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_fill_1
XFILLER_34_835 VPWR VGND sg13g2_decap_8
XFILLER_33_367 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0933_ u_ppwm_u_ex__1061_/A u_ppwm_u_ex__0933_/C net352 u_ppwm_u_ex__0933_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_14_1007 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0864_ VGND VPWR u_ppwm_u_ex__0882_/B u_ppwm_u_ex__0863_/Y u_ppwm_u_ex__0864_/Y
+ net358 sg13g2_a21oi_1
Xu_ppwm_u_pwm__249_ net198 VGND VPWR u_ppwm_u_pwm__249_/D net2 clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__0795_ u_ppwm_u_ex__0794_/Y VPWR u_ppwm_u_ex__0795_/Y VGND net378 u_ppwm_u_ex__0792_/Y
+ sg13g2_o21ai_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
Xhold19 hold19/A VPWR VGND net217 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1214__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_45_18 VPWR VGND sg13g2_decap_8
XFILLER_37_640 VPWR VGND sg13g2_decap_8
XFILLER_25_813 VPWR VGND sg13g2_decap_8
XFILLER_40_838 VPWR VGND sg13g2_decap_8
XFILLER_33_890 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1104__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_0_901 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_decap_4
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_47_459 VPWR VGND sg13g2_decap_8
XFILLER_28_673 VPWR VGND sg13g2_decap_8
XFILLER_43_643 VPWR VGND sg13g2_decap_8
XFILLER_15_334 VPWR VGND sg13g2_decap_8
XFILLER_16_846 VPWR VGND sg13g2_decap_8
XFILLER_37_1018 VPWR VGND sg13g2_decap_8
XFILLER_31_849 VPWR VGND sg13g2_decap_8
XFILLER_7_500 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0930_ net512 VPWR u_ppwm_u_mem__0930_/Y VGND net425 hold177/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0861_ VGND VPWR net424 u_ppwm_u_mem__0724_/Y hold230/A u_ppwm_u_mem__0860_/Y
+ sg13g2_a21oi_1
XFILLER_11_595 VPWR VGND sg13g2_decap_8
XFILLER_7_577 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0580_ VPWR u_ppwm_u_ex__0781_/A u_ppwm/instr\[0\] VGND sg13g2_inv_1
Xu_ppwm_u_mem__0792_ net475 u_ppwm_u_mem__0785_/Y u_ppwm_u_mem__0787_/Y u_ppwm_u_mem__0791_/Y
+ u_ppwm_u_mem__0789_/Y net393 u_ppwm_u_mem__0792_/X VPWR VGND sg13g2_mux4_1
XFILLER_3_772 VPWR VGND sg13g2_decap_8
XFILLER_39_927 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__121_ net507 VGND VPWR net623 hold254/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1063_ u_ppwm_u_ex__1063_/A u_ppwm_u_ex__1061_/Y u_ppwm_u_ex__1121_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_19_673 VPWR VGND sg13g2_decap_8
XFILLER_34_632 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0916_ net491 VPWR u_ppwm_u_ex__0917_/A VGND net458 net352 sg13g2_o21ai_1
XFILLER_30_882 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0847_ VPWR u_ppwm_u_ex__0847_/Y u_ppwm_u_ex__0847_/A VGND sg13g2_inv_1
Xu_ppwm_u_ex__0778_ u_ppwm_u_ex__0778_/Y net365 net575 net366 net445 VPWR VGND sg13g2_a22oi_1
XFILLER_45_919 VPWR VGND sg13g2_decap_8
XFILLER_44_407 VPWR VGND sg13g2_decap_8
XFILLER_25_610 VPWR VGND sg13g2_decap_8
XFILLER_37_470 VPWR VGND sg13g2_fill_1
XFILLER_40_635 VPWR VGND sg13g2_decap_8
XFILLER_25_687 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_fill_1
XFILLER_4_547 VPWR VGND sg13g2_decap_8
XFILLER_43_1000 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
XFILLER_48_768 VPWR VGND sg13g2_decap_8
XFILLER_47_256 VPWR VGND sg13g2_decap_8
XFILLER_46_61 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1060_ net500 VPWR u_ppwm_u_mem__1060_/Y VGND net406 hold60/A sg13g2_o21ai_1
XFILLER_16_643 VPWR VGND sg13g2_decap_8
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_43_440 VPWR VGND sg13g2_decap_8
XFILLER_31_646 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__236__195 VPWR VGND net195 sg13g2_tiehi
XFILLER_7_11 VPWR VGND sg13g2_decap_4
XFILLER_12_860 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0913_ VGND VPWR net435 u_ppwm_u_mem__0698_/Y u_ppwm_u_mem__1133_/D
+ u_ppwm_u_mem__0912_/Y sg13g2_a21oi_1
XFILLER_8_842 VPWR VGND sg13g2_decap_8
XFILLER_11_381 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0701_ hold313/A u_ppwm_u_ex__1020_/B2 u_ppwm_u_ex__0701_/Y VPWR VGND
+ sg13g2_nor2b_1
Xhold308 hold308/A VPWR VGND net676 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0632_ u_ppwm_u_ex__0626_/Y VPWR u_ppwm_u_ex__0634_/A VGND u_ppwm_u_ex__0628_/A
+ u_ppwm_u_ex__0628_/B sg13g2_o21ai_1
Xu_ppwm_u_mem__0844_ hold147/A hold128/A net476 u_ppwm_u_mem__0845_/B VPWR VGND sg13g2_mux2_1
Xhold319 hold319/A VPWR VGND net687 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0775_ hold60/A hold92/A net477 u_ppwm_u_mem__0776_/B VPWR VGND sg13g2_mux2_1
XFILLER_39_724 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__104_ VGND VPWR u_ppwm_u_global_counter__058_/Y u_ppwm_u_global_counter__101_/Y
+ hold253/A u_ppwm_u_global_counter__105_/B sg13g2_a21oi_1
Xu_ppwm_u_ex__1115_ net42 VGND VPWR u_ppwm_u_ex__1115_/D hold292/A clknet_5_18__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1046_ net351 u_ppwm_u_ex__1046_/C u_ppwm_u_ex__1046_/A u_ppwm_u_ex__1046_/Y
+ VPWR VGND u_ppwm_u_ex__1046_/D sg13g2_nand4_1
XFILLER_19_470 VPWR VGND sg13g2_decap_8
XFILLER_35_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1189_ net59 VGND VPWR net327 hold212/A clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_10_808 VPWR VGND sg13g2_decap_8
XFILLER_21_123 VPWR VGND sg13g2_decap_8
XFILLER_22_668 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_212 VPWR VGND sg13g2_decap_8
XFILLER_45_716 VPWR VGND sg13g2_decap_8
XFILLER_26_974 VPWR VGND sg13g2_decap_8
XFILLER_41_922 VPWR VGND sg13g2_decap_8
XFILLER_13_668 VPWR VGND sg13g2_decap_8
XFILLER_41_999 VPWR VGND sg13g2_decap_8
XFILLER_9_628 VPWR VGND sg13g2_decap_8
XFILLER_5_801 VPWR VGND sg13g2_decap_8
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_0_572 VPWR VGND sg13g2_decap_8
XFILLER_48_565 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1112_ net138 VGND VPWR u_ppwm_u_mem__1112_/D hold79/A clknet_5_22__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1043_ VGND VPWR net405 u_ppwm_u_mem__0633_/Y u_ppwm_u_mem__1198_/D
+ u_ppwm_u_mem__1042_/Y sg13g2_a21oi_1
XFILLER_44_771 VPWR VGND sg13g2_decap_8
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_43_281 VPWR VGND sg13g2_decap_4
XFILLER_32_955 VPWR VGND sg13g2_decap_8
Xhold105 hold105/A VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold116 hold116/A VPWR VGND net314 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0615_ u_ppwm_u_ex__0614_/Y VPWR u_ppwm_u_ex__0615_/Y VGND net473 net483
+ sg13g2_o21ai_1
Xhold149 hold149/A VPWR VGND net347 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0827_ u_ppwm_u_mem__0826_/Y u_ppwm_u_mem__0825_/Y u_ppwm_u_mem__0816_/Y
+ fanout383/A VPWR VGND sg13g2_a21o_2
Xhold127 hold127/A VPWR VGND net325 sg13g2_dlygate4sd3_1
Xhold138 hold138/A VPWR VGND net336 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0758_ hold103/A hold109/A net477 u_ppwm_u_mem__0758_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0689_ VPWR u_ppwm_u_mem__0689_/Y net220 VGND sg13g2_inv_1
XFILLER_39_521 VPWR VGND sg13g2_decap_8
XFILLER_26_226 VPWR VGND sg13g2_fill_2
XFILLER_39_598 VPWR VGND sg13g2_decap_8
XFILLER_42_719 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1029_ u_ppwm_u_ex__1028_/Y VPWR u_ppwm_u_ex__1029_/Y VGND u_ppwm_u_ex__1006_/A
+ u_ppwm_u_ex__1027_/X sg13g2_o21ai_1
XFILLER_26_248 VPWR VGND sg13g2_decap_4
XFILLER_23_944 VPWR VGND sg13g2_decap_8
XFILLER_10_605 VPWR VGND sg13g2_decap_8
XFILLER_22_465 VPWR VGND sg13g2_decap_8
XFILLER_45_513 VPWR VGND sg13g2_decap_8
XFILLER_33_708 VPWR VGND sg13g2_decap_8
XFILLER_26_771 VPWR VGND sg13g2_decap_8
XFILLER_14_944 VPWR VGND sg13g2_decap_8
XFILLER_41_796 VPWR VGND sg13g2_decap_8
XFILLER_5_675 VPWR VGND sg13g2_decap_8
XFILLER_49_830 VPWR VGND sg13g2_decap_8
XFILLER_48_362 VPWR VGND sg13g2_decap_8
XFILLER_36_557 VPWR VGND sg13g2_decap_8
XFILLER_17_782 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1026_ net494 VPWR u_ppwm_u_mem__1026_/Y VGND net404 net326 sg13g2_o21ai_1
Xu_ppwm_u_mem__1169__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_16_281 VPWR VGND sg13g2_fill_1
XFILLER_32_752 VPWR VGND sg13g2_decap_8
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_914 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_fill_1
XFILLER_9_992 VPWR VGND sg13g2_decap_8
Xfanout404 net405 net404 VPWR VGND sg13g2_buf_8
Xfanout415 net416 net415 VPWR VGND sg13g2_buf_8
Xfanout448 net671 net448 VPWR VGND sg13g2_buf_8
Xfanout426 net438 net426 VPWR VGND sg13g2_buf_8
Xfanout437 net438 net437 VPWR VGND sg13g2_buf_2
Xfanout459 hold301/A net459 VPWR VGND sg13g2_buf_1
Xu_ppwm_u_mem__1191__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_15_719 VPWR VGND sg13g2_decap_8
XFILLER_27_557 VPWR VGND sg13g2_decap_8
XFILLER_42_516 VPWR VGND sg13g2_decap_8
XFILLER_23_741 VPWR VGND sg13g2_decap_8
XFILLER_11_903 VPWR VGND sg13g2_decap_8
XFILLER_2_667 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_46_811 VPWR VGND sg13g2_decap_8
XFILLER_38_51 VPWR VGND sg13g2_fill_1
XFILLER_45_310 VPWR VGND sg13g2_decap_8
XFILLER_18_568 VPWR VGND sg13g2_decap_8
XFILLER_46_888 VPWR VGND sg13g2_decap_8
XFILLER_45_387 VPWR VGND sg13g2_decap_8
XFILLER_14_741 VPWR VGND sg13g2_decap_8
XFILLER_41_593 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0880_ u_ppwm_u_ex__0880_/Y net460 net372 VPWR VGND sg13g2_nand2_1
XFILLER_13_273 VPWR VGND sg13g2_fill_1
XFILLER_6_940 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__196_ u_ppwm_u_pwm__195_/Y VPWR u_ppwm_u_pwm__196_/Y VGND u_ppwm_u_pwm__202_/A
+ u_ppwm_u_pwm__202_/B sg13g2_o21ai_1
XFILLER_5_472 VPWR VGND sg13g2_decap_8
XFILLER_36_310 VPWR VGND sg13g2_fill_2
XFILLER_37_822 VPWR VGND sg13g2_decap_8
XFILLER_37_899 VPWR VGND sg13g2_decap_8
XFILLER_24_549 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1009_ VGND VPWR net409 u_ppwm_u_mem__0650_/Y u_ppwm_u_mem__1181_/D
+ u_ppwm_u_mem__1008_/Y sg13g2_a21oi_1
XFILLER_20_711 VPWR VGND sg13g2_decap_8
Xclkload8 clknet_5_24__leaf_clk clkload8/X VPWR VGND sg13g2_buf_1
XFILLER_20_788 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1223__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_43_825 VPWR VGND sg13g2_decap_8
XFILLER_15_516 VPWR VGND sg13g2_decap_8
XFILLER_27_387 VPWR VGND sg13g2_fill_1
XFILLER_11_700 VPWR VGND sg13g2_decap_8
XFILLER_10_210 VPWR VGND sg13g2_fill_1
XFILLER_7_759 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_fill_1
XFILLER_11_777 VPWR VGND sg13g2_decap_8
XFILLER_3_954 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_855 VPWR VGND sg13g2_decap_8
XFILLER_46_685 VPWR VGND sg13g2_decap_8
XFILLER_18_365 VPWR VGND sg13g2_decap_8
XFILLER_34_814 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1133__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_21_519 VPWR VGND sg13g2_decap_8
XFILLER_42_880 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0932_ VGND VPWR net448 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0933_/C u_ppwm_u_ex__0931_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0863_ VGND VPWR u_ppwm_u_ex__0849_/Y u_ppwm_u_ex__0851_/X u_ppwm_u_ex__0863_/Y
+ u_ppwm_u_ex__0850_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0794_ u_ppwm_u_ex__0794_/Y net379 u_ppwm_u_ex__0866_/C VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_pwm__248_ net184 VGND VPWR net595 hold274/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__179_ VGND VPWR hold268/A u_ppwm_u_pwm__180_/C hold179/A net546 sg13g2_a21oi_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_24_313 VPWR VGND sg13g2_decap_8
XFILLER_25_869 VPWR VGND sg13g2_decap_8
XFILLER_37_696 VPWR VGND sg13g2_decap_8
XFILLER_40_817 VPWR VGND sg13g2_decap_8
XFILLER_20_585 VPWR VGND sg13g2_decap_8
XFILLER_4_729 VPWR VGND sg13g2_decap_8
XFILLER_0_957 VPWR VGND sg13g2_decap_8
XFILLER_47_438 VPWR VGND sg13g2_decap_8
XFILLER_19_107 VPWR VGND sg13g2_fill_2
XFILLER_19_129 VPWR VGND sg13g2_fill_1
XFILLER_28_652 VPWR VGND sg13g2_decap_8
XFILLER_15_302 VPWR VGND sg13g2_decap_8
XFILLER_16_825 VPWR VGND sg13g2_decap_8
XFILLER_43_622 VPWR VGND sg13g2_decap_8
XFILLER_27_195 VPWR VGND sg13g2_fill_1
XFILLER_43_699 VPWR VGND sg13g2_decap_8
XFILLER_31_828 VPWR VGND sg13g2_decap_8
XFILLER_11_574 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0860_ net513 VPWR u_ppwm_u_mem__0860_/Y VGND net423 net597 sg13g2_o21ai_1
XFILLER_7_556 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0791_ u_ppwm_u_mem__0790_/Y VPWR u_ppwm_u_mem__0791_/Y VGND u_ppwm_u_mem__0723_/Y
+ net484 sg13g2_o21ai_1
XFILLER_3_751 VPWR VGND sg13g2_decap_8
XFILLER_2_261 VPWR VGND sg13g2_fill_1
XFILLER_39_906 VPWR VGND sg13g2_decap_8
XFILLER_2_294 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__120_ net507 VGND VPWR net610 hold240/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1062_ net505 VPWR u_ppwm_u_ex__1063_/A VGND net448 net349 sg13g2_o21ai_1
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_18_151 VPWR VGND sg13g2_fill_1
XFILLER_19_652 VPWR VGND sg13g2_decap_8
XFILLER_46_482 VPWR VGND sg13g2_decap_8
XFILLER_34_611 VPWR VGND sg13g2_decap_8
XFILLER_33_132 VPWR VGND sg13g2_fill_2
XFILLER_15_880 VPWR VGND sg13g2_decap_8
XFILLER_33_165 VPWR VGND sg13g2_fill_1
XFILLER_34_688 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0915_ u_ppwm_u_ex__0915_/B u_ppwm_u_ex__1046_/A net353 u_ppwm_u_ex__0915_/Y
+ VPWR VGND u_ppwm_u_ex__0915_/D sg13g2_nand4_1
XFILLER_30_861 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0846_ u_ppwm_u_ex__0845_/Y VPWR u_ppwm_u_ex__0847_/A VGND net378 u_ppwm_u_ex__0812_/X
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0989_ VGND VPWR net416 u_ppwm_u_mem__0660_/Y hold106/A u_ppwm_u_mem__0988_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0777_ net366 net364 net359 u_ppwm_u_ex__0831_/B VPWR VGND sg13g2_nor3_2
XFILLER_29_416 VPWR VGND sg13g2_fill_1
XFILLER_25_666 VPWR VGND sg13g2_decap_8
XFILLER_40_614 VPWR VGND sg13g2_decap_8
XFILLER_12_316 VPWR VGND sg13g2_decap_4
XFILLER_21_883 VPWR VGND sg13g2_decap_8
XFILLER_4_526 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1179__99 VPWR VGND net99 sg13g2_tiehi
XFILLER_0_754 VPWR VGND sg13g2_decap_8
XFILLER_48_747 VPWR VGND sg13g2_decap_8
XFILLER_47_235 VPWR VGND sg13g2_decap_8
XFILLER_16_622 VPWR VGND sg13g2_decap_8
XFILLER_29_994 VPWR VGND sg13g2_decap_8
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_43_496 VPWR VGND sg13g2_decap_8
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_16_699 VPWR VGND sg13g2_decap_8
XFILLER_31_625 VPWR VGND sg13g2_decap_8
XFILLER_8_821 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0700_ net452 net440 u_ppwm_u_ex__0700_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0912_ net511 VPWR u_ppwm_u_mem__0912_/Y VGND net435 net336 sg13g2_o21ai_1
XFILLER_8_898 VPWR VGND sg13g2_decap_8
XFILLER_7_78 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0631_ u_ppwm_u_ex__0991_/A net674 u_ppwm_u_ex__1101_/D VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0843_ u_ppwm_u_mem__0842_/Y VPWR fanout380/A VGND u_ppwm_u_mem__0835_/Y
+ u_ppwm_u_mem__0836_/Y sg13g2_o21ai_1
Xhold309 hold309/A VPWR VGND net677 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0774_ u_ppwm_u_mem__0773_/X u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0764_/Y
+ u_ppwm/instr\[1\] VPWR VGND sg13g2_a21o_2
XFILLER_30_4 VPWR VGND sg13g2_fill_1
XFILLER_39_703 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__103_ net620 net392 u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__103_/D
+ u_ppwm_u_global_counter__105_/B VPWR VGND sg13g2_and4_1
Xu_ppwm_u_ex__1114_ net46 VGND VPWR u_ppwm_u_ex__1114_/D hold307/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_38_213 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__1045_ u_ppwm_u_ex__1044_/Y u_ppwm_u_ex__1043_/Y net359 u_ppwm_u_ex__1046_/D
+ VPWR VGND sg13g2_a21o_1
XFILLER_35_920 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1188_ net63 VGND VPWR u_ppwm_u_mem__1188_/D hold121/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_997 VPWR VGND sg13g2_decap_8
XFILLER_22_647 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0829_ u_ppwm_u_ex__0996_/A u_ppwm_u_ex__0829_/C net354 u_ppwm_u_ex__0833_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_44_205 VPWR VGND sg13g2_fill_2
XFILLER_41_901 VPWR VGND sg13g2_decap_8
XFILLER_26_953 VPWR VGND sg13g2_decap_8
XFILLER_9_607 VPWR VGND sg13g2_decap_8
XFILLER_12_135 VPWR VGND sg13g2_decap_4
XFILLER_13_647 VPWR VGND sg13g2_decap_8
XFILLER_41_978 VPWR VGND sg13g2_decap_8
XFILLER_40_488 VPWR VGND sg13g2_decap_8
XFILLER_8_128 VPWR VGND sg13g2_fill_2
XFILLER_21_680 VPWR VGND sg13g2_decap_8
XFILLER_5_857 VPWR VGND sg13g2_decap_8
XFILLER_10_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_551 VPWR VGND sg13g2_decap_8
XFILLER_48_544 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1111_ net140 VGND VPWR u_ppwm_u_mem__1111_/D hold44/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_29_791 VPWR VGND sg13g2_decap_8
XFILLER_36_739 VPWR VGND sg13g2_decap_8
XFILLER_44_750 VPWR VGND sg13g2_decap_8
XFILLER_17_964 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1042_ net495 VPWR u_ppwm_u_mem__1042_/Y VGND net405 net205 sg13g2_o21ai_1
XFILLER_32_934 VPWR VGND sg13g2_decap_8
XFILLER_16_496 VPWR VGND sg13g2_decap_8
Xhold106 hold106/A VPWR VGND net304 sg13g2_dlygate4sd3_1
Xhold117 hold117/A VPWR VGND net315 sg13g2_dlygate4sd3_1
XFILLER_8_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0614_ net447 VPWR u_ppwm_u_ex__0614_/Y VGND u_ppwm_u_ex__0622_/B u_ppwm_u_ex__0623_/B
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0826_ VGND VPWR u_ppwm_u_mem__0818_/Y u_ppwm_u_mem__0820_/Y u_ppwm_u_mem__0826_/Y
+ net467 sg13g2_a21oi_1
Xhold139 hold139/A VPWR VGND net337 sg13g2_dlygate4sd3_1
Xhold128 hold128/A VPWR VGND net326 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0757_ u_ppwm_u_mem__0756_/Y u_ppwm_u_mem__0751_/Y u_ppwm_u_mem__0749_/Y
+ u_ppwm/instr\[0\] VPWR VGND sg13g2_a21o_2
XFILLER_4_890 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0688_ VPWR u_ppwm_u_mem__0688_/Y net337 VGND sg13g2_inv_1
XFILLER_39_500 VPWR VGND sg13g2_decap_8
XFILLER_39_577 VPWR VGND sg13g2_decap_8
XFILLER_27_739 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1028_ net376 VPWR u_ppwm_u_ex__1028_/Y VGND net450 net451 sg13g2_o21ai_1
XFILLER_23_923 VPWR VGND sg13g2_decap_8
XFILLER_22_411 VPWR VGND sg13g2_fill_1
XFILLER_22_444 VPWR VGND sg13g2_decap_8
XFILLER_35_794 VPWR VGND sg13g2_decap_8
XFILLER_2_849 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_fill_1
XFILLER_45_569 VPWR VGND sg13g2_decap_8
XFILLER_26_750 VPWR VGND sg13g2_decap_8
XFILLER_14_923 VPWR VGND sg13g2_decap_8
XFILLER_41_775 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_fill_1
XFILLER_5_654 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_fill_2
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_49_886 VPWR VGND sg13g2_decap_8
XFILLER_48_341 VPWR VGND sg13g2_decap_8
XFILLER_36_536 VPWR VGND sg13g2_decap_8
XFILLER_17_761 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1025_ VGND VPWR net410 u_ppwm_u_mem__0642_/Y hold129/A u_ppwm_u_mem__1024_/Y
+ sg13g2_a21oi_1
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
XFILLER_32_731 VPWR VGND sg13g2_decap_8
XFILLER_9_971 VPWR VGND sg13g2_decap_8
XFILLER_8_492 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0809_ u_ppwm_u_mem__0808_/Y u_ppwm_u_mem__0806_/Y u_ppwm_u_mem__0802_/Y
+ fanout387/A VPWR VGND sg13g2_a21o_1
Xfanout405 net406 net405 VPWR VGND sg13g2_buf_8
Xfanout416 net422 net416 VPWR VGND sg13g2_buf_2
Xfanout427 net431 net427 VPWR VGND sg13g2_buf_8
Xfanout438 fanout438/A net438 VPWR VGND sg13g2_buf_1
Xfanout449 net682 net449 VPWR VGND sg13g2_buf_8
XFILLER_27_536 VPWR VGND sg13g2_decap_8
XFILLER_23_720 VPWR VGND sg13g2_decap_8
XFILLER_35_591 VPWR VGND sg13g2_decap_8
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_fill_2
XFILLER_23_797 VPWR VGND sg13g2_decap_8
XFILLER_6_407 VPWR VGND sg13g2_fill_1
XFILLER_6_429 VPWR VGND sg13g2_decap_4
XFILLER_2_646 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_46_867 VPWR VGND sg13g2_decap_8
XFILLER_18_547 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1145__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_45_366 VPWR VGND sg13g2_decap_8
XFILLER_14_720 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_decap_8
XFILLER_9_201 VPWR VGND sg13g2_decap_4
XFILLER_14_797 VPWR VGND sg13g2_decap_8
XFILLER_9_245 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__195_ u_ppwm_u_pwm__195_/Y hold165/A hold283/A VPWR VGND sg13g2_nand2b_1
XFILLER_6_996 VPWR VGND sg13g2_decap_8
XFILLER_5_451 VPWR VGND sg13g2_decap_8
XFILLER_23_1021 VPWR VGND sg13g2_decap_8
XFILLER_37_801 VPWR VGND sg13g2_decap_8
XFILLER_49_683 VPWR VGND sg13g2_decap_8
XFILLER_24_528 VPWR VGND sg13g2_decap_8
XFILLER_37_878 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1008_ net496 VPWR u_ppwm_u_mem__1008_/Y VGND net409 net244 sg13g2_o21ai_1
XFILLER_20_767 VPWR VGND sg13g2_decap_8
Xclkload9 clknet_5_31__leaf_clk clkload9/X VPWR VGND sg13g2_buf_1
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_43_804 VPWR VGND sg13g2_decap_8
XFILLER_42_369 VPWR VGND sg13g2_fill_1
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_23_594 VPWR VGND sg13g2_decap_8
XFILLER_7_738 VPWR VGND sg13g2_decap_8
XFILLER_3_933 VPWR VGND sg13g2_decap_8
XFILLER_46_1021 VPWR VGND sg13g2_decap_8
XFILLER_2_443 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_19_834 VPWR VGND sg13g2_decap_8
XFILLER_18_311 VPWR VGND sg13g2_fill_2
XFILLER_46_664 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0931_ net361 u_ppwm_u_ex__0931_/B u_ppwm_u_ex__0931_/Y VPWR VGND sg13g2_nor2_1
XFILLER_14_594 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0862_ u_ppwm_u_ex__0882_/B net462 net374 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__0793_ net463 net451 net386 u_ppwm_u_ex__0866_/C VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_pwm__247_ net194 VGND VPWR u_ppwm_u_pwm__247_/D hold276/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__178_ u_ppwm_u_pwm__188_/A u_ppwm_u_pwm__178_/B u_ppwm_u_pwm__244_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_793 VPWR VGND sg13g2_decap_8
XFILLER_29_609 VPWR VGND sg13g2_decap_8
XFILLER_49_480 VPWR VGND sg13g2_decap_8
XFILLER_36_130 VPWR VGND sg13g2_fill_2
XFILLER_37_675 VPWR VGND sg13g2_decap_8
XFILLER_25_848 VPWR VGND sg13g2_decap_8
XFILLER_20_564 VPWR VGND sg13g2_decap_8
XFILLER_4_708 VPWR VGND sg13g2_decap_8
XFILLER_0_936 VPWR VGND sg13g2_decap_8
XFILLER_48_929 VPWR VGND sg13g2_decap_8
XFILLER_47_417 VPWR VGND sg13g2_decap_8
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_43_601 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_42_111 VPWR VGND sg13g2_fill_1
XFILLER_43_678 VPWR VGND sg13g2_decap_8
XFILLER_42_122 VPWR VGND sg13g2_fill_1
XFILLER_31_807 VPWR VGND sg13g2_decap_8
XFILLER_24_892 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_553 VPWR VGND sg13g2_decap_8
XFILLER_7_535 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0790_ u_ppwm_u_mem__0790_/Y hold193/A net484 VPWR VGND sg13g2_nand2_1
XFILLER_3_730 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1061_ net349 u_ppwm_u_ex__1061_/C u_ppwm_u_ex__1061_/A u_ppwm_u_ex__1061_/Y
+ VPWR VGND u_ppwm_u_ex__1061_/D sg13g2_nand4_1
XFILLER_19_631 VPWR VGND sg13g2_decap_8
XFILLER_47_984 VPWR VGND sg13g2_decap_8
XFILLER_46_461 VPWR VGND sg13g2_decap_8
XFILLER_18_196 VPWR VGND sg13g2_fill_2
XFILLER_34_667 VPWR VGND sg13g2_decap_8
XFILLER_22_829 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0914_ VGND VPWR hold299/A u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0915_/D
+ u_ppwm_u_ex__0913_/Y sg13g2_a21oi_1
XFILLER_21_339 VPWR VGND sg13g2_fill_1
XFILLER_30_840 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0845_ u_ppwm_u_ex__0845_/Y net378 u_ppwm_u_ex__0845_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0988_ net498 VPWR u_ppwm_u_mem__0988_/Y VGND net415 net251 sg13g2_o21ai_1
Xu_ppwm_u_ex__0776_ fanout361/A net388 u_ppwm_u_ex__0805_/C VPWR VGND sg13g2_nand2_2
XFILLER_6_590 VPWR VGND sg13g2_decap_8
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
XFILLER_38_984 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_fill_2
XFILLER_25_645 VPWR VGND sg13g2_decap_8
XFILLER_12_306 VPWR VGND sg13g2_fill_1
XFILLER_13_829 VPWR VGND sg13g2_decap_8
XFILLER_21_862 VPWR VGND sg13g2_decap_8
XFILLER_20_372 VPWR VGND sg13g2_fill_2
XFILLER_4_505 VPWR VGND sg13g2_decap_8
XFILLER_0_733 VPWR VGND sg13g2_decap_8
XFILLER_48_726 VPWR VGND sg13g2_decap_8
XFILLER_47_214 VPWR VGND sg13g2_decap_8
XFILLER_29_973 VPWR VGND sg13g2_decap_8
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_16_601 VPWR VGND sg13g2_decap_8
XFILLER_43_475 VPWR VGND sg13g2_decap_8
XFILLER_16_678 VPWR VGND sg13g2_decap_8
XFILLER_31_604 VPWR VGND sg13g2_decap_8
XFILLER_15_199 VPWR VGND sg13g2_fill_2
XFILLER_30_114 VPWR VGND sg13g2_fill_2
XFILLER_8_800 VPWR VGND sg13g2_decap_8
XFILLER_30_169 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0911_ VGND VPWR net436 u_ppwm_u_mem__0699_/Y u_ppwm_u_mem__1132_/D
+ u_ppwm_u_mem__0910_/Y sg13g2_a21oi_1
XFILLER_11_372 VPWR VGND sg13g2_decap_8
XFILLER_12_895 VPWR VGND sg13g2_decap_8
XFILLER_8_877 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0630_ u_ppwm_u_ex__0629_/Y VPWR hold306/A VGND net447 net469 sg13g2_o21ai_1
Xu_ppwm_u_mem__0842_ u_ppwm_u_mem__0842_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0842_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0773_ net475 u_ppwm_u_mem__0766_/Y u_ppwm_u_mem__0768_/Y u_ppwm_u_mem__0772_/Y
+ u_ppwm_u_mem__0770_/Y net393 u_ppwm_u_mem__0773_/X VPWR VGND sg13g2_mux4_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__102_ hold278/A u_ppwm_u_global_counter__103_/D u_ppwm_u_global_counter__099_/B
+ u_ppwm_u_global_counter__098_/Y u_ppwm_u_global_counter__057_/Y VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_ex__1113_ net50 VGND VPWR u_ppwm_u_ex__1113_/D hold304/A clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_759 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1044_ u_ppwm_u_ex__1044_/Y fanout356/A hold259/A net362 net459 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_47_781 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1187_ net67 VGND VPWR u_ppwm_u_mem__1187_/D hold38/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_22_626 VPWR VGND sg13g2_decap_8
XFILLER_21_158 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1109__144 VPWR VGND net144 sg13g2_tiehi
Xu_ppwm_u_ex__0828_ u_ppwm_u_ex__0827_/Y VPWR u_ppwm_u_ex__0829_/C VGND u_ppwm_u_ex__0782_/Y
+ u_ppwm_u_ex__0826_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__0759_ hold236/A net456 u_ppwm_u_ex__0760_/D VPWR VGND sg13g2_xor2_1
XFILLER_27_1019 VPWR VGND sg13g2_decap_8
XFILLER_17_409 VPWR VGND sg13g2_decap_4
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_26_932 VPWR VGND sg13g2_decap_8
XFILLER_38_781 VPWR VGND sg13g2_decap_8
XFILLER_37_291 VPWR VGND sg13g2_decap_4
XFILLER_13_626 VPWR VGND sg13g2_decap_8
XFILLER_41_957 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_40_467 VPWR VGND sg13g2_decap_8
XFILLER_20_191 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1162__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_5_836 VPWR VGND sg13g2_decap_8
XFILLER_0_530 VPWR VGND sg13g2_decap_8
XFILLER_48_523 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1110_ net142 VGND VPWR net243 hold143/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_718 VPWR VGND sg13g2_decap_8
XFILLER_29_770 VPWR VGND sg13g2_decap_8
XFILLER_17_943 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1041_ VGND VPWR net405 u_ppwm_u_mem__0634_/Y hold8/A u_ppwm_u_mem__1040_/Y
+ sg13g2_a21oi_1
XFILLER_32_913 VPWR VGND sg13g2_decap_8
XFILLER_8_674 VPWR VGND sg13g2_decap_8
XFILLER_12_692 VPWR VGND sg13g2_decap_8
XFILLER_7_151 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0613_ u_ppwm_u_ex__0991_/A u_ppwm_u_ex__0613_/B u_ppwm_u_ex__1099_/D
+ VPWR VGND sg13g2_nor2_1
Xhold107 hold107/A VPWR VGND net305 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0825_ u_ppwm_u_mem__0825_/Y u_ppwm_u_mem__0825_/B u_ppwm_u_mem__0822_/Y
+ VPWR VGND sg13g2_nand2b_1
Xhold118 hold118/A VPWR VGND net316 sg13g2_dlygate4sd3_1
Xhold129 hold129/A VPWR VGND net327 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0756_ VGND VPWR u_ppwm_u_mem__0754_/Y u_ppwm_u_mem__0755_/Y u_ppwm_u_mem__0756_/Y
+ net467 sg13g2_a21oi_1
Xu_ppwm_u_mem__0687_ VPWR u_ppwm_u_mem__0687_/Y net320 VGND sg13g2_inv_1
XFILLER_27_718 VPWR VGND sg13g2_decap_8
XFILLER_39_556 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1027_ VGND VPWR u_ppwm_u_ex__1027_/X u_ppwm_u_ex__1027_/B u_ppwm_u_ex__1027_/A
+ sg13g2_or2_1
XFILLER_23_902 VPWR VGND sg13g2_decap_8
XFILLER_35_773 VPWR VGND sg13g2_decap_8
XFILLER_34_272 VPWR VGND sg13g2_fill_1
XFILLER_23_979 VPWR VGND sg13g2_decap_8
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1226__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_2_828 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_729 VPWR VGND sg13g2_decap_8
XFILLER_45_548 VPWR VGND sg13g2_decap_8
XFILLER_14_902 VPWR VGND sg13g2_decap_8
XFILLER_41_754 VPWR VGND sg13g2_decap_8
XFILLER_14_979 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_fill_2
XFILLER_22_990 VPWR VGND sg13g2_decap_8
XFILLER_5_633 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_4_36 VPWR VGND sg13g2_fill_2
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_48_320 VPWR VGND sg13g2_decap_8
XFILLER_49_865 VPWR VGND sg13g2_decap_8
XFILLER_48_397 VPWR VGND sg13g2_decap_8
XFILLER_17_740 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1024_ net495 VPWR u_ppwm_u_mem__1024_/Y VGND net410 hold212/A sg13g2_o21ai_1
XFILLER_32_710 VPWR VGND sg13g2_decap_8
XFILLER_16_294 VPWR VGND sg13g2_fill_2
XFILLER_13_990 VPWR VGND sg13g2_decap_8
XFILLER_20_949 VPWR VGND sg13g2_decap_8
XFILLER_32_787 VPWR VGND sg13g2_decap_8
XFILLER_9_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0808_ VGND VPWR net393 u_ppwm_u_mem__0807_/X u_ppwm_u_mem__0808_/Y
+ net467 sg13g2_a21oi_1
Xu_ppwm_u_mem__0739_ net488 net333 net1 u_ppwm_u_mem__0739_/Y VPWR VGND sg13g2_nand3_1
Xfanout428 net431 net428 VPWR VGND sg13g2_buf_1
Xfanout439 net654 net439 VPWR VGND sg13g2_buf_8
Xfanout406 net422 net406 VPWR VGND sg13g2_buf_8
Xfanout417 net418 net417 VPWR VGND sg13g2_buf_8
XFILLER_27_515 VPWR VGND sg13g2_decap_8
XFILLER_35_570 VPWR VGND sg13g2_decap_8
XFILLER_23_776 VPWR VGND sg13g2_decap_8
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_22_297 VPWR VGND sg13g2_fill_1
XFILLER_2_625 VPWR VGND sg13g2_decap_8
XFILLER_18_526 VPWR VGND sg13g2_decap_8
XFILLER_46_846 VPWR VGND sg13g2_decap_8
XFILLER_45_345 VPWR VGND sg13g2_decap_8
XFILLER_41_551 VPWR VGND sg13g2_decap_8
XFILLER_13_220 VPWR VGND sg13g2_decap_8
XFILLER_13_264 VPWR VGND sg13g2_decap_8
XFILLER_14_776 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1125__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_5_430 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__194_ hold283/A hold165/A u_ppwm_u_pwm__202_/C VPWR VGND sg13g2_nor2b_1
XFILLER_6_975 VPWR VGND sg13g2_decap_8
XFILLER_23_1000 VPWR VGND sg13g2_decap_8
XFILLER_49_662 VPWR VGND sg13g2_decap_8
XFILLER_48_194 VPWR VGND sg13g2_decap_8
XFILLER_37_857 VPWR VGND sg13g2_decap_8
XFILLER_24_507 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1007_ VGND VPWR net412 u_ppwm_u_mem__0651_/Y u_ppwm_u_mem__1180_/D
+ u_ppwm_u_mem__1006_/Y sg13g2_a21oi_1
XFILLER_32_584 VPWR VGND sg13g2_decap_8
XFILLER_20_746 VPWR VGND sg13g2_decap_8
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_301 VPWR VGND sg13g2_fill_1
XFILLER_28_813 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_fill_2
XFILLER_23_573 VPWR VGND sg13g2_decap_8
XFILLER_11_735 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_fill_2
XFILLER_10_256 VPWR VGND sg13g2_decap_4
XFILLER_7_717 VPWR VGND sg13g2_decap_8
XFILLER_3_912 VPWR VGND sg13g2_decap_8
XFILLER_46_1000 VPWR VGND sg13g2_decap_8
XFILLER_2_422 VPWR VGND sg13g2_decap_8
XFILLER_3_989 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
Xhold290 hold290/A VPWR VGND net658 sg13g2_dlygate4sd3_1
XFILLER_2_499 VPWR VGND sg13g2_decap_8
XFILLER_19_813 VPWR VGND sg13g2_decap_8
XFILLER_46_643 VPWR VGND sg13g2_decap_8
XFILLER_45_164 VPWR VGND sg13g2_fill_2
XFILLER_34_849 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0930_ u_ppwm_u_ex__0931_/B net365 net439 net367 hold236/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_14_573 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0861_ u_ppwm_u_ex__0861_/A u_ppwm_u_ex__0859_/Y u_ppwm_u_ex__1107_/D
+ VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_ex__0792_ u_ppwm_u_ex__0791_/X VPWR u_ppwm_u_ex__0792_/Y VGND net453 u_ppwm_u_ex__0979_/A
+ sg13g2_o21ai_1
Xu_ppwm_u_pwm__246_ net180 VGND VPWR u_ppwm_u_pwm__246_/D hold225/A clknet_5_1__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__177_ u_ppwm_u_pwm__178_/B net636 u_ppwm_u_pwm__180_/C VPWR VGND sg13g2_xnor2_1
XFILLER_6_772 VPWR VGND sg13g2_decap_8
XFILLER_37_654 VPWR VGND sg13g2_decap_8
XFILLER_18_890 VPWR VGND sg13g2_decap_8
XFILLER_25_827 VPWR VGND sg13g2_decap_8
XFILLER_20_543 VPWR VGND sg13g2_decap_8
XFILLER_0_915 VPWR VGND sg13g2_decap_8
XFILLER_48_908 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1119__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_28_610 VPWR VGND sg13g2_decap_8
XFILLER_28_687 VPWR VGND sg13g2_decap_8
XFILLER_43_657 VPWR VGND sg13g2_decap_8
XFILLER_15_359 VPWR VGND sg13g2_fill_2
XFILLER_24_871 VPWR VGND sg13g2_decap_8
XFILLER_11_532 VPWR VGND sg13g2_decap_8
XFILLER_7_514 VPWR VGND sg13g2_decap_8
XFILLER_3_786 VPWR VGND sg13g2_decap_8
XFILLER_2_296 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1060_ u_ppwm_u_ex__1059_/Y u_ppwm_u_ex__1058_/Y net359 u_ppwm_u_ex__1061_/D
+ VPWR VGND sg13g2_a21o_1
XFILLER_19_610 VPWR VGND sg13g2_decap_8
XFILLER_47_963 VPWR VGND sg13g2_decap_8
XFILLER_46_440 VPWR VGND sg13g2_decap_8
XFILLER_19_687 VPWR VGND sg13g2_decap_8
XFILLER_22_808 VPWR VGND sg13g2_decap_8
XFILLER_33_134 VPWR VGND sg13g2_fill_1
XFILLER_34_646 VPWR VGND sg13g2_decap_8
XFILLER_21_307 VPWR VGND sg13g2_fill_2
XFILLER_33_156 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0913_ net359 u_ppwm_u_ex__0913_/B u_ppwm_u_ex__0913_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0844_ net456 net448 net384 u_ppwm_u_ex__0845_/B VPWR VGND sg13g2_mux2_1
XFILLER_30_896 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0987_ VGND VPWR net420 u_ppwm_u_mem__0661_/Y hold54/A u_ppwm_u_mem__0986_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__229_ net187 VGND VPWR net216 hold17/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__0775_ net388 u_ppwm_u_ex__0805_/C u_ppwm_u_ex__0784_/A VPWR VGND sg13g2_and2_1
Xu_ppwm_u_ex__1101__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_44_0 VPWR VGND sg13g2_decap_4
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_37_451 VPWR VGND sg13g2_fill_1
XFILLER_38_963 VPWR VGND sg13g2_decap_8
XFILLER_25_624 VPWR VGND sg13g2_decap_8
XFILLER_13_808 VPWR VGND sg13g2_decap_8
XFILLER_40_649 VPWR VGND sg13g2_decap_8
XFILLER_21_841 VPWR VGND sg13g2_decap_8
XFILLER_0_712 VPWR VGND sg13g2_decap_8
XFILLER_43_1014 VPWR VGND sg13g2_decap_8
XFILLER_48_705 VPWR VGND sg13g2_decap_8
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_16_657 VPWR VGND sg13g2_decap_8
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_43_454 VPWR VGND sg13g2_decap_8
XFILLER_12_874 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0910_ net515 VPWR u_ppwm_u_mem__0910_/Y VGND net436 net262 sg13g2_o21ai_1
XFILLER_8_856 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0841_ net474 u_ppwm_u_mem__0837_/X u_ppwm_u_mem__0838_/X u_ppwm_u_mem__0840_/X
+ u_ppwm_u_mem__0839_/X net393 u_ppwm_u_mem__0842_/B VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0772_ u_ppwm_u_mem__0771_/Y VPWR u_ppwm_u_mem__0772_/Y VGND u_ppwm_u_mem__0724_/Y
+ net484 sg13g2_o21ai_1
XFILLER_3_583 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__101_ u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__103_/D
+ net392 u_ppwm_u_global_counter__101_/Y VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__1112_ net27 VGND VPWR u_ppwm_u_ex__1112_/D hold296/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_39_738 VPWR VGND sg13g2_decap_8
XFILLER_47_760 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1043_ u_ppwm_u_ex__1043_/Y hold254/A fanout355/A VPWR VGND sg13g2_nand2_1
XFILLER_19_440 VPWR VGND sg13g2_decap_8
XFILLER_19_484 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1186_ net71 VGND VPWR net237 hold51/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_955 VPWR VGND sg13g2_decap_8
XFILLER_22_605 VPWR VGND sg13g2_decap_8
XFILLER_21_137 VPWR VGND sg13g2_fill_2
XFILLER_21_148 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0827_ VGND VPWR u_ppwm_u_ex__0782_/Y u_ppwm_u_ex__0826_/Y u_ppwm_u_ex__0827_/Y
+ net358 sg13g2_a21oi_1
XFILLER_30_693 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0758_ u_ppwm_u_ex__0758_/A hold259/A u_ppwm_u_ex__0760_/C VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_ex__0689_ net381 net385 u_ppwm_u_ex__0983_/B VPWR VGND sg13g2_nor2_1
XFILLER_26_911 VPWR VGND sg13g2_decap_8
XFILLER_38_760 VPWR VGND sg13g2_decap_8
XFILLER_13_605 VPWR VGND sg13g2_decap_8
XFILLER_26_988 VPWR VGND sg13g2_decap_8
XFILLER_41_936 VPWR VGND sg13g2_decap_8
XFILLER_25_498 VPWR VGND sg13g2_decap_8
XFILLER_40_446 VPWR VGND sg13g2_decap_8
XFILLER_5_815 VPWR VGND sg13g2_decap_8
XFILLER_4_303 VPWR VGND sg13g2_decap_8
XFILLER_48_502 VPWR VGND sg13g2_decap_8
XFILLER_0_586 VPWR VGND sg13g2_decap_8
XFILLER_48_579 VPWR VGND sg13g2_decap_8
XFILLER_17_922 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1040_ net500 VPWR u_ppwm_u_mem__1040_/Y VGND net405 hold59/A sg13g2_o21ai_1
XFILLER_28_281 VPWR VGND sg13g2_decap_8
XFILLER_44_785 VPWR VGND sg13g2_decap_8
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_31_457 VPWR VGND sg13g2_fill_2
XFILLER_32_969 VPWR VGND sg13g2_decap_8
XFILLER_12_671 VPWR VGND sg13g2_decap_8
XFILLER_8_653 VPWR VGND sg13g2_decap_8
Xhold108 hold108/A VPWR VGND net306 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0612_ u_ppwm_u_ex__0612_/B net483 u_ppwm_u_ex__0613_/B VPWR VGND sg13g2_xor2_1
Xu_ppwm_u_mem__0824_ VGND VPWR net396 u_ppwm_u_mem__0823_/X u_ppwm_u_mem__0825_/B
+ net393 sg13g2_a21oi_1
Xhold119 hold119/A VPWR VGND net317 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0755_ VGND VPWR net473 u_ppwm_u_mem__0752_/X u_ppwm_u_mem__0755_/Y
+ net393 sg13g2_a21oi_1
Xu_ppwm_u_mem__0686_ VPWR u_ppwm_u_mem__0686_/Y net335 VGND sg13g2_inv_1
XFILLER_39_535 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1026_ net373 net449 u_ppwm_u_ex__1054_/A VPWR VGND sg13g2_xor2_1
Xu_ppwm_u_mem__1169_ net139 VGND VPWR net268 hold224/A clknet_5_15__leaf_clk sg13g2_dfrbpq_2
XFILLER_35_752 VPWR VGND sg13g2_decap_8
XFILLER_23_958 VPWR VGND sg13g2_decap_8
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
XFILLER_10_619 VPWR VGND sg13g2_decap_8
XFILLER_22_479 VPWR VGND sg13g2_decap_8
XFILLER_2_807 VPWR VGND sg13g2_decap_8
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
XFILLER_18_708 VPWR VGND sg13g2_decap_8
XFILLER_45_527 VPWR VGND sg13g2_decap_8
XFILLER_17_207 VPWR VGND sg13g2_fill_1
XFILLER_41_733 VPWR VGND sg13g2_decap_8
XFILLER_14_958 VPWR VGND sg13g2_decap_8
XFILLER_26_785 VPWR VGND sg13g2_decap_8
XFILLER_25_295 VPWR VGND sg13g2_fill_1
XFILLER_43_87 VPWR VGND sg13g2_decap_4
XFILLER_5_612 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__233__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_5_689 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_49_844 VPWR VGND sg13g2_decap_8
XFILLER_0_383 VPWR VGND sg13g2_decap_8
XFILLER_48_376 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1023_ VGND VPWR net409 u_ppwm_u_mem__0643_/Y u_ppwm_u_mem__1188_/D
+ u_ppwm_u_mem__1022_/Y sg13g2_a21oi_1
XFILLER_16_240 VPWR VGND sg13g2_decap_8
XFILLER_44_582 VPWR VGND sg13g2_decap_8
XFILLER_17_796 VPWR VGND sg13g2_decap_8
XFILLER_32_766 VPWR VGND sg13g2_decap_8
XFILLER_20_928 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0807_ net397 u_ppwm_u_mem__0708_/Y u_ppwm_u_mem__0722_/Y u_ppwm_u_mem__0701_/Y
+ u_ppwm_u_mem__0715_/Y net485 u_ppwm_u_mem__0807_/X VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0738_ u_ppwm_u_mem__0731_/Y net625 u_ppwm_u_mem__0737_/Y hold258/A
+ VPWR VGND sg13g2_a21o_1
Xfanout429 net431 net429 VPWR VGND sg13g2_buf_8
Xfanout407 net408 net407 VPWR VGND sg13g2_buf_8
Xfanout418 net421 net418 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0669_ VPWR u_ppwm_u_mem__0669_/Y net286 VGND sg13g2_inv_1
Xu_ppwm_u_ex__1009_ u_ppwm_u_ex__1010_/B net355 net440 net362 hold312/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_22_243 VPWR VGND sg13g2_fill_2
XFILLER_23_755 VPWR VGND sg13g2_decap_8
XFILLER_11_917 VPWR VGND sg13g2_decap_8
XFILLER_13_13 VPWR VGND sg13g2_fill_1
XFILLER_13_68 VPWR VGND sg13g2_decap_4
XFILLER_2_604 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_46_825 VPWR VGND sg13g2_decap_8
XFILLER_18_505 VPWR VGND sg13g2_decap_8
XFILLER_26_582 VPWR VGND sg13g2_decap_8
XFILLER_41_530 VPWR VGND sg13g2_decap_8
XFILLER_14_755 VPWR VGND sg13g2_decap_8
XFILLER_9_225 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1129__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_9_247 VPWR VGND sg13g2_fill_1
XFILLER_6_954 VPWR VGND sg13g2_decap_8
XFILLER_10_983 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__193_ hold165/A hold283/A u_ppwm_u_pwm__202_/B VPWR VGND sg13g2_nor2b_1
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_decap_8
XFILLER_49_641 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_191 VPWR VGND sg13g2_fill_2
XFILLER_48_173 VPWR VGND sg13g2_decap_8
XFILLER_37_836 VPWR VGND sg13g2_decap_8
XFILLER_45_891 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1006_ net497 VPWR u_ppwm_u_mem__1006_/Y VGND net412 net234 sg13g2_o21ai_1
XFILLER_17_593 VPWR VGND sg13g2_decap_8
XFILLER_20_725 VPWR VGND sg13g2_decap_8
XFILLER_32_563 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_313 VPWR VGND sg13g2_fill_2
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_43_839 VPWR VGND sg13g2_decap_8
XFILLER_11_714 VPWR VGND sg13g2_decap_8
XFILLER_23_552 VPWR VGND sg13g2_decap_8
XFILLER_6_206 VPWR VGND sg13g2_fill_1
XFILLER_2_401 VPWR VGND sg13g2_decap_8
XFILLER_3_968 VPWR VGND sg13g2_decap_8
Xhold280 hold280/A VPWR VGND net648 sg13g2_dlygate4sd3_1
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_2_478 VPWR VGND sg13g2_decap_8
Xhold291 hold291/A VPWR VGND net659 sg13g2_dlygate4sd3_1
XFILLER_46_622 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_869 VPWR VGND sg13g2_decap_8
XFILLER_46_699 VPWR VGND sg13g2_decap_8
XFILLER_18_379 VPWR VGND sg13g2_decap_4
XFILLER_33_316 VPWR VGND sg13g2_decap_4
XFILLER_34_828 VPWR VGND sg13g2_decap_8
XFILLER_14_552 VPWR VGND sg13g2_decap_8
XFILLER_42_894 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0860_ net508 VPWR u_ppwm_u_ex__0861_/A VGND net463 net354 sg13g2_o21ai_1
Xu_ppwm_u_ex__0791_ VGND VPWR u_ppwm_u_ex__0791_/X net386 net464 sg13g2_or2_1
Xu_ppwm_u_pwm__245_ net188 VGND VPWR net548 hold178/A clknet_5_1__leaf_clk sg13g2_dfrbpq_2
XFILLER_10_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__176_ u_ppwm_u_pwm__188_/A net602 u_ppwm_u_pwm__180_/C hold235/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_6_751 VPWR VGND sg13g2_decap_8
XFILLER_37_633 VPWR VGND sg13g2_decap_8
XFILLER_25_806 VPWR VGND sg13g2_decap_8
XFILLER_24_327 VPWR VGND sg13g2_fill_1
XFILLER_33_883 VPWR VGND sg13g2_decap_8
XFILLER_20_522 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0989_ u_ppwm_u_ex__0989_/B net350 u_ppwm_u_ex__0989_/A u_ppwm_u_ex__0989_/Y
+ VPWR VGND u_ppwm_u_ex__0989_/D sg13g2_nand4_1
XFILLER_20_599 VPWR VGND sg13g2_decap_8
XFILLER_27_132 VPWR VGND sg13g2_decap_8
XFILLER_28_666 VPWR VGND sg13g2_decap_8
XFILLER_16_839 VPWR VGND sg13g2_decap_8
XFILLER_43_636 VPWR VGND sg13g2_decap_8
XFILLER_24_850 VPWR VGND sg13g2_decap_8
XFILLER_11_511 VPWR VGND sg13g2_decap_8
XFILLER_11_588 VPWR VGND sg13g2_decap_8
XFILLER_13_1011 VPWR VGND sg13g2_decap_8
XFILLER_3_765 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1172__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_47_942 VPWR VGND sg13g2_decap_8
XFILLER_18_8 VPWR VGND sg13g2_fill_2
XFILLER_19_666 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_34_625 VPWR VGND sg13g2_decap_8
XFILLER_46_496 VPWR VGND sg13g2_decap_8
XFILLER_18_198 VPWR VGND sg13g2_fill_1
XFILLER_42_691 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0912_ u_ppwm_u_ex__0913_/B net365 hold254/A net367 hold259/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_15_894 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0843_ u_ppwm_u_ex__0843_/A u_ppwm_u_ex__0843_/B u_ppwm_u_ex__0867_/A
+ u_ppwm_u_ex__0843_/Y VPWR VGND sg13g2_nor3_1
XFILLER_30_875 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0986_ net503 VPWR u_ppwm_u_mem__0986_/Y VGND net420 hold69/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__228_ net190 VGND VPWR net200 hold1/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__0774_ VGND VPWR u_ppwm_u_ex__0578_/Y u_ppwm_u_ex__0772_/Y hold50/A u_ppwm_u_ex__0773_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1220__117 VPWR VGND net117 sg13g2_tiehi
Xu_ppwm_u_pwm__159_ net490 VPWR u_ppwm_u_pwm__159_/Y VGND net454 net391 sg13g2_o21ai_1
XFILLER_37_0 VPWR VGND sg13g2_fill_2
XFILLER_38_942 VPWR VGND sg13g2_decap_8
XFILLER_37_441 VPWR VGND sg13g2_fill_1
XFILLER_25_603 VPWR VGND sg13g2_decap_8
XFILLER_24_113 VPWR VGND sg13g2_decap_4
XFILLER_40_628 VPWR VGND sg13g2_decap_8
XFILLER_21_820 VPWR VGND sg13g2_decap_8
XFILLER_33_680 VPWR VGND sg13g2_decap_8
XFILLER_20_352 VPWR VGND sg13g2_decap_8
XFILLER_20_374 VPWR VGND sg13g2_fill_1
XFILLER_21_897 VPWR VGND sg13g2_decap_8
XFILLER_0_768 VPWR VGND sg13g2_decap_8
XFILLER_29_931 VPWR VGND sg13g2_decap_8
XFILLER_47_249 VPWR VGND sg13g2_decap_8
XFILLER_46_32 VPWR VGND sg13g2_fill_2
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_76 VPWR VGND sg13g2_fill_1
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_43_433 VPWR VGND sg13g2_decap_8
XFILLER_16_636 VPWR VGND sg13g2_decap_8
XFILLER_28_496 VPWR VGND sg13g2_fill_1
XFILLER_30_116 VPWR VGND sg13g2_fill_1
XFILLER_31_639 VPWR VGND sg13g2_decap_8
XFILLER_12_853 VPWR VGND sg13g2_decap_8
XFILLER_8_835 VPWR VGND sg13g2_decap_8
XFILLER_7_15 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0840_ hold79/A hold164/A net485 u_ppwm_u_mem__0840_/X VPWR VGND sg13g2_mux2_1
XFILLER_11_385 VPWR VGND sg13g2_decap_4
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0771_ u_ppwm_u_mem__0771_/Y hold100/A net484 VPWR VGND sg13g2_nand2_1
XFILLER_3_562 VPWR VGND sg13g2_decap_8
XFILLER_39_717 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__100_ net439 net645 u_ppwm_u_global_counter__103_/D VPWR
+ VGND sg13g2_and2_1
Xu_ppwm_u_ex__1111_ net29 VGND VPWR u_ppwm_u_ex__1111_/D hold309/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_38_227 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1042_ u_ppwm_u_ex__1041_/Y VPWR u_ppwm_u_ex__1046_/C VGND u_ppwm_u_ex__1038_/Y
+ u_ppwm_u_ex__1040_/Y sg13g2_o21ai_1
XFILLER_19_463 VPWR VGND sg13g2_decap_8
XFILLER_46_293 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1185_ net75 VGND VPWR net250 hold124/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_433 VPWR VGND sg13g2_decap_4
XFILLER_35_934 VPWR VGND sg13g2_decap_8
XFILLER_15_691 VPWR VGND sg13g2_decap_8
XFILLER_30_672 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0826_ u_ppwm_u_ex__0826_/Y net464 net379 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__0969_ VGND VPWR net420 u_ppwm_u_mem__0670_/Y u_ppwm_u_mem__1161_/D
+ u_ppwm_u_mem__0968_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0757_ u_ppwm_u_ex__0757_/A hold262/A u_ppwm_u_ex__0761_/C VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_ex__0688_ u_ppwm_u_ex__0688_/A u_ppwm_u_ex__0688_/B u_ppwm_u_ex__0688_/C
+ u_ppwm_u_ex__0688_/Y VPWR VGND sg13g2_nor3_1
XFILLER_45_709 VPWR VGND sg13g2_decap_8
XFILLER_26_967 VPWR VGND sg13g2_decap_8
XFILLER_41_915 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_fill_2
XFILLER_21_694 VPWR VGND sg13g2_decap_8
XFILLER_10_1025 VPWR VGND sg13g2_decap_4
XFILLER_0_565 VPWR VGND sg13g2_decap_8
XFILLER_48_558 VPWR VGND sg13g2_decap_8
XFILLER_17_901 VPWR VGND sg13g2_decap_8
XFILLER_28_271 VPWR VGND sg13g2_decap_4
XFILLER_44_764 VPWR VGND sg13g2_decap_8
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_43_285 VPWR VGND sg13g2_fill_1
XFILLER_32_948 VPWR VGND sg13g2_decap_8
XFILLER_12_650 VPWR VGND sg13g2_decap_8
XFILLER_40_992 VPWR VGND sg13g2_decap_8
XFILLER_8_632 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0611_ net446 VPWR u_ppwm_u_ex__0612_/B VGND net385 u_ppwm_u_ex__0636_/B
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0823_ hold191/A hold137/A net481 u_ppwm_u_mem__0823_/X VPWR VGND sg13g2_mux2_1
XFILLER_7_186 VPWR VGND sg13g2_fill_2
Xhold109 hold109/A VPWR VGND net307 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0754_ u_ppwm_u_mem__0754_/Y net397 u_ppwm_u_mem__0754_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0685_ VPWR u_ppwm_u_mem__0685_/Y net273 VGND sg13g2_inv_1
XFILLER_39_514 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1025_ u_ppwm_u_ex__1025_/A u_ppwm_u_ex__1049_/B u_ppwm_u_ex__1025_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_35_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1168_ net143 VGND VPWR u_ppwm_u_mem__1168_/D hold108/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_23_937 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1099_ u_ppwm_u_mem__1101_/B net618 net606 u_ppwm_u_mem__1102_/D VPWR
+ VGND sg13g2_and3_1
XFILLER_22_458 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0809_ net506 VPWR u_ppwm_u_ex__0809_/Y VGND net466 net354 sg13g2_o21ai_1
XFILLER_45_506 VPWR VGND sg13g2_decap_8
XFILLER_27_56 VPWR VGND sg13g2_fill_1
XFILLER_26_764 VPWR VGND sg13g2_decap_8
XFILLER_41_712 VPWR VGND sg13g2_decap_8
XFILLER_14_937 VPWR VGND sg13g2_decap_8
XFILLER_41_789 VPWR VGND sg13g2_decap_8
XFILLER_21_491 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_decap_8
XFILLER_49_823 VPWR VGND sg13g2_decap_8
XFILLER_0_362 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_48_355 VPWR VGND sg13g2_decap_8
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1022_ net496 VPWR u_ppwm_u_mem__1022_/Y VGND net409 net319 sg13g2_o21ai_1
XFILLER_44_561 VPWR VGND sg13g2_decap_8
XFILLER_17_775 VPWR VGND sg13g2_decap_8
XFILLER_20_907 VPWR VGND sg13g2_decap_8
XFILLER_32_745 VPWR VGND sg13g2_decap_8
XFILLER_9_985 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0806_ u_ppwm_u_mem__0805_/Y VPWR u_ppwm_u_mem__0806_/Y VGND net473
+ u_ppwm_u_mem__0803_/X sg13g2_o21ai_1
Xu_ppwm_u_mem__0737_ net618 u_ppwm_u_mem__0737_/B u_ppwm_u_mem__0737_/C u_ppwm_u_mem__0737_/D
+ u_ppwm_u_mem__0737_/Y VPWR VGND sg13g2_nor4_1
Xu_ppwm_u_mem__0668_ VPWR u_ppwm_u_mem__0668_/Y net531 VGND sg13g2_inv_1
Xfanout419 net420 net419 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_pwm__249__198 VPWR VGND net198 sg13g2_tiehi
Xfanout408 net422 net408 VPWR VGND sg13g2_buf_1
XFILLER_27_506 VPWR VGND sg13g2_decap_4
XFILLER_42_509 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1008_ u_ppwm_u_ex__1010_/A net443 fanout356/A VPWR VGND sg13g2_nand2_1
XFILLER_23_734 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_4
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_46_804 VPWR VGND sg13g2_decap_8
XFILLER_26_561 VPWR VGND sg13g2_decap_8
XFILLER_14_734 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1168__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_41_586 VPWR VGND sg13g2_decap_8
XFILLER_13_288 VPWR VGND sg13g2_decap_4
XFILLER_10_962 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__192_ hold5/A hold204/A u_ppwm_u_pwm__202_/A VPWR VGND sg13g2_nor2b_1
XFILLER_6_933 VPWR VGND sg13g2_decap_8
XFILLER_5_465 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_37_815 VPWR VGND sg13g2_decap_8
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_45_870 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1005_ VGND VPWR net412 u_ppwm_u_mem__0652_/Y hold37/A u_ppwm_u_mem__1004_/Y
+ sg13g2_a21oi_1
XFILLER_17_572 VPWR VGND sg13g2_decap_8
XFILLER_32_542 VPWR VGND sg13g2_decap_8
XFILLER_20_704 VPWR VGND sg13g2_decap_8
XFILLER_9_782 VPWR VGND sg13g2_decap_8
XFILLER_8_292 VPWR VGND sg13g2_decap_4
XFILLER_39_152 VPWR VGND sg13g2_fill_2
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_43_818 VPWR VGND sg13g2_decap_8
XFILLER_15_509 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1142__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_23_531 VPWR VGND sg13g2_decap_8
XFILLER_10_225 VPWR VGND sg13g2_decap_4
XFILLER_24_79 VPWR VGND sg13g2_fill_1
XFILLER_40_89 VPWR VGND sg13g2_decap_4
XFILLER_3_947 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_2_457 VPWR VGND sg13g2_decap_8
Xhold270 hold323/A VPWR VGND net638 sg13g2_dlygate4sd3_1
Xhold281 hold281/A VPWR VGND net649 sg13g2_dlygate4sd3_1
Xhold292 hold292/A VPWR VGND net660 sg13g2_dlygate4sd3_1
XFILLER_46_601 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_848 VPWR VGND sg13g2_decap_8
XFILLER_18_358 VPWR VGND sg13g2_decap_8
XFILLER_34_807 VPWR VGND sg13g2_decap_8
XFILLER_46_678 VPWR VGND sg13g2_decap_8
XFILLER_14_531 VPWR VGND sg13g2_decap_8
XFILLER_42_873 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0790_ u_ppwm_u_ex__0843_/A u_ppwm_u_ex__0789_/Y u_ppwm_u_ex__0790_/Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_6_730 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__244_ net192 VGND VPWR u_ppwm_u_pwm__244_/D hold268/A clknet_5_1__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__175_ u_ppwm_u_pwm__180_/C net601 net652 u_ppwm_u_pwm__175_/C VPWR VGND
+ sg13g2_and3_2
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_49_494 VPWR VGND sg13g2_decap_8
XFILLER_37_612 VPWR VGND sg13g2_decap_8
XFILLER_37_689 VPWR VGND sg13g2_decap_8
XFILLER_33_862 VPWR VGND sg13g2_decap_8
XFILLER_20_501 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0988_ u_ppwm_u_ex__0989_/D u_ppwm_u_ex__0987_/X u_ppwm_u_ex__0780_/X
+ u_ppwm_u_ex__0856_/B net383 VPWR VGND sg13g2_a22oi_1
XFILLER_32_394 VPWR VGND sg13g2_decap_4
XFILLER_20_578 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_fill_1
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_43_615 VPWR VGND sg13g2_decap_8
XFILLER_16_818 VPWR VGND sg13g2_decap_8
XFILLER_11_567 VPWR VGND sg13g2_decap_8
XFILLER_7_549 VPWR VGND sg13g2_decap_8
XFILLER_3_744 VPWR VGND sg13g2_decap_8
XFILLER_47_921 VPWR VGND sg13g2_decap_8
XFILLER_19_645 VPWR VGND sg13g2_decap_8
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1213__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_47_998 VPWR VGND sg13g2_decap_8
XFILLER_46_475 VPWR VGND sg13g2_decap_8
XFILLER_34_604 VPWR VGND sg13g2_decap_8
XFILLER_33_125 VPWR VGND sg13g2_decap_8
XFILLER_15_873 VPWR VGND sg13g2_decap_8
XFILLER_21_309 VPWR VGND sg13g2_fill_1
XFILLER_42_670 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0911_ VPWR VGND u_ppwm_u_ex__0797_/Y u_ppwm_u_ex__0907_/Y u_ppwm_u_ex__0910_/X
+ u_ppwm_u_ex__0790_/Y u_ppwm_u_ex__1046_/A u_ppwm_u_ex__0871_/X sg13g2_a221oi_1
Xu_ppwm_u_ex__0842_ u_ppwm_u_ex__0867_/A net381 u_ppwm_u_ex__0842_/B VPWR VGND sg13g2_nand2_1
XFILLER_30_854 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0985_ VGND VPWR net415 u_ppwm_u_mem__0662_/Y hold70/A u_ppwm_u_mem__0984_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__227_ u_ppwm_u_pwm__249_/D net489 u_ppwm_u_pwm__227_/B u_ppwm_u_pwm__227_/C
+ VPWR VGND sg13g2_and3_1
Xu_ppwm_u_ex__0773_ net492 VPWR u_ppwm_u_ex__0773_/Y VGND net384 u_ppwm_u_ex__0772_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_pwm__158_ VGND VPWR u_ppwm_u_pwm__218_/B net389 hold41/A u_ppwm_u_pwm__157_/Y
+ sg13g2_a21oi_1
XFILLER_38_921 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_38_998 VPWR VGND sg13g2_decap_8
XFILLER_25_659 VPWR VGND sg13g2_decap_8
XFILLER_40_607 VPWR VGND sg13g2_decap_8
XFILLER_36_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_876 VPWR VGND sg13g2_decap_8
XFILLER_4_519 VPWR VGND sg13g2_decap_8
XFILLER_21_47 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1100__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_0_747 VPWR VGND sg13g2_decap_8
XFILLER_47_228 VPWR VGND sg13g2_decap_8
XFILLER_29_910 VPWR VGND sg13g2_decap_8
XFILLER_16_615 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_decap_8
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_43_412 VPWR VGND sg13g2_decap_8
XFILLER_31_618 VPWR VGND sg13g2_decap_8
XFILLER_43_489 VPWR VGND sg13g2_decap_8
XFILLER_8_814 VPWR VGND sg13g2_decap_8
XFILLER_12_832 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0770_ u_ppwm_u_mem__0769_/Y VPWR u_ppwm_u_mem__0770_/Y VGND u_ppwm_u_mem__0710_/Y
+ net484 sg13g2_o21ai_1
XFILLER_3_541 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_ex__1110_ net31 VGND VPWR net670 hold301/A clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_217 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1041_ VGND VPWR u_ppwm_u_ex__1038_/Y u_ppwm_u_ex__1040_/Y u_ppwm_u_ex__1041_/Y
+ net358 sg13g2_a21oi_1
XFILLER_35_913 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1184_ net79 VGND VPWR net323 hold215/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_795 VPWR VGND sg13g2_decap_8
XFILLER_46_272 VPWR VGND sg13g2_decap_8
XFILLER_15_670 VPWR VGND sg13g2_decap_8
XFILLER_14_180 VPWR VGND sg13g2_fill_2
XFILLER_30_651 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0825_ u_ppwm_u_ex__0825_/Y net464 net379 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0968_ net502 VPWR u_ppwm_u_mem__0968_/Y VGND net420 net271 sg13g2_o21ai_1
Xu_ppwm_u_ex__0756_ VPWR VGND u_ppwm_u_ex__0754_/Y u_ppwm_u_ex__0755_/Y u_ppwm_u_ex__0752_/Y
+ u_ppwm_u_ex__0758_/A u_ppwm_u_ex__0760_/A hold259/A sg13g2_a221oi_1
Xu_ppwm_u_mem__0899_ VGND VPWR net435 u_ppwm_u_mem__0705_/Y hold134/A u_ppwm_u_mem__0898_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0687_ u_ppwm_u_ex__0686_/Y VPWR u_ppwm_u_ex__0688_/C VGND u_ppwm_u_ex__0757_/A
+ hold277/A sg13g2_o21ai_1
XFILLER_16_25 VPWR VGND sg13g2_decap_4
XFILLER_25_401 VPWR VGND sg13g2_fill_1
XFILLER_25_412 VPWR VGND sg13g2_fill_2
XFILLER_26_946 VPWR VGND sg13g2_decap_8
XFILLER_38_795 VPWR VGND sg13g2_decap_8
XFILLER_12_139 VPWR VGND sg13g2_fill_1
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_10_1004 VPWR VGND sg13g2_decap_8
XFILLER_0_544 VPWR VGND sg13g2_decap_8
XFILLER_48_537 VPWR VGND sg13g2_decap_8
XFILLER_28_250 VPWR VGND sg13g2_decap_8
XFILLER_17_957 VPWR VGND sg13g2_decap_8
XFILLER_29_784 VPWR VGND sg13g2_decap_8
XFILLER_44_743 VPWR VGND sg13g2_decap_8
XFILLER_16_489 VPWR VGND sg13g2_decap_8
XFILLER_32_927 VPWR VGND sg13g2_decap_8
XFILLER_40_971 VPWR VGND sg13g2_decap_8
XFILLER_8_611 VPWR VGND sg13g2_decap_8
XFILLER_8_688 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0610_ u_ppwm/instr\[0\] u_ppwm_u_ex__0610_/C fanout388/A u_ppwm_u_ex__0636_/B
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__0822_ VGND VPWR u_ppwm_u_mem__0672_/Y net482 u_ppwm_u_mem__0822_/Y
+ u_ppwm_u_mem__0821_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0753_ hold90/A hold177/A net483 u_ppwm_u_mem__0754_/B VPWR VGND sg13g2_mux2_1
XFILLER_4_883 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0684_ VPWR u_ppwm_u_mem__0684_/Y net596 VGND sg13g2_inv_1
XFILLER_21_4 VPWR VGND sg13g2_fill_2
XFILLER_47_592 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1024_ VGND VPWR u_ppwm_u_ex__0877_/C u_ppwm_u_ex__1022_/Y u_ppwm_u_ex__1118_/D
+ u_ppwm_u_ex__1023_/Y sg13g2_a21oi_1
XFILLER_35_710 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1167_ net147 VGND VPWR u_ppwm_u_mem__1167_/D hold66/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_23_916 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1098_ net618 u_ppwm_u_mem__1098_/B u_ppwm_u_mem__1100_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_35_787 VPWR VGND sg13g2_decap_8
XFILLER_22_437 VPWR VGND sg13g2_decap_8
XFILLER_31_982 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0808_ u_ppwm_u_ex__0989_/A net354 u_ppwm_u_ex__0808_/X VPWR VGND sg13g2_and2_1
Xu_ppwm_u_ex__0739_ u_ppwm_u_ex__0739_/Y u_ppwm_u_ex__0739_/A u_ppwm_u_ex__0739_/B
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_592 VPWR VGND sg13g2_decap_8
XFILLER_26_743 VPWR VGND sg13g2_decap_8
XFILLER_14_916 VPWR VGND sg13g2_decap_8
XFILLER_41_768 VPWR VGND sg13g2_decap_8
XFILLER_40_278 VPWR VGND sg13g2_fill_1
XFILLER_21_470 VPWR VGND sg13g2_decap_8
XFILLER_5_647 VPWR VGND sg13g2_decap_8
XFILLER_4_168 VPWR VGND sg13g2_fill_2
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_0_341 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_48_334 VPWR VGND sg13g2_decap_8
XFILLER_49_879 VPWR VGND sg13g2_decap_8
XFILLER_29_581 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_decap_8
XFILLER_44_540 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1021_ VGND VPWR net412 u_ppwm_u_mem__0644_/Y u_ppwm_u_mem__1187_/D
+ u_ppwm_u_mem__1020_/Y sg13g2_a21oi_1
XFILLER_17_754 VPWR VGND sg13g2_decap_8
XFILLER_32_724 VPWR VGND sg13g2_decap_8
XFILLER_9_964 VPWR VGND sg13g2_decap_8
XFILLER_8_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0805_ VGND VPWR net473 u_ppwm_u_mem__0804_/X u_ppwm_u_mem__0805_/Y
+ net393 sg13g2_a21oi_1
XFILLER_4_680 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0736_ u_ppwm_u_mem__0737_/D net400 net488 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0667_ VPWR u_ppwm_u_mem__0667_/Y net315 VGND sg13g2_inv_1
Xfanout409 net410 net409 VPWR VGND sg13g2_buf_2
XFILLER_3_190 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1139__84 VPWR VGND net84 sg13g2_tiehi
XFILLER_39_334 VPWR VGND sg13g2_fill_1
XFILLER_27_529 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1007_ VGND VPWR u_ppwm_u_ex__1006_/A u_ppwm_u_ex__1027_/A u_ppwm_u_ex__1007_/Y
+ net358 sg13g2_a21oi_1
Xu_ppwm_u_mem__1219_ net148 VGND VPWR u_ppwm_u_mem__1219_/D hold256/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_22_201 VPWR VGND sg13g2_decap_8
XFILLER_23_713 VPWR VGND sg13g2_decap_8
XFILLER_35_584 VPWR VGND sg13g2_decap_8
XFILLER_22_256 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__232__181 VPWR VGND net181 sg13g2_tiehi
Xu_ppwm_u_mem__1224__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_2_639 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_38_34 VPWR VGND sg13g2_fill_2
XFILLER_45_359 VPWR VGND sg13g2_decap_8
XFILLER_26_540 VPWR VGND sg13g2_decap_8
XFILLER_14_713 VPWR VGND sg13g2_decap_8
XFILLER_13_201 VPWR VGND sg13g2_decap_4
XFILLER_13_234 VPWR VGND sg13g2_decap_4
XFILLER_41_565 VPWR VGND sg13g2_decap_8
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
XFILLER_6_912 VPWR VGND sg13g2_decap_8
XFILLER_10_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__191_ net594 u_ppwm_u_pwm__191_/B u_ppwm_u_pwm__191_/C hold227/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_6_989 VPWR VGND sg13g2_decap_8
XFILLER_5_444 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1175__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_23_1014 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_decap_8
XFILLER_0_193 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1004_ net499 VPWR u_ppwm_u_mem__1004_/Y VGND net414 hold57/A sg13g2_o21ai_1
XFILLER_17_551 VPWR VGND sg13g2_decap_8
XFILLER_32_598 VPWR VGND sg13g2_decap_8
XFILLER_9_761 VPWR VGND sg13g2_decap_8
XFILLER_5_82 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0719_ VPWR u_ppwm_u_mem__0719_/Y net560 VGND sg13g2_inv_1
XFILLER_27_315 VPWR VGND sg13g2_fill_1
XFILLER_28_827 VPWR VGND sg13g2_decap_8
XFILLER_39_164 VPWR VGND sg13g2_fill_1
XFILLER_39_197 VPWR VGND sg13g2_fill_1
XFILLER_23_510 VPWR VGND sg13g2_decap_8
XFILLER_36_893 VPWR VGND sg13g2_decap_8
XFILLER_11_749 VPWR VGND sg13g2_decap_8
XFILLER_23_587 VPWR VGND sg13g2_decap_8
XFILLER_6_219 VPWR VGND sg13g2_decap_4
XFILLER_3_926 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1198__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_46_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_436 VPWR VGND sg13g2_decap_8
Xhold260 hold260/A VPWR VGND net628 sg13g2_dlygate4sd3_1
Xhold271 hold271/A VPWR VGND net639 sg13g2_dlygate4sd3_1
Xhold282 hold282/A VPWR VGND net650 sg13g2_dlygate4sd3_1
Xhold293 hold293/A VPWR VGND net661 sg13g2_dlygate4sd3_1
XFILLER_49_88 VPWR VGND sg13g2_decap_4
XFILLER_19_827 VPWR VGND sg13g2_decap_8
XFILLER_46_657 VPWR VGND sg13g2_decap_8
XFILLER_33_307 VPWR VGND sg13g2_fill_2
XFILLER_14_510 VPWR VGND sg13g2_decap_8
XFILLER_27_893 VPWR VGND sg13g2_decap_8
XFILLER_42_852 VPWR VGND sg13g2_decap_8
XFILLER_14_587 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__243_ net196 VGND VPWR net603 hold233/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__174_ VGND VPWR hold284/A u_ppwm_u_pwm__175_/C hold234/A net601 sg13g2_a21oi_1
XFILLER_6_786 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_fill_2
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
XFILLER_37_668 VPWR VGND sg13g2_decap_8
XFILLER_36_145 VPWR VGND sg13g2_fill_2
XFILLER_33_841 VPWR VGND sg13g2_decap_8
XFILLER_20_557 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0987_ fanout383/A hold292/A u_ppwm_u_ex__0987_/X VPWR VGND sg13g2_xor2_1
XFILLER_0_929 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1158__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_28_624 VPWR VGND sg13g2_decap_8
XFILLER_36_690 VPWR VGND sg13g2_decap_8
XFILLER_24_885 VPWR VGND sg13g2_decap_8
XFILLER_11_546 VPWR VGND sg13g2_decap_8
XFILLER_7_528 VPWR VGND sg13g2_decap_8
XFILLER_3_723 VPWR VGND sg13g2_decap_8
XFILLER_47_900 VPWR VGND sg13g2_decap_8
XFILLER_19_624 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_977 VPWR VGND sg13g2_decap_8
XFILLER_46_454 VPWR VGND sg13g2_decap_8
XFILLER_27_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0910_ u_ppwm_u_ex__0892_/Y u_ppwm_u_ex__0928_/B net377 u_ppwm_u_ex__0910_/X
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_852 VPWR VGND sg13g2_decap_8
XFILLER_14_373 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0841_ u_ppwm_u_ex__0843_/B u_ppwm_u_ex__0840_/Y u_ppwm_u_ex__0816_/B
+ u_ppwm_u_ex__0839_/Y u_ppwm_u_ex__0795_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_30_833 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0984_ net498 VPWR u_ppwm_u_mem__0984_/Y VGND net415 hold224/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0772_ net383 u_ppwm_u_ex__0772_/C net446 u_ppwm_u_ex__0772_/Y VPWR VGND
+ net369 sg13g2_nand4_1
Xu_ppwm_u_pwm__226_ net247 u_ppwm_u_pwm__226_/B u_ppwm_u_pwm__226_/C u_ppwm_u_pwm__227_/C
+ VPWR VGND sg13g2_or3_1
Xu_ppwm_u_pwm__157_ net490 VPWR u_ppwm_u_pwm__157_/Y VGND net455 net389 sg13g2_o21ai_1
XFILLER_6_583 VPWR VGND sg13g2_decap_8
XFILLER_37_2 VPWR VGND sg13g2_fill_1
XFILLER_38_900 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_25_638 VPWR VGND sg13g2_decap_8
XFILLER_24_159 VPWR VGND sg13g2_fill_2
XFILLER_21_855 VPWR VGND sg13g2_decap_8
XFILLER_20_343 VPWR VGND sg13g2_decap_4
XFILLER_0_726 VPWR VGND sg13g2_decap_8
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_719 VPWR VGND sg13g2_decap_8
XFILLER_47_207 VPWR VGND sg13g2_decap_8
XFILLER_29_966 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_43_468 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_fill_2
XFILLER_15_159 VPWR VGND sg13g2_decap_8
XFILLER_12_811 VPWR VGND sg13g2_decap_8
XFILLER_24_682 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_fill_2
XFILLER_11_354 VPWR VGND sg13g2_fill_2
XFILLER_12_888 VPWR VGND sg13g2_decap_8
XFILLER_3_520 VPWR VGND sg13g2_decap_8
XFILLER_3_597 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1040_ u_ppwm_u_ex__1040_/Y hold299/A net373 VPWR VGND sg13g2_xnor2_1
XFILLER_47_774 VPWR VGND sg13g2_decap_8
XFILLER_46_251 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1183_ net83 VGND VPWR net584 hold147/A clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_498 VPWR VGND sg13g2_decap_8
XFILLER_35_969 VPWR VGND sg13g2_decap_8
XFILLER_22_619 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0824_ u_ppwm_u_ex__0996_/A net379 u_ppwm_u_ex__0856_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0967_ VGND VPWR net428 u_ppwm_u_mem__0671_/Y hold74/A u_ppwm_u_mem__0966_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0755_ net461 u_ppwm_u_ex__0755_/B u_ppwm_u_ex__0755_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0686_ u_ppwm_u_ex__0686_/Y net454 hold217/A VPWR VGND sg13g2_nand2b_1
XFILLER_7_892 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__209_ u_ppwm_u_pwm__209_/B u_ppwm_u_pwm__209_/C u_ppwm_u_pwm__209_/A
+ u_ppwm_u_pwm__216_/A VPWR VGND u_ppwm_u_pwm__209_/D sg13g2_nand4_1
Xu_ppwm_u_mem__0898_ net511 VPWR u_ppwm_u_mem__0898_/Y VGND net432 hold161/A sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_38_774 VPWR VGND sg13g2_decap_8
XFILLER_26_925 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__089_ u_ppwm_u_global_counter__089_/A hold266/A u_ppwm_u_global_counter__118_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_37_295 VPWR VGND sg13g2_fill_2
XFILLER_40_427 VPWR VGND sg13g2_fill_2
XFILLER_13_619 VPWR VGND sg13g2_decap_8
XFILLER_21_652 VPWR VGND sg13g2_decap_8
XFILLER_5_829 VPWR VGND sg13g2_decap_8
XFILLER_4_317 VPWR VGND sg13g2_fill_2
XFILLER_0_523 VPWR VGND sg13g2_decap_8
XFILLER_48_516 VPWR VGND sg13g2_decap_8
XFILLER_29_763 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1190__55 VPWR VGND net55 sg13g2_tiehi
XFILLER_44_722 VPWR VGND sg13g2_decap_8
XFILLER_17_936 VPWR VGND sg13g2_decap_8
XFILLER_28_295 VPWR VGND sg13g2_fill_2
XFILLER_32_906 VPWR VGND sg13g2_decap_8
XFILLER_44_799 VPWR VGND sg13g2_decap_8
XFILLER_40_950 VPWR VGND sg13g2_decap_8
XFILLER_11_162 VPWR VGND sg13g2_fill_2
XFILLER_12_685 VPWR VGND sg13g2_decap_8
XFILLER_8_667 VPWR VGND sg13g2_decap_8
XFILLER_7_144 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0821_ net474 VPWR u_ppwm_u_mem__0821_/Y VGND hold174/A net482 sg13g2_o21ai_1
XFILLER_7_188 VPWR VGND sg13g2_fill_1
XFILLER_7_177 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0752_ hold188/A hold111/A net486 u_ppwm_u_mem__0752_/X VPWR VGND sg13g2_mux2_1
XFILLER_4_862 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0683_ VPWR u_ppwm_u_mem__0683_/Y net556 VGND sg13g2_inv_1
XFILLER_26_1023 VPWR VGND sg13g2_decap_4
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_39_549 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1023_ net506 VPWR u_ppwm_u_ex__1023_/Y VGND net450 net350 sg13g2_o21ai_1
XFILLER_47_571 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1166_ net149 VGND VPWR u_ppwm_u_mem__1166_/D hold26/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1097_ u_ppwm_u_mem__1103_/A net607 u_ppwm_u_mem__1098_/B u_ppwm_u_mem__1222_/D
+ VPWR VGND sg13g2_nor3_1
XFILLER_31_961 VPWR VGND sg13g2_decap_8
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
XFILLER_8_82 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0807_ u_ppwm_u_ex__0807_/A u_ppwm_u_ex__0803_/X fanout354/A VPWR VGND
+ sg13g2_nor2b_2
Xu_ppwm_u_ex__0738_ VPWR VGND hold294/A u_ppwm_u_ex__0737_/Y u_ppwm_u_ex__0757_/A
+ hold295/A u_ppwm_u_ex__0739_/B u_ppwm_u_ex__0954_/A sg13g2_a221oi_1
Xu_ppwm_u_ex__0669_ u_ppwm_u_ex__0669_/Y net464 u_ppwm_u_ex__0998_/B2 VPWR VGND sg13g2_nand2b_1
XFILLER_26_722 VPWR VGND sg13g2_decap_8
XFILLER_38_571 VPWR VGND sg13g2_decap_8
XFILLER_26_799 VPWR VGND sg13g2_decap_8
XFILLER_41_747 VPWR VGND sg13g2_decap_8
XFILLER_40_235 VPWR VGND sg13g2_decap_4
XFILLER_40_213 VPWR VGND sg13g2_decap_4
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_22_983 VPWR VGND sg13g2_decap_8
XFILLER_5_626 VPWR VGND sg13g2_decap_8
XFILLER_49_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_0_320 VPWR VGND sg13g2_decap_8
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_49_858 VPWR VGND sg13g2_decap_8
XFILLER_48_313 VPWR VGND sg13g2_decap_8
XFILLER_0_397 VPWR VGND sg13g2_decap_8
XFILLER_29_560 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1020_ net496 VPWR u_ppwm_u_mem__1020_/Y VGND net412 net236 sg13g2_o21ai_1
XFILLER_17_733 VPWR VGND sg13g2_decap_8
XFILLER_17_80 VPWR VGND sg13g2_fill_2
XFILLER_32_703 VPWR VGND sg13g2_decap_8
XFILLER_44_596 VPWR VGND sg13g2_decap_8
XFILLER_9_943 VPWR VGND sg13g2_decap_8
XFILLER_13_983 VPWR VGND sg13g2_decap_8
XFILLER_8_442 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0804_ hold80/A hold168/A net482 u_ppwm_u_mem__0804_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0735_ net618 u_ppwm_u_mem__0737_/B u_ppwm_u_mem__0737_/C hold251/A
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__0666_ VPWR u_ppwm_u_mem__0666_/Y net224 VGND sg13g2_inv_1
XFILLER_48_880 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1006_ VGND VPWR u_ppwm_u_ex__1017_/B u_ppwm_u_ex__1027_/A u_ppwm_u_ex__1006_/A
+ sg13g2_or2_1
Xu_ppwm_u_mem__1218_ net164 VGND VPWR u_ppwm_u_mem__1218_/D hold167/A clknet_5_3__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_563 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1149_ net64 VGND VPWR net523 hold188/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_769 VPWR VGND sg13g2_decap_8
XFILLER_2_618 VPWR VGND sg13g2_decap_8
XFILLER_46_839 VPWR VGND sg13g2_decap_8
XFILLER_18_519 VPWR VGND sg13g2_decap_8
XFILLER_45_338 VPWR VGND sg13g2_decap_8
XFILLER_13_213 VPWR VGND sg13g2_decap_8
XFILLER_26_596 VPWR VGND sg13g2_decap_8
XFILLER_41_544 VPWR VGND sg13g2_decap_8
XFILLER_13_257 VPWR VGND sg13g2_decap_8
XFILLER_14_769 VPWR VGND sg13g2_decap_8
XFILLER_16_1000 VPWR VGND sg13g2_decap_8
XFILLER_10_920 VPWR VGND sg13g2_decap_8
XFILLER_22_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__190_ hold284/A hold283/A hold233/A u_ppwm_u_pwm__191_/C VPWR VGND net572
+ sg13g2_nand4_1
XFILLER_10_997 VPWR VGND sg13g2_decap_8
XFILLER_6_968 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_172 VPWR VGND sg13g2_fill_1
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_655 VPWR VGND sg13g2_decap_8
XFILLER_48_187 VPWR VGND sg13g2_decap_8
XFILLER_17_530 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1003_ VGND VPWR net415 u_ppwm_u_mem__0653_/Y hold58/A u_ppwm_u_mem__1002_/Y
+ sg13g2_a21oi_1
XFILLER_44_393 VPWR VGND sg13g2_decap_8
XFILLER_44_360 VPWR VGND sg13g2_fill_1
XFILLER_13_780 VPWR VGND sg13g2_decap_8
XFILLER_20_739 VPWR VGND sg13g2_decap_8
XFILLER_32_577 VPWR VGND sg13g2_decap_8
XFILLER_9_740 VPWR VGND sg13g2_decap_8
XFILLER_12_290 VPWR VGND sg13g2_decap_8
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_272 VPWR VGND sg13g2_decap_4
XFILLER_5_990 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0718_ VPWR u_ppwm_u_mem__0718_/Y net284 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0649_ VPWR u_ppwm_u_mem__0649_/Y net345 VGND sg13g2_inv_1
XFILLER_28_806 VPWR VGND sg13g2_decap_8
XFILLER_39_1011 VPWR VGND sg13g2_decap_8
XFILLER_36_872 VPWR VGND sg13g2_decap_8
XFILLER_23_566 VPWR VGND sg13g2_decap_8
XFILLER_11_728 VPWR VGND sg13g2_decap_8
XFILLER_40_36 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1122__28 VPWR VGND net28 sg13g2_tiehi
XFILLER_3_905 VPWR VGND sg13g2_decap_8
XFILLER_2_415 VPWR VGND sg13g2_decap_8
Xhold261 hold261/A VPWR VGND net629 sg13g2_dlygate4sd3_1
Xhold250 hold250/A VPWR VGND net618 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1205__81 VPWR VGND net81 sg13g2_tiehi
Xhold294 hold294/A VPWR VGND net662 sg13g2_dlygate4sd3_1
Xhold283 hold283/A VPWR VGND net651 sg13g2_dlygate4sd3_1
Xhold272 hold272/A VPWR VGND net640 sg13g2_dlygate4sd3_1
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_19_806 VPWR VGND sg13g2_decap_8
XFILLER_46_636 VPWR VGND sg13g2_decap_8
XFILLER_27_872 VPWR VGND sg13g2_decap_8
XFILLER_42_831 VPWR VGND sg13g2_decap_8
XFILLER_41_341 VPWR VGND sg13g2_decap_4
XFILLER_14_566 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1141__80 VPWR VGND net80 sg13g2_tiehi
Xu_ppwm_u_pwm__242_ net178 VGND VPWR u_ppwm_u_pwm__242_/D hold284/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_10_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__173_ u_ppwm_u_pwm__188_/A u_ppwm_u_pwm__173_/B u_ppwm_u_pwm__242_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_765 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1222__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_2_982 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_37_647 VPWR VGND sg13g2_decap_8
XFILLER_18_883 VPWR VGND sg13g2_decap_8
XFILLER_33_820 VPWR VGND sg13g2_decap_8
XFILLER_33_897 VPWR VGND sg13g2_decap_8
XFILLER_20_536 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0986_ hold292/A net383 u_ppwm_u_ex__0994_/A VPWR VGND sg13g2_and2_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
XFILLER_28_603 VPWR VGND sg13g2_decap_8
XFILLER_23_341 VPWR VGND sg13g2_fill_2
XFILLER_24_864 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_525 VPWR VGND sg13g2_decap_8
XFILLER_23_385 VPWR VGND sg13g2_fill_2
XFILLER_7_507 VPWR VGND sg13g2_decap_8
XFILLER_13_1025 VPWR VGND sg13g2_decap_4
XFILLER_3_702 VPWR VGND sg13g2_decap_8
XFILLER_3_779 VPWR VGND sg13g2_decap_8
XFILLER_19_603 VPWR VGND sg13g2_decap_8
XFILLER_47_956 VPWR VGND sg13g2_decap_8
XFILLER_46_433 VPWR VGND sg13g2_decap_8
XFILLER_15_831 VPWR VGND sg13g2_decap_8
XFILLER_34_639 VPWR VGND sg13g2_decap_8
XFILLER_14_363 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0840_ net375 fanout370/A u_ppwm_u_ex__0840_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0983_ VGND VPWR net409 u_ppwm_u_mem__0663_/Y u_ppwm_u_mem__1168_/D
+ u_ppwm_u_mem__0982_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0771_ VGND VPWR u_ppwm_u_ex__0768_/Y u_ppwm_u_ex__0769_/Y hold282/A
+ net649 sg13g2_a21oi_1
XFILLER_30_889 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__225_ net247 VPWR u_ppwm_u_pwm__227_/B VGND u_ppwm_u_pwm__226_/B u_ppwm_u_pwm__226_/C
+ sg13g2_o21ai_1
XFILLER_6_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__156_ VGND VPWR u_ppwm_u_pwm__128_/Y net391 hold14/A u_ppwm_u_pwm__155_/Y
+ sg13g2_a21oi_1
XFILLER_10_591 VPWR VGND sg13g2_decap_8
XFILLER_44_4 VPWR VGND sg13g2_fill_1
XFILLER_38_956 VPWR VGND sg13g2_decap_8
XFILLER_18_680 VPWR VGND sg13g2_decap_8
XFILLER_25_617 VPWR VGND sg13g2_decap_8
XFILLER_21_834 VPWR VGND sg13g2_decap_8
XFILLER_33_694 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0969_ VGND VPWR u_ppwm_u_ex__0967_/Y u_ppwm_u_ex__0968_/Y u_ppwm_u_ex__0969_/Y
+ net357 sg13g2_a21oi_1
XFILLER_0_705 VPWR VGND sg13g2_decap_8
XFILLER_43_1007 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__229__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_29_945 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_43_447 VPWR VGND sg13g2_decap_8
XFILLER_15_127 VPWR VGND sg13g2_fill_1
XFILLER_24_661 VPWR VGND sg13g2_decap_8
XFILLER_12_867 VPWR VGND sg13g2_decap_8
XFILLER_8_849 VPWR VGND sg13g2_decap_8
XFILLER_3_576 VPWR VGND sg13g2_decap_8
XFILLER_4_1023 VPWR VGND sg13g2_decap_4
Xfanout390 net391 net390 VPWR VGND sg13g2_buf_8
XFILLER_19_411 VPWR VGND sg13g2_decap_8
XFILLER_19_433 VPWR VGND sg13g2_decap_8
XFILLER_47_753 VPWR VGND sg13g2_decap_8
XFILLER_46_230 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1182_ net87 VGND VPWR net346 hold172/A clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_477 VPWR VGND sg13g2_decap_8
XFILLER_35_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0823_ u_ppwm_u_ex__1000_/A u_ppwm_u_ex__0823_/A u_ppwm_u_ex__0823_/B
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_686 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0966_ net511 VPWR u_ppwm_u_mem__0966_/Y VGND net428 hold185/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__208_ u_ppwm_u_pwm__209_/D hold13/A hold178/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_ex__0754_ u_ppwm_u_ex__0754_/Y net443 u_ppwm_u_ex__0753_/Y u_ppwm_u_ex__0755_/B
+ net461 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_ex__0685_ u_ppwm_u_ex__0954_/A hold252/A u_ppwm_u_ex__0688_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_7_871 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0897_ VGND VPWR net436 u_ppwm_u_mem__0706_/Y hold162/A u_ppwm_u_mem__0896_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__139_ hold178/A hold268/A hold233/A hold284/A u_ppwm_u_pwm__140_/C VPWR
+ VGND sg13g2_nor4_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
XFILLER_26_904 VPWR VGND sg13g2_decap_8
XFILLER_38_753 VPWR VGND sg13g2_decap_8
XFILLER_37_285 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_global_counter__088_ net398 net392 net633 hold266/A VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__1099_ net52 VGND VPWR u_ppwm_u_ex__1099_/D fanout487/A clknet_5_24__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_41_929 VPWR VGND sg13g2_decap_8
XFILLER_21_631 VPWR VGND sg13g2_decap_8
XFILLER_20_152 VPWR VGND sg13g2_decap_8
XFILLER_5_808 VPWR VGND sg13g2_decap_8
XFILLER_0_502 VPWR VGND sg13g2_decap_8
XFILLER_0_579 VPWR VGND sg13g2_decap_8
XFILLER_28_241 VPWR VGND sg13g2_decap_4
XFILLER_29_742 VPWR VGND sg13g2_decap_8
XFILLER_44_701 VPWR VGND sg13g2_decap_8
XFILLER_17_915 VPWR VGND sg13g2_decap_8
XFILLER_44_778 VPWR VGND sg13g2_decap_8
XFILLER_25_981 VPWR VGND sg13g2_decap_8
XFILLER_12_664 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0820_ VGND VPWR net397 u_ppwm_u_mem__0819_/X u_ppwm_u_mem__0820_/Y
+ net469 sg13g2_a21oi_1
XFILLER_11_196 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0751_ u_ppwm_u_mem__0751_/Y fanout394/A u_ppwm_u_mem__0750_/X VPWR
+ VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1178__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_4_841 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0682_ VPWR u_ppwm_u_mem__0682_/Y net522 VGND sg13g2_inv_1
XFILLER_3_373 VPWR VGND sg13g2_decap_8
XFILLER_26_1002 VPWR VGND sg13g2_decap_8
XFILLER_21_6 VPWR VGND sg13g2_fill_1
XFILLER_39_528 VPWR VGND sg13g2_decap_8
XFILLER_47_550 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1022_ VGND VPWR u_ppwm_u_ex__1017_/Y u_ppwm_u_ex__1018_/Y u_ppwm_u_ex__1022_/Y
+ u_ppwm_u_ex__1021_/Y sg13g2_a21oi_1
XFILLER_19_263 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1165_ net151 VGND VPWR net225 hold117/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_285 VPWR VGND sg13g2_decap_4
XFILLER_35_745 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1096_ net606 u_ppwm_u_mem__1102_/D u_ppwm_u_mem__1098_/B VPWR VGND
+ sg13g2_and2_1
XFILLER_15_480 VPWR VGND sg13g2_fill_2
XFILLER_15_491 VPWR VGND sg13g2_fill_2
XFILLER_31_940 VPWR VGND sg13g2_decap_8
XFILLER_30_450 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0806_ net446 VPWR u_ppwm_u_ex__0807_/A VGND u_ppwm_u_ex__0784_/A u_ppwm_u_ex__0805_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0949_ VGND VPWR net429 u_ppwm_u_mem__0680_/Y hold81/A u_ppwm_u_mem__0948_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0737_ u_ppwm_u_ex__0973_/A net454 u_ppwm_u_ex__0737_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0668_ u_ppwm_u_ex__0673_/C VPWR u_ppwm_u_ex__0668_/Y VGND u_ppwm_u_ex__0850_/A
+ net440 sg13g2_o21ai_1
Xu_ppwm_u_ex__0599_ u_ppwm_u_ex__0715_/B net369 u_ppwm_u_ex__0772_/C u_ppwm_u_ex__0601_/C
+ VPWR VGND sg13g2_nand3_1
XFILLER_26_701 VPWR VGND sg13g2_decap_8
XFILLER_38_550 VPWR VGND sg13g2_decap_8
XFILLER_25_211 VPWR VGND sg13g2_fill_1
XFILLER_25_266 VPWR VGND sg13g2_fill_2
XFILLER_26_778 VPWR VGND sg13g2_decap_8
XFILLER_41_726 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_4
XFILLER_22_962 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_8
XFILLER_0_376 VPWR VGND sg13g2_decap_8
XFILLER_48_369 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_decap_8
XFILLER_16_222 VPWR VGND sg13g2_fill_2
XFILLER_44_575 VPWR VGND sg13g2_decap_8
XFILLER_17_789 VPWR VGND sg13g2_decap_8
XFILLER_16_277 VPWR VGND sg13g2_decap_4
XFILLER_13_962 VPWR VGND sg13g2_decap_8
XFILLER_32_759 VPWR VGND sg13g2_decap_8
XFILLER_9_922 VPWR VGND sg13g2_decap_8
XFILLER_9_999 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0803_ u_ppwm_u_mem__0694_/Y u_ppwm_u_mem__0687_/Y net482 u_ppwm_u_mem__0803_/X
+ VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0734_ hold323/A net617 net611 u_ppwm_u_mem__0737_/C VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__0665_ VPWR u_ppwm_u_mem__0665_/Y net264 VGND sg13g2_inv_1
Xu_ppwm_u_ex__1005_ u_ppwm_u_ex__1027_/A net451 net376 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__1217_ net61 VGND VPWR u_ppwm_u_mem__1217_/D hold97/A clknet_5_9__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1148_ net66 VGND VPWR net557 hold228/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_748 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1079_ VGND VPWR net403 u_ppwm_u_mem__0615_/Y hold98/A u_ppwm_u_mem__1078_/Y
+ sg13g2_a21oi_1
XFILLER_46_818 VPWR VGND sg13g2_decap_8
XFILLER_45_317 VPWR VGND sg13g2_decap_4
XFILLER_39_892 VPWR VGND sg13g2_decap_8
XFILLER_41_523 VPWR VGND sg13g2_decap_8
XFILLER_14_748 VPWR VGND sg13g2_decap_8
XFILLER_26_575 VPWR VGND sg13g2_decap_8
XFILLER_10_976 VPWR VGND sg13g2_decap_8
XFILLER_6_947 VPWR VGND sg13g2_decap_8
XFILLER_5_479 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_49_634 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_0_184 VPWR VGND sg13g2_decap_8
XFILLER_48_166 VPWR VGND sg13g2_decap_8
XFILLER_48_155 VPWR VGND sg13g2_fill_2
XFILLER_37_829 VPWR VGND sg13g2_decap_8
XFILLER_29_391 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1002_ net498 VPWR u_ppwm_u_mem__1002_/Y VGND net415 hold67/A sg13g2_o21ai_1
XFILLER_45_884 VPWR VGND sg13g2_decap_8
XFILLER_44_383 VPWR VGND sg13g2_decap_4
XFILLER_17_586 VPWR VGND sg13g2_decap_8
XFILLER_32_556 VPWR VGND sg13g2_decap_8
XFILLER_20_718 VPWR VGND sg13g2_decap_8
XFILLER_9_796 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0717_ VPWR u_ppwm_u_mem__0717_/Y net298 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0648_ VPWR u_ppwm_u_mem__0648_/Y net583 VGND sg13g2_inv_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
XFILLER_27_306 VPWR VGND sg13g2_decap_8
XFILLER_36_851 VPWR VGND sg13g2_decap_8
XFILLER_11_707 VPWR VGND sg13g2_decap_8
XFILLER_23_545 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1107__37 VPWR VGND net37 sg13g2_tiehi
Xhold240 hold240/A VPWR VGND net608 sg13g2_dlygate4sd3_1
Xhold262 hold262/A VPWR VGND net630 sg13g2_dlygate4sd3_1
Xhold251 hold251/A VPWR VGND net619 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
Xhold284 hold284/A VPWR VGND net652 sg13g2_dlygate4sd3_1
Xhold295 hold295/A VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold273 hold273/A VPWR VGND net641 sg13g2_dlygate4sd3_1
XFILLER_46_615 VPWR VGND sg13g2_decap_8
XFILLER_45_125 VPWR VGND sg13g2_decap_4
XFILLER_27_851 VPWR VGND sg13g2_decap_8
XFILLER_42_810 VPWR VGND sg13g2_decap_8
XFILLER_14_545 VPWR VGND sg13g2_decap_8
XFILLER_42_887 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__239__189 VPWR VGND net189 sg13g2_tiehi
Xu_ppwm_u_pwm__241_ net182 VGND VPWR u_ppwm_u_pwm__241_/D hold283/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_6_744 VPWR VGND sg13g2_decap_8
XFILLER_10_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__172_ u_ppwm_u_pwm__173_/B net652 u_ppwm_u_pwm__175_/C VPWR VGND sg13g2_xnor2_1
XFILLER_2_961 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_4
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_37_626 VPWR VGND sg13g2_decap_8
XFILLER_18_862 VPWR VGND sg13g2_decap_8
XFILLER_45_681 VPWR VGND sg13g2_decap_8
XFILLER_32_320 VPWR VGND sg13g2_decap_4
XFILLER_20_515 VPWR VGND sg13g2_decap_8
XFILLER_33_876 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0985_ u_ppwm_u_ex__0985_/A net446 fanout351/A VPWR VGND sg13g2_nor2b_1
XFILLER_9_593 VPWR VGND sg13g2_decap_8
XFILLER_28_659 VPWR VGND sg13g2_decap_8
XFILLER_43_629 VPWR VGND sg13g2_decap_8
XFILLER_15_309 VPWR VGND sg13g2_fill_1
XFILLER_23_320 VPWR VGND sg13g2_decap_8
XFILLER_24_843 VPWR VGND sg13g2_decap_8
XFILLER_11_504 VPWR VGND sg13g2_decap_8
XFILLER_13_1004 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_3_758 VPWR VGND sg13g2_decap_8
XFILLER_47_935 VPWR VGND sg13g2_decap_8
XFILLER_46_412 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_659 VPWR VGND sg13g2_decap_8
XFILLER_46_489 VPWR VGND sg13g2_decap_8
XFILLER_15_810 VPWR VGND sg13g2_decap_8
XFILLER_34_618 VPWR VGND sg13g2_decap_8
XFILLER_15_887 VPWR VGND sg13g2_decap_8
XFILLER_42_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0982_ net496 VPWR u_ppwm_u_mem__0982_/Y VGND net409 net306 sg13g2_o21ai_1
Xu_ppwm_u_ex__0770_ net492 VPWR hold281/A VGND net648 u_ppwm_u_ex__0718_/X sg13g2_o21ai_1
XFILLER_30_868 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__224_ u_ppwm_u_pwm__223_/Y VPWR u_ppwm_u_pwm__226_/C VGND u_ppwm_u_pwm__221_/A
+ u_ppwm_u_pwm__219_/Y sg13g2_o21ai_1
XFILLER_10_570 VPWR VGND sg13g2_decap_8
XFILLER_6_541 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__155_ net490 VPWR u_ppwm_u_pwm__155_/Y VGND hold296/A net389 sg13g2_o21ai_1
XFILLER_29_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_935 VPWR VGND sg13g2_decap_8
XFILLER_24_106 VPWR VGND sg13g2_fill_2
XFILLER_17_180 VPWR VGND sg13g2_fill_2
XFILLER_21_813 VPWR VGND sg13g2_decap_8
XFILLER_33_673 VPWR VGND sg13g2_decap_8
XFILLER_36_1026 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0968_ u_ppwm_u_ex__0968_/Y net454 net374 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__0899_ net505 VPWR u_ppwm_u_ex__0900_/A VGND net460 net353 sg13g2_o21ai_1
Xu_ppwm_u_mem__1171__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_924 VPWR VGND sg13g2_decap_8
XFILLER_43_426 VPWR VGND sg13g2_decap_8
XFILLER_16_629 VPWR VGND sg13g2_decap_8
XFILLER_37_990 VPWR VGND sg13g2_decap_8
XFILLER_24_640 VPWR VGND sg13g2_decap_8
XFILLER_12_846 VPWR VGND sg13g2_decap_8
XFILLER_8_828 VPWR VGND sg13g2_decap_8
XFILLER_11_345 VPWR VGND sg13g2_decap_4
XFILLER_7_316 VPWR VGND sg13g2_fill_2
XFILLER_11_389 VPWR VGND sg13g2_fill_2
XFILLER_3_555 VPWR VGND sg13g2_decap_8
XFILLER_47_732 VPWR VGND sg13g2_decap_8
Xfanout391 fanout391/A net391 VPWR VGND sg13g2_buf_8
XFILLER_4_1002 VPWR VGND sg13g2_decap_8
Xfanout380 fanout380/A net380 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1181_ net91 VGND VPWR u_ppwm_u_mem__1181_/D hold46/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_927 VPWR VGND sg13g2_decap_8
XFILLER_46_286 VPWR VGND sg13g2_decap_8
XFILLER_34_437 VPWR VGND sg13g2_fill_1
XFILLER_43_993 VPWR VGND sg13g2_decap_8
XFILLER_42_481 VPWR VGND sg13g2_decap_8
XFILLER_15_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0822_ u_ppwm_u_ex__0823_/B u_ppwm_u_ex__0821_/X u_ppwm_u_ex__0790_/Y
+ u_ppwm_u_ex__0814_/A u_ppwm_u_ex__0797_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_30_665 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0965_ VGND VPWR net428 u_ppwm_u_mem__0672_/Y u_ppwm_u_mem__1159_/D
+ u_ppwm_u_mem__0964_/Y sg13g2_a21oi_1
XFILLER_7_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__207_ u_ppwm_u_pwm__209_/C hold11/A hold268/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_ex__0753_ net463 u_ppwm_u_ex__0753_/B u_ppwm_u_ex__0753_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0684_ u_ppwm_u_ex__0683_/Y VPWR u_ppwm_u_ex__0688_/A VGND net455 u_ppwm_u_ex__0585_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0896_ net515 VPWR u_ppwm_u_mem__0896_/Y VGND net436 hold190/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__138_ hold276/A hold225/A u_ppwm_u_pwm__140_/B VPWR VGND sg13g2_nor2_1
XFILLER_38_732 VPWR VGND sg13g2_decap_8
XFILLER_41_908 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1098_ VGND VPWR u_ppwm_u_ex__1092_/Y u_ppwm_u_ex__1096_/Y hold290/A
+ u_ppwm_u_ex__1097_/Y sg13g2_a21oi_1
Xu_ppwm_u_global_counter__087_ VGND VPWR net398 net392 u_ppwm_u_global_counter__089_/A
+ net440 sg13g2_a21oi_1
XFILLER_40_429 VPWR VGND sg13g2_fill_1
XFILLER_21_610 VPWR VGND sg13g2_decap_8
XFILLER_34_982 VPWR VGND sg13g2_decap_8
XFILLER_21_687 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_fill_1
XFILLER_10_1018 VPWR VGND sg13g2_decap_8
XFILLER_0_558 VPWR VGND sg13g2_decap_8
XFILLER_29_721 VPWR VGND sg13g2_decap_8
XFILLER_28_264 VPWR VGND sg13g2_decap_8
XFILLER_28_275 VPWR VGND sg13g2_fill_2
XFILLER_29_798 VPWR VGND sg13g2_decap_8
XFILLER_44_757 VPWR VGND sg13g2_decap_8
XFILLER_25_960 VPWR VGND sg13g2_decap_8
XFILLER_12_643 VPWR VGND sg13g2_decap_8
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_8_625 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_fill_1
XFILLER_7_179 VPWR VGND sg13g2_fill_1
XFILLER_4_820 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0750_ net484 hold229/A hold86/A hold77/A hold149/A net475 u_ppwm_u_mem__0750_/X
+ VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0681_ VPWR u_ppwm_u_mem__0681_/Y net310 VGND sg13g2_inv_1
XFILLER_4_897 VPWR VGND sg13g2_decap_8
XFILLER_39_507 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1021_ net351 VPWR u_ppwm_u_ex__1021_/Y VGND net360 u_ppwm_u_ex__1020_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__1164_ net153 VGND VPWR net316 hold163/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1115__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_35_724 VPWR VGND sg13g2_decap_8
XFILLER_34_234 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1095_ net606 u_ppwm_u_mem__1102_/D hold239/A VPWR VGND sg13g2_nor2_1
XFILLER_22_407 VPWR VGND sg13g2_decap_4
XFILLER_43_790 VPWR VGND sg13g2_decap_8
XFILLER_16_993 VPWR VGND sg13g2_decap_8
XFILLER_31_996 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0805_ net388 net385 u_ppwm_u_ex__0805_/C u_ppwm_u_ex__0805_/Y VPWR VGND
+ sg13g2_nor3_1
Xu_ppwm_u_mem__0948_ net511 VPWR u_ppwm_u_mem__0948_/Y VGND net430 hold112/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0736_ u_ppwm_u_ex__0739_/A net455 u_ppwm_u_ex__0711_/A net454 u_ppwm_u_ex__0973_/A
+ VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_ex__0667_ u_ppwm_u_ex__0673_/C net462 u_ppwm_u_ex__1020_/B2 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0879_ VGND VPWR net434 u_ppwm_u_mem__0715_/Y u_ppwm_u_mem__1116_/D
+ u_ppwm_u_mem__0878_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0598_ net375 net378 fanout369/A VPWR VGND sg13g2_nor2_1
XFILLER_26_757 VPWR VGND sg13g2_decap_8
XFILLER_41_705 VPWR VGND sg13g2_decap_8
XFILLER_43_48 VPWR VGND sg13g2_fill_2
XFILLER_22_941 VPWR VGND sg13g2_decap_8
XFILLER_21_484 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_0_355 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_48_348 VPWR VGND sg13g2_decap_8
XFILLER_29_595 VPWR VGND sg13g2_decap_8
XFILLER_44_554 VPWR VGND sg13g2_decap_8
XFILLER_16_234 VPWR VGND sg13g2_fill_2
XFILLER_17_82 VPWR VGND sg13g2_fill_1
XFILLER_17_768 VPWR VGND sg13g2_decap_8
XFILLER_32_738 VPWR VGND sg13g2_decap_8
XFILLER_9_901 VPWR VGND sg13g2_decap_8
XFILLER_13_941 VPWR VGND sg13g2_decap_8
XFILLER_31_237 VPWR VGND sg13g2_fill_2
XFILLER_40_782 VPWR VGND sg13g2_decap_8
XFILLER_9_978 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0802_ VPWR VGND u_ppwm_u_mem__0801_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0799_/Y
+ u_ppwm_u_mem__0795_/Y u_ppwm_u_mem__0802_/Y u_ppwm_u_mem__0797_/Y sg13g2_a221oi_1
XFILLER_8_499 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0733_ net587 net606 net565 u_ppwm_u_mem__0737_/B VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__0664_ VPWR u_ppwm_u_mem__0664_/Y net306 VGND sg13g2_inv_1
XFILLER_4_694 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1004_ u_ppwm_u_ex__1017_/A net451 net376 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1216_ net77 VGND VPWR net296 hold159/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1147_ net68 VGND VPWR u_ppwm_u_mem__1147_/D hold75/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_23_727 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1078_ net494 VPWR u_ppwm_u_mem__1078_/Y VGND net403 hold159/A sg13g2_o21ai_1
XFILLER_35_598 VPWR VGND sg13g2_decap_8
XFILLER_16_790 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_fill_2
XFILLER_31_793 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0719_ u_ppwm_u_ex__1049_/A net457 u_ppwm_u_ex__0719_/Y VPWR VGND sg13g2_nor2_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_39_871 VPWR VGND sg13g2_decap_8
XFILLER_26_554 VPWR VGND sg13g2_decap_8
XFILLER_41_502 VPWR VGND sg13g2_decap_8
XFILLER_14_727 VPWR VGND sg13g2_decap_8
XFILLER_41_579 VPWR VGND sg13g2_decap_8
XFILLER_10_955 VPWR VGND sg13g2_decap_8
XFILLER_6_926 VPWR VGND sg13g2_decap_8
XFILLER_5_458 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_48_101 VPWR VGND sg13g2_fill_1
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_808 VPWR VGND sg13g2_decap_8
XFILLER_45_863 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1001_ VGND VPWR net414 u_ppwm_u_mem__0654_/Y hold68/A u_ppwm_u_mem__1000_/Y
+ sg13g2_a21oi_1
XFILLER_17_565 VPWR VGND sg13g2_decap_8
XFILLER_32_535 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1116__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_12_281 VPWR VGND sg13g2_fill_1
XFILLER_9_775 VPWR VGND sg13g2_decap_8
XFILLER_8_285 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0716_ VPWR u_ppwm_u_mem__0716_/Y net561 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0647_ VPWR u_ppwm_u_mem__0647_/Y net322 VGND sg13g2_inv_1
XFILLER_4_491 VPWR VGND sg13g2_decap_8
XFILLER_39_123 VPWR VGND sg13g2_fill_1
XFILLER_36_830 VPWR VGND sg13g2_decap_8
XFILLER_23_524 VPWR VGND sg13g2_decap_8
XFILLER_10_229 VPWR VGND sg13g2_fill_1
XFILLER_31_590 VPWR VGND sg13g2_decap_8
Xhold252 hold252/A VPWR VGND net620 sg13g2_dlygate4sd3_1
Xhold241 hold241/A VPWR VGND net609 sg13g2_dlygate4sd3_1
Xhold230 hold230/A VPWR VGND net598 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_8 VPWR VGND sg13g2_decap_8
Xhold296 hold296/A VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold263 hold263/A VPWR VGND net631 sg13g2_dlygate4sd3_1
Xhold285 hold285/A VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold274 hold274/A VPWR VGND net642 sg13g2_dlygate4sd3_1
XFILLER_18_307 VPWR VGND sg13g2_decap_4
XFILLER_27_830 VPWR VGND sg13g2_decap_8
XFILLER_42_866 VPWR VGND sg13g2_decap_8
XFILLER_14_524 VPWR VGND sg13g2_decap_8
XFILLER_41_387 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__240_ net186 VGND VPWR net574 hold204/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
XFILLER_14_72 VPWR VGND sg13g2_decap_4
XFILLER_10_752 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__171_ u_ppwm_u_pwm__188_/A u_ppwm_u_pwm__171_/B u_ppwm_u_pwm__175_/C
+ u_ppwm_u_pwm__241_/D VPWR VGND sg13g2_nor3_1
XFILLER_6_723 VPWR VGND sg13g2_decap_8
XFILLER_5_222 VPWR VGND sg13g2_decap_8
XFILLER_5_211 VPWR VGND sg13g2_decap_4
XFILLER_5_288 VPWR VGND sg13g2_decap_4
XFILLER_2_940 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_37_605 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_18_841 VPWR VGND sg13g2_decap_8
XFILLER_45_660 VPWR VGND sg13g2_decap_8
XFILLER_17_351 VPWR VGND sg13g2_decap_4
XFILLER_44_181 VPWR VGND sg13g2_fill_1
XFILLER_33_855 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0984_ u_ppwm_u_ex__0985_/A u_ppwm_u_ex__0983_/Y u_ppwm_u_ex__0784_/A
+ u_ppwm_u_ex__0804_/Y net385 VPWR VGND sg13g2_a22oi_1
XFILLER_32_398 VPWR VGND sg13g2_fill_1
XFILLER_9_572 VPWR VGND sg13g2_decap_8
XFILLER_28_638 VPWR VGND sg13g2_decap_8
XFILLER_43_608 VPWR VGND sg13g2_decap_8
XFILLER_24_822 VPWR VGND sg13g2_decap_8
XFILLER_23_343 VPWR VGND sg13g2_fill_1
XFILLER_23_387 VPWR VGND sg13g2_fill_1
XFILLER_24_899 VPWR VGND sg13g2_decap_8
XFILLER_3_737 VPWR VGND sg13g2_decap_8
XFILLER_2_247 VPWR VGND sg13g2_fill_1
XFILLER_47_914 VPWR VGND sg13g2_decap_8
XFILLER_19_638 VPWR VGND sg13g2_decap_8
XFILLER_46_468 VPWR VGND sg13g2_decap_8
XFILLER_42_663 VPWR VGND sg13g2_decap_8
XFILLER_14_343 VPWR VGND sg13g2_fill_1
XFILLER_15_866 VPWR VGND sg13g2_decap_8
XFILLER_41_184 VPWR VGND sg13g2_fill_1
XFILLER_41_162 VPWR VGND sg13g2_fill_1
XFILLER_14_398 VPWR VGND sg13g2_decap_4
XFILLER_30_847 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0981_ VGND VPWR net409 u_ppwm_u_mem__0664_/Y u_ppwm_u_mem__1167_/D
+ u_ppwm_u_mem__0980_/Y sg13g2_a21oi_1
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_pwm__223_ u_ppwm_u_pwm__223_/Y net644 u_ppwm_u_pwm__223_/B VPWR VGND sg13g2_nand2_1
XFILLER_6_520 VPWR VGND sg13g2_decap_8
XFILLER_41_81 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__154_ VGND VPWR u_ppwm_u_pwm__129_/Y net391 hold12/A u_ppwm_u_pwm__153_/Y
+ sg13g2_a21oi_1
XFILLER_6_597 VPWR VGND sg13g2_decap_8
XFILLER_29_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_fill_1
XFILLER_38_914 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_2_75 VPWR VGND sg13g2_decap_4
XFILLER_33_652 VPWR VGND sg13g2_decap_8
XFILLER_36_1005 VPWR VGND sg13g2_decap_8
XFILLER_32_173 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0967_ VGND VPWR u_ppwm_u_ex__0953_/Y u_ppwm_u_ex__0955_/X u_ppwm_u_ex__0967_/Y
+ u_ppwm_u_ex__0954_/Y sg13g2_a21oi_1
XFILLER_21_869 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1125__112 VPWR VGND net112 sg13g2_tiehi
Xu_ppwm_u_ex__0898_ u_ppwm_u_ex__0898_/B u_ppwm_u_ex__1035_/A net352 u_ppwm_u_ex__0898_/Y
+ VPWR VGND u_ppwm_u_ex__0898_/D sg13g2_nand4_1
XFILLER_29_903 VPWR VGND sg13g2_decap_8
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_43_405 VPWR VGND sg13g2_decap_8
XFILLER_16_608 VPWR VGND sg13g2_decap_8
XFILLER_12_825 VPWR VGND sg13g2_decap_8
XFILLER_24_696 VPWR VGND sg13g2_decap_8
XFILLER_8_807 VPWR VGND sg13g2_decap_8
XFILLER_11_379 VPWR VGND sg13g2_fill_2
XFILLER_3_534 VPWR VGND sg13g2_decap_8
XFILLER_47_711 VPWR VGND sg13g2_decap_8
Xfanout392 fanout392/A net392 VPWR VGND sg13g2_buf_2
Xfanout370 fanout370/A net370 VPWR VGND sg13g2_buf_8
XFILLER_19_402 VPWR VGND sg13g2_decap_4
Xfanout381 net383 net381 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1180_ net95 VGND VPWR u_ppwm_u_mem__1180_/D hold36/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_906 VPWR VGND sg13g2_decap_8
XFILLER_47_788 VPWR VGND sg13g2_decap_8
XFILLER_46_265 VPWR VGND sg13g2_decap_8
XFILLER_43_972 VPWR VGND sg13g2_decap_8
XFILLER_15_663 VPWR VGND sg13g2_decap_8
XFILLER_42_460 VPWR VGND sg13g2_decap_8
XFILLER_14_195 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0821_ u_ppwm_u_ex__0866_/C u_ppwm_u_ex__0800_/X net378 u_ppwm_u_ex__0821_/X
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_644 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0964_ net510 VPWR u_ppwm_u_mem__0964_/Y VGND net427 net536 sg13g2_o21ai_1
Xu_ppwm_u_ex__0752_ u_ppwm_u_ex__0751_/Y VPWR u_ppwm_u_ex__0752_/Y VGND u_ppwm_u_ex__0748_/Y
+ u_ppwm_u_ex__0750_/Y sg13g2_o21ai_1
Xu_ppwm_u_pwm__206_ u_ppwm_u_pwm__206_/Y u_ppwm_u_pwm__209_/A u_ppwm_u_pwm__209_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__0683_ u_ppwm_u_ex__0683_/Y u_ppwm_u_ex__0683_/A hold217/A VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0895_ VGND VPWR net436 u_ppwm_u_mem__0707_/Y u_ppwm_u_mem__1124_/D
+ u_ppwm_u_mem__0894_/Y sg13g2_a21oi_1
XFILLER_6_394 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__137_ hold283/A hold204/A hold181/A hold279/A u_ppwm_u_pwm__140_/A VPWR
+ VGND sg13g2_nor4_1
XFILLER_42_1020 VPWR VGND sg13g2_decap_8
XFILLER_38_711 VPWR VGND sg13g2_decap_8
XFILLER_26_939 VPWR VGND sg13g2_decap_8
XFILLER_38_788 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1097_ net491 VPWR u_ppwm_u_ex__1097_/Y VGND net657 net349 sg13g2_o21ai_1
XFILLER_16_18 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__086_ hold273/A fanout392/A net398 net640 u_ppwm_u_global_counter__054_/Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_25_427 VPWR VGND sg13g2_fill_1
XFILLER_34_961 VPWR VGND sg13g2_decap_8
XFILLER_21_666 VPWR VGND sg13g2_decap_8
XFILLER_20_198 VPWR VGND sg13g2_decap_4
XFILLER_0_537 VPWR VGND sg13g2_decap_8
XFILLER_29_700 VPWR VGND sg13g2_decap_8
XFILLER_29_777 VPWR VGND sg13g2_decap_8
XFILLER_44_736 VPWR VGND sg13g2_decap_8
XFILLER_12_622 VPWR VGND sg13g2_decap_8
XFILLER_31_419 VPWR VGND sg13g2_fill_1
XFILLER_40_964 VPWR VGND sg13g2_decap_8
XFILLER_8_604 VPWR VGND sg13g2_decap_8
XFILLER_24_493 VPWR VGND sg13g2_decap_8
XFILLER_12_699 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0680_ VPWR u_ppwm_u_mem__0680_/Y net278 VGND sg13g2_inv_1
XFILLER_4_876 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1020_ VPWR VGND u_ppwm_u_ex__1020_/B2 u_ppwm_u_ex__1019_/Y net355 net692
+ u_ppwm_u_ex__1020_/Y net362 sg13g2_a221oi_1
Xu_ppwm_u_mem__1163_ net155 VGND VPWR u_ppwm_u_mem__1163_/D hold88/A clknet_5_15__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_703 VPWR VGND sg13g2_decap_8
XFILLER_47_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1094_ u_ppwm_u_mem__1094_/A net612 u_ppwm_u_mem__1102_/D hold245/A
+ VPWR VGND sg13g2_nor3_1
XFILLER_23_909 VPWR VGND sg13g2_decap_8
XFILLER_34_257 VPWR VGND sg13g2_fill_1
XFILLER_16_972 VPWR VGND sg13g2_decap_8
XFILLER_31_975 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0804_ net388 u_ppwm_u_ex__0805_/C u_ppwm_u_ex__0804_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0735_ u_ppwm_u_ex__0735_/Y u_ppwm_u_ex__0735_/A hold296/A VPWR VGND
+ sg13g2_nand2_1
XFILLER_8_96 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0947_ VGND VPWR net429 u_ppwm_u_mem__0681_/Y hold113/A u_ppwm_u_mem__0946_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0666_ u_ppwm_u_ex__0666_/Y net466 hold207/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0878_ net514 VPWR u_ppwm_u_mem__0878_/Y VGND net434 net561 sg13g2_o21ai_1
XFILLER_40_0 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0597_ net381 net384 u_ppwm_u_ex__0715_/B VPWR VGND sg13g2_nor2b_2
XFILLER_26_736 VPWR VGND sg13g2_decap_8
XFILLER_38_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__069_ net599 net590 net659 u_ppwm_u_global_counter__085_/A
+ VPWR VGND net627 sg13g2_nand4_1
XFILLER_14_909 VPWR VGND sg13g2_decap_8
XFILLER_22_920 VPWR VGND sg13g2_decap_8
XFILLER_25_268 VPWR VGND sg13g2_fill_1
XFILLER_21_463 VPWR VGND sg13g2_decap_8
XFILLER_22_997 VPWR VGND sg13g2_decap_8
XFILLER_4_139 VPWR VGND sg13g2_fill_1
XFILLER_49_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_301 VPWR VGND sg13g2_fill_1
XFILLER_0_334 VPWR VGND sg13g2_decap_8
XFILLER_1_868 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1148__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_48_327 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_44_533 VPWR VGND sg13g2_decap_8
XFILLER_16_224 VPWR VGND sg13g2_fill_1
XFILLER_17_747 VPWR VGND sg13g2_decap_8
XFILLER_29_574 VPWR VGND sg13g2_decap_8
XFILLER_13_920 VPWR VGND sg13g2_decap_8
XFILLER_17_94 VPWR VGND sg13g2_fill_1
XFILLER_31_205 VPWR VGND sg13g2_decap_4
XFILLER_32_717 VPWR VGND sg13g2_decap_8
XFILLER_40_761 VPWR VGND sg13g2_decap_8
XFILLER_9_957 VPWR VGND sg13g2_decap_8
XFILLER_13_997 VPWR VGND sg13g2_decap_8
XFILLER_8_467 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0801_ VGND VPWR net395 u_ppwm_u_mem__0800_/X u_ppwm_u_mem__0801_/Y
+ net470 sg13g2_a21oi_1
Xu_ppwm_u_mem__0732_ VGND VPWR u_ppwm_u_mem__0726_/Y u_ppwm_u_mem__0731_/Y hold136/A
+ u_ppwm_u_mem__0730_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0663_ VPWR u_ppwm_u_mem__0663_/Y net592 VGND sg13g2_inv_1
XFILLER_4_673 VPWR VGND sg13g2_decap_8
XFILLER_3_183 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_4
Xhold1 hold1/A VPWR VGND net199 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__1003_ VGND VPWR u_ppwm_u_ex__0994_/A u_ppwm_u_ex__0994_/B u_ppwm_u_ex__1006_/A
+ u_ppwm_u_ex__0992_/X sg13g2_a21oi_1
Xu_ppwm_u_mem__1215_ net93 VGND VPWR u_ppwm_u_mem__1215_/D hold24/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_48_894 VPWR VGND sg13g2_decap_8
XFILLER_47_382 VPWR VGND sg13g2_decap_8
XFILLER_23_706 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1146_ net70 VGND VPWR net274 hold137/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1077_ VGND VPWR net404 u_ppwm_u_mem__0616_/Y u_ppwm_u_mem__1215_/D
+ u_ppwm_u_mem__1076_/Y sg13g2_a21oi_1
XFILLER_35_577 VPWR VGND sg13g2_decap_8
XFILLER_31_772 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0718_ net446 net388 u_ppwm_u_ex__0781_/A u_ppwm/instr\[1\] u_ppwm_u_ex__0718_/X
+ VPWR VGND sg13g2_and4_1
Xu_ppwm_u_ex__0649_ u_ppwm_u_ex__0649_/Y u_ppwm_u_ex__1019_/B net450 u_ppwm_u_ex__0755_/B
+ net449 VPWR VGND sg13g2_a22oi_1
XFILLER_39_850 VPWR VGND sg13g2_decap_8
XFILLER_14_706 VPWR VGND sg13g2_decap_8
XFILLER_26_533 VPWR VGND sg13g2_decap_8
XFILLER_13_205 VPWR VGND sg13g2_fill_2
XFILLER_41_558 VPWR VGND sg13g2_decap_8
XFILLER_13_227 VPWR VGND sg13g2_decap_8
XFILLER_13_238 VPWR VGND sg13g2_fill_1
XFILLER_13_249 VPWR VGND sg13g2_fill_2
XFILLER_16_1014 VPWR VGND sg13g2_decap_8
XFILLER_10_934 VPWR VGND sg13g2_decap_8
XFILLER_22_794 VPWR VGND sg13g2_decap_8
XFILLER_6_905 VPWR VGND sg13g2_decap_8
XFILLER_5_437 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_23_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_669 VPWR VGND sg13g2_decap_8
XFILLER_45_842 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1000_ net498 VPWR u_ppwm_u_mem__1000_/Y VGND net414 hold150/A sg13g2_o21ai_1
XFILLER_17_544 VPWR VGND sg13g2_decap_8
XFILLER_9_754 VPWR VGND sg13g2_decap_8
XFILLER_13_794 VPWR VGND sg13g2_decap_8
XFILLER_4_470 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0715_ VPWR u_ppwm_u_mem__0715_/Y net563 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0646_ VPWR u_ppwm_u_mem__0646_/Y net249 VGND sg13g2_inv_1
XFILLER_48_691 VPWR VGND sg13g2_decap_8
XFILLER_39_1025 VPWR VGND sg13g2_decap_4
XFILLER_23_503 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1129_ net104 VGND VPWR net525 hold84/A clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_886 VPWR VGND sg13g2_decap_8
XFILLER_3_919 VPWR VGND sg13g2_decap_8
Xhold220 hold220/A VPWR VGND net588 sg13g2_dlygate4sd3_1
Xhold253 hold253/A VPWR VGND net621 sg13g2_dlygate4sd3_1
XFILLER_2_429 VPWR VGND sg13g2_decap_8
Xhold242 hold242/A VPWR VGND net610 sg13g2_dlygate4sd3_1
Xhold231 hold231/A VPWR VGND net599 sg13g2_dlygate4sd3_1
XFILLER_46_1007 VPWR VGND sg13g2_decap_8
Xhold286 hold286/A VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold264 hold264/A VPWR VGND net632 sg13g2_dlygate4sd3_1
Xhold275 hold275/A VPWR VGND net643 sg13g2_dlygate4sd3_1
Xhold297 hold297/A VPWR VGND net665 sg13g2_dlygate4sd3_1
XFILLER_45_149 VPWR VGND sg13g2_fill_2
XFILLER_45_138 VPWR VGND sg13g2_fill_2
XFILLER_26_352 VPWR VGND sg13g2_decap_8
XFILLER_26_363 VPWR VGND sg13g2_fill_1
XFILLER_27_886 VPWR VGND sg13g2_decap_8
XFILLER_42_845 VPWR VGND sg13g2_decap_8
XFILLER_6_702 VPWR VGND sg13g2_decap_8
XFILLER_10_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__170_ net651 u_ppwm_u_pwm__170_/B u_ppwm_u_pwm__175_/C VPWR VGND sg13g2_and2_1
XFILLER_22_591 VPWR VGND sg13g2_decap_8
XFILLER_5_201 VPWR VGND sg13g2_fill_1
XFILLER_6_779 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_2_996 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_fill_2
XFILLER_18_820 VPWR VGND sg13g2_decap_8
XFILLER_18_897 VPWR VGND sg13g2_decap_8
XFILLER_33_834 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0983_ net379 u_ppwm_u_ex__0983_/B u_ppwm_u_ex__0983_/Y VPWR VGND sg13g2_nor2_1
XFILLER_9_551 VPWR VGND sg13g2_decap_8
XFILLER_13_591 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0629_ VPWR u_ppwm_u_mem__0629_/Y net213 VGND sg13g2_inv_1
XFILLER_28_617 VPWR VGND sg13g2_decap_8
XFILLER_24_801 VPWR VGND sg13g2_decap_8
XFILLER_35_160 VPWR VGND sg13g2_decap_4
XFILLER_36_683 VPWR VGND sg13g2_decap_8
XFILLER_24_878 VPWR VGND sg13g2_decap_8
XFILLER_11_539 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__238__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_3_716 VPWR VGND sg13g2_decap_8
XFILLER_19_617 VPWR VGND sg13g2_decap_8
XFILLER_46_447 VPWR VGND sg13g2_decap_8
XFILLER_15_845 VPWR VGND sg13g2_decap_8
XFILLER_26_182 VPWR VGND sg13g2_decap_8
XFILLER_27_683 VPWR VGND sg13g2_decap_8
XFILLER_42_642 VPWR VGND sg13g2_decap_8
XFILLER_30_826 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0980_ net496 VPWR u_ppwm_u_mem__0980_/Y VGND net412 net264 sg13g2_o21ai_1
Xu_ppwm_u_pwm__222_ u_ppwm_u_pwm__222_/A u_ppwm_u_pwm__222_/B u_ppwm_u_pwm__226_/B
+ VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_pwm__153_ net490 VPWR u_ppwm_u_pwm__153_/Y VGND net456 net389 sg13g2_o21ai_1
XFILLER_6_576 VPWR VGND sg13g2_decap_8
XFILLER_2_793 VPWR VGND sg13g2_decap_8
XFILLER_1_292 VPWR VGND sg13g2_fill_2
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_2_65 VPWR VGND sg13g2_fill_2
XFILLER_37_403 VPWR VGND sg13g2_fill_2
XFILLER_18_694 VPWR VGND sg13g2_decap_8
XFILLER_33_631 VPWR VGND sg13g2_decap_8
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0966_ u_ppwm_u_ex__0966_/A u_ppwm_u_ex__0964_/Y u_ppwm_u_ex__1113_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_20_336 VPWR VGND sg13g2_decap_8
XFILLER_20_347 VPWR VGND sg13g2_fill_1
XFILLER_21_848 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0897_ VGND VPWR net449 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0898_/D u_ppwm_u_ex__0896_/Y
+ sg13g2_a21oi_1
XFILLER_0_719 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_959 VPWR VGND sg13g2_decap_8
XFILLER_44_918 VPWR VGND sg13g2_decap_8
XFILLER_15_108 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1212__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_12_804 VPWR VGND sg13g2_decap_8
XFILLER_24_675 VPWR VGND sg13g2_decap_8
XFILLER_7_318 VPWR VGND sg13g2_fill_1
XFILLER_3_513 VPWR VGND sg13g2_decap_8
Xfanout371 net372 net371 VPWR VGND sg13g2_buf_8
Xfanout382 net383 net382 VPWR VGND sg13g2_buf_1
Xfanout360 fanout361/A net360 VPWR VGND sg13g2_buf_1
Xfanout393 net394 net393 VPWR VGND sg13g2_buf_8
XFILLER_46_211 VPWR VGND sg13g2_fill_2
XFILLER_19_447 VPWR VGND sg13g2_fill_2
XFILLER_47_767 VPWR VGND sg13g2_decap_8
XFILLER_46_244 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_34_417 VPWR VGND sg13g2_fill_2
XFILLER_43_951 VPWR VGND sg13g2_decap_8
XFILLER_15_642 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_fill_1
XFILLER_30_623 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0820_ u_ppwm_u_ex__0820_/B u_ppwm_u_ex__0820_/C net369 u_ppwm_u_ex__0823_/A
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__0751_ u_ppwm_u_ex__0751_/Y net443 u_ppwm_u_ex__0850_/A hold231/A u_ppwm_u_ex__0576_/Y
+ VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__0963_ VGND VPWR net430 u_ppwm_u_mem__0673_/Y u_ppwm_u_mem__1158_/D
+ u_ppwm_u_mem__0962_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__205_ u_ppwm_u_pwm__209_/B hold268/A hold11/A VPWR VGND sg13g2_nand2b_1
XFILLER_10_380 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0682_ u_ppwm_u_ex__0681_/Y VPWR u_ppwm_u_ex__0682_/Y VGND u_ppwm_u_ex__0664_/Y
+ u_ppwm_u_ex__0680_/Y sg13g2_o21ai_1
XFILLER_7_885 VPWR VGND sg13g2_decap_8
XFILLER_6_351 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__136_ u_ppwm_u_pwm__188_/A net489 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0894_ net515 VPWR u_ppwm_u_mem__0894_/Y VGND net436 net543 sg13g2_o21ai_1
XFILLER_6_384 VPWR VGND sg13g2_fill_1
XFILLER_2_590 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__228__190 VPWR VGND net190 sg13g2_tiehi
Xu_ppwm_u_global_counter__085_ u_ppwm_u_global_counter__085_/A hold298/A u_ppwm_u_global_counter__085_/C
+ fanout392/A VPWR VGND sg13g2_nor3_1
XFILLER_26_918 VPWR VGND sg13g2_decap_8
XFILLER_38_767 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1096_ VGND VPWR u_ppwm_u_ex__0820_/C u_ppwm_u_ex__0972_/Y u_ppwm_u_ex__1096_/Y
+ u_ppwm_u_ex__1095_/Y sg13g2_a21oi_1
XFILLER_19_981 VPWR VGND sg13g2_decap_8
XFILLER_18_491 VPWR VGND sg13g2_decap_8
XFILLER_34_940 VPWR VGND sg13g2_decap_8
XFILLER_33_461 VPWR VGND sg13g2_fill_1
XFILLER_21_645 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0949_ VGND VPWR u_ppwm_u_ex__0940_/Y u_ppwm_u_ex__0947_/X u_ppwm_u_ex__1112_/D
+ u_ppwm_u_ex__0948_/Y sg13g2_a21oi_1
XFILLER_0_516 VPWR VGND sg13g2_decap_8
XFILLER_48_509 VPWR VGND sg13g2_decap_8
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_29_756 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_decap_8
XFILLER_17_929 VPWR VGND sg13g2_decap_8
XFILLER_28_288 VPWR VGND sg13g2_decap_8
XFILLER_43_269 VPWR VGND sg13g2_fill_2
XFILLER_12_601 VPWR VGND sg13g2_decap_8
XFILLER_19_1023 VPWR VGND sg13g2_decap_4
XFILLER_24_472 VPWR VGND sg13g2_decap_8
XFILLER_25_995 VPWR VGND sg13g2_decap_8
XFILLER_40_943 VPWR VGND sg13g2_decap_8
XFILLER_12_678 VPWR VGND sg13g2_decap_8
XFILLER_4_855 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1016 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_564 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1162_ net157 VGND VPWR net287 hold119/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_244 VPWR VGND sg13g2_fill_2
XFILLER_16_951 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1093_ net611 net691 net624 net400 u_ppwm_u_mem__1102_/D VPWR VGND sg13g2_and4_1
XFILLER_35_759 VPWR VGND sg13g2_decap_8
XFILLER_31_954 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0803_ u_ppwm_u_ex__0983_/B net364 net361 u_ppwm_u_ex__0803_/X VPWR VGND
+ sg13g2_or3_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0734_ u_ppwm_u_ex__0733_/Y u_ppwm_u_ex__0731_/Y u_ppwm_u_ex__0719_/Y
+ u_ppwm_u_ex__0734_/X VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_mem__0946_ net511 VPWR u_ppwm_u_mem__0946_/Y VGND net429 hold154/A sg13g2_o21ai_1
XFILLER_7_682 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0665_ net464 u_ppwm_u_ex__0998_/B2 u_ppwm_u_ex__0665_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0877_ VGND VPWR net424 u_ppwm_u_mem__0716_/Y hold194/A u_ppwm_u_mem__0876_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0596_ net388 u_ppwm/instr\[0\] u_ppwm/instr\[1\] u_ppwm_u_ex__0772_/C
+ VPWR VGND sg13g2_nor3_1
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_38_564 VPWR VGND sg13g2_decap_8
XFILLER_26_715 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__068_ u_ppwm_u_global_counter__068_/B net590 hold223/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__1079_ u_ppwm_u_ex__1079_/Y hold295/A net371 VPWR VGND sg13g2_nand2_1
XFILLER_25_225 VPWR VGND sg13g2_fill_1
XFILLER_40_239 VPWR VGND sg13g2_fill_2
XFILLER_22_976 VPWR VGND sg13g2_decap_8
XFILLER_5_619 VPWR VGND sg13g2_decap_8
XFILLER_49_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_313 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_48_306 VPWR VGND sg13g2_decap_8
XFILLER_29_553 VPWR VGND sg13g2_decap_8
XFILLER_44_512 VPWR VGND sg13g2_decap_8
XFILLER_17_40 VPWR VGND sg13g2_fill_1
XFILLER_17_726 VPWR VGND sg13g2_decap_8
XFILLER_16_247 VPWR VGND sg13g2_fill_2
XFILLER_44_589 VPWR VGND sg13g2_decap_8
XFILLER_25_792 VPWR VGND sg13g2_decap_8
XFILLER_40_740 VPWR VGND sg13g2_decap_8
XFILLER_9_936 VPWR VGND sg13g2_decap_8
XFILLER_13_976 VPWR VGND sg13g2_decap_8
XFILLER_33_83 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0800_ hold26/A hold30/A net478 u_ppwm_u_mem__0800_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0731_ net1 u_ppwm_u_mem__1094_/A u_ppwm_u_mem__0731_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0662_ VPWR u_ppwm_u_mem__0662_/Y net267 VGND sg13g2_inv_1
XFILLER_4_652 VPWR VGND sg13g2_decap_8
XFILLER_0_880 VPWR VGND sg13g2_decap_8
Xhold2 hold2/A VPWR VGND net200 sg13g2_dlygate4sd3_1
XFILLER_48_873 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1002_ u_ppwm_u_ex__1002_/A u_ppwm_u_ex__1002_/B hold311/A VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_mem__1214_ net109 VGND VPWR net223 hold92/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_361 VPWR VGND sg13g2_decap_8
XFILLER_35_556 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1145_ net72 VGND VPWR u_ppwm_u_mem__1145_/D hold122/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1119__26 VPWR VGND net26 sg13g2_tiehi
Xu_ppwm_u_mem__1076_ net495 VPWR u_ppwm_u_mem__1076_/Y VGND net404 net222 sg13g2_o21ai_1
XFILLER_22_228 VPWR VGND sg13g2_fill_2
XFILLER_31_751 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0717_ VPWR VGND u_ppwm_u_ex__0708_/Y u_ppwm_u_ex__0716_/Y u_ppwm_u_ex__0714_/Y
+ u_ppwm_u_ex__0714_/A u_ppwm_u_ex__0769_/C u_ppwm_u_ex__0712_/Y sg13g2_a221oi_1
Xu_ppwm_u_mem__0929_ VGND VPWR net417 u_ppwm_u_mem__0690_/Y u_ppwm_u_mem__1141_/D
+ u_ppwm_u_mem__0928_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0648_ u_ppwm_u_ex__0647_/Y VPWR u_ppwm_u_ex__0648_/Y VGND net452 u_ppwm_u_ex__0591_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__0579_ net506 u_ppwm_u_ex__0991_/A VPWR VGND sg13g2_inv_4
XFILLER_26_589 VPWR VGND sg13g2_decap_8
XFILLER_41_537 VPWR VGND sg13g2_decap_8
XFILLER_10_913 VPWR VGND sg13g2_decap_8
XFILLER_22_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1209__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_648 VPWR VGND sg13g2_decap_8
XFILLER_48_136 VPWR VGND sg13g2_fill_2
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_17_523 VPWR VGND sg13g2_decap_8
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_4
XFILLER_9_733 VPWR VGND sg13g2_decap_8
XFILLER_13_773 VPWR VGND sg13g2_decap_8
XFILLER_5_983 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0714_ VPWR u_ppwm_u_mem__0714_/Y net280 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0645_ VPWR u_ppwm_u_mem__0645_/Y net236 VGND sg13g2_inv_1
XFILLER_39_103 VPWR VGND sg13g2_fill_2
XFILLER_48_670 VPWR VGND sg13g2_decap_8
XFILLER_39_1004 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1128_ net106 VGND VPWR net283 hold149/A clknet_5_23__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1135__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_36_865 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1150__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_23_559 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1059_ VGND VPWR net402 u_ppwm_u_mem__0625_/Y hold61/A u_ppwm_u_mem__1058_/Y
+ sg13g2_a21oi_1
Xhold210 hold210/A VPWR VGND net578 sg13g2_dlygate4sd3_1
XFILLER_2_408 VPWR VGND sg13g2_decap_8
Xhold232 hold232/A VPWR VGND net600 sg13g2_dlygate4sd3_1
Xhold221 hold221/A VPWR VGND net589 sg13g2_dlygate4sd3_1
Xhold243 hold243/A VPWR VGND net611 sg13g2_dlygate4sd3_1
Xhold276 hold276/A VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold254 hold254/A VPWR VGND net622 sg13g2_dlygate4sd3_1
Xhold287 hold291/A VPWR VGND net655 sg13g2_dlygate4sd3_1
Xhold265 hold265/A VPWR VGND net633 sg13g2_dlygate4sd3_1
XFILLER_49_49 VPWR VGND sg13g2_decap_8
Xhold298 hold298/A VPWR VGND net666 sg13g2_dlygate4sd3_1
XFILLER_46_629 VPWR VGND sg13g2_decap_8
XFILLER_27_865 VPWR VGND sg13g2_decap_8
XFILLER_42_824 VPWR VGND sg13g2_decap_8
XFILLER_14_559 VPWR VGND sg13g2_decap_8
XFILLER_10_710 VPWR VGND sg13g2_decap_8
XFILLER_22_570 VPWR VGND sg13g2_decap_8
XFILLER_10_787 VPWR VGND sg13g2_decap_8
XFILLER_6_758 VPWR VGND sg13g2_decap_8
XFILLER_30_40 VPWR VGND sg13g2_fill_1
XFILLER_2_975 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_17_320 VPWR VGND sg13g2_decap_4
XFILLER_18_876 VPWR VGND sg13g2_decap_8
XFILLER_33_813 VPWR VGND sg13g2_decap_8
XFILLER_45_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0982_ u_ppwm_u_ex__0981_/Y u_ppwm_u_ex__0980_/Y net360 u_ppwm_u_ex__0989_/B
+ VPWR VGND sg13g2_a21o_1
XFILLER_13_570 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_decap_8
XFILLER_9_530 VPWR VGND sg13g2_decap_8
XFILLER_5_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0628_ VPWR u_ppwm_u_mem__0628_/Y net328 VGND sg13g2_inv_1
XFILLER_36_662 VPWR VGND sg13g2_decap_8
XFILLER_23_334 VPWR VGND sg13g2_fill_2
XFILLER_24_857 VPWR VGND sg13g2_decap_8
XFILLER_35_194 VPWR VGND sg13g2_fill_2
XFILLER_11_518 VPWR VGND sg13g2_decap_8
XFILLER_13_1018 VPWR VGND sg13g2_decap_8
XFILLER_47_949 VPWR VGND sg13g2_decap_8
XFILLER_46_426 VPWR VGND sg13g2_decap_8
XFILLER_27_662 VPWR VGND sg13g2_decap_8
XFILLER_42_621 VPWR VGND sg13g2_decap_8
XFILLER_15_824 VPWR VGND sg13g2_decap_8
XFILLER_30_805 VPWR VGND sg13g2_decap_8
XFILLER_42_698 VPWR VGND sg13g2_decap_8
XFILLER_25_84 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__221_ u_ppwm_u_pwm__222_/B u_ppwm_u_pwm__221_/A u_ppwm_u_pwm__221_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_pwm__152_ VGND VPWR u_ppwm_u_pwm__214_/B net389 hold63/A u_ppwm_u_pwm__151_/Y
+ sg13g2_a21oi_1
XFILLER_10_584 VPWR VGND sg13g2_decap_8
XFILLER_6_555 VPWR VGND sg13g2_decap_8
XFILLER_2_772 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_38_949 VPWR VGND sg13g2_decap_8
XFILLER_46_993 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_decap_8
XFILLER_18_673 VPWR VGND sg13g2_decap_8
XFILLER_33_610 VPWR VGND sg13g2_decap_8
XFILLER_45_492 VPWR VGND sg13g2_decap_8
XFILLER_20_304 VPWR VGND sg13g2_decap_4
XFILLER_20_315 VPWR VGND sg13g2_fill_2
XFILLER_21_827 VPWR VGND sg13g2_decap_8
XFILLER_33_687 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0965_ net490 VPWR u_ppwm_u_ex__0966_/A VGND net455 net352 sg13g2_o21ai_1
XFILLER_32_175 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0896_ net359 u_ppwm_u_ex__0896_/B u_ppwm_u_ex__0896_/Y VPWR VGND sg13g2_nor2_1
XFILLER_29_938 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_4
XFILLER_24_654 VPWR VGND sg13g2_decap_8
XFILLER_23_142 VPWR VGND sg13g2_decap_4
XFILLER_20_893 VPWR VGND sg13g2_decap_8
XFILLER_3_569 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xfanout350 net351 net350 VPWR VGND sg13g2_buf_8
Xfanout372 net374 net372 VPWR VGND sg13g2_buf_2
XFILLER_4_1016 VPWR VGND sg13g2_decap_8
Xfanout361 fanout361/A net361 VPWR VGND sg13g2_buf_8
Xfanout383 fanout383/A net383 VPWR VGND sg13g2_buf_8
XFILLER_47_746 VPWR VGND sg13g2_decap_8
XFILLER_46_223 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
Xfanout394 fanout394/A net394 VPWR VGND sg13g2_buf_8
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_43_930 VPWR VGND sg13g2_decap_8
XFILLER_15_621 VPWR VGND sg13g2_decap_8
XFILLER_14_153 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_42_495 VPWR VGND sg13g2_decap_8
XFILLER_15_698 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0750_ VGND VPWR u_ppwm_u_ex__0746_/Y u_ppwm_u_ex__0749_/Y u_ppwm_u_ex__0750_/Y
+ u_ppwm_u_ex__0745_/Y sg13g2_a21oi_1
XFILLER_30_679 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0962_ net512 VPWR u_ppwm_u_mem__0962_/Y VGND net429 net245 sg13g2_o21ai_1
Xu_ppwm_u_pwm__204_ u_ppwm_u_pwm__209_/A hold178/A hold13/A VPWR VGND sg13g2_nand2b_1
XFILLER_11_882 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0681_ u_ppwm_u_ex__0681_/Y u_ppwm_u_ex__0757_/A hold277/A VPWR VGND
+ sg13g2_nand2_1
XFILLER_7_864 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__135_ VPWR u_ppwm_u_pwm__135_/Y net199 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0893_ VGND VPWR net433 u_ppwm_u_mem__0708_/Y hold176/A u_ppwm_u_mem__0892_/Y
+ sg13g2_a21oi_1
XFILLER_35_4 VPWR VGND sg13g2_fill_2
XFILLER_38_746 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1184__79 VPWR VGND net79 sg13g2_tiehi
Xu_ppwm_u_ex__1095_ net350 VPWR u_ppwm_u_ex__1095_/Y VGND net361 u_ppwm_u_ex__1094_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_global_counter__084_ net639 net575 net442 u_ppwm_u_global_counter__085_/C
+ VPWR VGND u_ppwm_u_ex__0998_/B2 sg13g2_nand4_1
XFILLER_19_960 VPWR VGND sg13g2_decap_8
XFILLER_46_790 VPWR VGND sg13g2_decap_8
XFILLER_34_996 VPWR VGND sg13g2_decap_8
XFILLER_21_624 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0948_ net491 VPWR u_ppwm_u_ex__0948_/Y VGND net664 net352 sg13g2_o21ai_1
Xu_ppwm_u_ex__0879_ u_ppwm_u_ex__0991_/A u_ppwm_u_ex__0879_/B u_ppwm_u_ex__1108_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_29_735 VPWR VGND sg13g2_decap_8
XFILLER_17_908 VPWR VGND sg13g2_decap_8
XFILLER_19_1002 VPWR VGND sg13g2_decap_8
XFILLER_40_922 VPWR VGND sg13g2_decap_8
XFILLER_25_974 VPWR VGND sg13g2_decap_8
XFILLER_11_134 VPWR VGND sg13g2_fill_1
XFILLER_12_657 VPWR VGND sg13g2_decap_8
XFILLER_40_999 VPWR VGND sg13g2_decap_8
XFILLER_8_639 VPWR VGND sg13g2_decap_8
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_fill_1
XFILLER_4_834 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1219__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_47_543 VPWR VGND sg13g2_decap_8
XFILLER_47_60 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1161_ net159 VGND VPWR u_ppwm_u_mem__1161_/D hold73/A clknet_5_27__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1154__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_19_234 VPWR VGND sg13g2_decap_4
XFILLER_35_738 VPWR VGND sg13g2_decap_8
XFILLER_16_930 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1092_ VGND VPWR net611 u_ppwm_u_mem__1085_/B hold244/A u_ppwm_u_mem__1091_/C
+ sg13g2_a21oi_1
XFILLER_31_933 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0802_ u_ppwm_u_ex__0989_/A u_ppwm_u_ex__0797_/Y u_ppwm_u_ex__0801_/X
+ u_ppwm_u_ex__0795_/Y u_ppwm_u_ex__0790_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_30_465 VPWR VGND sg13g2_decap_4
XFILLER_7_661 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0733_ VPWR VGND u_ppwm_u_ex__0651_/A u_ppwm_u_ex__0732_/Y net458 u_ppwm_u_ex__1049_/A
+ u_ppwm_u_ex__0733_/Y net457 sg13g2_a221oi_1
Xu_ppwm_u_mem__0945_ VGND VPWR net429 u_ppwm_u_mem__0682_/Y hold155/A u_ppwm_u_mem__0944_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0664_ net439 net456 u_ppwm_u_ex__0664_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0876_ net514 VPWR u_ppwm_u_mem__0876_/Y VGND net424 net298 sg13g2_o21ai_1
Xu_ppwm_u_ex__0595_ u_ppwm/instr\[0\] u_ppwm/instr\[1\] u_ppwm_u_ex__0805_/C VPWR
+ VGND sg13g2_nor2_2
XFILLER_38_543 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1078_ VGND VPWR u_ppwm_u_ex__1077_/Y u_ppwm_u_ex__1078_/Y u_ppwm_u_ex__1075_/Y
+ u_ppwm_u_ex__1029_/Y sg13g2_a21oi_2
Xu_ppwm_u_global_counter__067_ hold232/A net599 u_ppwm_u_global_counter__067_/B VPWR
+ VGND sg13g2_xnor2_1
XFILLER_41_719 VPWR VGND sg13g2_decap_8
XFILLER_40_207 VPWR VGND sg13g2_fill_1
XFILLER_34_793 VPWR VGND sg13g2_decap_8
XFILLER_22_955 VPWR VGND sg13g2_decap_8
XFILLER_21_498 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_0_369 VPWR VGND sg13g2_decap_8
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_29_532 VPWR VGND sg13g2_decap_8
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_16_204 VPWR VGND sg13g2_fill_1
XFILLER_44_568 VPWR VGND sg13g2_decap_8
XFILLER_25_771 VPWR VGND sg13g2_decap_8
XFILLER_24_270 VPWR VGND sg13g2_fill_2
XFILLER_9_915 VPWR VGND sg13g2_decap_8
XFILLER_13_955 VPWR VGND sg13g2_decap_8
XFILLER_33_51 VPWR VGND sg13g2_fill_2
XFILLER_40_796 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0730_ u_ppwm_u_mem__0730_/A u_ppwm_u_mem__1094_/A hold257/A u_ppwm_u_mem__0730_/Y
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__0661_ VPWR u_ppwm_u_mem__0661_/Y net251 VGND sg13g2_inv_1
XFILLER_4_631 VPWR VGND sg13g2_decap_8
Xhold3 hold3/A VPWR VGND net201 sg13g2_dlygate4sd3_1
XFILLER_48_852 VPWR VGND sg13g2_decap_8
XFILLER_47_340 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1001_ net506 VPWR u_ppwm_u_ex__1002_/B VGND net453 net350 sg13g2_o21ai_1
Xu_ppwm_u_mem__1213_ net125 VGND VPWR net291 hold109/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1144_ net74 VGND VPWR net321 hold139/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_535 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1075_ VGND VPWR net404 u_ppwm_u_mem__0617_/Y hold25/A u_ppwm_u_mem__1074_/Y
+ sg13g2_a21oi_1
XFILLER_15_270 VPWR VGND sg13g2_decap_4
XFILLER_31_730 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_ex__0716_ VPWR u_ppwm_u_ex__0716_/Y net364 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1217__61 VPWR VGND net61 sg13g2_tiehi
Xu_ppwm_u_mem__0928_ net504 VPWR u_ppwm_u_mem__0928_/Y VGND net417 net314 sg13g2_o21ai_1
Xu_ppwm_u_ex__0647_ u_ppwm_u_ex__0647_/Y hold231/A net450 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0859_ u_ppwm_u_mem__0858_/Y u_ppwm_u_mem__0856_/Y u_ppwm_u_mem__0852_/Y
+ fanout376/A VPWR VGND sg13g2_a21o_2
Xu_ppwm_u_ex__0578_ VPWR u_ppwm_u_ex__0578_/Y net247 VGND sg13g2_inv_1
XFILLER_39_885 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__119_ net507 VGND VPWR net635 u_ppwm_u_ex__1020_/B2 clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_41_516 VPWR VGND sg13g2_decap_8
XFILLER_26_568 VPWR VGND sg13g2_decap_8
XFILLER_22_752 VPWR VGND sg13g2_decap_8
XFILLER_34_590 VPWR VGND sg13g2_decap_8
XFILLER_21_240 VPWR VGND sg13g2_decap_4
XFILLER_21_273 VPWR VGND sg13g2_decap_8
XFILLER_10_969 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_8
XFILLER_0_177 VPWR VGND sg13g2_decap_8
XFILLER_48_148 VPWR VGND sg13g2_decap_8
XFILLER_0_199 VPWR VGND sg13g2_decap_8
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_17_502 VPWR VGND sg13g2_decap_8
XFILLER_28_84 VPWR VGND sg13g2_decap_4
XFILLER_29_384 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_decap_8
XFILLER_17_579 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1112__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_44_387 VPWR VGND sg13g2_fill_2
XFILLER_32_549 VPWR VGND sg13g2_decap_8
XFILLER_13_752 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_4
XFILLER_9_712 VPWR VGND sg13g2_decap_8
XFILLER_12_251 VPWR VGND sg13g2_fill_1
XFILLER_12_262 VPWR VGND sg13g2_decap_4
XFILLER_40_593 VPWR VGND sg13g2_decap_8
XFILLER_8_266 VPWR VGND sg13g2_fill_2
XFILLER_9_789 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0713_ VPWR u_ppwm_u_mem__0713_/Y net532 VGND sg13g2_inv_1
XFILLER_5_962 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0644_ VPWR u_ppwm_u_mem__0644_/Y net319 VGND sg13g2_inv_1
XFILLER_36_844 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1127_ net108 VGND VPWR u_ppwm_u_mem__1127_/D hold133/A clknet_5_18__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_343 VPWR VGND sg13g2_fill_1
XFILLER_23_538 VPWR VGND sg13g2_decap_8
XFILLER_35_376 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1058_ net488 VPWR u_ppwm_u_mem__1058_/Y VGND net402 hold103/A sg13g2_o21ai_1
Xhold211 hold211/A VPWR VGND net579 sg13g2_dlygate4sd3_1
Xhold200 hold200/A VPWR VGND net568 sg13g2_dlygate4sd3_1
Xhold233 hold233/A VPWR VGND net601 sg13g2_dlygate4sd3_1
Xhold222 hold222/A VPWR VGND net590 sg13g2_dlygate4sd3_1
Xhold244 hold244/A VPWR VGND net612 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
Xhold255 hold255/A VPWR VGND net623 sg13g2_dlygate4sd3_1
Xhold277 hold277/A VPWR VGND net645 sg13g2_dlygate4sd3_1
Xhold266 hold266/A VPWR VGND net634 sg13g2_dlygate4sd3_1
Xhold299 hold299/A VPWR VGND net667 sg13g2_dlygate4sd3_1
Xhold288 hold288/A VPWR VGND net656 sg13g2_dlygate4sd3_1
XFILLER_46_608 VPWR VGND sg13g2_decap_8
XFILLER_26_310 VPWR VGND sg13g2_fill_2
XFILLER_27_844 VPWR VGND sg13g2_decap_8
XFILLER_39_682 VPWR VGND sg13g2_decap_8
XFILLER_42_803 VPWR VGND sg13g2_decap_8
XFILLER_14_538 VPWR VGND sg13g2_decap_8
XFILLER_10_766 VPWR VGND sg13g2_decap_8
XFILLER_6_737 VPWR VGND sg13g2_decap_8
XFILLER_2_954 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_37_619 VPWR VGND sg13g2_decap_8
XFILLER_18_855 VPWR VGND sg13g2_decap_8
XFILLER_45_674 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0981_ u_ppwm_u_ex__0981_/Y net356 net445 net362 fanout466/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_33_869 VPWR VGND sg13g2_decap_8
XFILLER_41_880 VPWR VGND sg13g2_decap_8
XFILLER_20_508 VPWR VGND sg13g2_decap_8
XFILLER_9_586 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0627_ VPWR u_ppwm_u_mem__0627_/Y net312 VGND sg13g2_inv_1
XFILLER_49_991 VPWR VGND sg13g2_decap_8
XFILLER_36_641 VPWR VGND sg13g2_decap_8
XFILLER_23_313 VPWR VGND sg13g2_decap_8
XFILLER_24_836 VPWR VGND sg13g2_decap_8
XFILLER_35_173 VPWR VGND sg13g2_fill_1
XFILLER_2_217 VPWR VGND sg13g2_fill_2
Xfanout510 net511 net510 VPWR VGND sg13g2_buf_8
XFILLER_47_928 VPWR VGND sg13g2_decap_8
XFILLER_46_405 VPWR VGND sg13g2_decap_8
XFILLER_15_803 VPWR VGND sg13g2_decap_8
XFILLER_27_641 VPWR VGND sg13g2_decap_8
XFILLER_42_600 VPWR VGND sg13g2_decap_8
XFILLER_14_313 VPWR VGND sg13g2_decap_8
XFILLER_42_677 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__220_ VGND VPWR u_ppwm_u_pwm__183_/A hold40/A u_ppwm_u_pwm__221_/B u_ppwm_u_pwm__219_/Y
+ sg13g2_a21oi_1
XFILLER_22_390 VPWR VGND sg13g2_decap_8
XFILLER_41_73 VPWR VGND sg13g2_fill_2
XFILLER_41_62 VPWR VGND sg13g2_fill_1
XFILLER_6_534 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__151_ net490 VPWR u_ppwm_u_pwm__151_/Y VGND net458 net389 sg13g2_o21ai_1
XFILLER_10_563 VPWR VGND sg13g2_decap_8
XFILLER_29_1015 VPWR VGND sg13g2_decap_8
XFILLER_2_751 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_38_928 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_46_972 VPWR VGND sg13g2_decap_8
XFILLER_18_652 VPWR VGND sg13g2_decap_8
XFILLER_45_471 VPWR VGND sg13g2_decap_8
XFILLER_17_195 VPWR VGND sg13g2_fill_2
XFILLER_21_806 VPWR VGND sg13g2_decap_8
XFILLER_32_154 VPWR VGND sg13g2_decap_8
XFILLER_33_666 VPWR VGND sg13g2_decap_8
XFILLER_36_1019 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0964_ u_ppwm_u_ex__0964_/B u_ppwm_u_ex__1086_/A net352 u_ppwm_u_ex__0964_/Y
+ VPWR VGND u_ppwm_u_ex__0964_/D sg13g2_nand4_1
Xu_ppwm_u_mem__1164__153 VPWR VGND net153 sg13g2_tiehi
Xu_ppwm_u_ex__0895_ u_ppwm_u_ex__0896_/B net365 hold240/A net367 hold222/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_9_383 VPWR VGND sg13g2_fill_1
XFILLER_29_917 VPWR VGND sg13g2_decap_8
XFILLER_43_419 VPWR VGND sg13g2_decap_8
XFILLER_37_983 VPWR VGND sg13g2_decap_8
XFILLER_23_110 VPWR VGND sg13g2_decap_8
XFILLER_24_633 VPWR VGND sg13g2_decap_8
XFILLER_11_338 VPWR VGND sg13g2_decap_8
XFILLER_12_839 VPWR VGND sg13g2_decap_8
XFILLER_7_309 VPWR VGND sg13g2_decap_8
XFILLER_20_872 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_fill_1
XFILLER_3_548 VPWR VGND sg13g2_decap_8
Xfanout362 net363 net362 VPWR VGND sg13g2_buf_8
Xfanout373 net374 net373 VPWR VGND sg13g2_buf_8
Xfanout384 net385 net384 VPWR VGND sg13g2_buf_8
Xfanout351 fanout351/A net351 VPWR VGND sg13g2_buf_8
XFILLER_47_725 VPWR VGND sg13g2_decap_8
Xfanout395 net396 net395 VPWR VGND sg13g2_buf_2
XFILLER_19_449 VPWR VGND sg13g2_fill_1
XFILLER_46_279 VPWR VGND sg13g2_decap_8
XFILLER_15_600 VPWR VGND sg13g2_decap_8
XFILLER_34_419 VPWR VGND sg13g2_fill_1
XFILLER_27_482 VPWR VGND sg13g2_fill_1
XFILLER_43_986 VPWR VGND sg13g2_decap_8
XFILLER_15_677 VPWR VGND sg13g2_decap_8
XFILLER_42_474 VPWR VGND sg13g2_decap_8
XFILLER_14_187 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0961_ VGND VPWR net430 u_ppwm_u_mem__0674_/Y hold48/A u_ppwm_u_mem__0960_/Y
+ sg13g2_a21oi_1
XFILLER_11_861 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_decap_8
XFILLER_7_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__203_ u_ppwm_u_pwm__196_/Y VPWR u_ppwm_u_pwm__203_/Y VGND u_ppwm_u_pwm__200_/Y
+ u_ppwm_u_pwm__202_/X sg13g2_o21ai_1
Xu_ppwm_u_mem__0892_ net516 VPWR u_ppwm_u_mem__0892_/Y VGND net435 hold183/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0680_ VPWR VGND u_ppwm_u_ex__0672_/Y u_ppwm_u_ex__0679_/Y u_ppwm_u_ex__0678_/Y
+ u_ppwm_u_ex__0678_/B u_ppwm_u_ex__0680_/Y u_ppwm_u_ex__0676_/Y sg13g2_a221oi_1
Xu_ppwm_u_pwm__134_ VPWR u_ppwm_u_pwm__134_/Y net215 VGND sg13g2_inv_1
XFILLER_28_4 VPWR VGND sg13g2_fill_2
XFILLER_37_202 VPWR VGND sg13g2_decap_4
XFILLER_38_725 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1094_ VPWR VGND hold217/A u_ppwm_u_ex__1093_/Y net355 net441 u_ppwm_u_ex__1094_/Y
+ net356 sg13g2_a221oi_1
Xu_ppwm_u_global_counter__083_ hold208/A net575 u_ppwm_u_global_counter__083_/B VPWR
+ VGND sg13g2_xnor2_1
XFILLER_25_408 VPWR VGND sg13g2_decap_4
XFILLER_37_268 VPWR VGND sg13g2_fill_2
XFILLER_21_603 VPWR VGND sg13g2_decap_8
XFILLER_34_975 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0947_ u_ppwm_u_ex__0947_/X net352 u_ppwm_u_ex__1071_/A u_ppwm_u_ex__0947_/C
+ VPWR VGND sg13g2_and3_1
Xu_ppwm_u_ex__0878_ u_ppwm_u_ex__0877_/Y VPWR u_ppwm_u_ex__0879_/B VGND net462 net354
+ sg13g2_o21ai_1
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_714 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__242__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_28_257 VPWR VGND sg13g2_decap_8
XFILLER_37_780 VPWR VGND sg13g2_decap_8
XFILLER_24_430 VPWR VGND sg13g2_fill_2
XFILLER_25_953 VPWR VGND sg13g2_decap_8
XFILLER_40_901 VPWR VGND sg13g2_decap_8
XFILLER_12_636 VPWR VGND sg13g2_decap_8
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_8_618 VPWR VGND sg13g2_decap_8
XFILLER_4_813 VPWR VGND sg13g2_decap_8
XFILLER_3_334 VPWR VGND sg13g2_fill_2
XFILLER_47_522 VPWR VGND sg13g2_decap_8
XFILLER_19_213 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1160_ net161 VGND VPWR net272 hold185/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1091_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1091_/B u_ppwm_u_mem__1091_/C
+ u_ppwm_u_mem__1220_/D VPWR VGND sg13g2_nor3_1
XFILLER_35_717 VPWR VGND sg13g2_decap_8
XFILLER_16_986 VPWR VGND sg13g2_decap_8
XFILLER_31_912 VPWR VGND sg13g2_decap_8
XFILLER_43_783 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0801_ u_ppwm_u_ex__0799_/A u_ppwm_u_ex__0800_/X net370 u_ppwm_u_ex__0801_/X
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_989 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0732_ net449 u_ppwm_u_ex__0732_/B u_ppwm_u_ex__0732_/C u_ppwm_u_ex__0732_/Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_7_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0944_ net511 VPWR u_ppwm_u_mem__0944_/Y VGND net429 hold188/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0663_ net370 u_ppwm_u_ex__0715_/B u_ppwm_u_ex__0663_/C u_ppwm_u_ex__0663_/D
+ u_ppwm_u_ex__0769_/A VPWR VGND sg13g2_and4_1
Xu_ppwm_u_mem__0875_ VGND VPWR net423 u_ppwm_u_mem__0717_/Y u_ppwm_u_mem__1114_/D
+ u_ppwm_u_mem__0874_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__1122__118 VPWR VGND net118 sg13g2_tiehi
Xu_ppwm_u_ex__0594_ net469 u_ppwm_u_ex__0622_/B net468 u_ppwm_u_ex__0636_/A VPWR VGND
+ sg13g2_nand3_1
XFILLER_38_522 VPWR VGND sg13g2_decap_8
XFILLER_19_0 VPWR VGND sg13g2_fill_1
XFILLER_38_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1077_ u_ppwm_u_ex__1077_/Y u_ppwm_u_ex__1077_/B u_ppwm_u_ex__1052_/Y
+ VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_global_counter__066_ u_ppwm_u_global_counter__066_/A u_ppwm_u_global_counter__067_/B
+ u_ppwm_u_global_counter__068_/B VPWR VGND sg13g2_nor2_1
XFILLER_22_934 VPWR VGND sg13g2_decap_8
XFILLER_34_772 VPWR VGND sg13g2_decap_8
XFILLER_21_477 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_0_348 VPWR VGND sg13g2_decap_8
XFILLER_29_588 VPWR VGND sg13g2_decap_8
XFILLER_44_547 VPWR VGND sg13g2_decap_8
XFILLER_25_750 VPWR VGND sg13g2_decap_8
XFILLER_13_934 VPWR VGND sg13g2_decap_8
XFILLER_40_775 VPWR VGND sg13g2_decap_8
XFILLER_32_1011 VPWR VGND sg13g2_decap_8
XFILLER_33_63 VPWR VGND sg13g2_fill_2
XFILLER_4_610 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1225__175 VPWR VGND net175 sg13g2_tiehi
Xu_ppwm_u_mem__0660_ VPWR u_ppwm_u_mem__0660_/Y net303 VGND sg13g2_inv_1
XFILLER_3_142 VPWR VGND sg13g2_decap_8
XFILLER_4_687 VPWR VGND sg13g2_decap_8
Xhold4 hold4/A VPWR VGND net202 sg13g2_dlygate4sd3_1
XFILLER_48_831 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1000_ u_ppwm_u_ex__1000_/A u_ppwm_u_ex__1000_/B u_ppwm_u_ex__1000_/C
+ u_ppwm_u_ex__1000_/D u_ppwm_u_ex__1002_/A VPWR VGND sg13g2_nor4_1
Xu_ppwm_u_mem__1212_ net141 VGND VPWR net308 hold145/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1143_ net76 VGND VPWR net338 hold22/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_396 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1074_ net494 VPWR u_ppwm_u_mem__1074_/Y VGND net403 hold92/A sg13g2_o21ai_1
XFILLER_43_580 VPWR VGND sg13g2_decap_8
XFILLER_16_783 VPWR VGND sg13g2_decap_8
XFILLER_15_282 VPWR VGND sg13g2_fill_1
XFILLER_31_786 VPWR VGND sg13g2_decap_8
XFILLER_8_982 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0715_ net377 u_ppwm_u_ex__0715_/B fanout365/A VPWR VGND sg13g2_and2_1
Xu_ppwm_u_mem__0927_ VGND VPWR net417 u_ppwm_u_mem__0691_/Y u_ppwm_u_mem__1140_/D
+ u_ppwm_u_mem__0926_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0646_ VPWR VGND u_ppwm_u_ex__0644_/Y u_ppwm_u_ex__0645_/Y u_ppwm_u_ex__0643_/Y
+ net451 u_ppwm_u_ex__0646_/Y u_ppwm_u_ex__0591_/Y sg13g2_a221oi_1
Xu_ppwm_u_mem__0858_ VGND VPWR net393 u_ppwm_u_mem__0857_/X u_ppwm_u_mem__0858_/Y
+ net467 sg13g2_a21oi_1
Xu_ppwm_u_ex__0577_ net463 u_ppwm_u_ex__0850_/A VPWR VGND sg13g2_inv_4
Xu_ppwm_u_mem__0789_ u_ppwm_u_mem__0788_/Y VPWR u_ppwm_u_mem__0789_/Y VGND u_ppwm_u_mem__0709_/Y
+ net485 sg13g2_o21ai_1
XFILLER_39_864 VPWR VGND sg13g2_decap_8
XFILLER_38_363 VPWR VGND sg13g2_fill_2
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__118_ net509 VGND VPWR u_ppwm_u_global_counter__118_/D hold265/A
+ clknet_5_17__leaf_clk sg13g2_dfrbpq_2
XFILLER_26_547 VPWR VGND sg13g2_decap_8
XFILLER_22_731 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_919 VPWR VGND sg13g2_decap_8
XFILLER_10_948 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_49_606 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__248__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_48_138 VPWR VGND sg13g2_fill_1
XFILLER_45_856 VPWR VGND sg13g2_decap_8
XFILLER_17_558 VPWR VGND sg13g2_decap_8
XFILLER_13_731 VPWR VGND sg13g2_decap_8
XFILLER_40_572 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1124__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_9_768 VPWR VGND sg13g2_decap_8
XFILLER_5_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0712_ VPWR u_ppwm_u_mem__0712_/Y net293 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0643_ VPWR u_ppwm_u_mem__0643_/Y net580 VGND sg13g2_inv_1
XFILLER_5_78 VPWR VGND sg13g2_decap_4
XFILLER_4_484 VPWR VGND sg13g2_decap_8
XFILLER_36_823 VPWR VGND sg13g2_decap_8
XFILLER_47_193 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1126_ net110 VGND VPWR net332 hold161/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_517 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1057_ VGND VPWR net402 u_ppwm_u_mem__0626_/Y hold104/A u_ppwm_u_mem__1056_/Y
+ sg13g2_a21oi_1
XFILLER_16_580 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1115__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_31_583 VPWR VGND sg13g2_decap_8
Xhold201 hold201/A VPWR VGND net569 sg13g2_dlygate4sd3_1
Xhold212 hold212/A VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold223 hold223/A VPWR VGND net591 sg13g2_dlygate4sd3_1
Xhold234 hold234/A VPWR VGND net602 sg13g2_dlygate4sd3_1
Xhold278 hold278/A VPWR VGND net646 sg13g2_dlygate4sd3_1
Xhold267 hold267/A VPWR VGND net635 sg13g2_dlygate4sd3_1
Xhold245 hold245/A VPWR VGND net613 sg13g2_dlygate4sd3_1
Xhold256 hold256/A VPWR VGND net624 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0629_ u_ppwm_u_ex__0624_/Y VPWR u_ppwm_u_ex__0629_/Y VGND u_ppwm_u_ex__0636_/B
+ u_ppwm_u_ex__0628_/Y sg13g2_o21ai_1
Xhold289 hold289/A VPWR VGND net657 sg13g2_dlygate4sd3_1
XFILLER_39_661 VPWR VGND sg13g2_decap_8
XFILLER_27_823 VPWR VGND sg13g2_decap_8
XFILLER_14_517 VPWR VGND sg13g2_decap_8
XFILLER_42_859 VPWR VGND sg13g2_decap_8
XFILLER_10_745 VPWR VGND sg13g2_decap_8
XFILLER_14_65 VPWR VGND sg13g2_decap_8
XFILLER_6_716 VPWR VGND sg13g2_decap_8
XFILLER_5_215 VPWR VGND sg13g2_fill_1
XFILLER_2_933 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_18_834 VPWR VGND sg13g2_decap_8
XFILLER_45_653 VPWR VGND sg13g2_decap_8
XFILLER_17_355 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0980_ u_ppwm_u_ex__0980_/Y hold207/A net355 VPWR VGND sg13g2_nand2_1
XFILLER_33_848 VPWR VGND sg13g2_decap_8
XFILLER_32_369 VPWR VGND sg13g2_fill_1
XFILLER_9_565 VPWR VGND sg13g2_decap_8
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0626_ VPWR u_ppwm_u_mem__0626_/Y net301 VGND sg13g2_inv_1
XFILLER_49_970 VPWR VGND sg13g2_decap_8
XFILLER_36_620 VPWR VGND sg13g2_decap_8
XFILLER_24_815 VPWR VGND sg13g2_decap_8
XFILLER_36_697 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1109_ net144 VGND VPWR net342 hold209/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_892 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1103__45 VPWR VGND net45 sg13g2_tiehi
Xfanout500 net504 net500 VPWR VGND sg13g2_buf_8
Xfanout511 net512 net511 VPWR VGND sg13g2_buf_8
XFILLER_47_907 VPWR VGND sg13g2_decap_8
XFILLER_27_620 VPWR VGND sg13g2_decap_8
XFILLER_27_697 VPWR VGND sg13g2_decap_8
XFILLER_42_656 VPWR VGND sg13g2_decap_8
XFILLER_15_859 VPWR VGND sg13g2_decap_8
XFILLER_25_42 VPWR VGND sg13g2_fill_2
XFILLER_26_196 VPWR VGND sg13g2_decap_4
XFILLER_23_881 VPWR VGND sg13g2_decap_8
XFILLER_41_41 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__150_ VGND VPWR u_ppwm_u_pwm__213_/B net389 hold10/A u_ppwm_u_pwm__149_/Y
+ sg13g2_a21oi_1
XFILLER_10_542 VPWR VGND sg13g2_decap_8
XFILLER_6_513 VPWR VGND sg13g2_decap_8
XFILLER_2_730 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_38_907 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_46_951 VPWR VGND sg13g2_decap_8
XFILLER_18_631 VPWR VGND sg13g2_decap_8
XFILLER_45_450 VPWR VGND sg13g2_decap_8
XFILLER_32_122 VPWR VGND sg13g2_fill_2
XFILLER_33_645 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0963_ VGND VPWR net663 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0964_/D u_ppwm_u_ex__0962_/Y
+ sg13g2_a21oi_1
XFILLER_14_881 VPWR VGND sg13g2_decap_8
XFILLER_32_166 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0894_ VPWR VGND u_ppwm_u_ex__0797_/Y u_ppwm_u_ex__0890_/Y u_ppwm_u_ex__0893_/X
+ u_ppwm_u_ex__0790_/Y u_ppwm_u_ex__1035_/A u_ppwm_u_ex__0847_/A sg13g2_a221oi_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1187__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_37_962 VPWR VGND sg13g2_decap_8
XFILLER_24_612 VPWR VGND sg13g2_decap_8
XFILLER_36_472 VPWR VGND sg13g2_fill_1
XFILLER_12_818 VPWR VGND sg13g2_decap_8
XFILLER_24_689 VPWR VGND sg13g2_decap_8
XFILLER_11_317 VPWR VGND sg13g2_fill_2
XFILLER_20_851 VPWR VGND sg13g2_decap_8
XFILLER_3_527 VPWR VGND sg13g2_decap_8
XFILLER_11_77 VPWR VGND sg13g2_fill_2
XFILLER_47_704 VPWR VGND sg13g2_decap_8
Xfanout352 net353 net352 VPWR VGND sg13g2_buf_8
Xfanout363 fanout363/A net363 VPWR VGND sg13g2_buf_8
Xfanout374 fanout376/A net374 VPWR VGND sg13g2_buf_8
XFILLER_19_406 VPWR VGND sg13g2_fill_1
Xfanout385 net387 net385 VPWR VGND sg13g2_buf_8
Xfanout396 net397 net396 VPWR VGND sg13g2_buf_1
XFILLER_46_258 VPWR VGND sg13g2_decap_8
XFILLER_27_472 VPWR VGND sg13g2_fill_2
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_34_409 VPWR VGND sg13g2_fill_1
XFILLER_43_965 VPWR VGND sg13g2_decap_8
XFILLER_42_453 VPWR VGND sg13g2_decap_8
XFILLER_15_656 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0960_ net511 VPWR u_ppwm_u_mem__0960_/Y VGND net430 hold173/A sg13g2_o21ai_1
XFILLER_11_840 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__202_ u_ppwm_u_pwm__202_/A u_ppwm_u_pwm__202_/B u_ppwm_u_pwm__202_/C
+ u_ppwm_u_pwm__202_/D u_ppwm_u_pwm__202_/X VPWR VGND sg13g2_or4_1
XFILLER_7_822 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0891_ VGND VPWR net434 u_ppwm_u_mem__0709_/Y hold184/A u_ppwm_u_mem__0890_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__133_ VPWR u_ppwm_u_pwm__133_/Y net203 VGND sg13g2_inv_1
XFILLER_7_899 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_fill_2
XFILLER_42_1013 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1194__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_38_704 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1093_ VGND VPWR net381 net370 u_ppwm_u_ex__1093_/Y u_ppwm_u_ex__0683_/A
+ sg13g2_a21oi_1
Xu_ppwm_u_global_counter__082_ net639 net575 net201 hold272/A VPWR VGND u_ppwm_u_global_counter__082_/D
+ sg13g2_nand4_1
XFILLER_37_247 VPWR VGND sg13g2_fill_2
XFILLER_19_995 VPWR VGND sg13g2_decap_8
XFILLER_33_420 VPWR VGND sg13g2_fill_2
XFILLER_34_954 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0946_ u_ppwm_u_ex__0945_/Y u_ppwm_u_ex__0944_/Y net361 u_ppwm_u_ex__0947_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_21_659 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__235__197 VPWR VGND net197 sg13g2_tiehi
Xu_ppwm_u_ex__0877_ u_ppwm_u_ex__0877_/B u_ppwm_u_ex__0877_/C fanout354/A u_ppwm_u_ex__0877_/Y
+ VPWR VGND u_ppwm_u_ex__0877_/D sg13g2_nand4_1
XFILLER_44_729 VPWR VGND sg13g2_decap_8
XFILLER_43_228 VPWR VGND sg13g2_decap_4
XFILLER_25_932 VPWR VGND sg13g2_decap_8
XFILLER_24_442 VPWR VGND sg13g2_fill_1
XFILLER_12_615 VPWR VGND sg13g2_decap_8
XFILLER_24_486 VPWR VGND sg13g2_decap_8
XFILLER_40_957 VPWR VGND sg13g2_decap_8
XFILLER_7_129 VPWR VGND sg13g2_decap_4
XFILLER_4_869 VPWR VGND sg13g2_decap_8
XFILLER_3_313 VPWR VGND sg13g2_decap_4
XFILLER_47_501 VPWR VGND sg13g2_decap_8
XFILLER_47_578 VPWR VGND sg13g2_decap_8
XFILLER_47_95 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1090_ net638 u_ppwm_u_mem__1090_/B u_ppwm_u_mem__1091_/C VPWR VGND
+ sg13g2_and2_1
XFILLER_34_206 VPWR VGND sg13g2_fill_1
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_43_762 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_16_965 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0800_ net462 net450 net386 u_ppwm_u_ex__0800_/X VPWR VGND sg13g2_mux2_1
XFILLER_31_968 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0943_ VGND VPWR net427 u_ppwm_u_mem__0683_/Y hold189/A u_ppwm_u_mem__0942_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0731_ u_ppwm_u_ex__0730_/Y VPWR u_ppwm_u_ex__0731_/Y VGND u_ppwm_u_ex__0723_/Y
+ u_ppwm_u_ex__0725_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__0662_ VGND VPWR u_ppwm_u_ex__0973_/A net441 u_ppwm_u_ex__0663_/D u_ppwm_u_ex__0658_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0874_ net513 VPWR u_ppwm_u_mem__0874_/Y VGND net423 net284 sg13g2_o21ai_1
XFILLER_7_696 VPWR VGND sg13g2_decap_8
XFILLER_6_184 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0593_ net473 net480 u_ppwm_u_ex__0622_/B VPWR VGND sg13g2_and2_1
XFILLER_40_4 VPWR VGND sg13g2_fill_1
XFILLER_3_891 VPWR VGND sg13g2_decap_8
XFILLER_38_501 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__065_ hold288/A net443 u_ppwm_u_global_counter__070_/A VPWR
+ VGND sg13g2_xnor2_1
XFILLER_26_729 VPWR VGND sg13g2_decap_8
XFILLER_38_578 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1076_ net373 VPWR u_ppwm_u_ex__1077_/B VGND hold294/A net448 sg13g2_o21ai_1
XFILLER_19_792 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1180__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_34_751 VPWR VGND sg13g2_decap_8
XFILLER_22_913 VPWR VGND sg13g2_decap_8
XFILLER_21_423 VPWR VGND sg13g2_decap_8
XFILLER_33_294 VPWR VGND sg13g2_fill_2
XFILLER_21_456 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0929_ VPWR VGND u_ppwm_u_ex__0797_/Y u_ppwm_u_ex__0927_/Y u_ppwm_u_ex__0928_/X
+ u_ppwm_u_ex__0790_/Y u_ppwm_u_ex__1061_/A u_ppwm_u_ex__0893_/X sg13g2_a221oi_1
XFILLER_49_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_327 VPWR VGND sg13g2_decap_8
XFILLER_29_567 VPWR VGND sg13g2_decap_8
XFILLER_44_526 VPWR VGND sg13g2_decap_8
XFILLER_17_65 VPWR VGND sg13g2_fill_2
XFILLER_17_87 VPWR VGND sg13g2_decap_8
XFILLER_13_913 VPWR VGND sg13g2_decap_8
XFILLER_31_209 VPWR VGND sg13g2_fill_2
XFILLER_40_754 VPWR VGND sg13g2_decap_8
XFILLER_4_666 VPWR VGND sg13g2_decap_8
XFILLER_48_810 VPWR VGND sg13g2_decap_8
XFILLER_0_894 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_1
Xhold5 hold5/A VPWR VGND net203 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1211_ net152 VGND VPWR net344 hold169/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_887 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1142_ net78 VGND VPWR net221 hold177/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_375 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1073_ VGND VPWR net406 u_ppwm_u_mem__0618_/Y hold93/A u_ppwm_u_mem__1072_/Y
+ sg13g2_a21oi_1
XFILLER_16_762 VPWR VGND sg13g2_decap_8
XFILLER_31_765 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0714_ u_ppwm_u_ex__0714_/A u_ppwm_u_ex__0714_/B u_ppwm_u_ex__0714_/C
+ u_ppwm_u_ex__0714_/Y VPWR VGND sg13g2_nor3_1
XFILLER_8_961 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0926_ net502 VPWR u_ppwm_u_mem__0926_/Y VGND net417 net226 sg13g2_o21ai_1
XFILLER_7_493 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0645_ net444 net453 u_ppwm_u_ex__0645_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0857_ net397 u_ppwm_u_mem__0705_/Y u_ppwm_u_mem__0719_/Y u_ppwm_u_mem__0698_/Y
+ u_ppwm_u_mem__0712_/Y net484 u_ppwm_u_mem__0857_/X VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_ex__0576_ VPWR u_ppwm_u_ex__0576_/Y net462 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0788_ u_ppwm_u_mem__0788_/Y hold156/A net485 VPWR VGND sg13g2_nand2_1
XFILLER_31_0 VPWR VGND sg13g2_fill_2
XFILLER_39_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__117_ net508 VGND VPWR net641 u_ppwm_u_ex__0998_/B2 clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_526 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1059_ u_ppwm_u_ex__1059_/Y fanout355/A hold286/A net362 net457 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_22_710 VPWR VGND sg13g2_decap_8
XFILLER_16_1007 VPWR VGND sg13g2_decap_8
XFILLER_21_220 VPWR VGND sg13g2_fill_1
XFILLER_10_927 VPWR VGND sg13g2_decap_8
XFILLER_22_787 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_4
XFILLER_45_835 VPWR VGND sg13g2_decap_8
XFILLER_17_537 VPWR VGND sg13g2_decap_8
XFILLER_29_386 VPWR VGND sg13g2_fill_1
XFILLER_44_356 VPWR VGND sg13g2_decap_4
XFILLER_13_710 VPWR VGND sg13g2_decap_8
XFILLER_40_551 VPWR VGND sg13g2_decap_8
XFILLER_13_787 VPWR VGND sg13g2_decap_8
XFILLER_9_747 VPWR VGND sg13g2_decap_8
XFILLER_12_297 VPWR VGND sg13g2_fill_1
XFILLER_5_920 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0711_ VPWR u_ppwm_u_mem__0711_/Y net275 VGND sg13g2_inv_1
XFILLER_5_997 VPWR VGND sg13g2_decap_8
XFILLER_4_463 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0642_ VPWR u_ppwm_u_mem__0642_/Y net326 VGND sg13g2_inv_1
XFILLER_0_691 VPWR VGND sg13g2_decap_8
XFILLER_36_802 VPWR VGND sg13g2_decap_8
XFILLER_48_684 VPWR VGND sg13g2_decap_8
XFILLER_39_1018 VPWR VGND sg13g2_decap_8
XFILLER_36_879 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1125_ net112 VGND VPWR net530 hold190/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1056_ net488 VPWR u_ppwm_u_mem__1056_/Y VGND net402 hold114/A sg13g2_o21ai_1
XFILLER_44_890 VPWR VGND sg13g2_decap_8
XFILLER_31_562 VPWR VGND sg13g2_decap_8
Xhold202 hold202/A VPWR VGND net570 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0909_ VGND VPWR net436 u_ppwm_u_mem__0700_/Y hold65/A u_ppwm_u_mem__0908_/Y
+ sg13g2_a21oi_1
Xhold224 hold224/A VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold235 hold235/A VPWR VGND net603 sg13g2_dlygate4sd3_1
Xhold213 hold213/A VPWR VGND net581 sg13g2_dlygate4sd3_1
Xhold268 hold268/A VPWR VGND net636 sg13g2_dlygate4sd3_1
Xhold257 hold257/A VPWR VGND net625 sg13g2_dlygate4sd3_1
Xhold246 hold246/A VPWR VGND net614 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0628_ u_ppwm_u_ex__0628_/Y u_ppwm_u_ex__0628_/A u_ppwm_u_ex__0628_/B
+ VPWR VGND sg13g2_xnor2_1
Xhold279 hold279/A VPWR VGND net647 sg13g2_dlygate4sd3_1
XFILLER_22_1011 VPWR VGND sg13g2_decap_8
XFILLER_27_802 VPWR VGND sg13g2_decap_8
XFILLER_39_640 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_fill_1
XFILLER_26_345 VPWR VGND sg13g2_decap_8
XFILLER_27_879 VPWR VGND sg13g2_decap_8
XFILLER_42_838 VPWR VGND sg13g2_decap_8
XFILLER_41_304 VPWR VGND sg13g2_fill_2
XFILLER_14_11 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1111__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_10_724 VPWR VGND sg13g2_decap_8
XFILLER_22_584 VPWR VGND sg13g2_decap_8
XFILLER_2_912 VPWR VGND sg13g2_decap_8
XFILLER_2_989 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_18_813 VPWR VGND sg13g2_decap_8
XFILLER_45_632 VPWR VGND sg13g2_decap_8
XFILLER_33_827 VPWR VGND sg13g2_decap_8
XFILLER_26_890 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1132__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_9_544 VPWR VGND sg13g2_decap_8
XFILLER_13_584 VPWR VGND sg13g2_decap_8
XFILLER_5_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0625_ VPWR u_ppwm_u_mem__0625_/Y net258 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1197__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_48_481 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1108_ net146 VGND VPWR net578 u_ppwm_u_mem__1108_/Q clknet_5_23__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_164 VPWR VGND sg13g2_fill_1
XFILLER_36_676 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1039_ VGND VPWR net407 u_ppwm_u_mem__0635_/Y u_ppwm_u_mem__1196_/D
+ u_ppwm_u_mem__1038_/Y sg13g2_a21oi_1
XFILLER_32_871 VPWR VGND sg13g2_decap_8
XFILLER_3_709 VPWR VGND sg13g2_decap_8
XFILLER_2_219 VPWR VGND sg13g2_fill_1
Xfanout501 net504 net501 VPWR VGND sg13g2_buf_8
Xfanout512 net518 net512 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_pwm__245__188 VPWR VGND net188 sg13g2_tiehi
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_142 VPWR VGND sg13g2_fill_2
XFILLER_27_676 VPWR VGND sg13g2_decap_8
XFILLER_42_635 VPWR VGND sg13g2_decap_8
XFILLER_15_838 VPWR VGND sg13g2_decap_8
XFILLER_26_175 VPWR VGND sg13g2_decap_8
XFILLER_14_359 VPWR VGND sg13g2_fill_1
XFILLER_23_860 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_8
XFILLER_10_521 VPWR VGND sg13g2_decap_8
XFILLER_41_75 VPWR VGND sg13g2_fill_1
XFILLER_6_569 VPWR VGND sg13g2_decap_8
XFILLER_10_598 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_2_786 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_2_58 VPWR VGND sg13g2_decap_8
XFILLER_18_610 VPWR VGND sg13g2_decap_8
XFILLER_46_930 VPWR VGND sg13g2_decap_8
XFILLER_17_153 VPWR VGND sg13g2_fill_2
XFILLER_18_687 VPWR VGND sg13g2_decap_8
XFILLER_32_101 VPWR VGND sg13g2_fill_2
XFILLER_33_624 VPWR VGND sg13g2_decap_8
XFILLER_14_860 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0962_ net361 u_ppwm_u_ex__0962_/B u_ppwm_u_ex__0962_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0893_ u_ppwm_u_ex__0870_/Y u_ppwm_u_ex__0892_/Y net377 u_ppwm_u_ex__0893_/X
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_591 VPWR VGND sg13g2_decap_8
XFILLER_37_941 VPWR VGND sg13g2_decap_8
XFILLER_24_668 VPWR VGND sg13g2_decap_8
XFILLER_20_830 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
XFILLER_3_506 VPWR VGND sg13g2_decap_8
Xfanout353 net354 net353 VPWR VGND sg13g2_buf_8
Xfanout364 fanout365/A net364 VPWR VGND sg13g2_buf_8
Xfanout375 fanout376/A net375 VPWR VGND sg13g2_buf_8
XFILLER_46_204 VPWR VGND sg13g2_decap_8
Xfanout386 net387 net386 VPWR VGND sg13g2_buf_8
XFILLER_19_418 VPWR VGND sg13g2_fill_2
Xfanout397 fanout397/A net397 VPWR VGND sg13g2_buf_8
XFILLER_46_237 VPWR VGND sg13g2_decap_8
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_43_944 VPWR VGND sg13g2_decap_8
XFILLER_14_101 VPWR VGND sg13g2_decap_8
XFILLER_15_635 VPWR VGND sg13g2_decap_8
XFILLER_42_432 VPWR VGND sg13g2_decap_8
XFILLER_30_616 VPWR VGND sg13g2_decap_8
XFILLER_7_801 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__201_ hold204/A hold5/A u_ppwm_u_pwm__202_/D VPWR VGND sg13g2_nor2b_1
XFILLER_6_300 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0890_ net514 VPWR u_ppwm_u_mem__0890_/Y VGND net434 hold196/A sg13g2_o21ai_1
XFILLER_6_344 VPWR VGND sg13g2_decap_8
XFILLER_10_373 VPWR VGND sg13g2_decap_8
XFILLER_10_384 VPWR VGND sg13g2_fill_1
XFILLER_11_896 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__132_ VPWR u_ppwm_u_pwm__132_/Y net533 VGND sg13g2_inv_1
XFILLER_7_878 VPWR VGND sg13g2_decap_8
XFILLER_2_583 VPWR VGND sg13g2_decap_8
XFILLER_28_6 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1092_ u_ppwm_u_ex__1091_/Y VPWR u_ppwm_u_ex__1092_/Y VGND u_ppwm_u_ex__1089_/Y
+ u_ppwm_u_ex__1090_/X sg13g2_o21ai_1
Xu_ppwm_u_global_counter__081_ u_ppwm_u_global_counter__083_/B u_ppwm_u_global_counter__081_/B
+ u_ppwm_u_global_counter__115_/D VPWR VGND sg13g2_and2_1
XFILLER_37_226 VPWR VGND sg13g2_fill_2
XFILLER_19_974 VPWR VGND sg13g2_decap_8
XFILLER_34_933 VPWR VGND sg13g2_decap_8
XFILLER_21_638 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0945_ u_ppwm_u_ex__0945_/Y net364 hold277/A net366 hold262/A VPWR VGND
+ sg13g2_a22oi_1
XFILLER_20_137 VPWR VGND sg13g2_fill_2
XFILLER_20_159 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0876_ VGND VPWR net450 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0877_/D u_ppwm_u_ex__0875_/Y
+ sg13g2_a21oi_1
XFILLER_0_509 VPWR VGND sg13g2_decap_8
XFILLER_29_749 VPWR VGND sg13g2_decap_8
XFILLER_44_708 VPWR VGND sg13g2_decap_8
XFILLER_25_911 VPWR VGND sg13g2_decap_8
XFILLER_19_1016 VPWR VGND sg13g2_decap_8
XFILLER_19_1027 VPWR VGND sg13g2_fill_2
XFILLER_24_432 VPWR VGND sg13g2_fill_1
XFILLER_40_936 VPWR VGND sg13g2_decap_8
XFILLER_24_465 VPWR VGND sg13g2_decap_8
XFILLER_25_988 VPWR VGND sg13g2_decap_8
XFILLER_22_33 VPWR VGND sg13g2_fill_1
XFILLER_4_848 VPWR VGND sg13g2_decap_8
XFILLER_26_1009 VPWR VGND sg13g2_decap_8
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_19_259 VPWR VGND sg13g2_decap_4
XFILLER_16_944 VPWR VGND sg13g2_decap_8
XFILLER_28_771 VPWR VGND sg13g2_decap_8
XFILLER_43_741 VPWR VGND sg13g2_decap_8
XFILLER_30_435 VPWR VGND sg13g2_fill_2
XFILLER_31_947 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0730_ u_ppwm_u_ex__0730_/A u_ppwm_u_ex__0732_/C u_ppwm_u_ex__0730_/C
+ u_ppwm_u_ex__0730_/D u_ppwm_u_ex__0730_/Y VPWR VGND sg13g2_nor4_1
XFILLER_30_457 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0942_ net510 VPWR u_ppwm_u_mem__0942_/Y VGND net427 hold228/A sg13g2_o21ai_1
XFILLER_11_693 VPWR VGND sg13g2_decap_8
XFILLER_10_192 VPWR VGND sg13g2_decap_8
XFILLER_10_181 VPWR VGND sg13g2_fill_2
XFILLER_7_675 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0661_ u_ppwm_u_ex__0660_/Y VPWR u_ppwm_u_ex__0663_/C VGND u_ppwm_u_ex__0652_/Y
+ u_ppwm_u_ex__0654_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__0873_ VGND VPWR net423 u_ppwm_u_mem__0718_/Y hold87/A u_ppwm_u_mem__0872_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0592_ net399 VPWR u_ppwm_u_ex__0592_/Y VGND net217 net614 sg13g2_o21ai_1
XFILLER_3_870 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1075_ u_ppwm_u_ex__1075_/A u_ppwm_u_ex__1075_/B u_ppwm_u_ex__1075_/C
+ u_ppwm_u_ex__1075_/Y VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_global_counter__064_ hold297/A net443 net445 u_ppwm_u_global_counter__067_/B
+ VPWR VGND net398 sg13g2_nand4_1
XFILLER_26_708 VPWR VGND sg13g2_decap_8
XFILLER_38_557 VPWR VGND sg13g2_decap_8
XFILLER_18_270 VPWR VGND sg13g2_fill_2
XFILLER_19_771 VPWR VGND sg13g2_decap_8
XFILLER_25_207 VPWR VGND sg13g2_decap_4
XFILLER_34_730 VPWR VGND sg13g2_decap_8
XFILLER_22_969 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0928_ net370 u_ppwm_u_ex__0928_/B u_ppwm_u_ex__0928_/X VPWR VGND sg13g2_and2_1
XFILLER_30_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0859_ u_ppwm_u_ex__1012_/A u_ppwm_u_ex__0859_/C net354 u_ppwm_u_ex__0859_/Y
+ VPWR VGND u_ppwm_u_ex__0859_/D sg13g2_nand4_1
XFILLER_0_306 VPWR VGND sg13g2_decap_8
XFILLER_29_546 VPWR VGND sg13g2_decap_8
XFILLER_44_505 VPWR VGND sg13g2_decap_8
XFILLER_17_11 VPWR VGND sg13g2_decap_8
XFILLER_17_719 VPWR VGND sg13g2_decap_8
XFILLER_25_785 VPWR VGND sg13g2_decap_8
XFILLER_40_733 VPWR VGND sg13g2_decap_8
XFILLER_13_969 VPWR VGND sg13g2_decap_8
XFILLER_9_929 VPWR VGND sg13g2_decap_8
XFILLER_4_645 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1121__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_0_873 VPWR VGND sg13g2_decap_8
Xhold6 hold6/A VPWR VGND net204 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1210_ net160 VGND VPWR u_ppwm_u_mem__1210_/D hold160/A clknet_5_9__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_48_866 VPWR VGND sg13g2_decap_8
XFILLER_47_354 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1141_ net80 VGND VPWR u_ppwm_u_mem__1141_/D hold116/A clknet_5_24__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_16_741 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1072_ net500 VPWR u_ppwm_u_mem__1072_/Y VGND net402 hold109/A sg13g2_o21ai_1
XFILLER_35_549 VPWR VGND sg13g2_decap_8
XFILLER_31_744 VPWR VGND sg13g2_decap_8
XFILLER_8_940 VPWR VGND sg13g2_decap_8
XFILLER_30_276 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0713_ u_ppwm_u_ex__0712_/Y VPWR u_ppwm_u_ex__0714_/C VGND u_ppwm_u_ex__0735_/A
+ hold277/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0925_ VGND VPWR net419 u_ppwm_u_mem__0692_/Y hold29/A u_ppwm_u_mem__0924_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0644_ net445 hold292/A u_ppwm_u_ex__0644_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__0856_ u_ppwm_u_mem__0855_/Y VPWR u_ppwm_u_mem__0856_/Y VGND net474
+ u_ppwm_u_mem__0853_/X sg13g2_o21ai_1
XFILLER_48_1020 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0787_ u_ppwm_u_mem__0786_/Y VPWR u_ppwm_u_mem__0787_/Y VGND u_ppwm_u_mem__0681_/Y
+ net482 sg13g2_o21ai_1
Xu_ppwm_u_ex__0575_ VPWR u_ppwm_u_ex__0732_/B net460 VGND sg13g2_inv_1
XFILLER_39_822 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__116_ net509 VGND VPWR net576 hold207/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_899 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1127_ net48 VGND VPWR net643 hold318/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1058_ u_ppwm_u_ex__1058_/Y hold236/A net356 VPWR VGND sg13g2_nand2_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_21_210 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1118__30 VPWR VGND net30 sg13g2_tiehi
XFILLER_10_906 VPWR VGND sg13g2_decap_8
XFILLER_22_766 VPWR VGND sg13g2_decap_8
XFILLER_21_265 VPWR VGND sg13g2_fill_2
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_48_129 VPWR VGND sg13g2_decap_8
XFILLER_45_814 VPWR VGND sg13g2_decap_8
XFILLER_17_516 VPWR VGND sg13g2_decap_8
XFILLER_29_398 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1144__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_40_530 VPWR VGND sg13g2_decap_8
XFILLER_25_582 VPWR VGND sg13g2_decap_8
XFILLER_9_726 VPWR VGND sg13g2_decap_8
XFILLER_13_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0710_ VPWR u_ppwm_u_mem__0710_/Y net564 VGND sg13g2_inv_1
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_4_442 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0641_ VPWR u_ppwm_u_mem__0641_/Y net571 VGND sg13g2_inv_1
XFILLER_0_670 VPWR VGND sg13g2_decap_8
XFILLER_48_663 VPWR VGND sg13g2_decap_8
XFILLER_47_151 VPWR VGND sg13g2_fill_2
XFILLER_35_302 VPWR VGND sg13g2_fill_1
XFILLER_36_858 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1124_ net114 VGND VPWR u_ppwm_u_mem__1124_/D hold175/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1055_ VGND VPWR net408 u_ppwm_u_mem__0627_/Y hold115/A u_ppwm_u_mem__1054_/Y
+ sg13g2_a21oi_1
XFILLER_31_541 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0908_ net515 VPWR u_ppwm_u_mem__0908_/Y VGND net436 hold213/A sg13g2_o21ai_1
Xhold225 hold225/A VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold203 hold203/A VPWR VGND net571 sg13g2_dlygate4sd3_1
Xhold214 hold214/A VPWR VGND net582 sg13g2_dlygate4sd3_1
Xhold236 hold236/A VPWR VGND net604 sg13g2_dlygate4sd3_1
Xhold269 hold269/A VPWR VGND net637 sg13g2_dlygate4sd3_1
Xhold258 hold258/A VPWR VGND net626 sg13g2_dlygate4sd3_1
Xhold247 hold247/A VPWR VGND net615 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0627_ u_ppwm_u_ex__0628_/B net469 net380 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__0839_ hold161/A hold138/A net485 u_ppwm_u_mem__0839_/X VPWR VGND sg13g2_mux2_1
XFILLER_39_696 VPWR VGND sg13g2_decap_8
XFILLER_27_858 VPWR VGND sg13g2_decap_8
XFILLER_42_817 VPWR VGND sg13g2_decap_8
XFILLER_10_703 VPWR VGND sg13g2_decap_8
XFILLER_22_563 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1121__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_5_239 VPWR VGND sg13g2_fill_1
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_2_968 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_45_611 VPWR VGND sg13g2_decap_8
XFILLER_17_313 VPWR VGND sg13g2_decap_8
XFILLER_18_869 VPWR VGND sg13g2_decap_8
XFILLER_29_173 VPWR VGND sg13g2_fill_2
XFILLER_45_688 VPWR VGND sg13g2_decap_8
XFILLER_33_806 VPWR VGND sg13g2_decap_8
XFILLER_41_894 VPWR VGND sg13g2_decap_8
XFILLER_9_523 VPWR VGND sg13g2_decap_8
XFILLER_13_563 VPWR VGND sg13g2_decap_8
XFILLER_40_382 VPWR VGND sg13g2_fill_2
XFILLER_5_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0624_ VPWR u_ppwm_u_mem__0624_/Y net253 VGND sg13g2_inv_1
XFILLER_48_460 VPWR VGND sg13g2_decap_8
XFILLER_36_655 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1107_ net174 VGND VPWR net598 hold229/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_880 VPWR VGND sg13g2_decap_8
XFILLER_23_327 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1038_ net501 VPWR u_ppwm_u_mem__1038_/Y VGND net407 net232 sg13g2_o21ai_1
XFILLER_32_850 VPWR VGND sg13g2_decap_8
XFILLER_31_371 VPWR VGND sg13g2_decap_8
Xfanout502 net503 net502 VPWR VGND sg13g2_buf_8
Xfanout513 net517 net513 VPWR VGND sg13g2_buf_8
XFILLER_46_419 VPWR VGND sg13g2_decap_8
XFILLER_39_493 VPWR VGND sg13g2_decap_8
XFILLER_15_817 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_27_655 VPWR VGND sg13g2_decap_8
XFILLER_42_614 VPWR VGND sg13g2_decap_8
XFILLER_25_22 VPWR VGND sg13g2_decap_8
XFILLER_41_124 VPWR VGND sg13g2_fill_1
XFILLER_10_577 VPWR VGND sg13g2_decap_8
XFILLER_6_548 VPWR VGND sg13g2_decap_8
XFILLER_2_765 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_fill_1
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_46_986 VPWR VGND sg13g2_decap_8
XFILLER_17_132 VPWR VGND sg13g2_decap_4
XFILLER_18_666 VPWR VGND sg13g2_decap_8
XFILLER_33_603 VPWR VGND sg13g2_decap_8
XFILLER_45_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0961_ u_ppwm_u_ex__0962_/B net364 hold252/A net366 net442 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_20_308 VPWR VGND sg13g2_fill_2
XFILLER_41_691 VPWR VGND sg13g2_decap_8
XFILLER_9_331 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0892_ VGND VPWR u_ppwm_u_ex__0711_/A net384 u_ppwm_u_ex__0892_/Y u_ppwm_u_ex__0891_/Y
+ sg13g2_a21oi_1
XFILLER_12_1000 VPWR VGND sg13g2_decap_8
XFILLER_5_570 VPWR VGND sg13g2_decap_8
XFILLER_37_920 VPWR VGND sg13g2_decap_8
XFILLER_37_997 VPWR VGND sg13g2_decap_8
XFILLER_23_135 VPWR VGND sg13g2_decap_8
XFILLER_23_146 VPWR VGND sg13g2_fill_1
XFILLER_24_647 VPWR VGND sg13g2_decap_8
XFILLER_20_886 VPWR VGND sg13g2_decap_8
XFILLER_11_79 VPWR VGND sg13g2_fill_1
Xfanout365 fanout365/A net365 VPWR VGND sg13g2_buf_8
Xfanout354 fanout354/A net354 VPWR VGND sg13g2_buf_8
XFILLER_47_739 VPWR VGND sg13g2_decap_8
XFILLER_4_1009 VPWR VGND sg13g2_decap_8
Xfanout398 net399 net398 VPWR VGND sg13g2_buf_8
Xfanout376 fanout376/A net376 VPWR VGND sg13g2_buf_1
Xfanout387 fanout387/A net387 VPWR VGND sg13g2_buf_8
XFILLER_46_216 VPWR VGND sg13g2_decap_8
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_43_923 VPWR VGND sg13g2_decap_8
XFILLER_42_411 VPWR VGND sg13g2_decap_8
XFILLER_15_614 VPWR VGND sg13g2_decap_8
XFILLER_42_488 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__200_ VGND VPWR u_ppwm_u_pwm__198_/Y u_ppwm_u_pwm__199_/Y u_ppwm_u_pwm__200_/Y
+ u_ppwm_u_pwm__197_/Y sg13g2_a21oi_1
XFILLER_11_875 VPWR VGND sg13g2_decap_8
XFILLER_7_857 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__131_ u_ppwm_u_pwm__213_/B net207 VPWR VGND sg13g2_inv_2
XFILLER_42_9 VPWR VGND sg13g2_fill_1
XFILLER_2_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1091_ VGND VPWR u_ppwm_u_ex__1089_/Y u_ppwm_u_ex__1090_/X u_ppwm_u_ex__1091_/Y
+ net357 sg13g2_a21oi_1
Xu_ppwm_u_global_counter__080_ u_ppwm_u_global_counter__082_/D net201 net441 u_ppwm_u_global_counter__081_/B
+ VPWR VGND sg13g2_a21o_1
XFILLER_38_739 VPWR VGND sg13g2_decap_8
XFILLER_19_953 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1131__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_46_783 VPWR VGND sg13g2_decap_8
XFILLER_45_260 VPWR VGND sg13g2_fill_2
XFILLER_34_912 VPWR VGND sg13g2_decap_8
XFILLER_45_282 VPWR VGND sg13g2_decap_8
XFILLER_21_617 VPWR VGND sg13g2_decap_8
XFILLER_34_989 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0944_ hold294/A VPWR u_ppwm_u_ex__0944_/Y VGND net381 net370 sg13g2_o21ai_1
Xu_ppwm_u_ex__0875_ net360 u_ppwm_u_ex__0875_/B u_ppwm_u_ex__0875_/Y VPWR VGND sg13g2_nor2_1
XFILLER_9_194 VPWR VGND sg13g2_decap_8
XFILLER_29_728 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1183__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_37_794 VPWR VGND sg13g2_decap_8
XFILLER_25_967 VPWR VGND sg13g2_decap_8
XFILLER_40_915 VPWR VGND sg13g2_decap_8
XFILLER_11_127 VPWR VGND sg13g2_decap_8
XFILLER_20_683 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1108__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_4_827 VPWR VGND sg13g2_decap_8
XFILLER_47_536 VPWR VGND sg13g2_decap_8
XFILLER_47_53 VPWR VGND sg13g2_decap_8
XFILLER_19_227 VPWR VGND sg13g2_decap_8
XFILLER_19_238 VPWR VGND sg13g2_fill_2
XFILLER_28_750 VPWR VGND sg13g2_decap_8
XFILLER_43_720 VPWR VGND sg13g2_decap_8
XFILLER_16_923 VPWR VGND sg13g2_decap_8
XFILLER_31_926 VPWR VGND sg13g2_decap_8
XFILLER_43_797 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0941_ VGND VPWR net417 u_ppwm_u_mem__0684_/Y u_ppwm_u_mem__1147_/D
+ u_ppwm_u_mem__0940_/Y sg13g2_a21oi_1
XFILLER_11_672 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0660_ u_ppwm_u_ex__0660_/A u_ppwm_u_ex__0660_/B u_ppwm_u_ex__0660_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_7_654 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0872_ net513 VPWR u_ppwm_u_mem__0872_/Y VGND net423 hold192/A sg13g2_o21ai_1
Xu_ppwm_u_mem__1161__159 VPWR VGND net159 sg13g2_tiehi
Xu_ppwm_u_ex__0591_ VPWR u_ppwm_u_ex__0591_/Y net443 VGND sg13g2_inv_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_536 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1074_ VGND VPWR u_ppwm_u_ex__1067_/Y u_ppwm_u_ex__1072_/Y u_ppwm_u_ex__1122_/D
+ u_ppwm_u_ex__1073_/Y sg13g2_a21oi_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_global_counter__063_ u_ppwm_u_global_counter__070_/A u_ppwm_u_global_counter__063_/B
+ u_ppwm_u_global_counter__107_/D VPWR VGND sg13g2_and2_1
XFILLER_19_750 VPWR VGND sg13g2_decap_8
XFILLER_46_580 VPWR VGND sg13g2_decap_8
XFILLER_34_786 VPWR VGND sg13g2_decap_8
XFILLER_22_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0927_ VGND VPWR u_ppwm_u_ex__0925_/Y u_ppwm_u_ex__0926_/Y u_ppwm_u_ex__0927_/Y
+ u_ppwm_u_ex__0819_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0858_ VGND VPWR net451 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0859_/D u_ppwm_u_ex__0857_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__0789_ net381 net375 u_ppwm_u_ex__0789_/Y VPWR VGND sg13g2_nor2_1
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_29_525 VPWR VGND sg13g2_decap_8
XFILLER_37_591 VPWR VGND sg13g2_decap_8
XFILLER_40_712 VPWR VGND sg13g2_decap_8
XFILLER_24_252 VPWR VGND sg13g2_decap_4
XFILLER_25_764 VPWR VGND sg13g2_decap_8
XFILLER_9_908 VPWR VGND sg13g2_decap_8
XFILLER_13_948 VPWR VGND sg13g2_decap_8
XFILLER_40_789 VPWR VGND sg13g2_decap_8
XFILLER_21_981 VPWR VGND sg13g2_decap_8
XFILLER_32_1025 VPWR VGND sg13g2_decap_4
XFILLER_20_480 VPWR VGND sg13g2_decap_8
XFILLER_4_624 VPWR VGND sg13g2_decap_8
XFILLER_3_101 VPWR VGND sg13g2_fill_2
XFILLER_3_156 VPWR VGND sg13g2_fill_2
XFILLER_0_852 VPWR VGND sg13g2_decap_8
XFILLER_48_845 VPWR VGND sg13g2_decap_8
Xhold7 hold7/A VPWR VGND net205 sg13g2_dlygate4sd3_1
XFILLER_47_333 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1140_ net82 VGND VPWR u_ppwm_u_mem__1140_/D hold28/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1071_ VGND VPWR net402 u_ppwm_u_mem__0619_/Y hold110/A u_ppwm_u_mem__1070_/Y
+ sg13g2_a21oi_1
XFILLER_35_528 VPWR VGND sg13g2_decap_8
XFILLER_16_720 VPWR VGND sg13g2_decap_8
XFILLER_43_594 VPWR VGND sg13g2_decap_8
XFILLER_16_797 VPWR VGND sg13g2_decap_8
XFILLER_30_222 VPWR VGND sg13g2_decap_8
XFILLER_31_723 VPWR VGND sg13g2_decap_8
XFILLER_30_244 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0712_ u_ppwm_u_ex__0712_/Y hold289/A hold217/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0924_ net502 VPWR u_ppwm_u_mem__0924_/Y VGND net419 hold191/A sg13g2_o21ai_1
XFILLER_8_996 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0643_ u_ppwm_u_ex__0643_/Y net444 net453 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0855_ VGND VPWR net474 u_ppwm_u_mem__0854_/X u_ppwm_u_mem__0855_/Y
+ net394 sg13g2_a21oi_1
Xu_ppwm_u_mem__0786_ u_ppwm_u_mem__0786_/Y hold47/A net482 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__0574_ VPWR u_ppwm_u_ex__0758_/A net458 VGND sg13g2_inv_1
XFILLER_39_801 VPWR VGND sg13g2_decap_8
XFILLER_39_878 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__115_ net509 VGND VPWR u_ppwm_u_global_counter__115_/D hold271/A
+ clknet_5_21__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1126_ net32 VGND VPWR net219 hold19/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1057_ u_ppwm_u_ex__1056_/Y VPWR u_ppwm_u_ex__1061_/C VGND u_ppwm_u_ex__1051_/A
+ u_ppwm_u_ex__1055_/X sg13g2_o21ai_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_41_509 VPWR VGND sg13g2_decap_8
XFILLER_22_745 VPWR VGND sg13g2_decap_8
XFILLER_34_583 VPWR VGND sg13g2_decap_8
XFILLER_21_233 VPWR VGND sg13g2_decap_8
XFILLER_21_244 VPWR VGND sg13g2_fill_1
XFILLER_9_90 VPWR VGND sg13g2_fill_2
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_fill_2
XFILLER_44_325 VPWR VGND sg13g2_decap_4
XFILLER_25_561 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_4
XFILLER_9_705 VPWR VGND sg13g2_decap_8
XFILLER_13_745 VPWR VGND sg13g2_decap_8
XFILLER_40_586 VPWR VGND sg13g2_decap_8
XFILLER_8_204 VPWR VGND sg13g2_fill_2
XFILLER_12_266 VPWR VGND sg13g2_fill_1
XFILLER_12_277 VPWR VGND sg13g2_decap_4
XFILLER_8_259 VPWR VGND sg13g2_decap_8
XFILLER_5_955 VPWR VGND sg13g2_decap_8
XFILLER_4_421 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0640_ VPWR u_ppwm_u_mem__0640_/Y net538 VGND sg13g2_inv_1
XFILLER_4_498 VPWR VGND sg13g2_decap_8
XFILLER_48_642 VPWR VGND sg13g2_decap_8
XFILLER_36_837 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1123_ net116 VGND VPWR net544 hold183/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1054_ net501 VPWR u_ppwm_u_mem__1054_/Y VGND net408 hold130/A sg13g2_o21ai_1
XFILLER_16_594 VPWR VGND sg13g2_decap_8
XFILLER_15_1020 VPWR VGND sg13g2_decap_8
XFILLER_31_597 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0907_ VGND VPWR net434 u_ppwm_u_mem__0701_/Y u_ppwm_u_mem__1130_/D
+ u_ppwm_u_mem__0906_/Y sg13g2_a21oi_1
XFILLER_8_793 VPWR VGND sg13g2_decap_8
Xhold226 hold226/A VPWR VGND net594 sg13g2_dlygate4sd3_1
Xhold204 hold204/A VPWR VGND net572 sg13g2_dlygate4sd3_1
Xhold215 hold215/A VPWR VGND net583 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0838_ hold71/A hold73/A net481 u_ppwm_u_mem__0838_/X VPWR VGND sg13g2_mux2_1
Xhold237 hold237/A VPWR VGND net605 sg13g2_dlygate4sd3_1
Xhold259 hold259/A VPWR VGND net627 sg13g2_dlygate4sd3_1
Xhold248 hold248/A VPWR VGND net616 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0626_ u_ppwm_u_ex__0626_/Y net469 net380 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0769_ u_ppwm_u_mem__0769_/Y hold84/A net484 VPWR VGND sg13g2_nand2_1
XFILLER_26_303 VPWR VGND sg13g2_fill_2
XFILLER_27_837 VPWR VGND sg13g2_decap_8
XFILLER_39_675 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1109_ net33 VGND VPWR u_ppwm_u_ex__1109_/D hold308/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_892 VPWR VGND sg13g2_decap_8
XFILLER_22_542 VPWR VGND sg13g2_decap_8
XFILLER_10_759 VPWR VGND sg13g2_decap_8
XFILLER_5_229 VPWR VGND sg13g2_fill_1
XFILLER_2_947 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_29_163 VPWR VGND sg13g2_fill_1
XFILLER_18_848 VPWR VGND sg13g2_decap_8
XFILLER_45_667 VPWR VGND sg13g2_decap_8
XFILLER_32_306 VPWR VGND sg13g2_fill_1
XFILLER_13_542 VPWR VGND sg13g2_decap_8
XFILLER_41_873 VPWR VGND sg13g2_decap_8
XFILLER_9_502 VPWR VGND sg13g2_decap_8
XFILLER_9_579 VPWR VGND sg13g2_decap_8
XFILLER_5_752 VPWR VGND sg13g2_decap_8
XFILLER_4_251 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0623_ VPWR u_ppwm_u_mem__0623_/Y net318 VGND sg13g2_inv_1
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
XFILLER_49_984 VPWR VGND sg13g2_decap_8
XFILLER_36_634 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1106_ net566 u_ppwm_u_mem__1105_/Y hold199/A VPWR VGND sg13g2_nor2b_1
XFILLER_24_829 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1037_ VGND VPWR net407 u_ppwm_u_mem__0636_/Y hold35/A u_ppwm_u_mem__1036_/Y
+ sg13g2_a21oi_1
XFILLER_8_590 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0609_ u_ppwm_u_ex__0623_/B net388 u_ppwm/instr\[0\] u_ppwm_u_ex__0610_/C
+ VPWR VGND sg13g2_and3_1
Xfanout514 net517 net514 VPWR VGND sg13g2_buf_1
Xfanout503 net504 net503 VPWR VGND sg13g2_buf_8
XFILLER_27_634 VPWR VGND sg13g2_decap_8
XFILLER_39_472 VPWR VGND sg13g2_decap_8
XFILLER_26_144 VPWR VGND sg13g2_fill_1
XFILLER_14_306 VPWR VGND sg13g2_decap_8
XFILLER_14_339 VPWR VGND sg13g2_decap_4
XFILLER_22_372 VPWR VGND sg13g2_decap_4
XFILLER_23_895 VPWR VGND sg13g2_decap_8
XFILLER_41_66 VPWR VGND sg13g2_fill_2
XFILLER_6_527 VPWR VGND sg13g2_decap_8
XFILLER_10_556 VPWR VGND sg13g2_decap_8
XFILLER_41_88 VPWR VGND sg13g2_fill_1
XFILLER_29_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_744 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1118__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_18_645 VPWR VGND sg13g2_decap_8
XFILLER_46_965 VPWR VGND sg13g2_decap_8
XFILLER_45_464 VPWR VGND sg13g2_decap_8
XFILLER_17_122 VPWR VGND sg13g2_fill_1
XFILLER_17_155 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0960_ u_ppwm_u_ex__1086_/A u_ppwm_u_ex__0959_/Y u_ppwm_u_ex__0820_/C
+ u_ppwm_u_ex__0928_/X u_ppwm_u_ex__0790_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_32_147 VPWR VGND sg13g2_fill_2
XFILLER_33_659 VPWR VGND sg13g2_decap_8
XFILLER_41_670 VPWR VGND sg13g2_decap_8
XFILLER_13_350 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0891_ net455 net384 u_ppwm_u_ex__0891_/Y VPWR VGND sg13g2_nor2_1
XFILLER_14_895 VPWR VGND sg13g2_decap_8
XFILLER_28_409 VPWR VGND sg13g2_fill_2
XFILLER_49_781 VPWR VGND sg13g2_decap_8
XFILLER_37_976 VPWR VGND sg13g2_decap_8
XFILLER_24_626 VPWR VGND sg13g2_decap_8
XFILLER_36_486 VPWR VGND sg13g2_fill_1
XFILLER_20_865 VPWR VGND sg13g2_decap_8
Xfanout355 fanout355/A net355 VPWR VGND sg13g2_buf_8
Xfanout366 fanout367/A net366 VPWR VGND sg13g2_buf_8
XFILLER_47_718 VPWR VGND sg13g2_decap_8
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
Xfanout377 net378 net377 VPWR VGND sg13g2_buf_8
Xfanout399 net642 net399 VPWR VGND sg13g2_buf_8
Xfanout388 fanout388/A net388 VPWR VGND sg13g2_buf_8
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_43_902 VPWR VGND sg13g2_decap_8
XFILLER_43_979 VPWR VGND sg13g2_decap_8
XFILLER_42_467 VPWR VGND sg13g2_decap_8
XFILLER_23_692 VPWR VGND sg13g2_decap_8
XFILLER_10_342 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__130_ VPWR u_ppwm_u_pwm__214_/B net260 VGND sg13g2_inv_1
XFILLER_11_854 VPWR VGND sg13g2_decap_8
XFILLER_7_836 VPWR VGND sg13g2_decap_8
XFILLER_2_541 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_718 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1090_ net374 net657 u_ppwm_u_ex__1090_/X VPWR VGND sg13g2_xor2_1
XFILLER_19_932 VPWR VGND sg13g2_decap_8
XFILLER_46_762 VPWR VGND sg13g2_decap_8
XFILLER_34_968 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0943_ u_ppwm_u_ex__1071_/A u_ppwm_u_ex__0942_/Y u_ppwm_u_ex__0820_/C
+ u_ppwm_u_ex__0910_/X u_ppwm_u_ex__0790_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_14_692 VPWR VGND sg13g2_decap_8
XFILLER_33_489 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0874_ u_ppwm_u_ex__0875_/B net365 u_ppwm_u_ex__1020_/B2 net367 hold231/A
+ VPWR VGND sg13g2_a22oi_1
XFILLER_9_184 VPWR VGND sg13g2_decap_4
XFILLER_6_891 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_fill_2
XFILLER_29_707 VPWR VGND sg13g2_decap_8
XFILLER_3_1010 VPWR VGND sg13g2_decap_8
XFILLER_37_773 VPWR VGND sg13g2_decap_8
XFILLER_24_423 VPWR VGND sg13g2_decap_8
XFILLER_25_946 VPWR VGND sg13g2_decap_8
XFILLER_12_629 VPWR VGND sg13g2_decap_8
XFILLER_20_662 VPWR VGND sg13g2_decap_8
XFILLER_4_806 VPWR VGND sg13g2_decap_8
XFILLER_3_349 VPWR VGND sg13g2_fill_2
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_515 VPWR VGND sg13g2_decap_8
XFILLER_16_902 VPWR VGND sg13g2_decap_8
XFILLER_43_776 VPWR VGND sg13g2_decap_8
XFILLER_16_979 VPWR VGND sg13g2_decap_8
XFILLER_30_404 VPWR VGND sg13g2_decap_4
XFILLER_31_905 VPWR VGND sg13g2_decap_8
XFILLER_24_990 VPWR VGND sg13g2_decap_8
XFILLER_11_651 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0940_ net502 VPWR u_ppwm_u_mem__0940_/Y VGND net417 net273 sg13g2_o21ai_1
XFILLER_7_633 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0871_ VGND VPWR net432 u_ppwm_u_mem__0719_/Y u_ppwm_u_mem__1112_/D
+ u_ppwm_u_mem__0870_/Y sg13g2_a21oi_1
XFILLER_10_183 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0590_ VPWR u_ppwm_u_ex__1019_/B hold231/A VGND sg13g2_inv_1
XFILLER_38_515 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1073_ net505 VPWR u_ppwm_u_ex__1073_/Y VGND net662 net349 sg13g2_o21ai_1
Xu_ppwm_u_global_counter__062_ net399 net445 net444 u_ppwm_u_global_counter__063_/B
+ VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_pwm__241__182 VPWR VGND net182 sg13g2_tiehi
XFILLER_22_927 VPWR VGND sg13g2_decap_8
XFILLER_34_765 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0926_ u_ppwm_u_ex__0926_/Y u_ppwm_u_ex__0838_/Y u_ppwm_u_ex__0801_/X
+ u_ppwm_u_ex__0838_/B u_ppwm_u_ex__0866_/C VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_ex__0857_ u_ppwm_u_ex__1012_/B VPWR u_ppwm_u_ex__0857_/Y VGND net359 u_ppwm_u_ex__0855_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__0788_ u_ppwm_u_ex__0843_/A u_ppwm/instr\[0\] u_ppwm_u_ex__0819_/C VPWR
+ VGND sg13g2_nand2_2
Xu_ppwm_u_mem__1218__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_37_570 VPWR VGND sg13g2_decap_8
XFILLER_25_743 VPWR VGND sg13g2_decap_8
XFILLER_13_927 VPWR VGND sg13g2_decap_8
XFILLER_40_768 VPWR VGND sg13g2_decap_8
XFILLER_32_1004 VPWR VGND sg13g2_decap_8
XFILLER_21_960 VPWR VGND sg13g2_decap_8
XFILLER_4_603 VPWR VGND sg13g2_decap_8
XFILLER_3_113 VPWR VGND sg13g2_fill_2
XFILLER_0_831 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_48_824 VPWR VGND sg13g2_decap_8
XFILLER_47_312 VPWR VGND sg13g2_decap_8
Xhold8 hold8/A VPWR VGND net206 sg13g2_dlygate4sd3_1
XFILLER_47_389 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1070_ net493 VPWR u_ppwm_u_mem__1070_/Y VGND net406 hold145/A sg13g2_o21ai_1
XFILLER_15_253 VPWR VGND sg13g2_decap_4
XFILLER_16_776 VPWR VGND sg13g2_decap_8
XFILLER_31_702 VPWR VGND sg13g2_decap_8
XFILLER_43_573 VPWR VGND sg13g2_decap_8
XFILLER_31_779 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0923_ VGND VPWR net427 u_ppwm_u_mem__0693_/Y u_ppwm_u_mem__1138_/D
+ u_ppwm_u_mem__0922_/Y sg13g2_a21oi_1
XFILLER_8_975 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0711_ u_ppwm_u_ex__0711_/A hold252/A u_ppwm_u_ex__0714_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_12_993 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0642_ u_ppwm_u_ex__0642_/Y hold222/A u_ppwm_u_ex__1025_/A hold259/A
+ u_ppwm_u_ex__0651_/A VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__0854_ hold42/A hold119/A net480 u_ppwm_u_mem__0854_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0573_ u_ppwm_u_ex__0757_/A hold296/A VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0785_ u_ppwm_u_mem__0784_/Y VPWR u_ppwm_u_mem__0785_/Y VGND u_ppwm_u_mem__0695_/Y
+ net486 sg13g2_o21ai_1
Xu_ppwm_u_global_counter__114_ net507 VGND VPWR net202 hold3/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1125_ net54 VGND VPWR net616 hold246/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_345 VPWR VGND sg13g2_fill_2
XFILLER_39_857 VPWR VGND sg13g2_decap_8
XFILLER_38_356 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1056_ VGND VPWR u_ppwm_u_ex__1051_/A u_ppwm_u_ex__1055_/X u_ppwm_u_ex__1056_/Y
+ net357 sg13g2_a21oi_1
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
XFILLER_34_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1199_ net129 VGND VPWR u_ppwm_u_mem__1199_/D hold158/A clknet_5_12__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_22_724 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0909_ VGND VPWR u_ppwm_u_ex__0973_/A net384 u_ppwm_u_ex__0928_/B u_ppwm_u_ex__0908_/Y
+ sg13g2_a21oi_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_25_540 VPWR VGND sg13g2_decap_8
XFILLER_13_724 VPWR VGND sg13g2_decap_8
XFILLER_40_565 VPWR VGND sg13g2_decap_8
XFILLER_5_934 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_477 VPWR VGND sg13g2_decap_8
XFILLER_48_621 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1122_ net118 VGND VPWR net552 hold196/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_816 VPWR VGND sg13g2_decap_8
XFILLER_48_698 VPWR VGND sg13g2_decap_8
XFILLER_47_186 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1053_ VGND VPWR net407 u_ppwm_u_mem__0628_/Y u_ppwm_u_mem__1203_/D
+ u_ppwm_u_mem__1052_/Y sg13g2_a21oi_1
XFILLER_16_573 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1128__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_31_576 VPWR VGND sg13g2_decap_8
XFILLER_12_790 VPWR VGND sg13g2_decap_8
XFILLER_8_772 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0906_ net513 VPWR u_ppwm_u_mem__0906_/Y VGND net434 net524 sg13g2_o21ai_1
XFILLER_7_271 VPWR VGND sg13g2_decap_4
Xhold205 hold205/A VPWR VGND net573 sg13g2_dlygate4sd3_1
Xhold216 hold216/A VPWR VGND net584 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0837_ hold28/A hold75/A net480 u_ppwm_u_mem__0837_/X VPWR VGND sg13g2_mux2_1
Xhold227 hold227/A VPWR VGND net595 sg13g2_dlygate4sd3_1
Xhold238 hold238/A VPWR VGND net606 sg13g2_dlygate4sd3_1
Xhold249 hold256/A VPWR VGND net617 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0625_ VGND VPWR net473 net383 u_ppwm_u_ex__0628_/A u_ppwm_u_ex__0619_/C
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0768_ u_ppwm_u_mem__0767_/Y VPWR u_ppwm_u_mem__0768_/Y VGND u_ppwm_u_mem__0682_/Y
+ net482 sg13g2_o21ai_1
Xu_ppwm_u_mem__0699_ VPWR u_ppwm_u_mem__0699_/Y net336 VGND sg13g2_inv_1
XFILLER_22_1025 VPWR VGND sg13g2_decap_4
XFILLER_39_654 VPWR VGND sg13g2_decap_8
XFILLER_27_816 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1108_ net35 VGND VPWR u_ppwm_u_ex__1108_/D hold324/A clknet_5_25__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_326 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__1039_ net373 hold299/A u_ppwm_u_ex__1054_/B VPWR VGND sg13g2_xor2_1
XFILLER_26_359 VPWR VGND sg13g2_decap_4
XFILLER_35_871 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_22_521 VPWR VGND sg13g2_decap_8
XFILLER_6_709 VPWR VGND sg13g2_decap_8
XFILLER_10_738 VPWR VGND sg13g2_decap_8
XFILLER_22_598 VPWR VGND sg13g2_decap_8
XFILLER_30_46 VPWR VGND sg13g2_fill_1
XFILLER_2_926 VPWR VGND sg13g2_decap_8
XFILLER_39_11 VPWR VGND sg13g2_fill_1
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_99 VPWR VGND sg13g2_decap_4
XFILLER_18_827 VPWR VGND sg13g2_decap_8
XFILLER_29_153 VPWR VGND sg13g2_fill_1
XFILLER_45_646 VPWR VGND sg13g2_decap_8
XFILLER_44_101 VPWR VGND sg13g2_fill_1
XFILLER_41_852 VPWR VGND sg13g2_decap_8
XFILLER_13_521 VPWR VGND sg13g2_decap_8
XFILLER_9_558 VPWR VGND sg13g2_decap_8
XFILLER_13_598 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1112__27 VPWR VGND net27 sg13g2_tiehi
XFILLER_5_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0622_ VPWR u_ppwm_u_mem__0622_/Y net528 VGND sg13g2_inv_1
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_963 VPWR VGND sg13g2_decap_8
XFILLER_48_495 VPWR VGND sg13g2_decap_8
XFILLER_36_613 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1105_ VGND VPWR net565 u_ppwm_u_mem__1103_/C u_ppwm_u_mem__1105_/Y
+ u_ppwm_u_mem__1094_/A sg13g2_a21oi_1
XFILLER_24_808 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1036_ net501 VPWR u_ppwm_u_mem__1036_/Y VGND net407 hold107/A sg13g2_o21ai_1
XFILLER_32_885 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0608_ u_ppwm_u_ex__0610_/C u_ppwm/instr\[1\] hold280/A VPWR VGND sg13g2_nand2b_1
Xfanout504 rst_n net504 VPWR VGND sg13g2_buf_8
Xfanout515 net517 net515 VPWR VGND sg13g2_buf_8
XFILLER_27_613 VPWR VGND sg13g2_decap_8
XFILLER_26_167 VPWR VGND sg13g2_decap_4
XFILLER_26_189 VPWR VGND sg13g2_decap_8
XFILLER_42_649 VPWR VGND sg13g2_decap_8
XFILLER_25_79 VPWR VGND sg13g2_fill_2
XFILLER_23_874 VPWR VGND sg13g2_decap_8
XFILLER_10_535 VPWR VGND sg13g2_decap_8
XFILLER_6_506 VPWR VGND sg13g2_decap_8
XFILLER_2_723 VPWR VGND sg13g2_decap_8
XFILLER_1_288 VPWR VGND sg13g2_decap_4
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_46_944 VPWR VGND sg13g2_decap_8
XFILLER_18_624 VPWR VGND sg13g2_decap_8
XFILLER_45_443 VPWR VGND sg13g2_decap_8
XFILLER_33_638 VPWR VGND sg13g2_decap_8
XFILLER_9_300 VPWR VGND sg13g2_decap_4
XFILLER_14_874 VPWR VGND sg13g2_decap_8
XFILLER_13_362 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0890_ u_ppwm_u_ex__0890_/A u_ppwm_u_ex__0890_/B u_ppwm_u_ex__0890_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_49_760 VPWR VGND sg13g2_decap_8
XFILLER_48_292 VPWR VGND sg13g2_decap_8
XFILLER_37_955 VPWR VGND sg13g2_decap_8
XFILLER_24_605 VPWR VGND sg13g2_decap_8
XFILLER_36_476 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1019_ VGND VPWR net414 u_ppwm_u_mem__0645_/Y hold39/A u_ppwm_u_mem__1018_/Y
+ sg13g2_a21oi_1
XFILLER_32_682 VPWR VGND sg13g2_decap_8
XFILLER_20_844 VPWR VGND sg13g2_decap_8
XFILLER_11_59 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1186__71 VPWR VGND net71 sg13g2_tiehi
Xfanout356 fanout356/A net356 VPWR VGND sg13g2_buf_8
Xfanout389 net391 net389 VPWR VGND sg13g2_buf_8
Xfanout367 fanout367/A net367 VPWR VGND sg13g2_buf_2
Xfanout378 net379 net378 VPWR VGND sg13g2_buf_8
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_fill_1
XFILLER_43_958 VPWR VGND sg13g2_decap_8
XFILLER_42_446 VPWR VGND sg13g2_decap_8
XFILLER_15_649 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_decap_8
XFILLER_23_671 VPWR VGND sg13g2_decap_8
XFILLER_10_321 VPWR VGND sg13g2_fill_1
XFILLER_7_815 VPWR VGND sg13g2_decap_8
XFILLER_6_314 VPWR VGND sg13g2_fill_2
XFILLER_2_520 VPWR VGND sg13g2_decap_8
XFILLER_42_1006 VPWR VGND sg13g2_decap_8
XFILLER_2_597 VPWR VGND sg13g2_decap_8
XFILLER_18_410 VPWR VGND sg13g2_decap_8
XFILLER_19_911 VPWR VGND sg13g2_decap_8
XFILLER_46_741 VPWR VGND sg13g2_decap_8
XFILLER_19_988 VPWR VGND sg13g2_decap_8
XFILLER_33_402 VPWR VGND sg13g2_decap_8
XFILLER_18_498 VPWR VGND sg13g2_decap_8
XFILLER_34_947 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0942_ u_ppwm_u_ex__0941_/Y VPWR u_ppwm_u_ex__0942_/Y VGND u_ppwm_u_ex__0814_/Y
+ u_ppwm_u_ex__0839_/Y sg13g2_o21ai_1
XFILLER_14_671 VPWR VGND sg13g2_decap_8
XFILLER_9_152 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0873_ u_ppwm_u_ex__0872_/Y u_ppwm_u_ex__0868_/Y u_ppwm_u_ex__0843_/A
+ u_ppwm_u_ex__0877_/C VPWR VGND sg13g2_a21o_1
XFILLER_6_870 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__189_ hold279/A net489 net549 u_ppwm_u_pwm__191_/B VPWR VGND sg13g2_nand3_1
XFILLER_37_752 VPWR VGND sg13g2_decap_8
XFILLER_25_925 VPWR VGND sg13g2_decap_8
XFILLER_12_608 VPWR VGND sg13g2_decap_8
XFILLER_24_479 VPWR VGND sg13g2_decap_8
XFILLER_20_641 VPWR VGND sg13g2_decap_8
XFILLER_3_317 VPWR VGND sg13g2_fill_2
XFILLER_3_306 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1193__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_42_210 VPWR VGND sg13g2_decap_4
XFILLER_16_958 VPWR VGND sg13g2_decap_8
XFILLER_43_755 VPWR VGND sg13g2_decap_8
XFILLER_42_232 VPWR VGND sg13g2_decap_4
XFILLER_11_630 VPWR VGND sg13g2_decap_8
XFILLER_7_612 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0870_ net515 VPWR u_ppwm_u_mem__0870_/Y VGND net432 net277 sg13g2_o21ai_1
XFILLER_6_122 VPWR VGND sg13g2_decap_4
XFILLER_7_689 VPWR VGND sg13g2_decap_8
XFILLER_3_884 VPWR VGND sg13g2_decap_8
XFILLER_2_394 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1072_ u_ppwm_u_ex__1072_/A u_ppwm_u_ex__1072_/B u_ppwm_u_ex__1072_/Y
+ VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_global_counter__061_ net444 net398 net445 u_ppwm_u_global_counter__070_/A
+ VPWR VGND sg13g2_nand3_1
XFILLER_19_785 VPWR VGND sg13g2_decap_8
XFILLER_33_221 VPWR VGND sg13g2_fill_1
XFILLER_34_744 VPWR VGND sg13g2_decap_8
XFILLER_22_906 VPWR VGND sg13g2_decap_8
XFILLER_21_416 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0925_ u_ppwm_u_ex__0925_/Y net368 u_ppwm_u_ex__0925_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__0856_ u_ppwm_u_ex__1012_/B net375 u_ppwm_u_ex__0856_/B VPWR VGND sg13g2_nand2_1
XFILLER_30_994 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0787_ VGND VPWR net660 u_ppwm_u_ex__0831_/B u_ppwm_u_ex__0787_/Y u_ppwm_u_ex__0786_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0999_ VGND VPWR net411 u_ppwm_u_mem__0655_/Y hold151/A u_ppwm_u_mem__0998_/Y
+ sg13g2_a21oi_1
XFILLER_25_1023 VPWR VGND sg13g2_decap_4
XFILLER_44_519 VPWR VGND sg13g2_decap_8
XFILLER_17_25 VPWR VGND sg13g2_fill_2
XFILLER_25_722 VPWR VGND sg13g2_decap_8
XFILLER_13_906 VPWR VGND sg13g2_decap_8
XFILLER_24_232 VPWR VGND sg13g2_fill_2
XFILLER_25_799 VPWR VGND sg13g2_decap_8
XFILLER_40_747 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1160__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_4_659 VPWR VGND sg13g2_decap_8
XFILLER_3_103 VPWR VGND sg13g2_fill_1
XFILLER_0_810 VPWR VGND sg13g2_decap_8
XFILLER_48_803 VPWR VGND sg13g2_decap_8
Xhold9 hold9/A VPWR VGND net207 sg13g2_dlygate4sd3_1
XFILLER_0_887 VPWR VGND sg13g2_decap_8
XFILLER_47_368 VPWR VGND sg13g2_decap_8
XFILLER_28_582 VPWR VGND sg13g2_decap_8
XFILLER_43_552 VPWR VGND sg13g2_decap_8
XFILLER_15_232 VPWR VGND sg13g2_decap_8
XFILLER_16_755 VPWR VGND sg13g2_decap_8
XFILLER_31_758 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0710_ u_ppwm_u_ex__0709_/Y VPWR u_ppwm_u_ex__0714_/A VGND hold295/A
+ u_ppwm_u_ex__0585_/Y sg13g2_o21ai_1
XFILLER_12_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0922_ net510 VPWR u_ppwm_u_mem__0922_/Y VGND net427 net324 sg13g2_o21ai_1
XFILLER_8_954 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0641_ u_ppwm_u_ex__0659_/B u_ppwm_u_ex__0711_/A net442 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0853_ u_ppwm_u_mem__0691_/Y u_ppwm_u_mem__0684_/Y net481 u_ppwm_u_mem__0853_/X
+ VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__0572_ u_ppwm_u_ex__0954_/A net455 VPWR VGND sg13g2_inv_2
XFILLER_7_486 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0784_ u_ppwm_u_mem__0784_/Y hold139/A net486 VPWR VGND sg13g2_nand2_1
XFILLER_3_681 VPWR VGND sg13g2_decap_8
XFILLER_39_836 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1124_ net53 VGND VPWR net658 hold289/A clknet_5_4__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__113_ net507 VGND VPWR net632 hold262/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_519 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1055_ u_ppwm_u_ex__1053_/X u_ppwm_u_ex__1029_/Y u_ppwm_u_ex__1052_/Y
+ u_ppwm_u_ex__1055_/X VPWR VGND sg13g2_a21o_1
XFILLER_19_582 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1198_ net137 VGND VPWR u_ppwm_u_mem__1198_/D hold7/A clknet_5_9__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_34_541 VPWR VGND sg13g2_decap_8
XFILLER_22_703 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0908_ hold307/A net384 u_ppwm_u_ex__0908_/Y VPWR VGND sg13g2_nor2_1
XFILLER_30_791 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0839_ u_ppwm_u_ex__0839_/Y u_ppwm_u_ex__0842_/B VPWR VGND net368 sg13g2_nand2b_2
XFILLER_45_828 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1109__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_13_703 VPWR VGND sg13g2_decap_8
XFILLER_40_544 VPWR VGND sg13g2_decap_8
XFILLER_25_596 VPWR VGND sg13g2_decap_8
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_fill_2
XFILLER_4_456 VPWR VGND sg13g2_decap_8
XFILLER_48_600 VPWR VGND sg13g2_decap_8
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_48_677 VPWR VGND sg13g2_decap_8
XFILLER_47_143 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1121_ net120 VGND VPWR u_ppwm_u_mem__1121_/D hold77/A clknet_5_23__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_16_552 VPWR VGND sg13g2_decap_8
XFILLER_18_90 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1052_ net501 VPWR u_ppwm_u_mem__1052_/Y VGND net407 net213 sg13g2_o21ai_1
XFILLER_44_883 VPWR VGND sg13g2_decap_8
XFILLER_31_555 VPWR VGND sg13g2_decap_8
XFILLER_8_751 VPWR VGND sg13g2_decap_8
XFILLER_7_250 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0905_ VGND VPWR net424 u_ppwm_u_mem__0702_/Y hold157/A u_ppwm_u_mem__0904_/Y
+ sg13g2_a21oi_1
XFILLER_7_283 VPWR VGND sg13g2_decap_4
Xhold217 hold217/A VPWR VGND net585 sg13g2_dlygate4sd3_1
Xhold206 hold206/A VPWR VGND net574 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0624_ u_ppwm_u_ex__0622_/X VPWR u_ppwm_u_ex__0624_/Y VGND u_ppwm_u_ex__0614_/Y
+ u_ppwm_u_ex__0623_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__0836_ net467 VPWR u_ppwm_u_mem__0836_/Y VGND u_ppwm_u_mem__0832_/Y
+ u_ppwm_u_mem__0833_/Y sg13g2_o21ai_1
Xhold239 hold239/A VPWR VGND net607 sg13g2_dlygate4sd3_1
Xhold228 hold228/A VPWR VGND net596 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0767_ u_ppwm_u_mem__0767_/Y hold173/A net482 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0698_ VPWR u_ppwm_u_mem__0698_/Y net570 VGND sg13g2_inv_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
XFILLER_22_1004 VPWR VGND sg13g2_decap_8
XFILLER_39_633 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1107_ net37 VGND VPWR u_ppwm_u_ex__1107_/D hold312/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_305 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__1038_ VGND VPWR u_ppwm_u_ex__1054_/A u_ppwm_u_ex__1029_/Y u_ppwm_u_ex__1038_/Y
+ u_ppwm_u_ex__1025_/Y sg13g2_a21oi_1
XFILLER_35_850 VPWR VGND sg13g2_decap_8
XFILLER_22_500 VPWR VGND sg13g2_decap_8
XFILLER_10_717 VPWR VGND sg13g2_decap_8
XFILLER_22_577 VPWR VGND sg13g2_decap_8
XFILLER_2_905 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_23 VPWR VGND sg13g2_fill_2
XFILLER_18_806 VPWR VGND sg13g2_decap_8
XFILLER_45_625 VPWR VGND sg13g2_decap_8
XFILLER_26_883 VPWR VGND sg13g2_decap_8
XFILLER_41_831 VPWR VGND sg13g2_decap_8
XFILLER_40_352 VPWR VGND sg13g2_fill_2
XFILLER_13_577 VPWR VGND sg13g2_decap_8
XFILLER_9_537 VPWR VGND sg13g2_decap_8
XFILLER_5_710 VPWR VGND sg13g2_decap_8
XFILLER_5_787 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0621_ VPWR u_ppwm_u_mem__0621_/Y net537 VGND sg13g2_inv_1
XFILLER_49_942 VPWR VGND sg13g2_decap_8
XFILLER_0_481 VPWR VGND sg13g2_decap_8
XFILLER_48_474 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1104_ VGND VPWR net565 u_ppwm_u_mem__1085_/B hold198/A u_ppwm_u_mem__1103_/C
+ sg13g2_a21oi_1
XFILLER_36_669 VPWR VGND sg13g2_decap_8
XFILLER_23_308 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1035_ VGND VPWR net418 u_ppwm_u_mem__0637_/Y u_ppwm_u_mem__1194_/D
+ u_ppwm_u_mem__1034_/Y sg13g2_a21oi_1
XFILLER_44_680 VPWR VGND sg13g2_decap_8
XFILLER_17_894 VPWR VGND sg13g2_decap_8
XFILLER_31_330 VPWR VGND sg13g2_fill_2
XFILLER_32_864 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0607_ VGND VPWR net218 u_ppwm_u_ex__0606_/Y hold21/A u_ppwm_u_ex__0991_/A
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0819_ hold44/A hold82/A net485 u_ppwm_u_mem__0819_/X VPWR VGND sg13g2_mux2_1
Xfanout505 net506 net505 VPWR VGND sg13g2_buf_8
Xfanout516 net517 net516 VPWR VGND sg13g2_buf_1
XFILLER_39_452 VPWR VGND sg13g2_decap_4
XFILLER_27_669 VPWR VGND sg13g2_decap_8
XFILLER_42_628 VPWR VGND sg13g2_decap_8
XFILLER_23_853 VPWR VGND sg13g2_decap_8
XFILLER_10_514 VPWR VGND sg13g2_decap_8
XFILLER_2_702 VPWR VGND sg13g2_decap_8
XFILLER_2_779 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_46_923 VPWR VGND sg13g2_decap_8
XFILLER_18_603 VPWR VGND sg13g2_decap_8
XFILLER_45_422 VPWR VGND sg13g2_decap_8
XFILLER_17_168 VPWR VGND sg13g2_fill_1
XFILLER_33_617 VPWR VGND sg13g2_decap_8
XFILLER_45_499 VPWR VGND sg13g2_decap_8
XFILLER_26_680 VPWR VGND sg13g2_decap_8
XFILLER_14_853 VPWR VGND sg13g2_decap_8
XFILLER_15_80 VPWR VGND sg13g2_fill_2
XFILLER_9_345 VPWR VGND sg13g2_fill_2
XFILLER_12_1014 VPWR VGND sg13g2_decap_8
XFILLER_5_584 VPWR VGND sg13g2_decap_8
XFILLER_48_271 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__244__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_37_934 VPWR VGND sg13g2_decap_8
XFILLER_17_691 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1018_ net499 VPWR u_ppwm_u_mem__1018_/Y VGND net414 hold51/A sg13g2_o21ai_1
XFILLER_20_823 VPWR VGND sg13g2_decap_8
XFILLER_32_661 VPWR VGND sg13g2_decap_8
Xfanout357 net358 net357 VPWR VGND sg13g2_buf_8
Xfanout368 net369 net368 VPWR VGND sg13g2_buf_8
Xfanout379 net380 net379 VPWR VGND sg13g2_buf_8
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_43_937 VPWR VGND sg13g2_decap_8
XFILLER_42_425 VPWR VGND sg13g2_decap_8
XFILLER_15_628 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1228__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_23_650 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_11_812 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_2_576 VPWR VGND sg13g2_decap_8
XFILLER_37_219 VPWR VGND sg13g2_decap_8
XFILLER_46_720 VPWR VGND sg13g2_decap_8
XFILLER_19_967 VPWR VGND sg13g2_decap_8
XFILLER_34_926 VPWR VGND sg13g2_decap_8
XFILLER_46_797 VPWR VGND sg13g2_decap_8
XFILLER_45_296 VPWR VGND sg13g2_fill_1
XFILLER_14_650 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0941_ u_ppwm_u_ex__0941_/Y u_ppwm_u_ex__0845_/B net368 u_ppwm_u_ex__0838_/B
+ u_ppwm_u_ex__0800_/X VPWR VGND sg13g2_a22oi_1
XFILLER_42_992 VPWR VGND sg13g2_decap_8
XFILLER_9_142 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0872_ u_ppwm_u_ex__0872_/Y u_ppwm_u_ex__0871_/X u_ppwm_u_ex__0796_/Y
+ u_ppwm_u_ex__0814_/A u_ppwm_u_ex__0789_/Y VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_pwm__188_ u_ppwm_u_pwm__188_/A u_ppwm_u_pwm__188_/B u_ppwm_u_pwm__247_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_83 VPWR VGND sg13g2_fill_1
XFILLER_37_731 VPWR VGND sg13g2_decap_8
XFILLER_25_904 VPWR VGND sg13g2_decap_8
XFILLER_19_1009 VPWR VGND sg13g2_decap_8
XFILLER_40_929 VPWR VGND sg13g2_decap_8
XFILLER_33_981 VPWR VGND sg13g2_decap_8
XFILLER_20_620 VPWR VGND sg13g2_decap_8
XFILLER_20_697 VPWR VGND sg13g2_decap_8
XFILLER_3_329 VPWR VGND sg13g2_fill_1
XFILLER_28_764 VPWR VGND sg13g2_decap_8
XFILLER_43_734 VPWR VGND sg13g2_decap_8
XFILLER_16_937 VPWR VGND sg13g2_decap_8
XFILLER_30_417 VPWR VGND sg13g2_fill_1
XFILLER_6_112 VPWR VGND sg13g2_decap_4
XFILLER_11_686 VPWR VGND sg13g2_decap_8
XFILLER_7_668 VPWR VGND sg13g2_decap_8
XFILLER_3_863 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1071_ u_ppwm_u_ex__1072_/B u_ppwm_u_ex__1071_/A net349 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_global_counter__060_ net398 net445 u_ppwm_u_global_counter__106_/D VPWR
+ VGND sg13g2_xor2_1
XFILLER_19_764 VPWR VGND sg13g2_decap_8
XFILLER_46_594 VPWR VGND sg13g2_decap_8
XFILLER_34_723 VPWR VGND sg13g2_decap_8
XFILLER_33_233 VPWR VGND sg13g2_decap_4
XFILLER_33_266 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0924_ u_ppwm_u_ex__0924_/B u_ppwm_u_ex__0924_/A u_ppwm_u_ex__0924_/X
+ VPWR VGND sg13g2_xor2_1
XFILLER_15_992 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0855_ u_ppwm_u_ex__0855_/Y net364 net440 net367 net443 VPWR VGND sg13g2_a22oi_1
XFILLER_30_973 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0998_ net498 VPWR u_ppwm_u_mem__0998_/Y VGND net411 hold211/A sg13g2_o21ai_1
Xu_ppwm_u_ex__0786_ u_ppwm_u_ex__0785_/Y VPWR u_ppwm_u_ex__0786_/Y VGND net359 u_ppwm_u_ex__0778_/Y
+ sg13g2_o21ai_1
XFILLER_25_1002 VPWR VGND sg13g2_decap_8
XFILLER_29_539 VPWR VGND sg13g2_decap_8
XFILLER_25_701 VPWR VGND sg13g2_decap_8
XFILLER_40_726 VPWR VGND sg13g2_decap_8
XFILLER_24_266 VPWR VGND sg13g2_decap_4
XFILLER_25_778 VPWR VGND sg13g2_decap_8
XFILLER_12_439 VPWR VGND sg13g2_fill_1
XFILLER_20_494 VPWR VGND sg13g2_decap_8
XFILLER_21_995 VPWR VGND sg13g2_decap_8
XFILLER_4_638 VPWR VGND sg13g2_decap_8
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_859 VPWR VGND sg13g2_decap_8
XFILLER_47_347 VPWR VGND sg13g2_decap_8
XFILLER_16_734 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_43_531 VPWR VGND sg13g2_decap_8
XFILLER_31_737 VPWR VGND sg13g2_decap_8
XFILLER_12_951 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0921_ VGND VPWR net426 u_ppwm_u_mem__0694_/Y hold127/A u_ppwm_u_mem__0920_/Y
+ sg13g2_a21oi_1
XFILLER_8_933 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0640_ u_ppwm_u_ex__0640_/A net684 hold317/A VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0852_ VPWR VGND u_ppwm_u_mem__0851_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0850_/Y
+ u_ppwm_u_mem__0845_/Y u_ppwm_u_mem__0852_/Y u_ppwm_u_mem__0847_/Y sg13g2_a221oi_1
Xu_ppwm_u_ex__0571_ VPWR u_ppwm_u_ex__0683_/A net454 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0783_ VPWR VGND u_ppwm_u_mem__0782_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0780_/Y
+ u_ppwm_u_mem__0776_/Y u_ppwm_u_mem__0783_/Y u_ppwm_u_mem__0778_/Y sg13g2_a221oi_1
XFILLER_48_1013 VPWR VGND sg13g2_decap_8
XFILLER_3_660 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_815 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__112_ net507 VGND VPWR net605 hold236/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1123_ net40 VGND VPWR u_ppwm_u_ex__1123_/D hold295/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_mem__1138__86 VPWR VGND net86 sg13g2_tiehi
Xu_ppwm_u_mem__1153__56 VPWR VGND net56 sg13g2_tiehi
Xu_ppwm_u_ex__1054_ u_ppwm_u_ex__1075_/B u_ppwm_u_ex__1054_/A u_ppwm_u_ex__1054_/B
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_561 VPWR VGND sg13g2_decap_8
XFILLER_46_391 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1197_ net145 VGND VPWR net206 hold59/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_22_759 VPWR VGND sg13g2_decap_8
XFILLER_34_597 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0907_ VGND VPWR net368 u_ppwm_u_ex__0799_/Y u_ppwm_u_ex__0907_/Y u_ppwm_u_ex__0906_/Y
+ sg13g2_a21oi_1
XFILLER_30_770 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1208__57 VPWR VGND net57 sg13g2_tiehi
Xu_ppwm_u_ex__0838_ net368 u_ppwm_u_ex__0838_/B u_ppwm_u_ex__0838_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0769_ u_ppwm_u_ex__0769_/A u_ppwm_u_ex__0769_/B u_ppwm_u_ex__0769_/C
+ u_ppwm_u_ex__0769_/D u_ppwm_u_ex__0769_/Y VPWR VGND sg13g2_nor4_1
XFILLER_45_807 VPWR VGND sg13g2_decap_8
XFILLER_17_509 VPWR VGND sg13g2_decap_8
XFILLER_37_380 VPWR VGND sg13g2_fill_1
XFILLER_25_575 VPWR VGND sg13g2_decap_8
XFILLER_40_523 VPWR VGND sg13g2_decap_8
XFILLER_13_759 VPWR VGND sg13g2_decap_8
XFILLER_9_719 VPWR VGND sg13g2_decap_8
XFILLER_21_792 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_pwm__231__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_4_435 VPWR VGND sg13g2_decap_8
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_48_656 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1120_ net122 VGND VPWR net276 hold95/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_531 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1051_ VGND VPWR net407 u_ppwm_u_mem__0629_/Y hold16/A u_ppwm_u_mem__1050_/Y
+ sg13g2_a21oi_1
XFILLER_28_380 VPWR VGND sg13g2_fill_2
XFILLER_35_339 VPWR VGND sg13g2_fill_1
XFILLER_44_862 VPWR VGND sg13g2_decap_8
XFILLER_31_534 VPWR VGND sg13g2_decap_8
XFILLER_8_730 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0904_ net514 VPWR u_ppwm_u_mem__0904_/Y VGND net424 net282 sg13g2_o21ai_1
Xhold207 hold207/A VPWR VGND net575 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0623_ net469 u_ppwm_u_ex__0623_/B u_ppwm_u_ex__0623_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0835_ net470 u_ppwm_u_mem__0835_/B u_ppwm_u_mem__0835_/Y VPWR VGND
+ sg13g2_nor2_1
Xhold218 hold218/A VPWR VGND net586 sg13g2_dlygate4sd3_1
Xhold229 hold229/A VPWR VGND net597 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0766_ u_ppwm_u_mem__0765_/Y VPWR u_ppwm_u_mem__0766_/Y VGND u_ppwm_u_mem__0696_/Y
+ net483 sg13g2_o21ai_1
Xu_ppwm_u_mem__0697_ VPWR u_ppwm_u_mem__0697_/Y net288 VGND sg13g2_inv_1
XFILLER_38_100 VPWR VGND sg13g2_decap_8
XFILLER_39_612 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1106_ net39 VGND VPWR net688 hold319/A clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_328 VPWR VGND sg13g2_fill_1
XFILLER_39_689 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1037_ u_ppwm_u_ex__1037_/A u_ppwm_u_ex__1035_/Y u_ppwm_u_ex__1119_/D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_22_556 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_45_604 VPWR VGND sg13g2_decap_8
XFILLER_17_306 VPWR VGND sg13g2_fill_2
XFILLER_41_810 VPWR VGND sg13g2_decap_8
XFILLER_26_862 VPWR VGND sg13g2_decap_8
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_9_516 VPWR VGND sg13g2_decap_8
XFILLER_13_556 VPWR VGND sg13g2_decap_8
XFILLER_41_887 VPWR VGND sg13g2_decap_8
XFILLER_5_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0620_ VPWR u_ppwm_u_mem__0620_/Y net343 VGND sg13g2_inv_1
XFILLER_49_921 VPWR VGND sg13g2_decap_8
XFILLER_0_460 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
XFILLER_48_453 VPWR VGND sg13g2_decap_8
XFILLER_49_998 VPWR VGND sg13g2_decap_8
Xhold90 hold90/A VPWR VGND net288 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1103_ u_ppwm_u_mem__1103_/A net588 u_ppwm_u_mem__1103_/C hold221/A
+ VPWR VGND sg13g2_nor3_1
XFILLER_36_648 VPWR VGND sg13g2_decap_8
XFILLER_17_873 VPWR VGND sg13g2_decap_8
XFILLER_35_169 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1034_ net501 VPWR u_ppwm_u_mem__1034_/Y VGND net418 net230 sg13g2_o21ai_1
XFILLER_32_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0606_ u_ppwm_u_ex__0772_/C u_ppwm_u_ex__0715_/B net446 u_ppwm_u_ex__0606_/Y
+ VPWR VGND net369 sg13g2_nand4_1
Xu_ppwm_u_mem__0818_ u_ppwm_u_mem__0818_/Y net475 u_ppwm_u_mem__0818_/B VPWR VGND
+ sg13g2_nand2_1
Xfanout506 net518 net506 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0749_ VPWR VGND u_ppwm_u_mem__0748_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0746_/Y
+ u_ppwm_u_mem__0743_/Y u_ppwm_u_mem__0749_/Y u_ppwm_u_mem__0744_/Y sg13g2_a221oi_1
Xfanout517 net518 net517 VPWR VGND sg13g2_buf_2
XFILLER_6_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_420 VPWR VGND sg13g2_decap_4
XFILLER_39_486 VPWR VGND sg13g2_decap_8
XFILLER_27_648 VPWR VGND sg13g2_decap_8
XFILLER_42_607 VPWR VGND sg13g2_decap_8
XFILLER_23_832 VPWR VGND sg13g2_decap_8
XFILLER_22_320 VPWR VGND sg13g2_fill_2
XFILLER_22_397 VPWR VGND sg13g2_fill_1
XFILLER_2_758 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1196__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_46_902 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1157__167 VPWR VGND net167 sg13g2_tiehi
XFILLER_45_401 VPWR VGND sg13g2_decap_8
XFILLER_18_659 VPWR VGND sg13g2_decap_8
XFILLER_46_979 VPWR VGND sg13g2_decap_8
XFILLER_45_478 VPWR VGND sg13g2_decap_8
XFILLER_14_832 VPWR VGND sg13g2_decap_8
XFILLER_32_128 VPWR VGND sg13g2_fill_2
XFILLER_41_684 VPWR VGND sg13g2_decap_8
XFILLER_9_324 VPWR VGND sg13g2_fill_1
XFILLER_5_563 VPWR VGND sg13g2_decap_8
XFILLER_0_290 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_49_795 VPWR VGND sg13g2_decap_8
XFILLER_48_250 VPWR VGND sg13g2_decap_8
XFILLER_37_913 VPWR VGND sg13g2_decap_8
XFILLER_17_670 VPWR VGND sg13g2_decap_8
XFILLER_23_117 VPWR VGND sg13g2_decap_8
XFILLER_23_128 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1017_ VGND VPWR net414 u_ppwm_u_mem__0646_/Y hold52/A u_ppwm_u_mem__1016_/Y
+ sg13g2_a21oi_1
XFILLER_32_640 VPWR VGND sg13g2_decap_8
XFILLER_20_802 VPWR VGND sg13g2_decap_8
XFILLER_9_880 VPWR VGND sg13g2_decap_8
XFILLER_20_879 VPWR VGND sg13g2_decap_8
Xfanout369 fanout369/A net369 VPWR VGND sg13g2_buf_1
Xfanout358 fanout358/A net358 VPWR VGND sg13g2_buf_8
XFILLER_39_250 VPWR VGND sg13g2_decap_4
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_43_916 VPWR VGND sg13g2_decap_8
XFILLER_15_607 VPWR VGND sg13g2_decap_8
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_6_316 VPWR VGND sg13g2_fill_1
XFILLER_11_868 VPWR VGND sg13g2_decap_8
XFILLER_2_555 VPWR VGND sg13g2_decap_8
XFILLER_19_946 VPWR VGND sg13g2_decap_8
XFILLER_46_776 VPWR VGND sg13g2_decap_8
XFILLER_45_253 VPWR VGND sg13g2_decap_8
XFILLER_34_905 VPWR VGND sg13g2_decap_8
XFILLER_45_275 VPWR VGND sg13g2_decap_8
XFILLER_33_437 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0940_ u_ppwm_u_ex__0939_/Y VPWR u_ppwm_u_ex__0940_/Y VGND u_ppwm_u_ex__0937_/Y
+ u_ppwm_u_ex__0950_/D sg13g2_o21ai_1
XFILLER_42_971 VPWR VGND sg13g2_decap_8
XFILLER_41_481 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0871_ u_ppwm_u_ex__0845_/B u_ppwm_u_ex__0870_/Y net377 u_ppwm_u_ex__0871_/X
+ VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_pwm__187_ u_ppwm_u_pwm__187_/B net644 u_ppwm_u_pwm__188_/B VPWR VGND sg13g2_xor2_1
XFILLER_37_710 VPWR VGND sg13g2_decap_8
XFILLER_49_592 VPWR VGND sg13g2_decap_8
XFILLER_3_1024 VPWR VGND sg13g2_decap_4
XFILLER_36_242 VPWR VGND sg13g2_decap_4
XFILLER_36_275 VPWR VGND sg13g2_fill_2
XFILLER_37_787 VPWR VGND sg13g2_decap_8
XFILLER_40_908 VPWR VGND sg13g2_decap_8
XFILLER_33_960 VPWR VGND sg13g2_decap_8
XFILLER_20_676 VPWR VGND sg13g2_decap_8
XFILLER_47_529 VPWR VGND sg13g2_decap_8
XFILLER_47_46 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_fill_2
XFILLER_28_743 VPWR VGND sg13g2_decap_8
XFILLER_16_916 VPWR VGND sg13g2_decap_8
XFILLER_43_713 VPWR VGND sg13g2_decap_8
XFILLER_15_426 VPWR VGND sg13g2_fill_2
XFILLER_31_919 VPWR VGND sg13g2_decap_8
XFILLER_10_131 VPWR VGND sg13g2_fill_2
XFILLER_11_665 VPWR VGND sg13g2_decap_8
XFILLER_10_153 VPWR VGND sg13g2_fill_2
XFILLER_7_647 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1202__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_3_842 VPWR VGND sg13g2_decap_8
XFILLER_38_529 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1070_ VGND VPWR u_ppwm_u_ex__1068_/Y u_ppwm_u_ex__1069_/Y u_ppwm_u_ex__1072_/A
+ net361 sg13g2_a21oi_1
XFILLER_18_220 VPWR VGND sg13g2_fill_2
XFILLER_19_743 VPWR VGND sg13g2_decap_8
XFILLER_34_702 VPWR VGND sg13g2_decap_8
XFILLER_46_573 VPWR VGND sg13g2_decap_8
XFILLER_15_971 VPWR VGND sg13g2_decap_8
XFILLER_34_779 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0923_ u_ppwm_u_ex__0952_/A VPWR u_ppwm_u_ex__0924_/B VGND u_ppwm_u_ex__0884_/Y
+ u_ppwm_u_ex__0950_/C sg13g2_o21ai_1
Xu_ppwm_u_ex__0854_ u_ppwm_u_ex__0851_/X u_ppwm_u_ex__0849_/Y u_ppwm_u_ex__0853_/Y
+ u_ppwm_u_ex__0859_/C VPWR VGND sg13g2_a21o_1
XFILLER_30_952 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0997_ VGND VPWR net410 u_ppwm_u_mem__0656_/Y u_ppwm_u_mem__1175_/D
+ u_ppwm_u_mem__0996_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__239_ net189 VGND VPWR net550 hold181/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__0785_ u_ppwm_u_ex__0785_/Y u_ppwm_u_ex__0856_/B net382 u_ppwm_u_ex__0783_/X
+ u_ppwm_u_ex__0780_/X VPWR VGND sg13g2_a22oi_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_5_190 VPWR VGND sg13g2_fill_2
XFILLER_29_518 VPWR VGND sg13g2_decap_8
XFILLER_37_584 VPWR VGND sg13g2_decap_8
XFILLER_24_234 VPWR VGND sg13g2_fill_1
XFILLER_24_245 VPWR VGND sg13g2_decap_8
XFILLER_25_757 VPWR VGND sg13g2_decap_8
XFILLER_40_705 VPWR VGND sg13g2_decap_8
XFILLER_21_974 VPWR VGND sg13g2_decap_8
XFILLER_32_1018 VPWR VGND sg13g2_decap_8
XFILLER_20_473 VPWR VGND sg13g2_decap_8
XFILLER_4_617 VPWR VGND sg13g2_decap_8
XFILLER_3_149 VPWR VGND sg13g2_decap_8
XFILLER_0_845 VPWR VGND sg13g2_decap_8
XFILLER_48_838 VPWR VGND sg13g2_decap_8
XFILLER_47_326 VPWR VGND sg13g2_decap_8
XFILLER_28_540 VPWR VGND sg13g2_decap_8
XFILLER_43_510 VPWR VGND sg13g2_decap_8
XFILLER_16_713 VPWR VGND sg13g2_decap_8
XFILLER_43_587 VPWR VGND sg13g2_decap_8
XFILLER_31_716 VPWR VGND sg13g2_decap_8
XFILLER_12_930 VPWR VGND sg13g2_decap_8
XFILLER_8_912 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0920_ net510 VPWR u_ppwm_u_mem__0920_/Y VGND net426 hold186/A sg13g2_o21ai_1
XFILLER_7_400 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0851_ VGND VPWR net395 u_ppwm_u_mem__0848_/X u_ppwm_u_mem__0851_/Y
+ net394 sg13g2_a21oi_1
XFILLER_8_989 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0570_ VPWR u_ppwm_u_ex__0570_/Y net451 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0782_ VGND VPWR net395 u_ppwm_u_mem__0781_/X u_ppwm_u_mem__0782_/Y
+ net470 sg13g2_a21oi_1
Xu_ppwm_u_ex__1122_ net28 VGND VPWR u_ppwm_u_ex__1122_/D hold294/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__111_ net507 VGND VPWR net629 hold259/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_17_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1053_ u_ppwm_u_ex__1054_/A u_ppwm_u_ex__1054_/B u_ppwm_u_ex__1053_/X
+ VPWR VGND sg13g2_and2_1
XFILLER_19_540 VPWR VGND sg13g2_decap_8
XFILLER_47_893 VPWR VGND sg13g2_decap_8
XFILLER_46_370 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_63 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1196_ net150 VGND VPWR u_ppwm_u_mem__1196_/D hold34/A clknet_5_13__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_34_576 VPWR VGND sg13g2_decap_8
XFILLER_22_738 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0906_ u_ppwm_u_ex__0905_/Y VPWR u_ppwm_u_ex__0906_/Y VGND u_ppwm_u_ex__0821_/X
+ u_ppwm_u_ex__0839_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__0837_ u_ppwm_u_ex__0842_/B net375 net377 VPWR VGND sg13g2_nand2_2
Xu_ppwm_u_ex__0768_ u_ppwm_u_ex__0767_/Y VPWR u_ppwm_u_ex__0768_/Y VGND u_ppwm_u_ex__0763_/Y
+ u_ppwm_u_ex__0765_/Y sg13g2_o21ai_1
XFILLER_1_609 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0699_ VGND VPWR u_ppwm_u_ex__0695_/Y u_ppwm_u_ex__0698_/Y u_ppwm_u_ex__0699_/Y
+ u_ppwm_u_ex__0694_/Y sg13g2_a21oi_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_28_48 VPWR VGND sg13g2_fill_2
XFILLER_38_893 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_44_36 VPWR VGND sg13g2_decap_4
XFILLER_40_502 VPWR VGND sg13g2_decap_8
XFILLER_25_554 VPWR VGND sg13g2_decap_8
XFILLER_13_738 VPWR VGND sg13g2_decap_8
XFILLER_40_579 VPWR VGND sg13g2_decap_8
XFILLER_21_771 VPWR VGND sg13g2_decap_8
XFILLER_20_281 VPWR VGND sg13g2_fill_2
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_0_642 VPWR VGND sg13g2_decap_8
XFILLER_48_635 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1050_ net501 VPWR u_ppwm_u_mem__1050_/Y VGND net408 hold141/A sg13g2_o21ai_1
XFILLER_29_882 VPWR VGND sg13g2_decap_8
XFILLER_44_841 VPWR VGND sg13g2_decap_8
XFILLER_16_510 VPWR VGND sg13g2_decap_8
XFILLER_16_587 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1167__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_15_1013 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0903_ VGND VPWR net424 u_ppwm_u_mem__0703_/Y hold85/A u_ppwm_u_mem__0902_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0834_ net478 hold108/A hold99/A hold172/A hold212/A net471 u_ppwm_u_mem__0835_/B
+ VPWR VGND sg13g2_mux4_1
XFILLER_8_786 VPWR VGND sg13g2_decap_8
Xhold208 hold208/A VPWR VGND net576 sg13g2_dlygate4sd3_1
Xu_ppwm_u_ex__0622_ VGND VPWR u_ppwm_u_ex__0622_/X u_ppwm_u_ex__0622_/B net469 sg13g2_or2_1
Xhold219 hold219/A VPWR VGND net587 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0765_ u_ppwm_u_mem__0765_/Y hold22/A net483 VPWR VGND sg13g2_nand2_1
XFILLER_4_981 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0696_ VPWR u_ppwm_u_mem__0696_/Y net329 VGND sg13g2_inv_1
Xu_ppwm_u_ex__1105_ net41 VGND VPWR net661 fanout466/A clknet_5_19__leaf_clk sg13g2_dfrbpq_2
XFILLER_39_668 VPWR VGND sg13g2_decap_8
XFILLER_47_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1036_ net505 VPWR u_ppwm_u_ex__1037_/A VGND net449 net349 sg13g2_o21ai_1
Xu_ppwm_u_mem__1179_ net99 VGND VPWR net235 hold57/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_35_885 VPWR VGND sg13g2_decap_8
XFILLER_22_535 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_26_841 VPWR VGND sg13g2_decap_8
XFILLER_38_690 VPWR VGND sg13g2_decap_8
XFILLER_13_535 VPWR VGND sg13g2_decap_8
XFILLER_25_373 VPWR VGND sg13g2_fill_1
XFILLER_41_866 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1140__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_40_354 VPWR VGND sg13g2_fill_1
XFILLER_5_745 VPWR VGND sg13g2_decap_8
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_49_900 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_49_977 VPWR VGND sg13g2_decap_8
XFILLER_48_432 VPWR VGND sg13g2_decap_8
Xhold80 hold80/A VPWR VGND net278 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1102_ net587 hold250/A hold238/A u_ppwm_u_mem__1102_/D u_ppwm_u_mem__1103_/C
+ VPWR VGND sg13g2_and4_1
Xhold91 hold91/A VPWR VGND net289 sg13g2_dlygate4sd3_1
XFILLER_36_627 VPWR VGND sg13g2_decap_8
XFILLER_17_852 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1033_ VGND VPWR net418 u_ppwm_u_mem__0638_/Y hold33/A u_ppwm_u_mem__1032_/Y
+ sg13g2_a21oi_1
XFILLER_32_822 VPWR VGND sg13g2_decap_8
XFILLER_32_899 VPWR VGND sg13g2_decap_8
XFILLER_8_583 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0605_ hold20/A u_ppwm_u_ex__0605_/A net217 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0817_ hold190/A hold64/A net485 u_ppwm_u_mem__0818_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0748_ VGND VPWR net472 u_ppwm_u_mem__0747_/X u_ppwm_u_mem__0748_/Y
+ net394 sg13g2_a21oi_1
Xu_ppwm_u_mem__0679_ VPWR u_ppwm_u_mem__0679_/Y net542 VGND sg13g2_inv_1
Xfanout507 net509 net507 VPWR VGND sg13g2_buf_8
Xfanout518 rst_n net518 VPWR VGND sg13g2_buf_8
XFILLER_27_627 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1019_ net387 u_ppwm_u_ex__1019_/B net362 u_ppwm_u_ex__1019_/Y VPWR VGND
+ sg13g2_nor3_1
XFILLER_26_148 VPWR VGND sg13g2_fill_2
XFILLER_22_310 VPWR VGND sg13g2_fill_1
XFILLER_23_811 VPWR VGND sg13g2_decap_8
XFILLER_25_38 VPWR VGND sg13g2_decap_4
XFILLER_35_682 VPWR VGND sg13g2_decap_8
XFILLER_22_365 VPWR VGND sg13g2_fill_2
XFILLER_22_376 VPWR VGND sg13g2_fill_1
XFILLER_23_888 VPWR VGND sg13g2_decap_8
XFILLER_10_549 VPWR VGND sg13g2_decap_8
XFILLER_2_737 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_46_958 VPWR VGND sg13g2_decap_8
XFILLER_18_638 VPWR VGND sg13g2_decap_8
XFILLER_45_457 VPWR VGND sg13g2_decap_8
XFILLER_14_811 VPWR VGND sg13g2_decap_8
XFILLER_13_343 VPWR VGND sg13g2_decap_8
XFILLER_41_663 VPWR VGND sg13g2_decap_8
XFILLER_14_888 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_fill_1
XFILLER_5_542 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_49_774 VPWR VGND sg13g2_decap_8
XFILLER_37_969 VPWR VGND sg13g2_decap_8
XFILLER_24_619 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1016_ net498 VPWR u_ppwm_u_mem__1016_/Y VGND net414 hold124/A sg13g2_o21ai_1
XFILLER_31_151 VPWR VGND sg13g2_fill_2
XFILLER_20_858 VPWR VGND sg13g2_decap_8
XFILLER_32_696 VPWR VGND sg13g2_decap_8
XFILLER_8_380 VPWR VGND sg13g2_fill_2
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
Xfanout359 fanout361/A net359 VPWR VGND sg13g2_buf_8
XFILLER_28_925 VPWR VGND sg13g2_decap_8
XFILLER_36_15 VPWR VGND sg13g2_decap_4
XFILLER_36_991 VPWR VGND sg13g2_decap_8
XFILLER_23_685 VPWR VGND sg13g2_decap_8
XFILLER_11_847 VPWR VGND sg13g2_decap_8
XFILLER_7_829 VPWR VGND sg13g2_decap_8
XFILLER_2_534 VPWR VGND sg13g2_decap_8
XFILLER_19_925 VPWR VGND sg13g2_decap_8
XFILLER_46_755 VPWR VGND sg13g2_decap_8
XFILLER_27_991 VPWR VGND sg13g2_decap_8
XFILLER_42_950 VPWR VGND sg13g2_decap_8
XFILLER_41_460 VPWR VGND sg13g2_decap_8
XFILLER_9_111 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0870_ VGND VPWR u_ppwm_u_ex__0735_/A net384 u_ppwm_u_ex__0870_/Y u_ppwm_u_ex__0869_/Y
+ sg13g2_a21oi_1
XFILLER_14_685 VPWR VGND sg13g2_decap_8
XFILLER_9_188 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__186_ net593 net546 hold276/A hold226/A VPWR VGND hold268/A sg13g2_nand4_1
XFILLER_6_884 VPWR VGND sg13g2_decap_8
XFILLER_3_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_37_766 VPWR VGND sg13g2_decap_8
XFILLER_24_405 VPWR VGND sg13g2_fill_1
XFILLER_25_939 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0999_ VGND VPWR u_ppwm_u_ex__0997_/Y u_ppwm_u_ex__0998_/Y u_ppwm_u_ex__1000_/D
+ net360 sg13g2_a21oi_1
XFILLER_20_655 VPWR VGND sg13g2_decap_8
XFILLER_47_508 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_41_1020 VPWR VGND sg13g2_decap_8
XFILLER_28_722 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_43_769 VPWR VGND sg13g2_decap_8
XFILLER_24_983 VPWR VGND sg13g2_decap_8
XFILLER_30_408 VPWR VGND sg13g2_fill_2
XFILLER_23_482 VPWR VGND sg13g2_decap_8
XFILLER_11_644 VPWR VGND sg13g2_decap_8
XFILLER_7_626 VPWR VGND sg13g2_decap_8
XFILLER_3_821 VPWR VGND sg13g2_decap_8
XFILLER_3_898 VPWR VGND sg13g2_decap_8
XFILLER_38_508 VPWR VGND sg13g2_decap_8
XFILLER_19_722 VPWR VGND sg13g2_decap_8
XFILLER_46_552 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_18_254 VPWR VGND sg13g2_fill_1
XFILLER_19_799 VPWR VGND sg13g2_decap_8
XFILLER_34_758 VPWR VGND sg13g2_decap_8
XFILLER_15_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0922_ u_ppwm_u_ex__0950_/C u_ppwm_u_ex__0922_/B u_ppwm_u_ex__0881_/Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_30_931 VPWR VGND sg13g2_decap_8
XFILLER_41_290 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0853_ u_ppwm_u_ex__0780_/X VPWR u_ppwm_u_ex__0853_/Y VGND u_ppwm_u_ex__0849_/Y
+ u_ppwm_u_ex__0851_/X sg13g2_o21ai_1
Xu_ppwm_u_pwm__238_ net191 VGND VPWR u_ppwm_u_pwm__238_/D hold279/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__0784_ u_ppwm_u_ex__0784_/A u_ppwm_u_ex__0819_/C u_ppwm_u_ex__0856_/B
+ VPWR VGND sg13g2_nor2_2
Xu_ppwm_u_mem__0996_ net496 VPWR u_ppwm_u_mem__0996_/Y VGND net410 net297 sg13g2_o21ai_1
XFILLER_6_681 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__169_ net651 u_ppwm_u_pwm__170_/B u_ppwm_u_pwm__171_/B VPWR VGND sg13g2_nor2_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_37_563 VPWR VGND sg13g2_decap_8
XFILLER_25_736 VPWR VGND sg13g2_decap_8
XFILLER_33_38 VPWR VGND sg13g2_fill_1
XFILLER_21_953 VPWR VGND sg13g2_decap_8
XFILLER_32_290 VPWR VGND sg13g2_fill_2
XFILLER_20_452 VPWR VGND sg13g2_decap_8
XFILLER_0_824 VPWR VGND sg13g2_decap_8
XFILLER_48_817 VPWR VGND sg13g2_decap_8
XFILLER_47_305 VPWR VGND sg13g2_decap_8
XFILLER_28_596 VPWR VGND sg13g2_decap_8
XFILLER_43_566 VPWR VGND sg13g2_decap_8
XFILLER_15_246 VPWR VGND sg13g2_decap_8
XFILLER_16_769 VPWR VGND sg13g2_decap_8
XFILLER_24_780 VPWR VGND sg13g2_decap_8
XFILLER_30_205 VPWR VGND sg13g2_decap_4
XFILLER_12_986 VPWR VGND sg13g2_decap_8
XFILLER_23_82 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0850_ u_ppwm_u_mem__0850_/Y net471 u_ppwm_u_mem__0850_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_8_968 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0781_ hold117/A hold105/A net478 u_ppwm_u_mem__0781_/X VPWR VGND sg13g2_mux2_1
XFILLER_3_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__110_ net507 VGND VPWR net591 hold222/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1121_ net36 VGND VPWR u_ppwm_u_ex__1121_/D hold303/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1052_ VGND VPWR u_ppwm_u_ex__0651_/A u_ppwm_u_ex__1025_/A u_ppwm_u_ex__1052_/Y
+ u_ppwm_u_ex__1049_/B sg13g2_a21oi_1
XFILLER_47_872 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1195_ net154 VGND VPWR net233 hold107/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_596 VPWR VGND sg13g2_decap_8
XFILLER_22_717 VPWR VGND sg13g2_decap_8
XFILLER_34_555 VPWR VGND sg13g2_decap_8
XFILLER_21_216 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0905_ VGND VPWR u_ppwm_u_ex__0792_/Y u_ppwm_u_ex__0838_/B u_ppwm_u_ex__0905_/Y
+ u_ppwm_u_ex__0819_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0836_ net375 net377 u_ppwm_u_ex__0838_/B VPWR VGND sg13g2_and2_1
Xu_ppwm_u_mem__0979_ VGND VPWR net413 u_ppwm_u_mem__0665_/Y u_ppwm_u_mem__1166_/D
+ u_ppwm_u_mem__0978_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0767_ net382 net386 net378 u_ppwm_u_ex__0767_/D u_ppwm_u_ex__0767_/Y
+ VPWR VGND sg13g2_nor4_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0698_ u_ppwm_u_ex__0698_/Y hold310/A u_ppwm_u_ex__0998_/B2 VPWR VGND
+ sg13g2_nand2b_1
XFILLER_9_1020 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_29_316 VPWR VGND sg13g2_fill_1
XFILLER_38_872 VPWR VGND sg13g2_decap_8
XFILLER_25_533 VPWR VGND sg13g2_decap_8
XFILLER_13_717 VPWR VGND sg13g2_decap_8
XFILLER_40_558 VPWR VGND sg13g2_decap_8
XFILLER_21_750 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
XFILLER_0_621 VPWR VGND sg13g2_decap_8
XFILLER_48_614 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_decap_8
XFILLER_36_809 VPWR VGND sg13g2_decap_8
XFILLER_47_179 VPWR VGND sg13g2_decap_8
XFILLER_29_861 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_decap_8
XFILLER_16_566 VPWR VGND sg13g2_decap_8
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_31_569 VPWR VGND sg13g2_decap_8
XFILLER_12_783 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0902_ net513 VPWR u_ppwm_u_mem__0902_/Y VGND net424 hold149/A sg13g2_o21ai_1
XFILLER_8_765 VPWR VGND sg13g2_decap_8
XFILLER_11_293 VPWR VGND sg13g2_decap_4
XFILLER_7_275 VPWR VGND sg13g2_fill_2
XFILLER_7_264 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0621_ VGND VPWR u_ppwm_u_ex__0615_/Y u_ppwm_u_ex__0619_/X u_ppwm_u_ex__1100_/D
+ u_ppwm_u_ex__0620_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0833_ net470 VPWR u_ppwm_u_mem__0833_/Y VGND u_ppwm_u_mem__0828_/Y
+ u_ppwm_u_mem__0829_/Y sg13g2_o21ai_1
Xhold209 hold209/A VPWR VGND net577 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0764_ VGND VPWR u_ppwm_u_mem__0760_/Y u_ppwm_u_mem__0761_/Y u_ppwm_u_mem__0764_/Y
+ u_ppwm_u_mem__0763_/Y sg13g2_a21oi_1
XFILLER_4_960 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0695_ VPWR u_ppwm_u_mem__0695_/Y net554 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1174__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_3_492 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1104_ net43 VGND VPWR net248 hold49/A clknet_5_7__leaf_clk sg13g2_dfrbpq_2
XFILLER_22_1018 VPWR VGND sg13g2_decap_8
XFILLER_27_809 VPWR VGND sg13g2_decap_8
XFILLER_39_647 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1035_ net351 u_ppwm_u_ex__1035_/C u_ppwm_u_ex__1035_/A u_ppwm_u_ex__1035_/Y
+ VPWR VGND u_ppwm_u_ex__1035_/D sg13g2_nand4_1
Xu_ppwm_u_mem__1178_ net103 VGND VPWR net256 hold67/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_352 VPWR VGND sg13g2_fill_2
XFILLER_35_864 VPWR VGND sg13g2_decap_8
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_22_514 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1106__39 VPWR VGND net39 sg13g2_tiehi
Xu_ppwm_u_ex__0819_ net381 u_ppwm_u_ex__0819_/C u_ppwm/instr\[0\] u_ppwm_u_ex__0819_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_2_919 VPWR VGND sg13g2_decap_8
XFILLER_39_48 VPWR VGND sg13g2_fill_1
XFILLER_45_639 VPWR VGND sg13g2_decap_8
XFILLER_26_820 VPWR VGND sg13g2_decap_8
XFILLER_25_341 VPWR VGND sg13g2_decap_4
XFILLER_13_514 VPWR VGND sg13g2_decap_8
XFILLER_25_363 VPWR VGND sg13g2_decap_4
XFILLER_26_897 VPWR VGND sg13g2_decap_8
XFILLER_41_845 VPWR VGND sg13g2_decap_8
XFILLER_5_724 VPWR VGND sg13g2_decap_8
XFILLER_4_223 VPWR VGND sg13g2_fill_2
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_48_411 VPWR VGND sg13g2_decap_8
XFILLER_49_956 VPWR VGND sg13g2_decap_8
XFILLER_0_495 VPWR VGND sg13g2_decap_8
Xhold81 hold81/A VPWR VGND net279 sg13g2_dlygate4sd3_1
Xhold70 hold70/A VPWR VGND net268 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1101_ net587 u_ppwm_u_mem__1101_/B hold220/A VPWR VGND sg13g2_nor2_1
Xhold92 hold92/A VPWR VGND net290 sg13g2_dlygate4sd3_1
XFILLER_36_606 VPWR VGND sg13g2_decap_8
XFILLER_48_488 VPWR VGND sg13g2_decap_8
XFILLER_17_831 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1032_ net503 VPWR u_ppwm_u_mem__1032_/Y VGND net418 hold200/A sg13g2_o21ai_1
XFILLER_44_694 VPWR VGND sg13g2_decap_8
XFILLER_43_160 VPWR VGND sg13g2_fill_1
XFILLER_32_801 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_fill_1
XFILLER_31_311 VPWR VGND sg13g2_fill_2
XFILLER_32_878 VPWR VGND sg13g2_decap_8
XFILLER_12_580 VPWR VGND sg13g2_decap_8
XFILLER_8_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0604_ net615 VPWR hold248/A VGND u_ppwm_u_ex__0636_/A u_ppwm_u_ex__0600_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0816_ VGND VPWR u_ppwm_u_mem__0811_/X u_ppwm_u_mem__0813_/Y u_ppwm_u_mem__0816_/Y
+ u_ppwm_u_mem__0815_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0747_ hold114/A hold145/A net477 u_ppwm_u_mem__0747_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0678_ VPWR u_ppwm_u_mem__0678_/Y net269 VGND sg13g2_inv_1
Xfanout508 net509 net508 VPWR VGND sg13g2_buf_8
XFILLER_20_0 VPWR VGND sg13g2_fill_1
XFILLER_27_606 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1018_ net358 u_ppwm_u_ex__1018_/B u_ppwm_u_ex__1018_/Y VPWR VGND sg13g2_nor2_1
XFILLER_35_661 VPWR VGND sg13g2_decap_8
XFILLER_22_322 VPWR VGND sg13g2_fill_1
XFILLER_23_867 VPWR VGND sg13g2_decap_8
XFILLER_10_528 VPWR VGND sg13g2_decap_8
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_fill_1
XFILLER_1_226 VPWR VGND sg13g2_fill_1
XFILLER_18_617 VPWR VGND sg13g2_decap_8
XFILLER_46_937 VPWR VGND sg13g2_decap_8
XFILLER_45_436 VPWR VGND sg13g2_decap_8
XFILLER_41_642 VPWR VGND sg13g2_decap_8
XFILLER_14_867 VPWR VGND sg13g2_decap_8
XFILLER_26_694 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_5_521 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_82 VPWR VGND sg13g2_fill_1
XFILLER_5_598 VPWR VGND sg13g2_decap_8
XFILLER_49_753 VPWR VGND sg13g2_decap_8
XFILLER_48_285 VPWR VGND sg13g2_decap_8
XFILLER_37_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1015_ VGND VPWR net414 u_ppwm_u_mem__0647_/Y hold125/A u_ppwm_u_mem__1014_/Y
+ sg13g2_a21oi_1
XFILLER_44_491 VPWR VGND sg13g2_decap_8
XFILLER_16_171 VPWR VGND sg13g2_decap_4
XFILLER_32_675 VPWR VGND sg13g2_decap_8
XFILLER_20_837 VPWR VGND sg13g2_decap_8
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
Xfanout349 net351 net349 VPWR VGND sg13g2_buf_8
XFILLER_28_904 VPWR VGND sg13g2_decap_8
XFILLER_14_108 VPWR VGND sg13g2_fill_2
XFILLER_36_970 VPWR VGND sg13g2_decap_8
XFILLER_42_439 VPWR VGND sg13g2_decap_8
XFILLER_23_664 VPWR VGND sg13g2_decap_8
XFILLER_10_314 VPWR VGND sg13g2_decap_8
XFILLER_11_826 VPWR VGND sg13g2_decap_8
XFILLER_7_808 VPWR VGND sg13g2_decap_8
XFILLER_6_307 VPWR VGND sg13g2_decap_8
XFILLER_2_513 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_fill_2
XFILLER_19_904 VPWR VGND sg13g2_decap_8
XFILLER_46_734 VPWR VGND sg13g2_decap_8
XFILLER_45_233 VPWR VGND sg13g2_decap_4
XFILLER_27_970 VPWR VGND sg13g2_decap_8
XFILLER_26_491 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1211__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_14_664 VPWR VGND sg13g2_decap_8
XFILLER_9_156 VPWR VGND sg13g2_fill_2
XFILLER_42_92 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_pwm__185_ VGND VPWR u_ppwm_u_pwm__183_/A net637 u_ppwm_u_pwm__246_/D u_ppwm_u_pwm__184_/Y
+ sg13g2_a21oi_1
XFILLER_6_863 VPWR VGND sg13g2_decap_8
XFILLER_10_892 VPWR VGND sg13g2_decap_8
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_37_745 VPWR VGND sg13g2_decap_8
XFILLER_18_981 VPWR VGND sg13g2_decap_8
XFILLER_25_918 VPWR VGND sg13g2_decap_8
XFILLER_36_277 VPWR VGND sg13g2_fill_1
XFILLER_20_634 VPWR VGND sg13g2_decap_8
XFILLER_33_995 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0998_ u_ppwm_u_ex__0998_/Y net355 u_ppwm_u_ex__0998_/B2 net362 net465
+ VPWR VGND sg13g2_a22oi_1
XFILLER_47_37 VPWR VGND sg13g2_fill_1
XFILLER_28_701 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_28_778 VPWR VGND sg13g2_decap_8
XFILLER_43_748 VPWR VGND sg13g2_decap_8
XFILLER_42_236 VPWR VGND sg13g2_fill_2
XFILLER_42_225 VPWR VGND sg13g2_decap_8
XFILLER_42_214 VPWR VGND sg13g2_fill_1
XFILLER_15_428 VPWR VGND sg13g2_fill_1
XFILLER_27_299 VPWR VGND sg13g2_fill_2
XFILLER_24_962 VPWR VGND sg13g2_decap_8
XFILLER_11_623 VPWR VGND sg13g2_decap_8
XFILLER_10_111 VPWR VGND sg13g2_fill_1
XFILLER_7_605 VPWR VGND sg13g2_decap_8
XFILLER_6_126 VPWR VGND sg13g2_fill_2
XFILLER_3_800 VPWR VGND sg13g2_decap_8
XFILLER_12_84 VPWR VGND sg13g2_decap_4
XFILLER_3_877 VPWR VGND sg13g2_decap_8
XFILLER_19_701 VPWR VGND sg13g2_decap_8
XFILLER_46_531 VPWR VGND sg13g2_decap_8
XFILLER_18_222 VPWR VGND sg13g2_fill_1
XFILLER_19_778 VPWR VGND sg13g2_decap_8
XFILLER_34_737 VPWR VGND sg13g2_decap_8
XFILLER_21_409 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0921_ net371 VPWR u_ppwm_u_ex__0952_/A VGND net458 net460 sg13g2_o21ai_1
XFILLER_14_472 VPWR VGND sg13g2_fill_2
XFILLER_18_1023 VPWR VGND sg13g2_decap_4
XFILLER_30_910 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0852_ u_ppwm_u_ex__0882_/A net463 net374 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__0995_ VGND VPWR net409 u_ppwm_u_mem__0657_/Y u_ppwm_u_mem__1174_/D
+ u_ppwm_u_mem__0994_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0783_ net383 net466 u_ppwm_u_ex__0783_/X VPWR VGND sg13g2_xor2_1
XFILLER_30_987 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__237_ net193 VGND VPWR net300 hold101/A clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_6_660 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1107__174 VPWR VGND net174 sg13g2_tiehi
Xu_ppwm_u_pwm__168_ u_ppwm_u_pwm__188_/A net573 u_ppwm_u_pwm__170_/B hold206/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_25_1016 VPWR VGND sg13g2_decap_8
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_18 VPWR VGND sg13g2_decap_8
XFILLER_37_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1114__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_25_715 VPWR VGND sg13g2_decap_8
XFILLER_21_932 VPWR VGND sg13g2_decap_8
XFILLER_33_792 VPWR VGND sg13g2_decap_8
XFILLER_0_803 VPWR VGND sg13g2_decap_8
XFILLER_28_575 VPWR VGND sg13g2_decap_8
XFILLER_16_748 VPWR VGND sg13g2_decap_8
XFILLER_43_545 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1127__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_12_965 VPWR VGND sg13g2_decap_8
XFILLER_8_947 VPWR VGND sg13g2_decap_8
XFILLER_23_50 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0780_ u_ppwm_u_mem__0780_/Y net471 u_ppwm_u_mem__0780_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_48_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_674 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1120_ net44 VGND VPWR u_ppwm_u_ex__1120_/D hold299/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_829 VPWR VGND sg13g2_decap_8
XFILLER_47_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1051_ VPWR u_ppwm_u_ex__1075_/A u_ppwm_u_ex__1051_/A VGND sg13g2_inv_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_19_575 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1194_ net158 VGND VPWR u_ppwm_u_mem__1194_/D hold32/A clknet_5_13__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_34_534 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_21_206 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0904_ u_ppwm_u_ex__0903_/Y VPWR u_ppwm_u_ex__0915_/B VGND u_ppwm_u_ex__0901_/Y
+ u_ppwm_u_ex__0922_/B sg13g2_o21ai_1
XFILLER_30_784 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0835_ u_ppwm_u_ex__0835_/A u_ppwm_u_ex__0835_/B hold320/A VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_mem__0978_ net497 VPWR u_ppwm_u_mem__0978_/Y VGND net413 net224 sg13g2_o21ai_1
Xu_ppwm_u_ex__0766_ net454 net441 u_ppwm_u_ex__0767_/D VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_ex__0697_ u_ppwm_u_ex__0696_/Y VPWR u_ppwm_u_ex__0697_/Y VGND u_ppwm_u_ex__0570_/Y
+ net440 sg13g2_o21ai_1
XFILLER_38_851 VPWR VGND sg13g2_decap_8
XFILLER_25_512 VPWR VGND sg13g2_decap_8
XFILLER_25_589 VPWR VGND sg13g2_decap_8
XFILLER_40_537 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_fill_2
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_20_283 VPWR VGND sg13g2_fill_1
XFILLER_4_449 VPWR VGND sg13g2_decap_8
XFILLER_0_600 VPWR VGND sg13g2_decap_8
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_47_136 VPWR VGND sg13g2_decap_8
XFILLER_47_114 VPWR VGND sg13g2_fill_2
XFILLER_29_840 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_fill_1
XFILLER_44_876 VPWR VGND sg13g2_decap_8
XFILLER_16_545 VPWR VGND sg13g2_decap_8
XFILLER_31_548 VPWR VGND sg13g2_decap_8
XFILLER_12_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0901_ VGND VPWR net423 u_ppwm_u_mem__0704_/Y u_ppwm_u_mem__1127_/D
+ u_ppwm_u_mem__0900_/Y sg13g2_a21oi_1
XFILLER_8_744 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1123__40 VPWR VGND net40 sg13g2_tiehi
XFILLER_11_261 VPWR VGND sg13g2_decap_8
XFILLER_11_272 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0620_ net512 VPWR u_ppwm_u_ex__0620_/Y VGND net447 net473 sg13g2_o21ai_1
Xu_ppwm_u_mem__0832_ VGND VPWR u_ppwm_u_mem__0830_/Y u_ppwm_u_mem__0831_/Y u_ppwm_u_mem__0832_/Y
+ net472 sg13g2_a21oi_1
Xu_ppwm_u_mem__0763_ net467 VPWR u_ppwm_u_mem__0763_/Y VGND net470 u_ppwm_u_mem__0762_/X
+ sg13g2_o21ai_1
XFILLER_3_471 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0694_ VPWR u_ppwm_u_mem__0694_/Y net324 VGND sg13g2_inv_1
XFILLER_39_626 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1103_ net45 VGND VPWR net650 hold280/A clknet_5_5__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1034_ u_ppwm_u_ex__1033_/Y u_ppwm_u_ex__1032_/Y net359 u_ppwm_u_ex__1035_/D
+ VPWR VGND sg13g2_a21o_1
XFILLER_35_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1177_ net107 VGND VPWR net266 hold150/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_375 VPWR VGND sg13g2_decap_4
XFILLER_30_581 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0818_ u_ppwm_u_ex__0820_/C u_ppwm/instr\[0\] net381 u_ppwm_u_ex__0819_/C
+ VPWR VGND sg13g2_and3_2
Xu_ppwm_u_ex__0749_ u_ppwm_u_ex__0749_/Y net464 net444 VPWR VGND sg13g2_nand2b_1
XFILLER_39_16 VPWR VGND sg13g2_decap_8
XFILLER_45_618 VPWR VGND sg13g2_decap_8
XFILLER_41_824 VPWR VGND sg13g2_decap_8
XFILLER_26_876 VPWR VGND sg13g2_decap_8
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_25_386 VPWR VGND sg13g2_fill_1
XFILLER_5_703 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_fill_2
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_49_935 VPWR VGND sg13g2_decap_8
XFILLER_0_474 VPWR VGND sg13g2_decap_8
XFILLER_48_467 VPWR VGND sg13g2_decap_8
Xhold71 hold71/A VPWR VGND net269 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1100_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1100_/B u_ppwm_u_mem__1101_/B
+ u_ppwm_u_mem__1223_/D VPWR VGND sg13g2_nor3_1
Xhold60 hold60/A VPWR VGND net258 sg13g2_dlygate4sd3_1
Xhold82 hold82/A VPWR VGND net280 sg13g2_dlygate4sd3_1
XFILLER_17_810 VPWR VGND sg13g2_decap_8
Xhold93 hold93/A VPWR VGND net291 sg13g2_dlygate4sd3_1
XFILLER_28_180 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1031_ VGND VPWR net411 u_ppwm_u_mem__0639_/Y hold201/A u_ppwm_u_mem__1030_/Y
+ sg13g2_a21oi_1
XFILLER_44_673 VPWR VGND sg13g2_decap_8
XFILLER_16_353 VPWR VGND sg13g2_decap_4
XFILLER_16_375 VPWR VGND sg13g2_decap_8
XFILLER_17_887 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_fill_1
XFILLER_32_857 VPWR VGND sg13g2_decap_8
XFILLER_31_378 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_8_541 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0603_ VGND VPWR u_ppwm_u_ex__0605_/A net614 hold247/A u_ppwm_u_ex__0991_/A
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0815_ net467 VPWR u_ppwm_u_mem__0815_/Y VGND net470 u_ppwm_u_mem__0814_/X
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0746_ u_ppwm_u_mem__0746_/Y net395 u_ppwm_u_mem__0746_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0677_ VPWR u_ppwm_u_mem__0677_/Y net240 VGND sg13g2_inv_1
Xfanout509 net518 net509 VPWR VGND sg13g2_buf_8
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__1017_ u_ppwm_u_ex__1017_/B u_ppwm_u_ex__1027_/B u_ppwm_u_ex__1017_/A
+ u_ppwm_u_ex__1017_/Y VPWR VGND sg13g2_nand3_1
XFILLER_35_640 VPWR VGND sg13g2_decap_8
XFILLER_25_29 VPWR VGND sg13g2_decap_4
XFILLER_23_846 VPWR VGND sg13g2_decap_8
XFILLER_10_507 VPWR VGND sg13g2_decap_8
XFILLER_22_367 VPWR VGND sg13g2_fill_1
XFILLER_46_916 VPWR VGND sg13g2_decap_8
XFILLER_45_415 VPWR VGND sg13g2_decap_8
XFILLER_39_990 VPWR VGND sg13g2_decap_8
XFILLER_26_673 VPWR VGND sg13g2_decap_8
XFILLER_41_621 VPWR VGND sg13g2_decap_8
XFILLER_14_846 VPWR VGND sg13g2_decap_8
XFILLER_9_316 VPWR VGND sg13g2_fill_2
XFILLER_41_698 VPWR VGND sg13g2_decap_8
XFILLER_9_338 VPWR VGND sg13g2_decap_8
XFILLER_12_1007 VPWR VGND sg13g2_decap_8
XFILLER_5_500 VPWR VGND sg13g2_decap_8
XFILLER_5_577 VPWR VGND sg13g2_decap_8
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_48_264 VPWR VGND sg13g2_decap_8
XFILLER_37_927 VPWR VGND sg13g2_decap_8
XFILLER_45_982 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1014_ net498 VPWR u_ppwm_u_mem__1014_/Y VGND net411 hold215/A sg13g2_o21ai_1
XFILLER_44_470 VPWR VGND sg13g2_decap_8
XFILLER_16_183 VPWR VGND sg13g2_fill_1
XFILLER_17_684 VPWR VGND sg13g2_decap_8
XFILLER_20_816 VPWR VGND sg13g2_decap_8
XFILLER_32_654 VPWR VGND sg13g2_decap_8
XFILLER_31_153 VPWR VGND sg13g2_fill_1
XFILLER_31_164 VPWR VGND sg13g2_decap_4
XFILLER_9_894 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0729_ net467 u_ppwm_u_mem__0842_/A VPWR VGND sg13g2_inv_4
XFILLER_42_418 VPWR VGND sg13g2_decap_8
XFILLER_11_805 VPWR VGND sg13g2_decap_8
XFILLER_23_643 VPWR VGND sg13g2_decap_8
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1124__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_2_569 VPWR VGND sg13g2_decap_8
XFILLER_46_713 VPWR VGND sg13g2_decap_8
XFILLER_18_426 VPWR VGND sg13g2_fill_2
XFILLER_45_212 VPWR VGND sg13g2_fill_1
XFILLER_34_919 VPWR VGND sg13g2_decap_8
XFILLER_45_289 VPWR VGND sg13g2_decap_8
XFILLER_14_643 VPWR VGND sg13g2_decap_8
XFILLER_42_985 VPWR VGND sg13g2_decap_8
XFILLER_42_60 VPWR VGND sg13g2_fill_1
XFILLER_41_495 VPWR VGND sg13g2_decap_8
XFILLER_9_146 VPWR VGND sg13g2_fill_2
XFILLER_10_871 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__184_ u_ppwm_u_pwm__184_/Y net489 u_ppwm_u_pwm__187_/B VPWR VGND sg13g2_nand2_1
XFILLER_6_842 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_37_724 VPWR VGND sg13g2_decap_8
XFILLER_36_234 VPWR VGND sg13g2_decap_4
XFILLER_18_960 VPWR VGND sg13g2_decap_8
XFILLER_17_481 VPWR VGND sg13g2_decap_8
XFILLER_33_974 VPWR VGND sg13g2_decap_8
XFILLER_20_613 VPWR VGND sg13g2_decap_8
XFILLER_32_462 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__0997_ u_ppwm_u_ex__0997_/Y net444 net356 VPWR VGND sg13g2_nand2_1
XFILLER_9_691 VPWR VGND sg13g2_decap_8
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_223 VPWR VGND sg13g2_decap_4
XFILLER_28_757 VPWR VGND sg13g2_decap_8
XFILLER_43_727 VPWR VGND sg13g2_decap_8
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_27_267 VPWR VGND sg13g2_fill_1
XFILLER_42_259 VPWR VGND sg13g2_fill_2
XFILLER_24_941 VPWR VGND sg13g2_decap_8
XFILLER_11_602 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_fill_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
XFILLER_11_679 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_4
XFILLER_3_856 VPWR VGND sg13g2_decap_8
XFILLER_2_377 VPWR VGND sg13g2_decap_8
Xhold190 hold190/A VPWR VGND net558 sg13g2_dlygate4sd3_1
XFILLER_46_510 VPWR VGND sg13g2_decap_8
XFILLER_19_757 VPWR VGND sg13g2_decap_8
XFILLER_34_716 VPWR VGND sg13g2_decap_8
XFILLER_46_587 VPWR VGND sg13g2_decap_8
XFILLER_33_226 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0920_ u_ppwm_u_ex__0950_/A u_ppwm_u_ex__0950_/B u_ppwm_u_ex__0924_/A
+ VPWR VGND sg13g2_nor2_1
XFILLER_18_1002 VPWR VGND sg13g2_decap_8
XFILLER_33_237 VPWR VGND sg13g2_fill_2
XFILLER_42_782 VPWR VGND sg13g2_decap_8
XFILLER_14_462 VPWR VGND sg13g2_fill_1
XFILLER_15_985 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0851_ net373 net463 u_ppwm_u_ex__0851_/X VPWR VGND sg13g2_xor2_1
XFILLER_30_966 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0994_ net496 VPWR u_ppwm_u_mem__0994_/Y VGND net412 net292 sg13g2_o21ai_1
Xu_ppwm_u_ex__0782_ u_ppwm_u_ex__0782_/Y net466 net382 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_pwm__236_ net195 VGND VPWR net239 hold40/A clknet_5_4__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__167_ net625 net572 net549 net647 u_ppwm_u_pwm__170_/B VPWR VGND sg13g2_and4_1
Xu_ppwm_u_mem__1177__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_37_521 VPWR VGND sg13g2_decap_8
XFILLER_37_598 VPWR VGND sg13g2_decap_8
XFILLER_40_719 VPWR VGND sg13g2_decap_8
XFILLER_21_911 VPWR VGND sg13g2_decap_8
XFILLER_33_771 VPWR VGND sg13g2_decap_8
XFILLER_32_292 VPWR VGND sg13g2_fill_1
XFILLER_21_988 VPWR VGND sg13g2_decap_8
XFILLER_20_487 VPWR VGND sg13g2_decap_8
XFILLER_0_859 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_20 VPWR VGND uo_out[2] sg13g2_tielo
Xu_ppwm_u_mem__1147__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_28_554 VPWR VGND sg13g2_decap_8
XFILLER_43_524 VPWR VGND sg13g2_decap_8
XFILLER_16_727 VPWR VGND sg13g2_decap_8
XFILLER_12_944 VPWR VGND sg13g2_decap_8
XFILLER_30_229 VPWR VGND sg13g2_fill_2
XFILLER_8_926 VPWR VGND sg13g2_decap_8
XFILLER_48_1006 VPWR VGND sg13g2_decap_8
XFILLER_3_653 VPWR VGND sg13g2_decap_8
XFILLER_2_141 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_808 VPWR VGND sg13g2_decap_8
XFILLER_47_830 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1050_ net373 net448 u_ppwm_u_ex__1051_/A VPWR VGND sg13g2_xor2_1
XFILLER_19_554 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1193_ net162 VGND VPWR net231 hold200/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_46_384 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_15_782 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0903_ VGND VPWR u_ppwm_u_ex__0901_/Y u_ppwm_u_ex__0922_/B u_ppwm_u_ex__0903_/Y
+ net357 sg13g2_a21oi_1
XFILLER_14_292 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__0834_ net508 VPWR u_ppwm_u_ex__0835_/B VGND net464 net354 sg13g2_o21ai_1
XFILLER_30_763 VPWR VGND sg13g2_decap_8
XFILLER_31_1010 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0977_ VGND VPWR net413 u_ppwm_u_mem__0666_/Y hold27/A u_ppwm_u_mem__0976_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__219_ net644 u_ppwm_u_pwm__223_/B u_ppwm_u_pwm__219_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__0765_ u_ppwm_u_ex__0764_/Y VPWR u_ppwm_u_ex__0765_/Y VGND u_ppwm_u_ex__0683_/A
+ net441 sg13g2_o21ai_1
Xu_ppwm_u_ex__0696_ u_ppwm_u_ex__0696_/Y net450 u_ppwm_u_ex__1020_/B2 VPWR VGND sg13g2_nand2b_1
XFILLER_43_0 VPWR VGND sg13g2_decap_4
XFILLER_38_830 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__099_ u_ppwm_u_global_counter__099_/B net439 u_ppwm_u_global_counter__122_/D
+ VPWR VGND sg13g2_xor2_1
XFILLER_25_568 VPWR VGND sg13g2_decap_8
XFILLER_40_516 VPWR VGND sg13g2_decap_8
XFILLER_20_273 VPWR VGND sg13g2_fill_2
XFILLER_21_785 VPWR VGND sg13g2_decap_8
XFILLER_20_295 VPWR VGND sg13g2_decap_4
XFILLER_4_428 VPWR VGND sg13g2_decap_8
XFILLER_0_656 VPWR VGND sg13g2_decap_8
XFILLER_48_649 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_decap_8
XFILLER_29_896 VPWR VGND sg13g2_decap_8
XFILLER_44_855 VPWR VGND sg13g2_decap_8
XFILLER_43_398 VPWR VGND sg13g2_decap_8
XFILLER_12_741 VPWR VGND sg13g2_decap_8
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0900_ net513 VPWR u_ppwm_u_mem__0900_/Y VGND net432 net331 sg13g2_o21ai_1
XFILLER_8_723 VPWR VGND sg13g2_decap_8
XFILLER_7_211 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0831_ u_ppwm_u_mem__0831_/Y hold34/A net480 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0762_ net478 hold163/A hold53/A hold67/A hold124/A net472 u_ppwm_u_mem__0762_/X
+ VPWR VGND sg13g2_mux4_1
XFILLER_4_995 VPWR VGND sg13g2_decap_8
XFILLER_3_450 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0693_ VPWR u_ppwm_u_mem__0693_/Y net559 VGND sg13g2_inv_1
Xu_ppwm_u_pwm__247__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_39_605 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1102_ net47 VGND VPWR net685 hold315/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__1033_ u_ppwm_u_ex__1033_/Y net355 hold240/A net362 net461 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_35_822 VPWR VGND sg13g2_decap_8
XFILLER_19_395 VPWR VGND sg13g2_decap_8
XFILLER_34_321 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1176_ net111 VGND VPWR net519 hold211/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_899 VPWR VGND sg13g2_decap_8
XFILLER_22_549 VPWR VGND sg13g2_decap_8
XFILLER_30_560 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0817_ u_ppwm_u_ex__0816_/Y VPWR u_ppwm_u_ex__0820_/B VGND net370 u_ppwm_u_ex__0792_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__0748_ u_ppwm_u_ex__0753_/B VPWR u_ppwm_u_ex__0748_/Y VGND u_ppwm_u_ex__0850_/A
+ net443 sg13g2_o21ai_1
Xu_ppwm_u_ex__0679_ net457 net439 u_ppwm_u_ex__0679_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_26_855 VPWR VGND sg13g2_decap_8
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_803 VPWR VGND sg13g2_decap_8
XFILLER_13_549 VPWR VGND sg13g2_decap_8
XFILLER_9_509 VPWR VGND sg13g2_decap_8
XFILLER_21_582 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1105__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_5_759 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1120__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_20_85 VPWR VGND sg13g2_fill_1
XFILLER_49_914 VPWR VGND sg13g2_decap_8
XFILLER_0_453 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
Xhold50 hold50/A VPWR VGND net248 sg13g2_dlygate4sd3_1
XFILLER_48_446 VPWR VGND sg13g2_decap_8
Xhold72 hold72/A VPWR VGND net270 sg13g2_dlygate4sd3_1
Xhold61 hold61/A VPWR VGND net259 sg13g2_dlygate4sd3_1
XFILLER_29_83 VPWR VGND sg13g2_fill_1
Xhold83 hold83/A VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold94 hold94/A VPWR VGND net292 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1030_ net495 VPWR u_ppwm_u_mem__1030_/Y VGND net411 net538 sg13g2_o21ai_1
XFILLER_16_321 VPWR VGND sg13g2_fill_1
XFILLER_17_866 VPWR VGND sg13g2_decap_8
XFILLER_29_693 VPWR VGND sg13g2_decap_8
XFILLER_44_652 VPWR VGND sg13g2_decap_8
XFILLER_31_313 VPWR VGND sg13g2_fill_1
XFILLER_32_836 VPWR VGND sg13g2_decap_8
XFILLER_40_880 VPWR VGND sg13g2_decap_8
XFILLER_8_520 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0814_ net478 hold66/A hold94/A hold46/A hold121/A net472 u_ppwm_u_mem__0814_/X
+ VPWR VGND sg13g2_mux4_1
XFILLER_8_597 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0602_ VGND VPWR u_ppwm_u_ex__0592_/Y u_ppwm_u_ex__0601_/Y hold275/A
+ u_ppwm_u_ex__0991_/A sg13g2_a21oi_1
XFILLER_6_98 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0745_ hold203/A hold7/A net477 u_ppwm_u_mem__0746_/B VPWR VGND sg13g2_mux2_1
XFILLER_4_792 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0676_ VPWR u_ppwm_u_mem__0676_/Y net309 VGND sg13g2_inv_1
XFILLER_6_1003 VPWR VGND sg13g2_decap_8
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_39_424 VPWR VGND sg13g2_fill_1
XFILLER_39_479 VPWR VGND sg13g2_decap_8
XFILLER_19_181 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__1016_ VGND VPWR u_ppwm_u_ex__1017_/A u_ppwm_u_ex__1017_/B u_ppwm_u_ex__1018_/B
+ u_ppwm_u_ex__1027_/B sg13g2_a21oi_1
Xu_ppwm_u_mem__1228_ net101 VGND VPWR u_ppwm_u_mem__1228_/D fanout438/A clknet_5_7__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_mem__1159_ net163 VGND VPWR u_ppwm_u_mem__1159_/D hold168/A clknet_5_27__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_23_825 VPWR VGND sg13g2_decap_8
XFILLER_35_696 VPWR VGND sg13g2_decap_8
XFILLER_31_891 VPWR VGND sg13g2_decap_8
XFILLER_38_490 VPWR VGND sg13g2_fill_1
XFILLER_41_600 VPWR VGND sg13g2_decap_8
XFILLER_26_652 VPWR VGND sg13g2_decap_8
XFILLER_14_825 VPWR VGND sg13g2_decap_8
XFILLER_41_677 VPWR VGND sg13g2_decap_8
XFILLER_13_368 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__237__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_5_556 VPWR VGND sg13g2_decap_8
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_48_243 VPWR VGND sg13g2_decap_8
XFILLER_0_283 VPWR VGND sg13g2_decap_8
XFILLER_37_906 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_8
XFILLER_36_405 VPWR VGND sg13g2_fill_1
XFILLER_29_490 VPWR VGND sg13g2_fill_1
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1013_ VGND VPWR net411 u_ppwm_u_mem__0648_/Y hold216/A u_ppwm_u_mem__1012_/Y
+ sg13g2_a21oi_1
XFILLER_32_633 VPWR VGND sg13g2_decap_8
XFILLER_31_198 VPWR VGND sg13g2_decap_8
XFILLER_9_873 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0728_ VPWR fanout394/A hold305/A VGND sg13g2_inv_1
Xu_ppwm_u_mem__0659_ VPWR u_ppwm_u_mem__0659_/Y net228 VGND sg13g2_inv_1
XFILLER_39_243 VPWR VGND sg13g2_decap_8
XFILLER_28_939 VPWR VGND sg13g2_decap_8
XFILLER_43_909 VPWR VGND sg13g2_decap_8
XFILLER_23_622 VPWR VGND sg13g2_decap_8
XFILLER_23_699 VPWR VGND sg13g2_decap_8
XFILLER_10_338 VPWR VGND sg13g2_decap_4
XFILLER_7_6 VPWR VGND sg13g2_fill_1
XFILLER_2_548 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_19_939 VPWR VGND sg13g2_decap_8
XFILLER_46_769 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1170__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_45_246 VPWR VGND sg13g2_decap_8
XFILLER_14_622 VPWR VGND sg13g2_decap_8
XFILLER_42_964 VPWR VGND sg13g2_decap_8
XFILLER_13_110 VPWR VGND sg13g2_fill_1
XFILLER_41_474 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_fill_2
XFILLER_14_699 VPWR VGND sg13g2_decap_8
XFILLER_6_821 VPWR VGND sg13g2_decap_8
XFILLER_10_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__183_ VGND VPWR u_ppwm_u_pwm__187_/B hold269/A u_ppwm_u_pwm__183_/A
+ sg13g2_or2_1
XFILLER_5_342 VPWR VGND sg13g2_fill_2
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_6_898 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
XFILLER_3_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_703 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_246 VPWR VGND sg13g2_fill_2
XFILLER_33_953 VPWR VGND sg13g2_decap_8
XFILLER_32_452 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__0996_ u_ppwm_u_ex__1000_/C u_ppwm_u_ex__0996_/A net350 VPWR VGND sg13g2_nand2_1
XFILLER_9_670 VPWR VGND sg13g2_decap_8
XFILLER_20_669 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_28_736 VPWR VGND sg13g2_decap_8
XFILLER_43_706 VPWR VGND sg13g2_decap_8
XFILLER_16_909 VPWR VGND sg13g2_decap_8
XFILLER_24_920 VPWR VGND sg13g2_decap_8
XFILLER_24_997 VPWR VGND sg13g2_decap_8
XFILLER_10_124 VPWR VGND sg13g2_decap_8
XFILLER_11_658 VPWR VGND sg13g2_decap_8
XFILLER_23_496 VPWR VGND sg13g2_decap_8
XFILLER_10_146 VPWR VGND sg13g2_decap_8
XFILLER_3_835 VPWR VGND sg13g2_decap_8
Xhold180 hold180/A VPWR VGND net548 sg13g2_dlygate4sd3_1
XFILLER_2_367 VPWR VGND sg13g2_fill_1
Xhold191 hold191/A VPWR VGND net559 sg13g2_dlygate4sd3_1
XFILLER_19_736 VPWR VGND sg13g2_decap_8
XFILLER_46_566 VPWR VGND sg13g2_decap_8
XFILLER_15_964 VPWR VGND sg13g2_decap_8
XFILLER_42_761 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0850_ u_ppwm_u_ex__0850_/A u_ppwm_u_ex__1049_/B u_ppwm_u_ex__0850_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_30_945 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0993_ VGND VPWR net413 u_ppwm_u_mem__0658_/Y u_ppwm_u_mem__1173_/D
+ u_ppwm_u_mem__0992_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0781_ fanout358/A u_ppwm_u_ex__0781_/A u_ppwm_u_ex__0819_/C VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_pwm__235_ net197 VGND VPWR net212 hold13/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__166_ VGND VPWR net549 u_ppwm_u_pwm__163_/A hold205/A net572 sg13g2_a21oi_1
XFILLER_6_695 VPWR VGND sg13g2_decap_8
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_37_577 VPWR VGND sg13g2_decap_8
XFILLER_33_750 VPWR VGND sg13g2_decap_8
XFILLER_20_466 VPWR VGND sg13g2_decap_8
XFILLER_21_967 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0979_ u_ppwm_u_ex__0979_/A net363 fanout355/A VPWR VGND sg13g2_nor2_2
XFILLER_0_838 VPWR VGND sg13g2_decap_8
XFILLER_47_319 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_10 VPWR VGND uio_oe[7] sg13g2_tielo
Xheichips25_ppwm_21 VPWR VGND uo_out[3] sg13g2_tielo
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_decap_8
XFILLER_43_503 VPWR VGND sg13g2_decap_8
XFILLER_31_709 VPWR VGND sg13g2_decap_8
XFILLER_12_923 VPWR VGND sg13g2_decap_8
XFILLER_8_905 VPWR VGND sg13g2_decap_8
XFILLER_24_794 VPWR VGND sg13g2_decap_8
XFILLER_3_632 VPWR VGND sg13g2_decap_8
XFILLER_2_120 VPWR VGND sg13g2_decap_8
Xfanout490 net492 net490 VPWR VGND sg13g2_buf_8
XFILLER_19_533 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1192_ net166 VGND VPWR net569 hold170/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_886 VPWR VGND sg13g2_decap_8
XFILLER_46_363 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_9_21 VPWR VGND sg13g2_fill_2
XFILLER_15_761 VPWR VGND sg13g2_decap_8
XFILLER_34_569 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0902_ net371 net458 u_ppwm_u_ex__0922_/B VPWR VGND sg13g2_xor2_1
Xu_ppwm_u_ex__0833_ u_ppwm_u_ex__1000_/A u_ppwm_u_ex__0833_/B u_ppwm_u_ex__0833_/C
+ u_ppwm_u_ex__0835_/A VPWR VGND sg13g2_nor3_1
XFILLER_30_742 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0976_ net496 VPWR u_ppwm_u_mem__0976_/Y VGND net412 hold117/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__218_ u_ppwm_u_pwm__221_/A hold225/A u_ppwm_u_pwm__218_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_ex__0764_ u_ppwm_u_ex__0764_/Y net455 net442 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_ex__0695_ u_ppwm_u_ex__0695_/Y hold292/A hold207/A VPWR VGND sg13g2_nand2b_1
XFILLER_6_492 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__149_ net490 VPWR u_ppwm_u_pwm__149_/Y VGND net460 net389 sg13g2_o21ai_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_38_886 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__098_ net392 u_ppwm_u_global_counter__103_/C net439 u_ppwm_u_global_counter__098_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_25_547 VPWR VGND sg13g2_decap_8
XFILLER_20_230 VPWR VGND sg13g2_decap_8
XFILLER_20_241 VPWR VGND sg13g2_fill_1
XFILLER_21_764 VPWR VGND sg13g2_decap_8
XFILLER_0_635 VPWR VGND sg13g2_decap_8
XFILLER_48_628 VPWR VGND sg13g2_decap_8
XFILLER_44_834 VPWR VGND sg13g2_decap_8
XFILLER_16_503 VPWR VGND sg13g2_decap_8
XFILLER_29_875 VPWR VGND sg13g2_decap_8
XFILLER_12_720 VPWR VGND sg13g2_decap_8
XFILLER_24_591 VPWR VGND sg13g2_decap_8
XFILLER_8_702 VPWR VGND sg13g2_decap_8
XFILLER_15_1006 VPWR VGND sg13g2_decap_8
XFILLER_34_84 VPWR VGND sg13g2_fill_2
XFILLER_12_797 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0830_ u_ppwm_u_mem__0830_/Y hold15/A net480 VPWR VGND sg13g2_nand2_1
XFILLER_8_779 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0761_ VGND VPWR net472 u_ppwm_u_mem__0758_/X u_ppwm_u_mem__0761_/Y
+ net394 sg13g2_a21oi_1
Xu_ppwm_u_mem__0692_ VPWR u_ppwm_u_mem__0692_/Y net226 VGND sg13g2_inv_1
XFILLER_4_974 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1101_ net49 VGND VPWR u_ppwm_u_ex__1101_/D hold305/A clknet_5_25__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1032_ u_ppwm_u_ex__1032_/Y hold222/A net356 VPWR VGND sg13g2_nand2_1
XFILLER_47_683 VPWR VGND sg13g2_decap_8
XFILLER_35_801 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1175_ net115 VGND VPWR u_ppwm_u_mem__1175_/D hold99/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1134__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_35_878 VPWR VGND sg13g2_decap_8
XFILLER_22_528 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0816_ u_ppwm_u_ex__0816_/Y net370 u_ppwm_u_ex__0816_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__0747_ u_ppwm_u_ex__0753_/B net462 hold231/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0959_ VGND VPWR net429 u_ppwm_u_mem__0675_/Y u_ppwm_u_mem__1156_/D
+ u_ppwm_u_mem__0958_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__0678_ u_ppwm_u_ex__0678_/A u_ppwm_u_ex__0678_/B u_ppwm_u_ex__0678_/C
+ u_ppwm_u_ex__0678_/Y VPWR VGND sg13g2_nor3_1
XFILLER_29_116 VPWR VGND sg13g2_fill_1
XFILLER_38_683 VPWR VGND sg13g2_decap_8
XFILLER_26_834 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_859 VPWR VGND sg13g2_decap_8
XFILLER_13_528 VPWR VGND sg13g2_decap_8
XFILLER_21_561 VPWR VGND sg13g2_decap_8
XFILLER_5_738 VPWR VGND sg13g2_decap_8
XFILLER_0_432 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
XFILLER_48_425 VPWR VGND sg13g2_decap_8
Xhold40 hold40/A VPWR VGND net238 sg13g2_dlygate4sd3_1
Xhold73 hold73/A VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold51 hold51/A VPWR VGND net249 sg13g2_dlygate4sd3_1
Xhold62 hold62/A VPWR VGND net260 sg13g2_dlygate4sd3_1
Xhold84 hold84/A VPWR VGND net282 sg13g2_dlygate4sd3_1
XFILLER_29_672 VPWR VGND sg13g2_decap_8
Xhold95 hold95/A VPWR VGND net293 sg13g2_dlygate4sd3_1
XFILLER_44_631 VPWR VGND sg13g2_decap_8
XFILLER_16_333 VPWR VGND sg13g2_fill_2
XFILLER_17_845 VPWR VGND sg13g2_decap_8
XFILLER_32_815 VPWR VGND sg13g2_decap_8
XFILLER_12_594 VPWR VGND sg13g2_decap_8
XFILLER_8_576 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__0601_ u_ppwm_u_ex__0636_/A u_ppwm_u_ex__0601_/C net446 u_ppwm_u_ex__0601_/Y
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__0813_ VGND VPWR net396 u_ppwm_u_mem__0812_/X u_ppwm_u_mem__0813_/Y
+ net394 sg13g2_a21oi_1
Xu_ppwm_u_mem__0744_ VGND VPWR net472 u_ppwm_u_mem__0741_/X u_ppwm_u_mem__0744_/Y
+ net470 sg13g2_a21oi_1
XFILLER_4_771 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0675_ VPWR u_ppwm_u_mem__0675_/Y net541 VGND sg13g2_inv_1
XFILLER_48_992 VPWR VGND sg13g2_decap_8
XFILLER_47_480 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1227_ net156 VGND VPWR net626 hold257/A clknet_5_3__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__1015_ u_ppwm_u_ex__1027_/B net450 net376 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__1158_ net165 VGND VPWR u_ppwm_u_mem__1158_/D hold47/A clknet_5_31__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_23_804 VPWR VGND sg13g2_decap_8
XFILLER_35_675 VPWR VGND sg13g2_decap_8
XFILLER_34_174 VPWR VGND sg13g2_decap_4
XFILLER_22_336 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1089_ net638 u_ppwm_u_mem__1090_/B u_ppwm_u_mem__1091_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_31_870 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__1099__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_26_631 VPWR VGND sg13g2_decap_8
XFILLER_14_804 VPWR VGND sg13g2_decap_8
XFILLER_41_656 VPWR VGND sg13g2_decap_8
XFILLER_40_144 VPWR VGND sg13g2_fill_1
XFILLER_22_892 VPWR VGND sg13g2_decap_8
XFILLER_5_535 VPWR VGND sg13g2_decap_8
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_262 VPWR VGND sg13g2_fill_2
XFILLER_49_767 VPWR VGND sg13g2_decap_8
XFILLER_48_222 VPWR VGND sg13g2_decap_8
XFILLER_48_299 VPWR VGND sg13g2_decap_8
XFILLER_45_940 VPWR VGND sg13g2_decap_8
XFILLER_36_439 VPWR VGND sg13g2_fill_1
XFILLER_17_642 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1012_ net494 VPWR u_ppwm_u_mem__1012_/Y VGND net411 net345 sg13g2_o21ai_1
XFILLER_32_612 VPWR VGND sg13g2_decap_8
XFILLER_32_689 VPWR VGND sg13g2_decap_8
XFILLER_9_852 VPWR VGND sg13g2_decap_8
XFILLER_13_892 VPWR VGND sg13g2_decap_8
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0727_ VPWR fanout397/A net475 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0658_ VPWR u_ppwm_u_mem__0658_/Y net292 VGND sg13g2_inv_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
.ends

