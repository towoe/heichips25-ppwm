magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755750214
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 9675 38408 9717 38417
rect 9675 38368 9676 38408
rect 9716 38368 9717 38408
rect 9675 38359 9717 38368
rect 9571 38240 9629 38241
rect 9571 38200 9580 38240
rect 9620 38200 9629 38240
rect 9571 38199 9629 38200
rect 9867 38240 9909 38249
rect 9867 38200 9868 38240
rect 9908 38200 9909 38240
rect 9867 38191 9909 38200
rect 10531 38240 10589 38241
rect 10531 38200 10540 38240
rect 10580 38200 10589 38240
rect 10531 38199 10589 38200
rect 10723 38240 10781 38241
rect 10723 38200 10732 38240
rect 10772 38200 10781 38240
rect 10723 38199 10781 38200
rect 11595 38240 11637 38249
rect 11595 38200 11596 38240
rect 11636 38200 11637 38240
rect 11595 38191 11637 38200
rect 11787 38240 11829 38249
rect 11787 38200 11788 38240
rect 11828 38200 11829 38240
rect 11787 38191 11829 38200
rect 11875 38240 11933 38241
rect 11875 38200 11884 38240
rect 11924 38200 11933 38240
rect 11875 38199 11933 38200
rect 8043 38072 8085 38081
rect 8043 38032 8044 38072
rect 8084 38032 8085 38072
rect 8043 38023 8085 38032
rect 11595 38072 11637 38081
rect 11595 38032 11596 38072
rect 11636 38032 11637 38072
rect 11595 38023 11637 38032
rect 12267 38072 12309 38081
rect 12267 38032 12268 38072
rect 12308 38032 12309 38072
rect 12267 38023 12309 38032
rect 11395 37988 11453 37989
rect 11395 37948 11404 37988
rect 11444 37948 11453 37988
rect 11395 37947 11453 37948
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 9859 37652 9917 37653
rect 9859 37612 9868 37652
rect 9908 37612 9917 37652
rect 9859 37611 9917 37612
rect 7075 37400 7133 37401
rect 7075 37360 7084 37400
rect 7124 37360 7133 37400
rect 7075 37359 7133 37360
rect 7843 37400 7901 37401
rect 7843 37360 7852 37400
rect 7892 37360 7901 37400
rect 7843 37359 7901 37360
rect 8707 37400 8765 37401
rect 8707 37360 8716 37400
rect 8756 37360 8765 37400
rect 8707 37359 8765 37360
rect 10051 37400 10109 37401
rect 10051 37360 10060 37400
rect 10100 37360 10109 37400
rect 10051 37359 10109 37360
rect 11587 37400 11645 37401
rect 11587 37360 11596 37400
rect 11636 37360 11645 37400
rect 11587 37359 11645 37360
rect 12451 37400 12509 37401
rect 12451 37360 12460 37400
rect 12500 37360 12509 37400
rect 12451 37359 12509 37360
rect 12843 37400 12885 37409
rect 12843 37360 12844 37400
rect 12884 37360 12885 37400
rect 12843 37351 12885 37360
rect 13987 37400 14045 37401
rect 13987 37360 13996 37400
rect 14036 37360 14045 37400
rect 13987 37359 14045 37360
rect 16387 37400 16445 37401
rect 16387 37360 16396 37400
rect 16436 37360 16445 37400
rect 16387 37359 16445 37360
rect 7467 37316 7509 37325
rect 7467 37276 7468 37316
rect 7508 37276 7509 37316
rect 7467 37267 7509 37276
rect 6987 37232 7029 37241
rect 6987 37192 6988 37232
rect 7028 37192 7029 37232
rect 6987 37183 7029 37192
rect 9859 37232 9917 37233
rect 9859 37192 9868 37232
rect 9908 37192 9917 37232
rect 9859 37191 9917 37192
rect 10155 37232 10197 37241
rect 10155 37192 10156 37232
rect 10196 37192 10197 37232
rect 10155 37183 10197 37192
rect 10435 37232 10493 37233
rect 10435 37192 10444 37232
rect 10484 37192 10493 37232
rect 10435 37191 10493 37192
rect 14659 37232 14717 37233
rect 14659 37192 14668 37232
rect 14708 37192 14717 37232
rect 14659 37191 14717 37192
rect 15715 37232 15773 37233
rect 15715 37192 15724 37232
rect 15764 37192 15773 37232
rect 15715 37191 15773 37192
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 9955 36896 10013 36897
rect 9955 36856 9964 36896
rect 10004 36856 10013 36896
rect 9955 36855 10013 36856
rect 15523 36896 15581 36897
rect 15523 36856 15532 36896
rect 15572 36856 15581 36896
rect 15523 36855 15581 36856
rect 16491 36812 16533 36821
rect 16491 36772 16492 36812
rect 16532 36772 16533 36812
rect 16491 36763 16533 36772
rect 6499 36728 6557 36729
rect 6499 36688 6508 36728
rect 6548 36688 6557 36728
rect 6499 36687 6557 36688
rect 7179 36728 7221 36737
rect 7179 36688 7180 36728
rect 7220 36688 7221 36728
rect 7179 36679 7221 36688
rect 7555 36728 7613 36729
rect 7555 36688 7564 36728
rect 7604 36688 7613 36728
rect 7555 36687 7613 36688
rect 8419 36728 8477 36729
rect 8419 36688 8428 36728
rect 8468 36688 8477 36728
rect 8419 36687 8477 36688
rect 10627 36728 10685 36729
rect 10627 36688 10636 36728
rect 10676 36688 10685 36728
rect 10627 36687 10685 36688
rect 11107 36728 11165 36729
rect 11107 36688 11116 36728
rect 11156 36688 11165 36728
rect 11107 36687 11165 36688
rect 11211 36728 11253 36737
rect 11211 36688 11212 36728
rect 11252 36688 11253 36728
rect 11211 36679 11253 36688
rect 11403 36728 11445 36737
rect 11403 36688 11404 36728
rect 11444 36688 11445 36728
rect 11403 36679 11445 36688
rect 11779 36728 11837 36729
rect 11779 36688 11788 36728
rect 11828 36688 11837 36728
rect 11779 36687 11837 36688
rect 14851 36728 14909 36729
rect 14851 36688 14860 36728
rect 14900 36688 14909 36728
rect 14851 36687 14909 36688
rect 14955 36728 14997 36737
rect 14955 36688 14956 36728
rect 14996 36688 14997 36728
rect 14955 36679 14997 36688
rect 15331 36728 15389 36729
rect 15331 36688 15340 36728
rect 15380 36688 15389 36728
rect 15331 36687 15389 36688
rect 15435 36728 15477 36737
rect 15435 36688 15436 36728
rect 15476 36688 15477 36728
rect 15435 36679 15477 36688
rect 15627 36728 15669 36737
rect 15627 36688 15628 36728
rect 15668 36688 15669 36728
rect 15627 36679 15669 36688
rect 15811 36728 15869 36729
rect 15811 36688 15820 36728
rect 15860 36688 15869 36728
rect 15811 36687 15869 36688
rect 16683 36728 16725 36737
rect 16683 36688 16684 36728
rect 16724 36688 16725 36728
rect 16683 36679 16725 36688
rect 16779 36728 16821 36737
rect 16779 36688 16780 36728
rect 16820 36688 16821 36728
rect 16779 36679 16821 36688
rect 16875 36728 16917 36737
rect 16875 36688 16876 36728
rect 16916 36688 16917 36728
rect 16875 36679 16917 36688
rect 16971 36728 17013 36737
rect 16971 36688 16972 36728
rect 17012 36688 17013 36728
rect 16971 36679 17013 36688
rect 17539 36728 17597 36729
rect 17539 36688 17548 36728
rect 17588 36688 17597 36728
rect 17539 36687 17597 36688
rect 6603 36644 6645 36653
rect 6603 36604 6604 36644
rect 6644 36604 6645 36644
rect 6603 36595 6645 36604
rect 9579 36644 9621 36653
rect 9579 36604 9580 36644
rect 9620 36604 9621 36644
rect 9579 36595 9621 36604
rect 4299 36560 4341 36569
rect 4299 36520 4300 36560
rect 4340 36520 4341 36560
rect 4299 36511 4341 36520
rect 4683 36560 4725 36569
rect 4683 36520 4684 36560
rect 4724 36520 4725 36560
rect 4683 36511 4725 36520
rect 6987 36560 7029 36569
rect 6987 36520 6988 36560
rect 7028 36520 7029 36560
rect 6987 36511 7029 36520
rect 11403 36560 11445 36569
rect 11403 36520 11404 36560
rect 11444 36520 11445 36560
rect 11403 36511 11445 36520
rect 12651 36560 12693 36569
rect 12651 36520 12652 36560
rect 12692 36520 12693 36560
rect 12651 36511 12693 36520
rect 17163 36560 17205 36569
rect 17163 36520 17164 36560
rect 17204 36520 17205 36560
rect 17163 36511 17205 36520
rect 9955 36476 10013 36477
rect 9955 36436 9964 36476
rect 10004 36436 10013 36476
rect 9955 36435 10013 36436
rect 12451 36476 12509 36477
rect 12451 36436 12460 36476
rect 12500 36436 12509 36476
rect 12451 36435 12509 36436
rect 17643 36476 17685 36485
rect 17643 36436 17644 36476
rect 17684 36436 17685 36476
rect 17643 36427 17685 36436
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 6891 36140 6933 36149
rect 6891 36100 6892 36140
rect 6932 36100 6933 36140
rect 6891 36091 6933 36100
rect 8331 36140 8373 36149
rect 8331 36100 8332 36140
rect 8372 36100 8373 36140
rect 8331 36091 8373 36100
rect 8523 36056 8565 36065
rect 8523 36016 8524 36056
rect 8564 36016 8565 36056
rect 8523 36007 8565 36016
rect 11107 36056 11165 36057
rect 11107 36016 11116 36056
rect 11156 36016 11165 36056
rect 11107 36015 11165 36016
rect 14563 36056 14621 36057
rect 14563 36016 14572 36056
rect 14612 36016 14621 36056
rect 14563 36015 14621 36016
rect 19179 36056 19221 36065
rect 19179 36016 19180 36056
rect 19220 36016 19221 36056
rect 19179 36007 19221 36016
rect 4291 35888 4349 35889
rect 4291 35848 4300 35888
rect 4340 35848 4349 35888
rect 4291 35847 4349 35848
rect 5155 35888 5213 35889
rect 5155 35848 5164 35888
rect 5204 35848 5213 35888
rect 5155 35847 5213 35848
rect 6595 35888 6653 35889
rect 6595 35848 6604 35888
rect 6644 35848 6653 35888
rect 6595 35847 6653 35848
rect 6699 35888 6741 35897
rect 6699 35848 6700 35888
rect 6740 35848 6741 35888
rect 6699 35839 6741 35848
rect 6891 35888 6933 35897
rect 6891 35848 6892 35888
rect 6932 35848 6933 35888
rect 6891 35839 6933 35848
rect 7747 35888 7805 35889
rect 7747 35848 7756 35888
rect 7796 35848 7805 35888
rect 7747 35847 7805 35848
rect 8035 35888 8093 35889
rect 8035 35848 8044 35888
rect 8084 35848 8093 35888
rect 8035 35847 8093 35848
rect 8139 35888 8181 35897
rect 8139 35848 8140 35888
rect 8180 35848 8181 35888
rect 8139 35839 8181 35848
rect 8331 35888 8373 35897
rect 8331 35848 8332 35888
rect 8372 35848 8373 35888
rect 8331 35839 8373 35848
rect 9003 35888 9045 35897
rect 9003 35848 9004 35888
rect 9044 35848 9045 35888
rect 9003 35839 9045 35848
rect 9099 35888 9141 35897
rect 9099 35848 9100 35888
rect 9140 35848 9141 35888
rect 9099 35839 9141 35848
rect 9195 35888 9237 35897
rect 9195 35848 9196 35888
rect 9236 35848 9237 35888
rect 9195 35839 9237 35848
rect 9387 35888 9429 35897
rect 9387 35848 9388 35888
rect 9428 35848 9429 35888
rect 9387 35839 9429 35848
rect 9483 35888 9525 35897
rect 9483 35848 9484 35888
rect 9524 35848 9525 35888
rect 9483 35839 9525 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9675 35888 9717 35897
rect 9675 35848 9676 35888
rect 9716 35848 9717 35888
rect 9675 35839 9717 35848
rect 9867 35888 9909 35897
rect 9867 35848 9868 35888
rect 9908 35848 9909 35888
rect 9867 35839 9909 35848
rect 9963 35888 10005 35897
rect 9963 35848 9964 35888
rect 10004 35848 10005 35888
rect 9963 35839 10005 35848
rect 10059 35888 10101 35897
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10155 35888 10197 35897
rect 10155 35848 10156 35888
rect 10196 35848 10197 35888
rect 10155 35839 10197 35848
rect 10435 35888 10493 35889
rect 10435 35848 10444 35888
rect 10484 35848 10493 35888
rect 10435 35847 10493 35848
rect 10731 35888 10773 35897
rect 10731 35848 10732 35888
rect 10772 35848 10773 35888
rect 10731 35839 10773 35848
rect 10827 35888 10869 35897
rect 10827 35848 10828 35888
rect 10868 35848 10869 35888
rect 10827 35839 10869 35848
rect 11587 35888 11645 35889
rect 11587 35848 11596 35888
rect 11636 35848 11645 35888
rect 11587 35847 11645 35848
rect 11779 35888 11837 35889
rect 11779 35848 11788 35888
rect 11828 35848 11837 35888
rect 11779 35847 11837 35848
rect 11979 35888 12021 35897
rect 11979 35848 11980 35888
rect 12020 35848 12021 35888
rect 11979 35839 12021 35848
rect 12355 35888 12413 35889
rect 12355 35848 12364 35888
rect 12404 35848 12413 35888
rect 12355 35847 12413 35848
rect 13219 35888 13277 35889
rect 13219 35848 13228 35888
rect 13268 35848 13277 35888
rect 13219 35847 13277 35848
rect 14859 35888 14901 35897
rect 14859 35848 14860 35888
rect 14900 35848 14901 35888
rect 14859 35839 14901 35848
rect 14955 35888 14997 35897
rect 14955 35848 14956 35888
rect 14996 35848 14997 35888
rect 14955 35839 14997 35848
rect 15235 35888 15293 35889
rect 15235 35848 15244 35888
rect 15284 35848 15293 35888
rect 15235 35847 15293 35848
rect 15627 35888 15669 35897
rect 15627 35848 15628 35888
rect 15668 35848 15669 35888
rect 15627 35839 15669 35848
rect 16003 35888 16061 35889
rect 16003 35848 16012 35888
rect 16052 35848 16061 35888
rect 16003 35847 16061 35848
rect 16867 35888 16925 35889
rect 16867 35848 16876 35888
rect 16916 35848 16925 35888
rect 16867 35847 16925 35848
rect 18307 35888 18365 35889
rect 18307 35848 18316 35888
rect 18356 35848 18365 35888
rect 18307 35847 18365 35848
rect 21091 35888 21149 35889
rect 21091 35848 21100 35888
rect 21140 35848 21149 35888
rect 21091 35847 21149 35848
rect 3915 35804 3957 35813
rect 3915 35764 3916 35804
rect 3956 35764 3957 35804
rect 3915 35755 3957 35764
rect 8907 35804 8949 35813
rect 8907 35764 8908 35804
rect 8948 35764 8949 35804
rect 8907 35755 8949 35764
rect 6307 35720 6365 35721
rect 6307 35680 6316 35720
rect 6356 35680 6365 35720
rect 6307 35679 6365 35680
rect 7075 35720 7133 35721
rect 7075 35680 7084 35720
rect 7124 35680 7133 35720
rect 7075 35679 7133 35680
rect 14371 35720 14429 35721
rect 14371 35680 14380 35720
rect 14420 35680 14429 35720
rect 14371 35679 14429 35680
rect 18019 35720 18077 35721
rect 18019 35680 18028 35720
rect 18068 35680 18077 35720
rect 18019 35679 18077 35680
rect 18979 35720 19037 35721
rect 18979 35680 18988 35720
rect 19028 35680 19037 35720
rect 18979 35679 19037 35680
rect 21195 35720 21237 35729
rect 21195 35680 21196 35720
rect 21236 35680 21237 35720
rect 21195 35671 21237 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 8523 35384 8565 35393
rect 8523 35344 8524 35384
rect 8564 35344 8565 35384
rect 8523 35335 8565 35344
rect 9195 35384 9237 35393
rect 9195 35344 9196 35384
rect 9236 35344 9237 35384
rect 9195 35335 9237 35344
rect 21091 35384 21149 35385
rect 21091 35344 21100 35384
rect 21140 35344 21149 35384
rect 21091 35343 21149 35344
rect 3435 35300 3477 35309
rect 3435 35260 3436 35300
rect 3476 35260 3477 35300
rect 3435 35251 3477 35260
rect 10923 35300 10965 35309
rect 10923 35260 10924 35300
rect 10964 35260 10965 35300
rect 10923 35251 10965 35260
rect 16875 35300 16917 35309
rect 16875 35260 16876 35300
rect 16916 35260 16917 35300
rect 16875 35251 16917 35260
rect 17163 35300 17205 35309
rect 17163 35260 17164 35300
rect 17204 35260 17205 35300
rect 17163 35251 17205 35260
rect 18219 35300 18261 35309
rect 18219 35260 18220 35300
rect 18260 35260 18261 35300
rect 18219 35251 18261 35260
rect 18411 35300 18453 35309
rect 18411 35260 18412 35300
rect 18452 35260 18453 35300
rect 18411 35251 18453 35260
rect 3235 35216 3293 35217
rect 3235 35176 3244 35216
rect 3284 35176 3293 35216
rect 3235 35175 3293 35176
rect 3339 35216 3381 35225
rect 3339 35176 3340 35216
rect 3380 35176 3381 35216
rect 3339 35167 3381 35176
rect 3531 35216 3573 35225
rect 3531 35176 3532 35216
rect 3572 35176 3573 35216
rect 3531 35167 3573 35176
rect 3723 35216 3765 35225
rect 3723 35176 3724 35216
rect 3764 35176 3765 35216
rect 3723 35167 3765 35176
rect 3819 35216 3861 35225
rect 3819 35176 3820 35216
rect 3860 35176 3861 35216
rect 3819 35167 3861 35176
rect 3915 35216 3957 35225
rect 3915 35176 3916 35216
rect 3956 35176 3957 35216
rect 3915 35167 3957 35176
rect 4011 35216 4053 35225
rect 4011 35176 4012 35216
rect 4052 35176 4053 35216
rect 4011 35167 4053 35176
rect 4203 35216 4245 35225
rect 4203 35176 4204 35216
rect 4244 35176 4245 35216
rect 4203 35167 4245 35176
rect 4579 35216 4637 35217
rect 4579 35176 4588 35216
rect 4628 35176 4637 35216
rect 4579 35175 4637 35176
rect 5443 35216 5501 35217
rect 5443 35176 5452 35216
rect 5492 35176 5501 35216
rect 5443 35175 5501 35176
rect 6787 35216 6845 35217
rect 6787 35176 6796 35216
rect 6836 35176 6845 35216
rect 6787 35175 6845 35176
rect 7651 35216 7709 35217
rect 7651 35176 7660 35216
rect 7700 35176 7709 35216
rect 7651 35175 7709 35176
rect 8035 35216 8093 35217
rect 8035 35176 8044 35216
rect 8084 35176 8093 35216
rect 8035 35175 8093 35176
rect 9579 35216 9621 35225
rect 9579 35176 9580 35216
rect 9620 35176 9621 35216
rect 9579 35167 9621 35176
rect 9675 35216 9717 35225
rect 9675 35176 9676 35216
rect 9716 35176 9717 35216
rect 9675 35167 9717 35176
rect 9771 35216 9813 35225
rect 9771 35176 9772 35216
rect 9812 35176 9813 35216
rect 9771 35167 9813 35176
rect 9867 35216 9909 35225
rect 9867 35176 9868 35216
rect 9908 35176 9909 35216
rect 9867 35167 9909 35176
rect 10723 35216 10781 35217
rect 10723 35176 10732 35216
rect 10772 35176 10781 35216
rect 10723 35175 10781 35176
rect 11019 35216 11061 35225
rect 11019 35176 11020 35216
rect 11060 35176 11061 35216
rect 11019 35167 11061 35176
rect 11115 35216 11157 35225
rect 11115 35176 11116 35216
rect 11156 35176 11157 35216
rect 11115 35167 11157 35176
rect 11211 35216 11253 35225
rect 11211 35176 11212 35216
rect 11252 35176 11253 35216
rect 11211 35167 11253 35176
rect 11395 35216 11453 35217
rect 11395 35176 11404 35216
rect 11444 35176 11453 35216
rect 11395 35175 11453 35176
rect 12355 35216 12413 35217
rect 12355 35176 12364 35216
rect 12404 35176 12413 35216
rect 12355 35175 12413 35176
rect 13411 35216 13469 35217
rect 13411 35176 13420 35216
rect 13460 35176 13469 35216
rect 13411 35175 13469 35176
rect 13603 35216 13661 35217
rect 13603 35176 13612 35216
rect 13652 35176 13661 35216
rect 13603 35175 13661 35176
rect 14083 35216 14141 35217
rect 14083 35176 14092 35216
rect 14132 35176 14141 35216
rect 14083 35175 14141 35176
rect 15339 35216 15381 35225
rect 15339 35176 15340 35216
rect 15380 35176 15381 35216
rect 15339 35167 15381 35176
rect 16195 35216 16253 35217
rect 16195 35176 16204 35216
rect 16244 35176 16253 35216
rect 16195 35175 16253 35176
rect 16587 35216 16629 35225
rect 16587 35176 16588 35216
rect 16628 35176 16629 35216
rect 16587 35167 16629 35176
rect 16683 35216 16725 35225
rect 16683 35176 16684 35216
rect 16724 35176 16725 35216
rect 16683 35167 16725 35176
rect 16779 35216 16821 35225
rect 16779 35176 16780 35216
rect 16820 35176 16821 35216
rect 16779 35167 16821 35176
rect 17067 35216 17109 35225
rect 17067 35176 17068 35216
rect 17108 35176 17109 35216
rect 17067 35167 17109 35176
rect 17259 35216 17301 35225
rect 17259 35176 17260 35216
rect 17300 35176 17301 35216
rect 17259 35167 17301 35176
rect 17347 35216 17405 35217
rect 17347 35176 17356 35216
rect 17396 35176 17405 35216
rect 17347 35175 17405 35176
rect 17539 35216 17597 35217
rect 17539 35176 17548 35216
rect 17588 35176 17597 35216
rect 17539 35175 17597 35176
rect 18787 35216 18845 35217
rect 18787 35176 18796 35216
rect 18836 35176 18845 35216
rect 18787 35175 18845 35176
rect 19651 35216 19709 35217
rect 19651 35176 19660 35216
rect 19700 35176 19709 35216
rect 19651 35175 19709 35176
rect 21763 35216 21821 35217
rect 21763 35176 21772 35216
rect 21812 35176 21821 35216
rect 21763 35175 21821 35176
rect 24067 35216 24125 35217
rect 24067 35176 24076 35216
rect 24116 35176 24125 35216
rect 24067 35175 24125 35176
rect 26467 35216 26525 35217
rect 26467 35176 26476 35216
rect 26516 35176 26525 35216
rect 26467 35175 26525 35176
rect 30211 35216 30269 35217
rect 30211 35176 30220 35216
rect 30260 35176 30269 35216
rect 30211 35175 30269 35176
rect 32131 35216 32189 35217
rect 32131 35176 32140 35216
rect 32180 35176 32189 35216
rect 32131 35175 32189 35176
rect 6603 35132 6645 35141
rect 6603 35092 6604 35132
rect 6644 35092 6645 35132
rect 6603 35083 6645 35092
rect 9379 35132 9437 35133
rect 9379 35092 9388 35132
rect 9428 35092 9437 35132
rect 9379 35091 9437 35092
rect 1995 35048 2037 35057
rect 1995 35008 1996 35048
rect 2036 35008 2037 35048
rect 1995 34999 2037 35008
rect 13227 35048 13269 35057
rect 13227 35008 13228 35048
rect 13268 35008 13269 35048
rect 13227 34999 13269 35008
rect 21963 35048 22005 35057
rect 21963 35008 21964 35048
rect 22004 35008 22005 35048
rect 21963 34999 22005 35008
rect 26667 35048 26709 35057
rect 26667 35008 26668 35048
rect 26708 35008 26709 35048
rect 26667 34999 26709 35008
rect 29355 35048 29397 35057
rect 29355 35008 29356 35048
rect 29396 35008 29397 35048
rect 29355 34999 29397 35008
rect 32715 35048 32757 35057
rect 32715 35008 32716 35048
rect 32756 35008 32757 35048
rect 32715 34999 32757 35008
rect 7459 34964 7517 34965
rect 7459 34924 7468 34964
rect 7508 34924 7517 34964
rect 7459 34923 7517 34924
rect 7755 34964 7797 34973
rect 7755 34924 7756 34964
rect 7796 34924 7797 34964
rect 7755 34915 7797 34924
rect 8715 34964 8757 34973
rect 8715 34924 8716 34964
rect 8756 34924 8757 34964
rect 8715 34915 8757 34924
rect 10051 34964 10109 34965
rect 10051 34924 10060 34964
rect 10100 34924 10109 34964
rect 10051 34923 10109 34924
rect 14755 34964 14813 34965
rect 14755 34924 14764 34964
rect 14804 34924 14813 34964
rect 14755 34923 14813 34924
rect 20803 34964 20861 34965
rect 20803 34924 20812 34964
rect 20852 34924 20861 34964
rect 20803 34923 20861 34924
rect 23395 34964 23453 34965
rect 23395 34924 23404 34964
rect 23444 34924 23453 34964
rect 23395 34923 23453 34924
rect 25795 34964 25853 34965
rect 25795 34924 25804 34964
rect 25844 34924 25853 34964
rect 25795 34923 25853 34924
rect 29539 34964 29597 34965
rect 29539 34924 29548 34964
rect 29588 34924 29597 34964
rect 29539 34923 29597 34924
rect 31459 34964 31517 34965
rect 31459 34924 31468 34964
rect 31508 34924 31517 34964
rect 31459 34923 31517 34924
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 5443 34628 5501 34629
rect 5443 34588 5452 34628
rect 5492 34588 5501 34628
rect 5443 34587 5501 34588
rect 6795 34628 6837 34637
rect 6795 34588 6796 34628
rect 6836 34588 6837 34628
rect 6795 34579 6837 34588
rect 10147 34628 10205 34629
rect 10147 34588 10156 34628
rect 10196 34588 10205 34628
rect 10147 34587 10205 34588
rect 13323 34628 13365 34637
rect 13323 34588 13324 34628
rect 13364 34588 13365 34628
rect 13323 34579 13365 34588
rect 31651 34628 31709 34629
rect 31651 34588 31660 34628
rect 31700 34588 31709 34628
rect 31651 34587 31709 34588
rect 1323 34544 1365 34553
rect 1323 34504 1324 34544
rect 1364 34504 1365 34544
rect 1323 34495 1365 34504
rect 10731 34544 10773 34553
rect 10731 34504 10732 34544
rect 10772 34504 10773 34544
rect 10731 34495 10773 34504
rect 18315 34544 18357 34553
rect 18315 34504 18316 34544
rect 18356 34504 18357 34544
rect 18315 34495 18357 34504
rect 18795 34544 18837 34553
rect 18795 34504 18796 34544
rect 18836 34504 18837 34544
rect 18795 34495 18837 34504
rect 24843 34544 24885 34553
rect 24843 34504 24844 34544
rect 24884 34504 24885 34544
rect 24843 34495 24885 34504
rect 35499 34544 35541 34553
rect 35499 34504 35500 34544
rect 35540 34504 35541 34544
rect 35499 34495 35541 34504
rect 37995 34544 38037 34553
rect 37995 34504 37996 34544
rect 38036 34504 38037 34544
rect 37995 34495 38037 34504
rect 5259 34421 5301 34430
rect 1891 34376 1949 34377
rect 1891 34336 1900 34376
rect 1940 34336 1949 34376
rect 1891 34335 1949 34336
rect 2755 34376 2813 34377
rect 2755 34336 2764 34376
rect 2804 34336 2813 34376
rect 2755 34335 2813 34336
rect 4491 34376 4533 34385
rect 4491 34336 4492 34376
rect 4532 34336 4533 34376
rect 4491 34327 4533 34336
rect 4587 34376 4629 34385
rect 4587 34336 4588 34376
rect 4628 34336 4629 34376
rect 4587 34327 4629 34336
rect 4683 34376 4725 34385
rect 4683 34336 4684 34376
rect 4724 34336 4725 34376
rect 4683 34327 4725 34336
rect 4779 34376 4821 34385
rect 4779 34336 4780 34376
rect 4820 34336 4821 34376
rect 4779 34327 4821 34336
rect 5067 34376 5109 34385
rect 5067 34336 5068 34376
rect 5108 34336 5109 34376
rect 5067 34327 5109 34336
rect 5163 34376 5205 34385
rect 5163 34336 5164 34376
rect 5204 34336 5205 34376
rect 5259 34381 5260 34421
rect 5300 34381 5301 34421
rect 5259 34372 5301 34381
rect 6115 34376 6173 34377
rect 5163 34327 5205 34336
rect 6115 34336 6124 34376
rect 6164 34336 6173 34376
rect 6115 34335 6173 34336
rect 6315 34376 6357 34385
rect 6315 34336 6316 34376
rect 6356 34336 6357 34376
rect 6315 34327 6357 34336
rect 6411 34376 6453 34385
rect 6411 34336 6412 34376
rect 6452 34336 6453 34376
rect 6411 34327 6453 34336
rect 6507 34376 6549 34385
rect 6507 34336 6508 34376
rect 6548 34336 6549 34376
rect 6507 34327 6549 34336
rect 6603 34376 6645 34385
rect 6603 34336 6604 34376
rect 6644 34336 6645 34376
rect 6603 34327 6645 34336
rect 6795 34376 6837 34385
rect 6795 34336 6796 34376
rect 6836 34336 6837 34376
rect 6795 34327 6837 34336
rect 6987 34376 7029 34385
rect 6987 34336 6988 34376
rect 7028 34336 7029 34376
rect 6987 34327 7029 34336
rect 7075 34376 7133 34377
rect 7075 34336 7084 34376
rect 7124 34336 7133 34376
rect 7075 34335 7133 34336
rect 7267 34376 7325 34377
rect 7267 34336 7276 34376
rect 7316 34336 7325 34376
rect 7267 34335 7325 34336
rect 7371 34376 7413 34385
rect 7371 34336 7372 34376
rect 7412 34336 7413 34376
rect 7371 34327 7413 34336
rect 7563 34376 7605 34385
rect 7563 34336 7564 34376
rect 7604 34336 7605 34376
rect 7563 34327 7605 34336
rect 8131 34376 8189 34377
rect 8131 34336 8140 34376
rect 8180 34336 8189 34376
rect 8131 34335 8189 34336
rect 8995 34376 9053 34377
rect 8995 34336 9004 34376
rect 9044 34336 9053 34376
rect 8995 34335 9053 34336
rect 10435 34376 10493 34377
rect 10435 34336 10444 34376
rect 10484 34336 10493 34376
rect 10435 34335 10493 34336
rect 10539 34376 10581 34385
rect 10539 34336 10540 34376
rect 10580 34336 10581 34376
rect 10539 34327 10581 34336
rect 10731 34376 10773 34385
rect 10731 34336 10732 34376
rect 10772 34336 10773 34376
rect 10731 34327 10773 34336
rect 10915 34376 10973 34377
rect 10915 34336 10924 34376
rect 10964 34336 10973 34376
rect 10915 34335 10973 34336
rect 11979 34376 12021 34385
rect 11979 34336 11980 34376
rect 12020 34336 12021 34376
rect 11979 34327 12021 34336
rect 13027 34376 13085 34377
rect 13027 34336 13036 34376
rect 13076 34336 13085 34376
rect 13027 34335 13085 34336
rect 13987 34376 14045 34377
rect 13987 34336 13996 34376
rect 14036 34336 14045 34376
rect 13987 34335 14045 34336
rect 14371 34376 14429 34377
rect 14371 34336 14380 34376
rect 14420 34336 14429 34376
rect 14371 34335 14429 34336
rect 14947 34376 15005 34377
rect 14947 34336 14956 34376
rect 14996 34336 15005 34376
rect 14947 34335 15005 34336
rect 15811 34376 15869 34377
rect 15811 34336 15820 34376
rect 15860 34336 15869 34376
rect 15811 34335 15869 34336
rect 17827 34376 17885 34377
rect 17827 34336 17836 34376
rect 17876 34336 17885 34376
rect 17827 34335 17885 34336
rect 18499 34376 18557 34377
rect 18499 34336 18508 34376
rect 18548 34336 18557 34376
rect 18499 34335 18557 34336
rect 18603 34376 18645 34385
rect 18603 34336 18604 34376
rect 18644 34336 18645 34376
rect 18603 34327 18645 34336
rect 18795 34376 18837 34385
rect 18795 34336 18796 34376
rect 18836 34336 18837 34376
rect 18795 34327 18837 34336
rect 19651 34376 19709 34377
rect 19651 34336 19660 34376
rect 19700 34336 19709 34376
rect 19651 34335 19709 34336
rect 19851 34376 19893 34385
rect 19851 34336 19852 34376
rect 19892 34336 19893 34376
rect 19851 34327 19893 34336
rect 19947 34376 19989 34385
rect 19947 34336 19948 34376
rect 19988 34336 19989 34376
rect 19947 34327 19989 34336
rect 20043 34376 20085 34385
rect 20043 34336 20044 34376
rect 20084 34336 20085 34376
rect 21187 34376 21245 34377
rect 20043 34327 20085 34336
rect 20139 34355 20181 34364
rect 20139 34315 20140 34355
rect 20180 34315 20181 34355
rect 21187 34336 21196 34376
rect 21236 34336 21245 34376
rect 21187 34335 21245 34336
rect 21763 34376 21821 34377
rect 21763 34336 21772 34376
rect 21812 34336 21821 34376
rect 21763 34335 21821 34336
rect 22627 34376 22685 34377
rect 22627 34336 22636 34376
rect 22676 34336 22685 34376
rect 22627 34335 22685 34336
rect 24643 34376 24701 34377
rect 24643 34336 24652 34376
rect 24692 34336 24701 34376
rect 24643 34335 24701 34336
rect 25603 34376 25661 34377
rect 25603 34336 25612 34376
rect 25652 34336 25661 34376
rect 25603 34335 25661 34336
rect 26179 34376 26237 34377
rect 26179 34336 26188 34376
rect 26228 34336 26237 34376
rect 26179 34335 26237 34336
rect 27043 34376 27101 34377
rect 27043 34336 27052 34376
rect 27092 34336 27101 34376
rect 27043 34335 27101 34336
rect 29059 34376 29117 34377
rect 29059 34336 29068 34376
rect 29108 34336 29117 34376
rect 29059 34335 29117 34336
rect 29259 34376 29301 34385
rect 29259 34336 29260 34376
rect 29300 34336 29301 34376
rect 29259 34327 29301 34336
rect 29635 34376 29693 34377
rect 29635 34336 29644 34376
rect 29684 34336 29693 34376
rect 29635 34335 29693 34336
rect 30499 34376 30557 34377
rect 30499 34336 30508 34376
rect 30548 34336 30557 34376
rect 30499 34335 30557 34336
rect 32611 34376 32669 34377
rect 32611 34336 32620 34376
rect 32660 34336 32669 34376
rect 32611 34335 32669 34336
rect 33475 34376 33533 34377
rect 33475 34336 33484 34376
rect 33524 34336 33533 34376
rect 33475 34335 33533 34336
rect 36355 34376 36413 34377
rect 36355 34336 36364 34376
rect 36404 34336 36413 34376
rect 36355 34335 36413 34336
rect 36555 34376 36597 34385
rect 36555 34336 36556 34376
rect 36596 34336 36597 34376
rect 36555 34327 36597 34336
rect 36651 34376 36693 34385
rect 36651 34336 36652 34376
rect 36692 34336 36693 34376
rect 36651 34327 36693 34336
rect 36747 34376 36789 34385
rect 36747 34336 36748 34376
rect 36788 34336 36789 34376
rect 36747 34327 36789 34336
rect 37027 34376 37085 34377
rect 37027 34336 37036 34376
rect 37076 34336 37085 34376
rect 37027 34335 37085 34336
rect 37227 34376 37269 34385
rect 37227 34336 37228 34376
rect 37268 34336 37269 34376
rect 37227 34327 37269 34336
rect 20139 34306 20181 34315
rect 1515 34292 1557 34301
rect 1515 34252 1516 34292
rect 1556 34252 1557 34292
rect 1515 34243 1557 34252
rect 7755 34292 7797 34301
rect 7755 34252 7756 34292
rect 7796 34252 7797 34292
rect 7755 34243 7797 34252
rect 14571 34292 14613 34301
rect 14571 34252 14572 34292
rect 14612 34252 14613 34292
rect 14571 34243 14613 34252
rect 21387 34292 21429 34301
rect 21387 34252 21388 34292
rect 21428 34252 21429 34292
rect 21387 34243 21429 34252
rect 25803 34292 25845 34301
rect 25803 34252 25804 34292
rect 25844 34252 25845 34292
rect 25803 34243 25845 34252
rect 32235 34292 32277 34301
rect 32235 34252 32236 34292
rect 32276 34252 32277 34292
rect 32235 34243 32277 34252
rect 37131 34292 37173 34301
rect 37131 34252 37132 34292
rect 37172 34252 37173 34292
rect 37131 34243 37173 34252
rect 3907 34208 3965 34209
rect 3907 34168 3916 34208
rect 3956 34168 3965 34208
rect 3907 34167 3965 34168
rect 4963 34208 5021 34209
rect 4963 34168 4972 34208
rect 5012 34168 5021 34208
rect 4963 34167 5021 34168
rect 7459 34208 7517 34209
rect 7459 34168 7468 34208
rect 7508 34168 7517 34208
rect 7459 34167 7517 34168
rect 10147 34208 10205 34209
rect 10147 34168 10156 34208
rect 10196 34168 10205 34208
rect 10147 34167 10205 34168
rect 11587 34208 11645 34209
rect 11587 34168 11596 34208
rect 11636 34168 11645 34208
rect 11587 34167 11645 34168
rect 12363 34208 12405 34217
rect 12363 34168 12364 34208
rect 12404 34168 12405 34208
rect 12363 34159 12405 34168
rect 14283 34208 14325 34217
rect 14283 34168 14284 34208
rect 14324 34168 14325 34208
rect 14283 34159 14325 34168
rect 16963 34208 17021 34209
rect 16963 34168 16972 34208
rect 17012 34168 17021 34208
rect 16963 34167 17021 34168
rect 17155 34208 17213 34209
rect 17155 34168 17164 34208
rect 17204 34168 17213 34208
rect 17155 34167 17213 34168
rect 18979 34208 19037 34209
rect 18979 34168 18988 34208
rect 19028 34168 19037 34208
rect 18979 34167 19037 34168
rect 20515 34208 20573 34209
rect 20515 34168 20524 34208
rect 20564 34168 20573 34208
rect 20515 34167 20573 34168
rect 23779 34208 23837 34209
rect 23779 34168 23788 34208
rect 23828 34168 23837 34208
rect 23779 34167 23837 34168
rect 23971 34208 24029 34209
rect 23971 34168 23980 34208
rect 24020 34168 24029 34208
rect 23971 34167 24029 34168
rect 25515 34208 25557 34217
rect 25515 34168 25516 34208
rect 25556 34168 25557 34208
rect 25515 34159 25557 34168
rect 28195 34208 28253 34209
rect 28195 34168 28204 34208
rect 28244 34168 28253 34208
rect 28195 34167 28253 34168
rect 28387 34208 28445 34209
rect 28387 34168 28396 34208
rect 28436 34168 28445 34208
rect 28387 34167 28445 34168
rect 34627 34208 34685 34209
rect 34627 34168 34636 34208
rect 34676 34168 34685 34208
rect 34627 34167 34685 34168
rect 35683 34208 35741 34209
rect 35683 34168 35692 34208
rect 35732 34168 35741 34208
rect 35683 34167 35741 34168
rect 36835 34208 36893 34209
rect 36835 34168 36844 34208
rect 36884 34168 36893 34208
rect 36835 34167 36893 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 6115 33872 6173 33873
rect 6115 33832 6124 33872
rect 6164 33832 6173 33872
rect 6115 33831 6173 33832
rect 9387 33872 9429 33881
rect 9387 33832 9388 33872
rect 9428 33832 9429 33872
rect 9387 33823 9429 33832
rect 13699 33872 13757 33873
rect 13699 33832 13708 33872
rect 13748 33832 13757 33872
rect 13699 33831 13757 33832
rect 14947 33872 15005 33873
rect 14947 33832 14956 33872
rect 14996 33832 15005 33872
rect 14947 33831 15005 33832
rect 18315 33872 18357 33881
rect 18315 33832 18316 33872
rect 18356 33832 18357 33872
rect 18315 33823 18357 33832
rect 21379 33872 21437 33873
rect 21379 33832 21388 33872
rect 21428 33832 21437 33872
rect 21379 33831 21437 33832
rect 22147 33872 22205 33873
rect 22147 33832 22156 33872
rect 22196 33832 22205 33872
rect 22147 33831 22205 33832
rect 23107 33872 23165 33873
rect 23107 33832 23116 33872
rect 23156 33832 23165 33872
rect 23107 33831 23165 33832
rect 26083 33872 26141 33873
rect 26083 33832 26092 33872
rect 26132 33832 26141 33872
rect 26083 33831 26141 33832
rect 28963 33872 29021 33873
rect 28963 33832 28972 33872
rect 29012 33832 29021 33872
rect 28963 33831 29021 33832
rect 30795 33872 30837 33881
rect 30795 33832 30796 33872
rect 30836 33832 30837 33872
rect 30795 33823 30837 33832
rect 32227 33872 32285 33873
rect 32227 33832 32236 33872
rect 32276 33832 32285 33872
rect 32227 33831 32285 33832
rect 37795 33872 37853 33873
rect 37795 33832 37804 33872
rect 37844 33832 37853 33872
rect 37795 33831 37853 33832
rect 8139 33788 8181 33797
rect 8139 33748 8140 33788
rect 8180 33748 8181 33788
rect 8139 33739 8181 33748
rect 11011 33788 11069 33789
rect 11011 33748 11020 33788
rect 11060 33748 11069 33788
rect 11011 33747 11069 33748
rect 11307 33788 11349 33797
rect 11307 33748 11308 33788
rect 11348 33748 11349 33788
rect 11307 33739 11349 33748
rect 16107 33788 16149 33797
rect 16107 33748 16108 33788
rect 16148 33748 16149 33788
rect 16107 33739 16149 33748
rect 18987 33788 19029 33797
rect 18987 33748 18988 33788
rect 19028 33748 19029 33788
rect 18987 33739 19029 33748
rect 23403 33788 23445 33797
rect 23403 33748 23404 33788
rect 23444 33748 23445 33788
rect 23403 33739 23445 33748
rect 27147 33788 27189 33797
rect 27147 33748 27148 33788
rect 27188 33748 27189 33788
rect 27147 33739 27189 33748
rect 35403 33788 35445 33797
rect 35403 33748 35404 33788
rect 35444 33748 35445 33788
rect 35403 33739 35445 33748
rect 6507 33724 6549 33733
rect 1227 33704 1269 33713
rect 1227 33664 1228 33704
rect 1268 33664 1269 33704
rect 1227 33655 1269 33664
rect 1603 33704 1661 33705
rect 1603 33664 1612 33704
rect 1652 33664 1661 33704
rect 1603 33663 1661 33664
rect 2467 33704 2525 33705
rect 2467 33664 2476 33704
rect 2516 33664 2525 33704
rect 2467 33663 2525 33664
rect 3819 33704 3861 33713
rect 3819 33664 3820 33704
rect 3860 33664 3861 33704
rect 3819 33655 3861 33664
rect 4011 33704 4053 33713
rect 4011 33664 4012 33704
rect 4052 33664 4053 33704
rect 4011 33655 4053 33664
rect 4099 33704 4157 33705
rect 4099 33664 4108 33704
rect 4148 33664 4157 33704
rect 4099 33663 4157 33664
rect 4299 33704 4341 33713
rect 4299 33664 4300 33704
rect 4340 33664 4341 33704
rect 4299 33655 4341 33664
rect 4491 33704 4533 33713
rect 4491 33664 4492 33704
rect 4532 33664 4533 33704
rect 4491 33655 4533 33664
rect 4579 33704 4637 33705
rect 4579 33664 4588 33704
rect 4628 33664 4637 33704
rect 4579 33663 4637 33664
rect 4779 33704 4821 33713
rect 4779 33664 4780 33704
rect 4820 33664 4821 33704
rect 4779 33655 4821 33664
rect 4875 33704 4917 33713
rect 4875 33664 4876 33704
rect 4916 33664 4917 33704
rect 4875 33655 4917 33664
rect 4971 33704 5013 33713
rect 4971 33664 4972 33704
rect 5012 33664 5013 33704
rect 4971 33655 5013 33664
rect 5067 33704 5109 33713
rect 5067 33664 5068 33704
rect 5108 33664 5109 33704
rect 5067 33655 5109 33664
rect 5443 33704 5501 33705
rect 5443 33664 5452 33704
rect 5492 33664 5501 33704
rect 5443 33663 5501 33664
rect 6411 33704 6453 33713
rect 6411 33664 6412 33704
rect 6452 33664 6453 33704
rect 6507 33684 6508 33724
rect 6548 33684 6549 33724
rect 6507 33675 6549 33684
rect 6891 33704 6933 33713
rect 6411 33655 6453 33664
rect 6891 33664 6892 33704
rect 6932 33664 6933 33704
rect 6891 33655 6933 33664
rect 6987 33704 7029 33713
rect 6987 33664 6988 33704
rect 7028 33664 7029 33704
rect 6987 33655 7029 33664
rect 7459 33704 7517 33705
rect 7459 33664 7468 33704
rect 7508 33664 7517 33704
rect 9475 33704 9533 33705
rect 7459 33663 7517 33664
rect 7947 33690 7989 33699
rect 7947 33650 7948 33690
rect 7988 33650 7989 33690
rect 9475 33664 9484 33704
rect 9524 33664 9533 33704
rect 9475 33663 9533 33664
rect 10147 33704 10205 33705
rect 10147 33664 10156 33704
rect 10196 33664 10205 33704
rect 10147 33663 10205 33664
rect 11683 33704 11741 33705
rect 11683 33664 11692 33704
rect 11732 33664 11741 33704
rect 11683 33663 11741 33664
rect 12547 33704 12605 33705
rect 12547 33664 12556 33704
rect 12596 33664 12605 33704
rect 12547 33663 12605 33664
rect 14755 33704 14813 33705
rect 14755 33664 14764 33704
rect 14804 33664 14813 33704
rect 14755 33663 14813 33664
rect 15619 33704 15677 33705
rect 15619 33664 15628 33704
rect 15668 33664 15677 33704
rect 16771 33704 16829 33705
rect 15619 33663 15677 33664
rect 7947 33641 7989 33650
rect 16251 33662 16293 33671
rect 16771 33664 16780 33704
rect 16820 33664 16829 33704
rect 16771 33663 16829 33664
rect 17355 33704 17397 33713
rect 17355 33664 17356 33704
rect 17396 33664 17397 33704
rect 3627 33620 3669 33629
rect 3627 33580 3628 33620
rect 3668 33580 3669 33620
rect 16251 33622 16252 33662
rect 16292 33622 16293 33662
rect 17355 33655 17397 33664
rect 17739 33704 17781 33713
rect 17739 33664 17740 33704
rect 17780 33664 17781 33704
rect 17739 33655 17781 33664
rect 17835 33704 17877 33713
rect 17835 33664 17836 33704
rect 17876 33664 17877 33704
rect 17835 33655 17877 33664
rect 18211 33704 18269 33705
rect 18211 33664 18220 33704
rect 18260 33664 18269 33704
rect 18211 33663 18269 33664
rect 18507 33704 18549 33713
rect 18507 33664 18508 33704
rect 18548 33664 18549 33704
rect 18507 33655 18549 33664
rect 18699 33704 18741 33713
rect 18699 33664 18700 33704
rect 18740 33664 18741 33704
rect 18699 33655 18741 33664
rect 18787 33704 18845 33705
rect 18787 33664 18796 33704
rect 18836 33664 18845 33704
rect 18787 33663 18845 33664
rect 19363 33704 19421 33705
rect 19363 33664 19372 33704
rect 19412 33664 19421 33704
rect 19363 33663 19421 33664
rect 20227 33704 20285 33705
rect 20227 33664 20236 33704
rect 20276 33664 20285 33704
rect 20227 33663 20285 33664
rect 21579 33704 21621 33713
rect 21579 33664 21580 33704
rect 21620 33664 21621 33704
rect 21579 33655 21621 33664
rect 21675 33704 21717 33713
rect 21675 33664 21676 33704
rect 21716 33664 21717 33704
rect 21675 33655 21717 33664
rect 21771 33704 21813 33713
rect 21771 33664 21772 33704
rect 21812 33664 21813 33704
rect 21771 33655 21813 33664
rect 21867 33704 21909 33713
rect 21867 33664 21868 33704
rect 21908 33664 21909 33704
rect 21867 33655 21909 33664
rect 22059 33704 22101 33713
rect 22059 33664 22060 33704
rect 22100 33664 22101 33704
rect 22059 33655 22101 33664
rect 22251 33704 22293 33713
rect 22251 33664 22252 33704
rect 22292 33664 22293 33704
rect 22251 33655 22293 33664
rect 22339 33704 22397 33705
rect 22339 33664 22348 33704
rect 22388 33664 22397 33704
rect 22339 33663 22397 33664
rect 22915 33704 22973 33705
rect 22915 33664 22924 33704
rect 22964 33664 22973 33704
rect 22915 33663 22973 33664
rect 23019 33704 23061 33713
rect 23019 33664 23020 33704
rect 23060 33664 23061 33704
rect 23019 33655 23061 33664
rect 23211 33704 23253 33713
rect 23211 33664 23212 33704
rect 23252 33664 23253 33704
rect 23211 33655 23253 33664
rect 23779 33704 23837 33705
rect 23779 33664 23788 33704
rect 23828 33664 23837 33704
rect 23779 33663 23837 33664
rect 24643 33704 24701 33705
rect 24643 33664 24652 33704
rect 24692 33664 24701 33704
rect 24643 33663 24701 33664
rect 25995 33704 26037 33713
rect 25995 33664 25996 33704
rect 26036 33664 26037 33704
rect 25995 33655 26037 33664
rect 26187 33704 26229 33713
rect 26187 33664 26188 33704
rect 26228 33664 26229 33704
rect 26187 33655 26229 33664
rect 26275 33704 26333 33705
rect 26275 33664 26284 33704
rect 26324 33664 26333 33704
rect 26275 33663 26333 33664
rect 26755 33704 26813 33705
rect 26755 33664 26764 33704
rect 26804 33664 26813 33704
rect 26755 33663 26813 33664
rect 27051 33704 27093 33713
rect 27051 33664 27052 33704
rect 27092 33664 27093 33704
rect 27051 33655 27093 33664
rect 28099 33704 28157 33705
rect 28099 33664 28108 33704
rect 28148 33664 28157 33704
rect 28099 33663 28157 33664
rect 28203 33704 28245 33713
rect 28203 33664 28204 33704
rect 28244 33664 28245 33704
rect 28203 33655 28245 33664
rect 28771 33704 28829 33705
rect 28771 33664 28780 33704
rect 28820 33664 28829 33704
rect 28771 33663 28829 33664
rect 28875 33704 28917 33713
rect 28875 33664 28876 33704
rect 28916 33664 28917 33704
rect 28875 33655 28917 33664
rect 29067 33704 29109 33713
rect 29067 33664 29068 33704
rect 29108 33664 29109 33704
rect 29067 33655 29109 33664
rect 29923 33704 29981 33705
rect 29923 33664 29932 33704
rect 29972 33664 29981 33704
rect 29923 33663 29981 33664
rect 30883 33704 30941 33705
rect 30883 33664 30892 33704
rect 30932 33664 30941 33704
rect 30883 33663 30941 33664
rect 31083 33704 31125 33713
rect 31083 33664 31084 33704
rect 31124 33664 31125 33704
rect 31083 33655 31125 33664
rect 31179 33704 31221 33713
rect 31179 33664 31180 33704
rect 31220 33664 31221 33704
rect 31179 33655 31221 33664
rect 31275 33704 31317 33713
rect 31275 33664 31276 33704
rect 31316 33664 31317 33704
rect 31275 33655 31317 33664
rect 31371 33704 31413 33713
rect 31371 33664 31372 33704
rect 31412 33664 31413 33704
rect 31371 33655 31413 33664
rect 31563 33704 31605 33713
rect 31563 33664 31564 33704
rect 31604 33664 31605 33704
rect 31563 33655 31605 33664
rect 31659 33704 31701 33713
rect 31659 33664 31660 33704
rect 31700 33664 31701 33704
rect 31659 33655 31701 33664
rect 31755 33704 31797 33713
rect 31755 33664 31756 33704
rect 31796 33664 31797 33704
rect 31755 33655 31797 33664
rect 31851 33704 31893 33713
rect 31851 33664 31852 33704
rect 31892 33664 31893 33704
rect 31851 33655 31893 33664
rect 32035 33704 32093 33705
rect 32035 33664 32044 33704
rect 32084 33664 32093 33704
rect 32035 33663 32093 33664
rect 32139 33704 32181 33713
rect 32139 33664 32140 33704
rect 32180 33664 32181 33704
rect 32139 33655 32181 33664
rect 32331 33704 32373 33713
rect 32331 33664 32332 33704
rect 32372 33664 32373 33704
rect 32331 33655 32373 33664
rect 32523 33704 32565 33713
rect 32523 33664 32524 33704
rect 32564 33664 32565 33704
rect 32523 33655 32565 33664
rect 32899 33704 32957 33705
rect 32899 33664 32908 33704
rect 32948 33664 32957 33704
rect 32899 33663 32957 33664
rect 33763 33704 33821 33705
rect 33763 33664 33772 33704
rect 33812 33664 33821 33704
rect 33763 33663 33821 33664
rect 35203 33704 35261 33705
rect 35203 33664 35212 33704
rect 35252 33664 35261 33704
rect 35203 33663 35261 33664
rect 35779 33704 35837 33705
rect 35779 33664 35788 33704
rect 35828 33664 35837 33704
rect 35779 33663 35837 33664
rect 36643 33704 36701 33705
rect 36643 33664 36652 33704
rect 36692 33664 36701 33704
rect 36643 33663 36701 33664
rect 37987 33704 38045 33705
rect 37987 33664 37996 33704
rect 38036 33664 38045 33704
rect 37987 33663 38045 33664
rect 16251 33613 16293 33622
rect 17259 33620 17301 33629
rect 3627 33571 3669 33580
rect 17259 33580 17260 33620
rect 17300 33580 17301 33620
rect 17259 33571 17301 33580
rect 25803 33620 25845 33629
rect 25803 33580 25804 33620
rect 25844 33580 25845 33620
rect 25803 33571 25845 33580
rect 9867 33536 9909 33545
rect 9867 33496 9868 33536
rect 9908 33496 9909 33536
rect 9867 33487 9909 33496
rect 28587 33536 28629 33545
rect 28587 33496 28588 33536
rect 28628 33496 28629 33536
rect 28587 33487 28629 33496
rect 3819 33452 3861 33461
rect 3819 33412 3820 33452
rect 3860 33412 3861 33452
rect 3819 33403 3861 33412
rect 4299 33452 4341 33461
rect 4299 33412 4300 33452
rect 4340 33412 4341 33452
rect 4299 33403 4341 33412
rect 6115 33452 6173 33453
rect 6115 33412 6124 33452
rect 6164 33412 6173 33452
rect 6115 33411 6173 33412
rect 14083 33452 14141 33453
rect 14083 33412 14092 33452
rect 14132 33412 14141 33452
rect 14083 33411 14141 33412
rect 18507 33452 18549 33461
rect 18507 33412 18508 33452
rect 18548 33412 18549 33452
rect 18507 33403 18549 33412
rect 21379 33452 21437 33453
rect 21379 33412 21388 33452
rect 21428 33412 21437 33452
rect 21379 33411 21437 33412
rect 27427 33452 27485 33453
rect 27427 33412 27436 33452
rect 27476 33412 27485 33452
rect 27427 33411 27485 33412
rect 29251 33452 29309 33453
rect 29251 33412 29260 33452
rect 29300 33412 29309 33452
rect 29251 33411 29309 33412
rect 34915 33452 34973 33453
rect 34915 33412 34924 33452
rect 34964 33412 34973 33452
rect 34915 33411 34973 33412
rect 35115 33452 35157 33461
rect 35115 33412 35116 33452
rect 35156 33412 35157 33452
rect 35115 33403 35157 33412
rect 38659 33452 38717 33453
rect 38659 33412 38668 33452
rect 38708 33412 38717 33452
rect 38659 33411 38717 33412
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 2379 33116 2421 33125
rect 2379 33076 2380 33116
rect 2420 33076 2421 33116
rect 2379 33067 2421 33076
rect 3243 33116 3285 33125
rect 3243 33076 3244 33116
rect 3284 33076 3285 33116
rect 3243 33067 3285 33076
rect 5643 33116 5685 33125
rect 5643 33076 5644 33116
rect 5684 33076 5685 33116
rect 5643 33067 5685 33076
rect 6219 33116 6261 33125
rect 6219 33076 6220 33116
rect 6260 33076 6261 33116
rect 6219 33067 6261 33076
rect 19851 33116 19893 33125
rect 19851 33076 19852 33116
rect 19892 33076 19893 33116
rect 19851 33067 19893 33076
rect 23499 33116 23541 33125
rect 23499 33076 23500 33116
rect 23540 33076 23541 33116
rect 23499 33067 23541 33076
rect 24843 33116 24885 33125
rect 24843 33076 24844 33116
rect 24884 33076 24885 33116
rect 24843 33067 24885 33076
rect 31947 33116 31989 33125
rect 31947 33076 31948 33116
rect 31988 33076 31989 33116
rect 31947 33067 31989 33076
rect 34155 33116 34197 33125
rect 34155 33076 34156 33116
rect 34196 33076 34197 33116
rect 34155 33067 34197 33076
rect 34339 33116 34397 33117
rect 34339 33076 34348 33116
rect 34388 33076 34397 33116
rect 34339 33075 34397 33076
rect 35203 33116 35261 33117
rect 35203 33076 35212 33116
rect 35252 33076 35261 33116
rect 35203 33075 35261 33076
rect 1611 33032 1653 33041
rect 1611 32992 1612 33032
rect 1652 32992 1653 33032
rect 1611 32983 1653 32992
rect 6699 33032 6741 33041
rect 6699 32992 6700 33032
rect 6740 32992 6741 33032
rect 6699 32983 6741 32992
rect 10627 33032 10685 33033
rect 10627 32992 10636 33032
rect 10676 32992 10685 33032
rect 10627 32991 10685 32992
rect 19659 33032 19701 33041
rect 19659 32992 19660 33032
rect 19700 32992 19701 33032
rect 19659 32983 19701 32992
rect 21283 33032 21341 33033
rect 21283 32992 21292 33032
rect 21332 32992 21341 33032
rect 21283 32991 21341 32992
rect 33003 33032 33045 33041
rect 33003 32992 33004 33032
rect 33044 32992 33045 33032
rect 33003 32983 33045 32992
rect 33675 33032 33717 33041
rect 33675 32992 33676 33032
rect 33716 32992 33717 33032
rect 33675 32983 33717 32992
rect 36459 33032 36501 33041
rect 36459 32992 36460 33032
rect 36500 32992 36501 33032
rect 36459 32983 36501 32992
rect 9291 32948 9333 32957
rect 9291 32908 9292 32948
rect 9332 32908 9333 32948
rect 9291 32899 9333 32908
rect 12739 32948 12797 32949
rect 12739 32908 12748 32948
rect 12788 32908 12797 32948
rect 12739 32907 12797 32908
rect 16395 32948 16437 32957
rect 16395 32908 16396 32948
rect 16436 32908 16437 32948
rect 16395 32899 16437 32908
rect 19275 32948 19317 32957
rect 19275 32908 19276 32948
rect 19316 32908 19317 32948
rect 19275 32899 19317 32908
rect 28587 32948 28629 32957
rect 28587 32908 28588 32948
rect 28628 32908 28629 32948
rect 28587 32899 28629 32908
rect 33475 32948 33533 32949
rect 33475 32908 33484 32948
rect 33524 32908 33533 32948
rect 33475 32907 33533 32908
rect 2467 32864 2525 32865
rect 2467 32824 2476 32864
rect 2516 32824 2525 32864
rect 2467 32823 2525 32824
rect 2667 32864 2709 32873
rect 2667 32824 2668 32864
rect 2708 32824 2709 32864
rect 2667 32815 2709 32824
rect 2755 32864 2813 32865
rect 2755 32824 2764 32864
rect 2804 32824 2813 32864
rect 2755 32823 2813 32824
rect 2947 32864 3005 32865
rect 2947 32824 2956 32864
rect 2996 32824 3005 32864
rect 2947 32823 3005 32824
rect 3051 32864 3093 32873
rect 3051 32824 3052 32864
rect 3092 32824 3093 32864
rect 3051 32815 3093 32824
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3523 32864 3581 32865
rect 3523 32824 3532 32864
rect 3572 32824 3581 32864
rect 3523 32823 3581 32824
rect 3715 32864 3773 32865
rect 3715 32824 3724 32864
rect 3764 32824 3773 32864
rect 3715 32823 3773 32824
rect 3907 32864 3965 32865
rect 3907 32824 3916 32864
rect 3956 32824 3965 32864
rect 3907 32823 3965 32824
rect 4771 32864 4829 32865
rect 4771 32824 4780 32864
rect 4820 32824 4829 32864
rect 4771 32823 4829 32824
rect 5643 32864 5685 32873
rect 5643 32824 5644 32864
rect 5684 32824 5685 32864
rect 5643 32815 5685 32824
rect 5835 32864 5877 32873
rect 5835 32824 5836 32864
rect 5876 32824 5877 32864
rect 5835 32815 5877 32824
rect 5923 32864 5981 32865
rect 5923 32824 5932 32864
rect 5972 32824 5981 32864
rect 5923 32823 5981 32824
rect 6115 32864 6173 32865
rect 6115 32824 6124 32864
rect 6164 32824 6173 32864
rect 6115 32823 6173 32824
rect 7267 32864 7325 32865
rect 7267 32824 7276 32864
rect 7316 32824 7325 32864
rect 7267 32823 7325 32824
rect 8131 32864 8189 32865
rect 8131 32824 8140 32864
rect 8180 32824 8189 32864
rect 8131 32823 8189 32824
rect 9955 32864 10013 32865
rect 9955 32824 9964 32864
rect 10004 32824 10013 32864
rect 9955 32823 10013 32824
rect 10251 32864 10293 32873
rect 10251 32824 10252 32864
rect 10292 32824 10293 32864
rect 10251 32815 10293 32824
rect 10347 32864 10389 32873
rect 10347 32824 10348 32864
rect 10388 32824 10389 32864
rect 10347 32815 10389 32824
rect 10819 32864 10877 32865
rect 10819 32824 10828 32864
rect 10868 32824 10877 32864
rect 10819 32823 10877 32824
rect 10923 32864 10965 32873
rect 10923 32824 10924 32864
rect 10964 32824 10965 32864
rect 10923 32815 10965 32824
rect 11115 32864 11157 32873
rect 11115 32824 11116 32864
rect 11156 32824 11157 32864
rect 11115 32815 11157 32824
rect 11403 32864 11445 32873
rect 11403 32824 11404 32864
rect 11444 32824 11445 32864
rect 11403 32815 11445 32824
rect 11499 32864 11541 32873
rect 11499 32824 11500 32864
rect 11540 32824 11541 32864
rect 11499 32815 11541 32824
rect 11595 32864 11637 32873
rect 11595 32824 11596 32864
rect 11636 32824 11637 32864
rect 11595 32815 11637 32824
rect 11691 32864 11733 32873
rect 11691 32824 11692 32864
rect 11732 32824 11733 32864
rect 11691 32815 11733 32824
rect 11883 32864 11925 32873
rect 11883 32824 11884 32864
rect 11924 32824 11925 32864
rect 11883 32815 11925 32824
rect 11979 32864 12021 32873
rect 11979 32824 11980 32864
rect 12020 32824 12021 32864
rect 11979 32815 12021 32824
rect 12075 32864 12117 32873
rect 12075 32824 12076 32864
rect 12116 32824 12117 32864
rect 12075 32815 12117 32824
rect 12171 32864 12213 32873
rect 12171 32824 12172 32864
rect 12212 32824 12213 32864
rect 12171 32815 12213 32824
rect 12547 32864 12605 32865
rect 12547 32824 12556 32864
rect 12596 32824 12605 32864
rect 12547 32823 12605 32824
rect 13795 32864 13853 32865
rect 13795 32824 13804 32864
rect 13844 32824 13853 32864
rect 13795 32823 13853 32824
rect 13995 32864 14037 32873
rect 13995 32824 13996 32864
rect 14036 32824 14037 32864
rect 13995 32815 14037 32824
rect 14371 32864 14429 32865
rect 14371 32824 14380 32864
rect 14420 32824 14429 32864
rect 14371 32823 14429 32824
rect 15235 32864 15293 32865
rect 15235 32824 15244 32864
rect 15284 32824 15293 32864
rect 15235 32823 15293 32824
rect 16683 32864 16725 32873
rect 16683 32824 16684 32864
rect 16724 32824 16725 32864
rect 16683 32815 16725 32824
rect 16779 32864 16821 32873
rect 16779 32824 16780 32864
rect 16820 32824 16821 32864
rect 16779 32815 16821 32824
rect 16875 32864 16917 32873
rect 16875 32824 16876 32864
rect 16916 32824 16917 32864
rect 16875 32815 16917 32824
rect 17547 32864 17589 32873
rect 17547 32824 17548 32864
rect 17588 32824 17589 32864
rect 17547 32815 17589 32824
rect 18403 32864 18461 32865
rect 18403 32824 18412 32864
rect 18452 32824 18461 32864
rect 18403 32823 18461 32824
rect 18595 32864 18653 32865
rect 18595 32824 18604 32864
rect 18644 32824 18653 32864
rect 18595 32823 18653 32824
rect 19939 32864 19997 32865
rect 19939 32824 19948 32864
rect 19988 32824 19997 32864
rect 19939 32823 19997 32824
rect 21579 32864 21621 32873
rect 21579 32824 21580 32864
rect 21620 32824 21621 32864
rect 21579 32815 21621 32824
rect 21675 32864 21717 32873
rect 21675 32824 21676 32864
rect 21716 32824 21717 32864
rect 21675 32815 21717 32824
rect 21955 32864 22013 32865
rect 21955 32824 21964 32864
rect 22004 32824 22013 32864
rect 21955 32823 22013 32824
rect 23587 32864 23645 32865
rect 23587 32824 23596 32864
rect 23636 32824 23645 32864
rect 23587 32823 23645 32824
rect 23787 32864 23829 32873
rect 23787 32824 23788 32864
rect 23828 32824 23829 32864
rect 23787 32815 23829 32824
rect 23883 32864 23925 32873
rect 23883 32824 23884 32864
rect 23924 32824 23925 32864
rect 23883 32815 23925 32824
rect 23979 32864 24021 32873
rect 23979 32824 23980 32864
rect 24020 32824 24021 32864
rect 23979 32815 24021 32824
rect 24075 32864 24117 32873
rect 24075 32824 24076 32864
rect 24116 32824 24117 32864
rect 24075 32815 24117 32824
rect 24355 32864 24413 32865
rect 24355 32824 24364 32864
rect 24404 32824 24413 32864
rect 24355 32823 24413 32824
rect 25315 32864 25373 32865
rect 25315 32824 25324 32864
rect 25364 32824 25373 32864
rect 25315 32823 25373 32824
rect 25707 32864 25749 32873
rect 25707 32824 25708 32864
rect 25748 32824 25749 32864
rect 25707 32815 25749 32824
rect 25803 32864 25845 32873
rect 25803 32824 25804 32864
rect 25844 32824 25845 32864
rect 25803 32815 25845 32824
rect 25899 32864 25941 32873
rect 25899 32824 25900 32864
rect 25940 32824 25941 32864
rect 25899 32815 25941 32824
rect 25995 32864 26037 32873
rect 25995 32824 25996 32864
rect 26036 32824 26037 32864
rect 25995 32815 26037 32824
rect 26563 32864 26621 32865
rect 26563 32824 26572 32864
rect 26612 32824 26621 32864
rect 26563 32823 26621 32824
rect 27427 32864 27485 32865
rect 27427 32824 27436 32864
rect 27476 32824 27485 32864
rect 27427 32823 27485 32824
rect 28779 32864 28821 32873
rect 28779 32824 28780 32864
rect 28820 32824 28821 32864
rect 28779 32815 28821 32824
rect 29155 32864 29213 32865
rect 29155 32824 29164 32864
rect 29204 32824 29213 32864
rect 29155 32823 29213 32824
rect 30019 32864 30077 32865
rect 30019 32824 30028 32864
rect 30068 32824 30077 32864
rect 30019 32823 30077 32824
rect 31651 32864 31709 32865
rect 31651 32824 31660 32864
rect 31700 32824 31709 32864
rect 31651 32823 31709 32824
rect 31755 32864 31797 32873
rect 31755 32824 31756 32864
rect 31796 32824 31797 32864
rect 31755 32815 31797 32824
rect 31947 32864 31989 32873
rect 31947 32824 31948 32864
rect 31988 32824 31989 32864
rect 31947 32815 31989 32824
rect 32131 32864 32189 32865
rect 32131 32824 32140 32864
rect 32180 32824 32189 32864
rect 32131 32823 32189 32824
rect 33859 32864 33917 32865
rect 33859 32824 33868 32864
rect 33908 32824 33917 32864
rect 33859 32823 33917 32824
rect 33963 32864 34005 32873
rect 33963 32824 33964 32864
rect 34004 32824 34005 32864
rect 33963 32815 34005 32824
rect 34155 32864 34197 32873
rect 34155 32824 34156 32864
rect 34196 32824 34197 32864
rect 34155 32815 34197 32824
rect 35011 32864 35069 32865
rect 35011 32824 35020 32864
rect 35060 32824 35069 32864
rect 35011 32823 35069 32824
rect 35875 32864 35933 32865
rect 35875 32824 35884 32864
rect 35924 32824 35933 32864
rect 35875 32823 35933 32824
rect 36163 32864 36221 32865
rect 36163 32824 36172 32864
rect 36212 32824 36221 32864
rect 36163 32823 36221 32824
rect 36267 32864 36309 32873
rect 36267 32824 36268 32864
rect 36308 32824 36309 32864
rect 36267 32815 36309 32824
rect 36459 32864 36501 32873
rect 36459 32824 36460 32864
rect 36500 32824 36501 32864
rect 36459 32815 36501 32824
rect 36643 32864 36701 32865
rect 36643 32824 36652 32864
rect 36692 32824 36701 32864
rect 36643 32823 36701 32824
rect 37891 32864 37949 32865
rect 37891 32824 37900 32864
rect 37940 32824 37949 32864
rect 37891 32823 37949 32824
rect 38755 32864 38813 32865
rect 38755 32824 38764 32864
rect 38804 32824 38813 32864
rect 38755 32823 38813 32824
rect 4587 32780 4629 32789
rect 4587 32740 4588 32780
rect 4628 32740 4629 32780
rect 4587 32731 4629 32740
rect 5451 32780 5493 32789
rect 5451 32740 5452 32780
rect 5492 32740 5493 32780
rect 5451 32731 5493 32740
rect 6891 32780 6933 32789
rect 6891 32740 6892 32780
rect 6932 32740 6933 32780
rect 6891 32731 6933 32740
rect 11019 32780 11061 32789
rect 11019 32740 11020 32780
rect 11060 32740 11061 32780
rect 11019 32731 11061 32740
rect 26187 32780 26229 32789
rect 26187 32740 26188 32780
rect 26228 32740 26229 32780
rect 26187 32731 26229 32740
rect 37323 32780 37365 32789
rect 37323 32740 37324 32780
rect 37364 32740 37365 32780
rect 37323 32731 37365 32740
rect 37515 32780 37557 32789
rect 37515 32740 37516 32780
rect 37556 32740 37557 32780
rect 37515 32731 37557 32740
rect 12459 32696 12501 32705
rect 12459 32656 12460 32696
rect 12500 32656 12501 32696
rect 12459 32647 12501 32656
rect 13123 32696 13181 32697
rect 13123 32656 13132 32696
rect 13172 32656 13181 32696
rect 13123 32655 13181 32656
rect 16579 32696 16637 32697
rect 16579 32656 16588 32696
rect 16628 32656 16637 32696
rect 16579 32655 16637 32656
rect 31171 32696 31229 32697
rect 31171 32656 31180 32696
rect 31220 32656 31229 32696
rect 31171 32655 31229 32656
rect 32803 32696 32861 32697
rect 32803 32656 32812 32696
rect 32852 32656 32861 32696
rect 32803 32655 32861 32656
rect 39907 32696 39965 32697
rect 39907 32656 39916 32696
rect 39956 32656 39965 32696
rect 39907 32655 39965 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 3715 32360 3773 32361
rect 3715 32320 3724 32360
rect 3764 32320 3773 32360
rect 3715 32319 3773 32320
rect 5259 32360 5301 32369
rect 5259 32320 5260 32360
rect 5300 32320 5301 32360
rect 5259 32311 5301 32320
rect 6411 32360 6453 32369
rect 6411 32320 6412 32360
rect 6452 32320 6453 32360
rect 6411 32311 6453 32320
rect 6795 32360 6837 32369
rect 6795 32320 6796 32360
rect 6836 32320 6837 32360
rect 6795 32311 6837 32320
rect 7267 32360 7325 32361
rect 7267 32320 7276 32360
rect 7316 32320 7325 32360
rect 7267 32319 7325 32320
rect 13603 32360 13661 32361
rect 13603 32320 13612 32360
rect 13652 32320 13661 32360
rect 13603 32319 13661 32320
rect 18115 32360 18173 32361
rect 18115 32320 18124 32360
rect 18164 32320 18173 32360
rect 18115 32319 18173 32320
rect 22155 32360 22197 32369
rect 22155 32320 22156 32360
rect 22196 32320 22197 32360
rect 22155 32311 22197 32320
rect 26371 32360 26429 32361
rect 26371 32320 26380 32360
rect 26420 32320 26429 32360
rect 26371 32319 26429 32320
rect 31939 32360 31997 32361
rect 31939 32320 31948 32360
rect 31988 32320 31997 32360
rect 31939 32319 31997 32320
rect 32427 32360 32469 32369
rect 32427 32320 32428 32360
rect 32468 32320 32469 32360
rect 32427 32311 32469 32320
rect 33195 32360 33237 32369
rect 33195 32320 33196 32360
rect 33236 32320 33237 32360
rect 33195 32311 33237 32320
rect 35787 32360 35829 32369
rect 35787 32320 35788 32360
rect 35828 32320 35829 32360
rect 35787 32311 35829 32320
rect 36259 32360 36317 32361
rect 36259 32320 36268 32360
rect 36308 32320 36317 32360
rect 36259 32319 36317 32320
rect 1131 32276 1173 32285
rect 1131 32236 1132 32276
rect 1172 32236 1173 32276
rect 1131 32227 1173 32236
rect 31467 32276 31509 32285
rect 31467 32236 31468 32276
rect 31508 32236 31509 32276
rect 31467 32227 31509 32236
rect 1507 32192 1565 32193
rect 1507 32152 1516 32192
rect 1556 32152 1565 32192
rect 1507 32151 1565 32152
rect 2371 32192 2429 32193
rect 2371 32152 2380 32192
rect 2420 32152 2429 32192
rect 2371 32151 2429 32152
rect 4387 32192 4445 32193
rect 4387 32152 4396 32192
rect 4436 32152 4445 32192
rect 4387 32151 4445 32152
rect 5731 32192 5789 32193
rect 5731 32152 5740 32192
rect 5780 32152 5789 32192
rect 5731 32151 5789 32152
rect 6115 32192 6173 32193
rect 6115 32152 6124 32192
rect 6164 32152 6173 32192
rect 6115 32151 6173 32152
rect 6307 32192 6365 32193
rect 6307 32152 6316 32192
rect 6356 32152 6365 32192
rect 6307 32151 6365 32152
rect 6691 32192 6749 32193
rect 6691 32152 6700 32192
rect 6740 32152 6749 32192
rect 6691 32151 6749 32152
rect 7179 32192 7221 32201
rect 7179 32152 7180 32192
rect 7220 32152 7221 32192
rect 7179 32143 7221 32152
rect 7371 32192 7413 32201
rect 7371 32152 7372 32192
rect 7412 32152 7413 32192
rect 7371 32143 7413 32152
rect 7459 32192 7517 32193
rect 7459 32152 7468 32192
rect 7508 32152 7517 32192
rect 7459 32151 7517 32152
rect 7947 32192 7989 32201
rect 7947 32152 7948 32192
rect 7988 32152 7989 32192
rect 7947 32143 7989 32152
rect 8043 32192 8085 32201
rect 8043 32152 8044 32192
rect 8084 32152 8085 32192
rect 8043 32143 8085 32152
rect 8139 32192 8181 32201
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8235 32192 8277 32201
rect 8235 32152 8236 32192
rect 8276 32152 8277 32192
rect 8235 32143 8277 32152
rect 9579 32192 9621 32201
rect 9579 32152 9580 32192
rect 9620 32152 9621 32192
rect 9579 32143 9621 32152
rect 10243 32192 10301 32193
rect 10243 32152 10252 32192
rect 10292 32152 10301 32192
rect 10243 32151 10301 32152
rect 11107 32192 11165 32193
rect 11107 32152 11116 32192
rect 11156 32152 11165 32192
rect 11107 32151 11165 32152
rect 11971 32192 12029 32193
rect 11971 32152 11980 32192
rect 12020 32152 12029 32192
rect 11971 32151 12029 32152
rect 12171 32192 12213 32201
rect 12171 32152 12172 32192
rect 12212 32152 12213 32192
rect 12171 32143 12213 32152
rect 12355 32192 12413 32193
rect 12355 32152 12364 32192
rect 12404 32152 12413 32192
rect 12355 32151 12413 32152
rect 12739 32192 12797 32193
rect 12739 32152 12748 32192
rect 12788 32152 12797 32192
rect 12739 32151 12797 32152
rect 13035 32192 13077 32201
rect 13035 32152 13036 32192
rect 13076 32152 13077 32192
rect 13035 32143 13077 32152
rect 13131 32192 13173 32201
rect 13131 32152 13132 32192
rect 13172 32152 13173 32192
rect 13131 32143 13173 32152
rect 14275 32192 14333 32193
rect 14275 32152 14284 32192
rect 14324 32152 14333 32192
rect 14275 32151 14333 32152
rect 14475 32192 14517 32201
rect 14475 32152 14476 32192
rect 14516 32152 14517 32192
rect 14475 32143 14517 32152
rect 14571 32192 14613 32201
rect 14571 32152 14572 32192
rect 14612 32152 14613 32192
rect 14571 32143 14613 32152
rect 14667 32192 14709 32201
rect 14667 32152 14668 32192
rect 14708 32152 14709 32192
rect 14667 32143 14709 32152
rect 14763 32192 14805 32201
rect 14763 32152 14764 32192
rect 14804 32152 14805 32192
rect 14763 32143 14805 32152
rect 16003 32192 16061 32193
rect 16003 32152 16012 32192
rect 16052 32152 16061 32192
rect 16003 32151 16061 32152
rect 16387 32192 16445 32193
rect 16387 32152 16396 32192
rect 16436 32152 16445 32192
rect 16387 32151 16445 32152
rect 16579 32192 16637 32193
rect 16579 32152 16588 32192
rect 16628 32152 16637 32192
rect 16579 32151 16637 32152
rect 17451 32192 17493 32201
rect 17451 32152 17452 32192
rect 17492 32152 17493 32192
rect 17451 32143 17493 32152
rect 17835 32192 17877 32201
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 17931 32192 17973 32201
rect 17931 32152 17932 32192
rect 17972 32152 17973 32192
rect 17931 32143 17973 32152
rect 18027 32192 18069 32201
rect 18027 32152 18028 32192
rect 18068 32152 18069 32192
rect 18027 32143 18069 32152
rect 18403 32192 18461 32193
rect 18403 32152 18412 32192
rect 18452 32152 18461 32192
rect 18403 32151 18461 32152
rect 19651 32192 19709 32193
rect 19651 32152 19660 32192
rect 19700 32152 19709 32192
rect 19651 32151 19709 32152
rect 20515 32192 20573 32193
rect 20515 32152 20524 32192
rect 20564 32152 20573 32192
rect 20515 32151 20573 32152
rect 20907 32192 20949 32201
rect 20907 32152 20908 32192
rect 20948 32152 20949 32192
rect 20907 32143 20949 32152
rect 22539 32192 22581 32201
rect 22539 32152 22540 32192
rect 22580 32152 22581 32192
rect 22539 32143 22581 32152
rect 23211 32192 23253 32201
rect 23211 32152 23212 32192
rect 23252 32152 23253 32192
rect 23211 32143 23253 32152
rect 25603 32192 25661 32193
rect 25603 32152 25612 32192
rect 25652 32152 25661 32192
rect 25603 32151 25661 32152
rect 25891 32192 25949 32193
rect 25891 32152 25900 32192
rect 25940 32152 25949 32192
rect 25891 32151 25949 32152
rect 25995 32192 26037 32201
rect 25995 32152 25996 32192
rect 26036 32152 26037 32192
rect 25995 32143 26037 32152
rect 26187 32192 26229 32201
rect 26187 32152 26188 32192
rect 26228 32152 26229 32192
rect 26187 32143 26229 32152
rect 27043 32192 27101 32193
rect 27043 32152 27052 32192
rect 27092 32152 27101 32192
rect 27043 32151 27101 32152
rect 27243 32192 27285 32201
rect 27243 32152 27244 32192
rect 27284 32152 27285 32192
rect 27243 32143 27285 32152
rect 27339 32192 27381 32201
rect 27339 32152 27340 32192
rect 27380 32152 27381 32192
rect 27339 32143 27381 32152
rect 27435 32192 27477 32201
rect 27435 32152 27436 32192
rect 27476 32152 27477 32192
rect 27435 32143 27477 32152
rect 27531 32192 27573 32201
rect 27531 32152 27532 32192
rect 27572 32152 27573 32192
rect 27531 32143 27573 32152
rect 28771 32192 28829 32193
rect 28771 32152 28780 32192
rect 28820 32152 28829 32192
rect 28771 32151 28829 32152
rect 28971 32192 29013 32201
rect 28971 32152 28972 32192
rect 29012 32152 29013 32192
rect 28971 32143 29013 32152
rect 29635 32192 29693 32193
rect 29635 32152 29644 32192
rect 29684 32152 29693 32192
rect 29635 32151 29693 32152
rect 30027 32192 30069 32201
rect 30027 32152 30028 32192
rect 30068 32152 30069 32192
rect 30027 32143 30069 32152
rect 30123 32192 30165 32201
rect 30123 32152 30124 32192
rect 30164 32152 30165 32192
rect 30123 32143 30165 32152
rect 30219 32192 30261 32201
rect 30219 32152 30220 32192
rect 30260 32152 30261 32192
rect 30219 32143 30261 32152
rect 30315 32192 30357 32201
rect 30315 32152 30316 32192
rect 30356 32152 30357 32192
rect 30315 32143 30357 32152
rect 30507 32192 30549 32201
rect 30507 32152 30508 32192
rect 30548 32152 30549 32192
rect 30507 32143 30549 32152
rect 30699 32192 30741 32201
rect 30699 32152 30700 32192
rect 30740 32152 30741 32192
rect 30699 32143 30741 32152
rect 30787 32192 30845 32193
rect 30787 32152 30796 32192
rect 30836 32152 30845 32192
rect 30787 32151 30845 32152
rect 31075 32192 31133 32193
rect 31075 32152 31084 32192
rect 31124 32152 31133 32192
rect 31075 32151 31133 32152
rect 31371 32192 31413 32201
rect 31371 32152 31372 32192
rect 31412 32152 31413 32192
rect 31371 32143 31413 32152
rect 32043 32192 32085 32201
rect 32043 32152 32044 32192
rect 32084 32152 32085 32192
rect 32043 32143 32085 32152
rect 32139 32192 32181 32201
rect 32139 32152 32140 32192
rect 32180 32152 32181 32192
rect 32139 32143 32181 32152
rect 32235 32192 32277 32201
rect 32235 32152 32236 32192
rect 32276 32152 32277 32192
rect 32235 32143 32277 32152
rect 32811 32192 32853 32201
rect 32811 32152 32812 32192
rect 32852 32152 32853 32192
rect 32811 32143 32853 32152
rect 32899 32192 32957 32193
rect 32899 32152 32908 32192
rect 32948 32152 32957 32192
rect 32899 32151 32957 32152
rect 33091 32192 33149 32193
rect 33091 32152 33100 32192
rect 33140 32152 33149 32192
rect 33091 32151 33149 32152
rect 33763 32192 33821 32193
rect 33763 32152 33772 32192
rect 33812 32152 33821 32192
rect 33763 32151 33821 32152
rect 34531 32192 34589 32193
rect 34531 32152 34540 32192
rect 34580 32152 34589 32192
rect 34531 32151 34589 32152
rect 35683 32192 35741 32193
rect 35683 32152 35692 32192
rect 35732 32152 35741 32192
rect 35683 32151 35741 32152
rect 35979 32192 36021 32201
rect 35979 32152 35980 32192
rect 36020 32152 36021 32192
rect 35979 32143 36021 32152
rect 36075 32192 36117 32201
rect 36075 32152 36076 32192
rect 36116 32152 36117 32192
rect 36075 32143 36117 32152
rect 36171 32192 36213 32201
rect 36171 32152 36172 32192
rect 36212 32152 36213 32192
rect 36171 32143 36213 32152
rect 36459 32192 36501 32201
rect 36459 32152 36460 32192
rect 36500 32152 36501 32192
rect 36459 32143 36501 32152
rect 36555 32192 36597 32201
rect 36555 32152 36556 32192
rect 36596 32152 36597 32192
rect 36555 32143 36597 32152
rect 36651 32192 36693 32201
rect 36651 32152 36652 32192
rect 36692 32152 36693 32192
rect 36651 32143 36693 32152
rect 36747 32192 36789 32201
rect 36747 32152 36748 32192
rect 36788 32152 36789 32192
rect 36747 32143 36789 32152
rect 36939 32192 36981 32201
rect 36939 32152 36940 32192
rect 36980 32152 36981 32192
rect 36939 32143 36981 32152
rect 37603 32192 37661 32193
rect 37603 32152 37612 32192
rect 37652 32152 37661 32192
rect 37603 32151 37661 32152
rect 38083 32192 38141 32193
rect 38083 32152 38092 32192
rect 38132 32152 38141 32192
rect 38083 32151 38141 32152
rect 39619 32192 39677 32193
rect 39619 32152 39628 32192
rect 39668 32152 39677 32192
rect 39619 32151 39677 32152
rect 40579 32192 40637 32193
rect 40579 32152 40588 32192
rect 40628 32152 40637 32192
rect 40579 32151 40637 32152
rect 32611 32108 32669 32109
rect 32611 32068 32620 32108
rect 32660 32068 32669 32108
rect 32611 32067 32669 32068
rect 39723 32108 39765 32117
rect 39723 32068 39724 32108
rect 39764 32068 39765 32108
rect 39723 32059 39765 32068
rect 6027 32024 6069 32033
rect 6027 31984 6028 32024
rect 6068 31984 6069 32024
rect 6027 31975 6069 31984
rect 9387 32024 9429 32033
rect 9387 31984 9388 32024
rect 9428 31984 9429 32024
rect 9387 31975 9429 31984
rect 14955 32024 14997 32033
rect 14955 31984 14956 32024
rect 14996 31984 14997 32024
rect 14955 31975 14997 31984
rect 24267 32024 24309 32033
rect 24267 31984 24268 32024
rect 24308 31984 24309 32024
rect 24267 31975 24309 31984
rect 26187 32024 26229 32033
rect 26187 31984 26188 32024
rect 26228 31984 26229 32024
rect 26187 31975 26229 31984
rect 27723 32024 27765 32033
rect 27723 31984 27724 32024
rect 27764 31984 27765 32024
rect 27723 31975 27765 31984
rect 34251 32024 34293 32033
rect 34251 31984 34252 32024
rect 34292 31984 34293 32024
rect 34251 31975 34293 31984
rect 34827 32024 34869 32033
rect 34827 31984 34828 32024
rect 34868 31984 34869 32024
rect 34827 31975 34869 31984
rect 38763 32024 38805 32033
rect 38763 31984 38764 32024
rect 38804 31984 38805 32024
rect 38763 31975 38805 31984
rect 39243 32024 39285 32033
rect 39243 31984 39244 32024
rect 39284 31984 39285 32024
rect 39243 31975 39285 31984
rect 3523 31940 3581 31941
rect 3523 31900 3532 31940
rect 3572 31900 3581 31940
rect 3523 31899 3581 31900
rect 10435 31940 10493 31941
rect 10435 31900 10444 31940
rect 10484 31900 10493 31940
rect 10435 31899 10493 31900
rect 11299 31940 11357 31941
rect 11299 31900 11308 31940
rect 11348 31900 11357 31940
rect 11299 31899 11357 31900
rect 12267 31940 12309 31949
rect 12267 31900 12268 31940
rect 12308 31900 12309 31940
rect 12267 31891 12309 31900
rect 13411 31940 13469 31941
rect 13411 31900 13420 31940
rect 13460 31900 13469 31940
rect 13411 31899 13469 31900
rect 15331 31940 15389 31941
rect 15331 31900 15340 31940
rect 15380 31900 15389 31940
rect 15331 31899 15389 31900
rect 16299 31940 16341 31949
rect 16299 31900 16300 31940
rect 16340 31900 16341 31940
rect 16299 31891 16341 31900
rect 23787 31940 23829 31949
rect 23787 31900 23788 31940
rect 23828 31900 23829 31940
rect 23787 31891 23829 31900
rect 24931 31940 24989 31941
rect 24931 31900 24940 31940
rect 24980 31900 24989 31940
rect 24931 31899 24989 31900
rect 28683 31940 28725 31949
rect 28683 31900 28684 31940
rect 28724 31900 28725 31940
rect 28683 31891 28725 31900
rect 30507 31940 30549 31949
rect 30507 31900 30508 31940
rect 30548 31900 30549 31940
rect 30507 31891 30549 31900
rect 31747 31940 31805 31941
rect 31747 31900 31756 31940
rect 31796 31900 31805 31940
rect 31747 31899 31805 31900
rect 33867 31940 33909 31949
rect 33867 31900 33868 31940
rect 33908 31900 33909 31940
rect 33867 31891 33909 31900
rect 38571 31940 38613 31949
rect 38571 31900 38572 31940
rect 38612 31900 38613 31940
rect 38571 31891 38613 31900
rect 39907 31940 39965 31941
rect 39907 31900 39916 31940
rect 39956 31900 39965 31940
rect 39907 31899 39965 31900
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 13995 31604 14037 31613
rect 13995 31564 13996 31604
rect 14036 31564 14037 31604
rect 13995 31555 14037 31564
rect 15147 31604 15189 31613
rect 15147 31564 15148 31604
rect 15188 31564 15189 31604
rect 15147 31555 15189 31564
rect 26179 31604 26237 31605
rect 26179 31564 26188 31604
rect 26228 31564 26237 31604
rect 26179 31563 26237 31564
rect 29643 31604 29685 31613
rect 29643 31564 29644 31604
rect 29684 31564 29685 31604
rect 29643 31555 29685 31564
rect 32427 31604 32469 31613
rect 32427 31564 32428 31604
rect 32468 31564 32469 31604
rect 32427 31555 32469 31564
rect 37123 31604 37181 31605
rect 37123 31564 37132 31604
rect 37172 31564 37181 31604
rect 37123 31563 37181 31564
rect 1323 31520 1365 31529
rect 1323 31480 1324 31520
rect 1364 31480 1365 31520
rect 1323 31471 1365 31480
rect 3907 31520 3965 31521
rect 3907 31480 3916 31520
rect 3956 31480 3965 31520
rect 3907 31479 3965 31480
rect 6315 31520 6357 31529
rect 6315 31480 6316 31520
rect 6356 31480 6357 31520
rect 6315 31471 6357 31480
rect 6891 31520 6933 31529
rect 6891 31480 6892 31520
rect 6932 31480 6933 31520
rect 6891 31471 6933 31480
rect 9771 31520 9813 31529
rect 9771 31480 9772 31520
rect 9812 31480 9813 31520
rect 9771 31471 9813 31480
rect 12355 31520 12413 31521
rect 12355 31480 12364 31520
rect 12404 31480 12413 31520
rect 12355 31479 12413 31480
rect 18219 31520 18261 31529
rect 18219 31480 18220 31520
rect 18260 31480 18261 31520
rect 18219 31471 18261 31480
rect 18411 31520 18453 31529
rect 18411 31480 18412 31520
rect 18452 31480 18453 31520
rect 18411 31471 18453 31480
rect 21675 31520 21717 31529
rect 21675 31480 21676 31520
rect 21716 31480 21717 31520
rect 21675 31471 21717 31480
rect 26475 31520 26517 31529
rect 26475 31480 26476 31520
rect 26516 31480 26517 31520
rect 26475 31471 26517 31480
rect 28299 31520 28341 31529
rect 28299 31480 28300 31520
rect 28340 31480 28341 31520
rect 28299 31471 28341 31480
rect 41931 31520 41973 31529
rect 41931 31480 41932 31520
rect 41972 31480 41973 31520
rect 41931 31471 41973 31480
rect 4875 31436 4917 31445
rect 4875 31396 4876 31436
rect 4916 31396 4917 31436
rect 4875 31387 4917 31396
rect 1891 31352 1949 31353
rect 1891 31312 1900 31352
rect 1940 31312 1949 31352
rect 1891 31311 1949 31312
rect 2755 31352 2813 31353
rect 2755 31312 2764 31352
rect 2804 31312 2813 31352
rect 2755 31311 2813 31312
rect 4395 31352 4437 31361
rect 4395 31312 4396 31352
rect 4436 31312 4437 31352
rect 4395 31303 4437 31312
rect 4491 31352 4533 31361
rect 4491 31312 4492 31352
rect 4532 31312 4533 31352
rect 4491 31303 4533 31312
rect 4971 31352 5013 31361
rect 5931 31357 5973 31366
rect 4971 31312 4972 31352
rect 5012 31312 5013 31352
rect 4971 31303 5013 31312
rect 5443 31352 5501 31353
rect 5443 31312 5452 31352
rect 5492 31312 5501 31352
rect 5443 31311 5501 31312
rect 5931 31317 5932 31357
rect 5972 31317 5973 31357
rect 5931 31308 5973 31317
rect 6403 31352 6461 31353
rect 6403 31312 6412 31352
rect 6452 31312 6461 31352
rect 6403 31311 6461 31312
rect 7083 31352 7125 31361
rect 7083 31312 7084 31352
rect 7124 31312 7125 31352
rect 7083 31303 7125 31312
rect 7747 31352 7805 31353
rect 7747 31312 7756 31352
rect 7796 31312 7805 31352
rect 7747 31311 7805 31312
rect 8811 31352 8853 31361
rect 8811 31312 8812 31352
rect 8852 31312 8853 31352
rect 8811 31303 8853 31312
rect 9667 31352 9725 31353
rect 9667 31312 9676 31352
rect 9716 31312 9725 31352
rect 9667 31311 9725 31312
rect 9963 31352 10005 31361
rect 9963 31312 9964 31352
rect 10004 31312 10005 31352
rect 9963 31303 10005 31312
rect 10339 31352 10397 31353
rect 10339 31312 10348 31352
rect 10388 31312 10397 31352
rect 10339 31311 10397 31312
rect 11203 31352 11261 31353
rect 11203 31312 11212 31352
rect 11252 31312 11261 31352
rect 11203 31311 11261 31312
rect 12555 31352 12597 31361
rect 12555 31312 12556 31352
rect 12596 31312 12597 31352
rect 12555 31303 12597 31312
rect 12651 31352 12693 31361
rect 12651 31312 12652 31352
rect 12692 31312 12693 31352
rect 12651 31303 12693 31312
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 13227 31352 13269 31361
rect 13227 31312 13228 31352
rect 13268 31312 13269 31352
rect 13227 31303 13269 31312
rect 13315 31352 13373 31353
rect 13315 31312 13324 31352
rect 13364 31312 13373 31352
rect 13315 31311 13373 31312
rect 13507 31352 13565 31353
rect 13507 31312 13516 31352
rect 13556 31312 13565 31352
rect 13507 31311 13565 31312
rect 13611 31352 13653 31361
rect 13611 31312 13612 31352
rect 13652 31312 13653 31352
rect 13611 31303 13653 31312
rect 13803 31352 13845 31361
rect 13803 31312 13804 31352
rect 13844 31312 13845 31352
rect 13803 31303 13845 31312
rect 13995 31352 14037 31361
rect 13995 31312 13996 31352
rect 14036 31312 14037 31352
rect 13995 31303 14037 31312
rect 14187 31352 14229 31361
rect 14187 31312 14188 31352
rect 14228 31312 14229 31352
rect 14187 31303 14229 31312
rect 14275 31352 14333 31353
rect 14275 31312 14284 31352
rect 14324 31312 14333 31352
rect 14275 31311 14333 31312
rect 14659 31352 14717 31353
rect 14659 31312 14668 31352
rect 14708 31312 14717 31352
rect 14659 31311 14717 31312
rect 14851 31352 14909 31353
rect 14851 31312 14860 31352
rect 14900 31312 14909 31352
rect 14851 31311 14909 31312
rect 14955 31352 14997 31361
rect 14955 31312 14956 31352
rect 14996 31312 14997 31352
rect 14955 31303 14997 31312
rect 15147 31352 15189 31361
rect 15147 31312 15148 31352
rect 15188 31312 15189 31352
rect 15147 31303 15189 31312
rect 15339 31352 15381 31361
rect 15339 31312 15340 31352
rect 15380 31312 15381 31352
rect 15339 31303 15381 31312
rect 15435 31352 15477 31361
rect 15435 31312 15436 31352
rect 15476 31312 15477 31352
rect 15435 31303 15477 31312
rect 15531 31352 15573 31361
rect 15531 31312 15532 31352
rect 15572 31312 15573 31352
rect 15531 31303 15573 31312
rect 15627 31352 15669 31361
rect 15627 31312 15628 31352
rect 15668 31312 15669 31352
rect 15627 31303 15669 31312
rect 15819 31352 15861 31361
rect 15819 31312 15820 31352
rect 15860 31312 15861 31352
rect 15819 31303 15861 31312
rect 16011 31352 16053 31361
rect 16011 31312 16012 31352
rect 16052 31312 16053 31352
rect 16011 31303 16053 31312
rect 16099 31352 16157 31353
rect 16099 31312 16108 31352
rect 16148 31312 16157 31352
rect 16099 31311 16157 31312
rect 16291 31352 16349 31353
rect 16291 31312 16300 31352
rect 16340 31312 16349 31352
rect 16291 31311 16349 31312
rect 17163 31352 17205 31361
rect 17163 31312 17164 31352
rect 17204 31312 17205 31352
rect 17163 31303 17205 31312
rect 17827 31352 17885 31353
rect 17827 31312 17836 31352
rect 17876 31312 17885 31352
rect 17827 31311 17885 31312
rect 20707 31352 20765 31353
rect 20707 31312 20716 31352
rect 20756 31312 20765 31352
rect 20707 31311 20765 31312
rect 20899 31352 20957 31353
rect 20899 31312 20908 31352
rect 20948 31312 20957 31352
rect 20899 31311 20957 31312
rect 22531 31352 22589 31353
rect 22531 31312 22540 31352
rect 22580 31312 22589 31352
rect 22531 31311 22589 31312
rect 22731 31352 22773 31361
rect 22731 31312 22732 31352
rect 22772 31312 22773 31352
rect 22731 31303 22773 31312
rect 22827 31352 22869 31361
rect 22827 31312 22828 31352
rect 22868 31312 22869 31352
rect 22827 31303 22869 31312
rect 22923 31352 22965 31361
rect 22923 31312 22924 31352
rect 22964 31312 22965 31352
rect 22923 31303 22965 31312
rect 24163 31352 24221 31353
rect 24163 31312 24172 31352
rect 24212 31312 24221 31352
rect 24163 31311 24221 31312
rect 25027 31352 25085 31353
rect 25027 31312 25036 31352
rect 25076 31312 25085 31352
rect 25027 31311 25085 31312
rect 26371 31352 26429 31353
rect 26371 31312 26380 31352
rect 26420 31312 26429 31352
rect 26371 31311 26429 31312
rect 28099 31352 28157 31353
rect 28099 31312 28108 31352
rect 28148 31312 28157 31352
rect 28099 31311 28157 31312
rect 29347 31352 29405 31353
rect 29347 31312 29356 31352
rect 29396 31312 29405 31352
rect 29347 31311 29405 31312
rect 29451 31352 29493 31361
rect 29451 31312 29452 31352
rect 29492 31312 29493 31352
rect 29451 31303 29493 31312
rect 29643 31352 29685 31361
rect 29643 31312 29644 31352
rect 29684 31312 29685 31352
rect 29643 31303 29685 31312
rect 30499 31352 30557 31353
rect 30499 31312 30508 31352
rect 30548 31312 30557 31352
rect 30499 31311 30557 31312
rect 30691 31352 30749 31353
rect 30691 31312 30700 31352
rect 30740 31312 30749 31352
rect 30691 31311 30749 31312
rect 31651 31352 31709 31353
rect 31651 31312 31660 31352
rect 31700 31312 31709 31352
rect 31651 31311 31709 31312
rect 31939 31352 31997 31353
rect 31939 31312 31948 31352
rect 31988 31312 31997 31352
rect 31939 31311 31997 31312
rect 32899 31352 32957 31353
rect 32899 31312 32908 31352
rect 32948 31312 32957 31352
rect 32899 31311 32957 31312
rect 33387 31352 33429 31361
rect 33387 31312 33388 31352
rect 33428 31312 33429 31352
rect 33387 31303 33429 31312
rect 35107 31352 35165 31353
rect 35107 31312 35116 31352
rect 35156 31312 35165 31352
rect 35107 31311 35165 31312
rect 35971 31352 36029 31353
rect 35971 31312 35980 31352
rect 36020 31312 36029 31352
rect 35971 31311 36029 31312
rect 38179 31352 38237 31353
rect 38179 31312 38188 31352
rect 38228 31312 38237 31352
rect 38179 31311 38237 31312
rect 38755 31352 38813 31353
rect 38755 31312 38764 31352
rect 38804 31312 38813 31352
rect 38755 31311 38813 31312
rect 39619 31352 39677 31353
rect 39619 31312 39628 31352
rect 39668 31312 39677 31352
rect 39619 31311 39677 31312
rect 43267 31352 43325 31353
rect 43267 31312 43276 31352
rect 43316 31312 43325 31352
rect 43267 31311 43325 31312
rect 1515 31268 1557 31277
rect 1515 31228 1516 31268
rect 1556 31228 1557 31268
rect 1515 31219 1557 31228
rect 8035 31268 8093 31269
rect 8035 31228 8044 31268
rect 8084 31228 8093 31268
rect 8035 31227 8093 31228
rect 13707 31268 13749 31277
rect 13707 31228 13708 31268
rect 13748 31228 13749 31268
rect 13707 31219 13749 31228
rect 15915 31268 15957 31277
rect 15915 31228 15916 31268
rect 15956 31228 15957 31268
rect 15915 31219 15957 31228
rect 23787 31268 23829 31277
rect 23787 31228 23788 31268
rect 23828 31228 23829 31268
rect 23787 31219 23829 31228
rect 34731 31268 34773 31277
rect 34731 31228 34732 31268
rect 34772 31228 34773 31268
rect 34731 31219 34773 31228
rect 38379 31268 38421 31277
rect 38379 31228 38380 31268
rect 38420 31228 38421 31268
rect 38379 31219 38421 31228
rect 6123 31184 6165 31193
rect 6123 31144 6124 31184
rect 6164 31144 6165 31184
rect 6123 31135 6165 31144
rect 12835 31184 12893 31185
rect 12835 31144 12844 31184
rect 12884 31144 12893 31184
rect 12835 31143 12893 31144
rect 14571 31184 14613 31193
rect 14571 31144 14572 31184
rect 14612 31144 14613 31184
rect 14571 31135 14613 31144
rect 16963 31184 17021 31185
rect 16963 31144 16972 31184
rect 17012 31144 17021 31184
rect 16963 31143 17021 31144
rect 21859 31184 21917 31185
rect 21859 31144 21868 31184
rect 21908 31144 21917 31184
rect 21859 31143 21917 31144
rect 23011 31184 23069 31185
rect 23011 31144 23020 31184
rect 23060 31144 23069 31184
rect 23011 31143 23069 31144
rect 27427 31184 27485 31185
rect 27427 31144 27436 31184
rect 27476 31144 27485 31184
rect 27427 31143 27485 31144
rect 29827 31184 29885 31185
rect 29827 31144 29836 31184
rect 29876 31144 29885 31184
rect 29827 31143 29885 31144
rect 33771 31184 33813 31193
rect 33771 31144 33772 31184
rect 33812 31144 33813 31184
rect 33771 31135 33813 31144
rect 37507 31184 37565 31185
rect 37507 31144 37516 31184
rect 37556 31144 37565 31184
rect 37507 31143 37565 31144
rect 40771 31184 40829 31185
rect 40771 31144 40780 31184
rect 40820 31144 40829 31184
rect 40771 31143 40829 31144
rect 43179 31184 43221 31193
rect 43179 31144 43180 31184
rect 43220 31144 43221 31184
rect 43179 31135 43221 31144
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 3907 30848 3965 30849
rect 3907 30808 3916 30848
rect 3956 30808 3965 30848
rect 3907 30807 3965 30808
rect 4771 30848 4829 30849
rect 4771 30808 4780 30848
rect 4820 30808 4829 30848
rect 4771 30807 4829 30808
rect 7555 30848 7613 30849
rect 7555 30808 7564 30848
rect 7604 30808 7613 30848
rect 7555 30807 7613 30808
rect 10915 30848 10973 30849
rect 10915 30808 10924 30848
rect 10964 30808 10973 30848
rect 10915 30807 10973 30808
rect 12835 30848 12893 30849
rect 12835 30808 12844 30848
rect 12884 30808 12893 30848
rect 12835 30807 12893 30808
rect 16483 30848 16541 30849
rect 16483 30808 16492 30848
rect 16532 30808 16541 30848
rect 16483 30807 16541 30808
rect 32227 30848 32285 30849
rect 32227 30808 32236 30848
rect 32276 30808 32285 30848
rect 32227 30807 32285 30808
rect 33291 30848 33333 30857
rect 33291 30808 33292 30848
rect 33332 30808 33333 30848
rect 33291 30799 33333 30808
rect 35587 30848 35645 30849
rect 35587 30808 35596 30848
rect 35636 30808 35645 30848
rect 35587 30807 35645 30808
rect 38947 30848 39005 30849
rect 38947 30808 38956 30848
rect 38996 30808 39005 30848
rect 38947 30807 39005 30808
rect 9963 30764 10005 30773
rect 9963 30724 9964 30764
rect 10004 30724 10005 30764
rect 9963 30715 10005 30724
rect 13515 30764 13557 30773
rect 13515 30724 13516 30764
rect 13556 30724 13557 30764
rect 13515 30715 13557 30724
rect 18891 30764 18933 30773
rect 18891 30724 18892 30764
rect 18932 30724 18933 30764
rect 18891 30715 18933 30724
rect 21387 30764 21429 30773
rect 21387 30724 21388 30764
rect 21428 30724 21429 30764
rect 21387 30715 21429 30724
rect 25995 30764 26037 30773
rect 25995 30724 25996 30764
rect 26036 30724 26037 30764
rect 25995 30715 26037 30724
rect 26763 30764 26805 30773
rect 26763 30724 26764 30764
rect 26804 30724 26805 30764
rect 26763 30715 26805 30724
rect 27435 30764 27477 30773
rect 27435 30724 27436 30764
rect 27476 30724 27477 30764
rect 27435 30715 27477 30724
rect 36651 30764 36693 30773
rect 36651 30724 36652 30764
rect 36692 30724 36693 30764
rect 36651 30715 36693 30724
rect 3715 30680 3773 30681
rect 3715 30640 3724 30680
rect 3764 30640 3773 30680
rect 3715 30639 3773 30640
rect 4579 30680 4637 30681
rect 4579 30640 4588 30680
rect 4628 30640 4637 30680
rect 4579 30639 4637 30640
rect 4875 30680 4917 30689
rect 4875 30640 4876 30680
rect 4916 30640 4917 30680
rect 4875 30631 4917 30640
rect 4971 30680 5013 30689
rect 4971 30640 4972 30680
rect 5012 30640 5013 30680
rect 4971 30631 5013 30640
rect 5067 30680 5109 30689
rect 5067 30640 5068 30680
rect 5108 30640 5109 30680
rect 5067 30631 5109 30640
rect 5827 30680 5885 30681
rect 5827 30640 5836 30680
rect 5876 30640 5885 30680
rect 5827 30639 5885 30640
rect 6019 30680 6077 30681
rect 6019 30640 6028 30680
rect 6068 30640 6077 30680
rect 6019 30639 6077 30640
rect 6219 30680 6261 30689
rect 6219 30640 6220 30680
rect 6260 30640 6261 30680
rect 6219 30631 6261 30640
rect 6315 30680 6357 30689
rect 6315 30640 6316 30680
rect 6356 30640 6357 30680
rect 6315 30631 6357 30640
rect 6411 30680 6453 30689
rect 6411 30640 6412 30680
rect 6452 30640 6453 30680
rect 6411 30631 6453 30640
rect 6507 30680 6549 30689
rect 6507 30640 6508 30680
rect 6548 30640 6549 30680
rect 6507 30631 6549 30640
rect 8707 30680 8765 30681
rect 8707 30640 8716 30680
rect 8756 30640 8765 30680
rect 8707 30639 8765 30640
rect 9571 30680 9629 30681
rect 9571 30640 9580 30680
rect 9620 30640 9629 30680
rect 9571 30639 9629 30640
rect 10723 30680 10781 30681
rect 10723 30640 10732 30680
rect 10772 30640 10781 30680
rect 10723 30639 10781 30640
rect 10827 30680 10869 30689
rect 10827 30640 10828 30680
rect 10868 30640 10869 30680
rect 10827 30631 10869 30640
rect 11019 30680 11061 30689
rect 11019 30640 11020 30680
rect 11060 30640 11061 30680
rect 11019 30631 11061 30640
rect 12075 30680 12117 30689
rect 12075 30640 12076 30680
rect 12116 30640 12117 30680
rect 12075 30631 12117 30640
rect 12555 30680 12597 30689
rect 12555 30640 12556 30680
rect 12596 30640 12597 30680
rect 12555 30631 12597 30640
rect 12651 30680 12693 30689
rect 12651 30640 12652 30680
rect 12692 30640 12693 30680
rect 12651 30631 12693 30640
rect 12747 30680 12789 30689
rect 12747 30640 12748 30680
rect 12788 30640 12789 30680
rect 12747 30631 12789 30640
rect 13123 30680 13181 30681
rect 13123 30640 13132 30680
rect 13172 30640 13181 30680
rect 13123 30639 13181 30640
rect 13419 30680 13461 30689
rect 13419 30640 13420 30680
rect 13460 30640 13461 30680
rect 13419 30631 13461 30640
rect 13987 30680 14045 30681
rect 13987 30640 13996 30680
rect 14036 30640 14045 30680
rect 13987 30639 14045 30640
rect 15523 30680 15581 30681
rect 15523 30640 15532 30680
rect 15572 30640 15581 30680
rect 15523 30639 15581 30640
rect 15819 30680 15861 30689
rect 15819 30640 15820 30680
rect 15860 30640 15861 30680
rect 15819 30631 15861 30640
rect 15915 30680 15957 30689
rect 15915 30640 15916 30680
rect 15956 30640 15957 30680
rect 15915 30631 15957 30640
rect 17635 30680 17693 30681
rect 17635 30640 17644 30680
rect 17684 30640 17693 30680
rect 17635 30639 17693 30640
rect 18499 30680 18557 30681
rect 18499 30640 18508 30680
rect 18548 30640 18557 30680
rect 18499 30639 18557 30640
rect 19083 30680 19125 30689
rect 19083 30640 19084 30680
rect 19124 30640 19125 30680
rect 19083 30631 19125 30640
rect 19179 30680 19221 30689
rect 19179 30640 19180 30680
rect 19220 30640 19221 30680
rect 19179 30631 19221 30640
rect 19275 30680 19317 30689
rect 19275 30640 19276 30680
rect 19316 30640 19317 30680
rect 19275 30631 19317 30640
rect 19371 30680 19413 30689
rect 19371 30640 19372 30680
rect 19412 30640 19413 30680
rect 19371 30631 19413 30640
rect 19659 30680 19701 30689
rect 19659 30640 19660 30680
rect 19700 30640 19701 30680
rect 19659 30631 19701 30640
rect 19755 30680 19797 30689
rect 19755 30640 19756 30680
rect 19796 30640 19797 30680
rect 19755 30631 19797 30640
rect 19851 30680 19893 30689
rect 19851 30640 19852 30680
rect 19892 30640 19893 30680
rect 20131 30680 20189 30681
rect 19851 30631 19893 30640
rect 19947 30635 19989 30644
rect 20131 30640 20140 30680
rect 20180 30640 20189 30680
rect 20131 30639 20189 30640
rect 21091 30680 21149 30681
rect 21091 30640 21100 30680
rect 21140 30640 21149 30680
rect 21091 30639 21149 30640
rect 21763 30680 21821 30681
rect 21763 30640 21772 30680
rect 21812 30640 21821 30680
rect 21763 30639 21821 30640
rect 22627 30680 22685 30681
rect 22627 30640 22636 30680
rect 22676 30640 22685 30680
rect 22627 30639 22685 30640
rect 25035 30680 25077 30689
rect 25035 30640 25036 30680
rect 25076 30640 25077 30680
rect 19947 30595 19948 30635
rect 19988 30595 19989 30635
rect 25035 30631 25077 30640
rect 25131 30680 25173 30689
rect 25131 30640 25132 30680
rect 25172 30640 25173 30680
rect 25131 30631 25173 30640
rect 25227 30680 25269 30689
rect 25227 30640 25228 30680
rect 25268 30640 25269 30680
rect 25227 30631 25269 30640
rect 25323 30680 25365 30689
rect 25323 30640 25324 30680
rect 25364 30640 25365 30680
rect 25323 30631 25365 30640
rect 25603 30680 25661 30681
rect 25603 30640 25612 30680
rect 25652 30640 25661 30680
rect 25603 30639 25661 30640
rect 25899 30680 25941 30689
rect 25899 30640 25900 30680
rect 25940 30640 25941 30680
rect 25899 30631 25941 30640
rect 26475 30680 26517 30689
rect 26475 30640 26476 30680
rect 26516 30640 26517 30680
rect 26475 30631 26517 30640
rect 26571 30680 26613 30689
rect 26571 30640 26572 30680
rect 26612 30640 26613 30680
rect 26571 30631 26613 30640
rect 26667 30680 26709 30689
rect 26667 30640 26668 30680
rect 26708 30640 26709 30680
rect 26667 30631 26709 30640
rect 26947 30680 27005 30681
rect 26947 30640 26956 30680
rect 26996 30640 27005 30680
rect 26947 30639 27005 30640
rect 27051 30680 27093 30689
rect 27051 30640 27052 30680
rect 27092 30640 27093 30680
rect 27051 30631 27093 30640
rect 27243 30680 27285 30689
rect 27243 30640 27244 30680
rect 27284 30640 27285 30680
rect 27243 30631 27285 30640
rect 27811 30680 27869 30681
rect 27811 30640 27820 30680
rect 27860 30640 27869 30680
rect 27811 30639 27869 30640
rect 28675 30680 28733 30681
rect 28675 30640 28684 30680
rect 28724 30640 28733 30680
rect 28675 30639 28733 30640
rect 30019 30680 30077 30681
rect 30019 30640 30028 30680
rect 30068 30640 30077 30680
rect 30019 30639 30077 30640
rect 31555 30680 31613 30681
rect 31555 30640 31564 30680
rect 31604 30640 31613 30680
rect 31555 30639 31613 30640
rect 31755 30680 31797 30689
rect 31755 30640 31756 30680
rect 31796 30640 31797 30680
rect 31755 30631 31797 30640
rect 31947 30680 31989 30689
rect 31947 30640 31948 30680
rect 31988 30640 31989 30680
rect 31947 30631 31989 30640
rect 32035 30680 32093 30681
rect 32035 30640 32044 30680
rect 32084 30640 32093 30680
rect 32035 30639 32093 30640
rect 32331 30680 32373 30689
rect 32331 30640 32332 30680
rect 32372 30640 32373 30680
rect 32331 30631 32373 30640
rect 32427 30680 32469 30689
rect 32427 30640 32428 30680
rect 32468 30640 32469 30680
rect 32427 30631 32469 30640
rect 32523 30680 32565 30689
rect 32523 30640 32524 30680
rect 32564 30640 32565 30680
rect 32523 30631 32565 30640
rect 33675 30680 33717 30689
rect 33675 30640 33676 30680
rect 33716 30640 33717 30680
rect 33675 30631 33717 30640
rect 34051 30680 34109 30681
rect 34051 30640 34060 30680
rect 34100 30640 34109 30680
rect 34051 30639 34109 30640
rect 34243 30680 34301 30681
rect 34243 30640 34252 30680
rect 34292 30640 34301 30680
rect 34243 30639 34301 30640
rect 34539 30680 34581 30689
rect 34539 30640 34540 30680
rect 34580 30640 34581 30680
rect 34539 30631 34581 30640
rect 34635 30680 34677 30689
rect 34635 30640 34636 30680
rect 34676 30640 34677 30680
rect 34635 30631 34677 30640
rect 34731 30680 34773 30689
rect 34731 30640 34732 30680
rect 34772 30640 34773 30680
rect 34731 30631 34773 30640
rect 34827 30680 34869 30689
rect 34827 30640 34828 30680
rect 34868 30640 34869 30680
rect 34827 30631 34869 30640
rect 35019 30680 35061 30689
rect 35019 30640 35020 30680
rect 35060 30640 35061 30680
rect 35019 30631 35061 30640
rect 35115 30680 35157 30689
rect 35115 30640 35116 30680
rect 35156 30640 35157 30680
rect 35115 30631 35157 30640
rect 35211 30680 35253 30689
rect 35211 30640 35212 30680
rect 35252 30640 35253 30680
rect 35211 30631 35253 30640
rect 35307 30680 35349 30689
rect 35307 30640 35308 30680
rect 35348 30640 35349 30680
rect 35307 30631 35349 30640
rect 35499 30680 35541 30689
rect 35499 30640 35500 30680
rect 35540 30640 35541 30680
rect 35499 30631 35541 30640
rect 35691 30680 35733 30689
rect 35691 30640 35692 30680
rect 35732 30640 35733 30680
rect 35691 30631 35733 30640
rect 35779 30680 35837 30681
rect 35779 30640 35788 30680
rect 35828 30640 35837 30680
rect 35779 30639 35837 30640
rect 36451 30680 36509 30681
rect 36451 30640 36460 30680
rect 36500 30640 36509 30680
rect 36451 30639 36509 30640
rect 36555 30680 36597 30689
rect 36555 30640 36556 30680
rect 36596 30640 36597 30680
rect 36555 30631 36597 30640
rect 36747 30680 36789 30689
rect 36747 30640 36748 30680
rect 36788 30640 36789 30680
rect 36747 30631 36789 30640
rect 36939 30680 36981 30689
rect 36939 30640 36940 30680
rect 36980 30640 36981 30680
rect 36939 30631 36981 30640
rect 37035 30680 37077 30689
rect 37035 30640 37036 30680
rect 37076 30640 37077 30680
rect 37035 30631 37077 30640
rect 37131 30680 37173 30689
rect 37131 30640 37132 30680
rect 37172 30640 37173 30680
rect 37131 30631 37173 30640
rect 37227 30680 37269 30689
rect 37227 30640 37228 30680
rect 37268 30640 37269 30680
rect 37227 30631 37269 30640
rect 37411 30680 37469 30681
rect 37411 30640 37420 30680
rect 37460 30640 37469 30680
rect 37411 30639 37469 30640
rect 38275 30680 38333 30681
rect 38275 30640 38284 30680
rect 38324 30640 38333 30680
rect 38275 30639 38333 30640
rect 39147 30680 39189 30689
rect 39147 30640 39148 30680
rect 39188 30640 39189 30680
rect 39147 30631 39189 30640
rect 39243 30680 39285 30689
rect 39243 30640 39244 30680
rect 39284 30640 39285 30680
rect 39243 30631 39285 30640
rect 39339 30680 39381 30689
rect 39339 30640 39340 30680
rect 39380 30640 39381 30680
rect 39339 30631 39381 30640
rect 39435 30680 39477 30689
rect 39435 30640 39436 30680
rect 39476 30640 39477 30680
rect 39435 30631 39477 30640
rect 40099 30680 40157 30681
rect 40099 30640 40108 30680
rect 40148 30640 40157 30680
rect 40099 30639 40157 30640
rect 41451 30680 41493 30689
rect 41451 30640 41452 30680
rect 41492 30640 41493 30680
rect 41451 30631 41493 30640
rect 41827 30680 41885 30681
rect 41827 30640 41836 30680
rect 41876 30640 41885 30680
rect 41827 30639 41885 30640
rect 42691 30680 42749 30681
rect 42691 30640 42700 30680
rect 42740 30640 42749 30680
rect 42691 30639 42749 30640
rect 44803 30680 44861 30681
rect 44803 30640 44812 30680
rect 44852 30640 44861 30680
rect 44803 30639 44861 30640
rect 45483 30680 45525 30689
rect 45483 30640 45484 30680
rect 45524 30640 45525 30680
rect 45483 30631 45525 30640
rect 45667 30680 45725 30681
rect 45667 30640 45676 30680
rect 45716 30640 45725 30680
rect 45667 30639 45725 30640
rect 19947 30586 19989 30595
rect 39619 30596 39677 30597
rect 39619 30556 39628 30596
rect 39668 30556 39677 30596
rect 39619 30555 39677 30556
rect 1803 30512 1845 30521
rect 1803 30472 1804 30512
rect 1844 30472 1845 30512
rect 1803 30463 1845 30472
rect 5355 30512 5397 30521
rect 5355 30472 5356 30512
rect 5396 30472 5397 30512
rect 5355 30463 5397 30472
rect 11499 30512 11541 30521
rect 11499 30472 11500 30512
rect 11540 30472 11541 30512
rect 11499 30463 11541 30472
rect 15051 30512 15093 30521
rect 15051 30472 15052 30512
rect 15092 30472 15093 30512
rect 15051 30463 15093 30472
rect 27243 30512 27285 30521
rect 27243 30472 27244 30512
rect 27284 30472 27285 30512
rect 27243 30463 27285 30472
rect 36171 30512 36213 30521
rect 36171 30472 36172 30512
rect 36212 30472 36213 30512
rect 36171 30463 36213 30472
rect 44427 30512 44469 30521
rect 44427 30472 44428 30512
rect 44468 30472 44469 30512
rect 44427 30463 44469 30472
rect 3043 30428 3101 30429
rect 3043 30388 3052 30428
rect 3092 30388 3101 30428
rect 3043 30387 3101 30388
rect 13795 30428 13853 30429
rect 13795 30388 13804 30428
rect 13844 30388 13853 30428
rect 13795 30387 13853 30388
rect 14659 30428 14717 30429
rect 14659 30388 14668 30428
rect 14708 30388 14717 30428
rect 14659 30387 14717 30388
rect 16195 30428 16253 30429
rect 16195 30388 16204 30428
rect 16244 30388 16253 30428
rect 16195 30387 16253 30388
rect 20619 30428 20661 30437
rect 20619 30388 20620 30428
rect 20660 30388 20661 30428
rect 20619 30379 20661 30388
rect 23779 30428 23837 30429
rect 23779 30388 23788 30428
rect 23828 30388 23837 30428
rect 23779 30387 23837 30388
rect 26275 30428 26333 30429
rect 26275 30388 26284 30428
rect 26324 30388 26333 30428
rect 26275 30387 26333 30388
rect 29827 30428 29885 30429
rect 29827 30388 29836 30428
rect 29876 30388 29885 30428
rect 29827 30387 29885 30388
rect 30691 30428 30749 30429
rect 30691 30388 30700 30428
rect 30740 30388 30749 30428
rect 30691 30387 30749 30388
rect 30883 30428 30941 30429
rect 30883 30388 30892 30428
rect 30932 30388 30941 30428
rect 30883 30387 30941 30388
rect 31755 30428 31797 30437
rect 31755 30388 31756 30428
rect 31796 30388 31797 30428
rect 31755 30379 31797 30388
rect 38083 30428 38141 30429
rect 38083 30388 38092 30428
rect 38132 30388 38141 30428
rect 38083 30387 38141 30388
rect 40011 30428 40053 30437
rect 40011 30388 40012 30428
rect 40052 30388 40053 30428
rect 40011 30379 40053 30388
rect 43843 30428 43901 30429
rect 43843 30388 43852 30428
rect 43892 30388 43901 30428
rect 43843 30387 43901 30388
rect 45771 30428 45813 30437
rect 45771 30388 45772 30428
rect 45812 30388 45813 30428
rect 45771 30379 45813 30388
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 3715 30092 3773 30093
rect 3715 30052 3724 30092
rect 3764 30052 3773 30092
rect 3715 30051 3773 30052
rect 4875 30092 4917 30101
rect 4875 30052 4876 30092
rect 4916 30052 4917 30092
rect 4875 30043 4917 30052
rect 6499 30092 6557 30093
rect 6499 30052 6508 30092
rect 6548 30052 6557 30092
rect 6499 30051 6557 30052
rect 12459 30092 12501 30101
rect 12459 30052 12460 30092
rect 12500 30052 12501 30092
rect 12459 30043 12501 30052
rect 13411 30092 13469 30093
rect 13411 30052 13420 30092
rect 13460 30052 13469 30092
rect 13411 30051 13469 30052
rect 16491 30092 16533 30101
rect 16491 30052 16492 30092
rect 16532 30052 16533 30092
rect 16491 30043 16533 30052
rect 22251 30092 22293 30101
rect 22251 30052 22252 30092
rect 22292 30052 22293 30092
rect 22251 30043 22293 30052
rect 26763 30092 26805 30101
rect 26763 30052 26764 30092
rect 26804 30052 26805 30092
rect 26763 30043 26805 30052
rect 36067 30092 36125 30093
rect 36067 30052 36076 30092
rect 36116 30052 36125 30092
rect 36067 30051 36125 30052
rect 41635 30092 41693 30093
rect 41635 30052 41644 30092
rect 41684 30052 41693 30092
rect 41635 30051 41693 30052
rect 7851 30008 7893 30017
rect 7851 29968 7852 30008
rect 7892 29968 7893 30008
rect 7851 29959 7893 29968
rect 9867 30008 9909 30017
rect 9867 29968 9868 30008
rect 9908 29968 9909 30008
rect 9867 29959 9909 29968
rect 20715 30008 20757 30017
rect 20715 29968 20716 30008
rect 20756 29968 20757 30008
rect 20715 29959 20757 29968
rect 27715 30008 27773 30009
rect 27715 29968 27724 30008
rect 27764 29968 27773 30008
rect 27715 29967 27773 29968
rect 29259 30008 29301 30017
rect 29259 29968 29260 30008
rect 29300 29968 29301 30008
rect 29259 29959 29301 29968
rect 33387 30008 33429 30017
rect 33387 29968 33388 30008
rect 33428 29968 33429 30008
rect 33387 29959 33429 29968
rect 40491 30008 40533 30017
rect 40491 29968 40492 30008
rect 40532 29968 40533 30008
rect 40491 29959 40533 29968
rect 46635 30008 46677 30017
rect 46635 29968 46636 30008
rect 46676 29968 46677 30008
rect 46635 29959 46677 29968
rect 37419 29924 37461 29933
rect 37419 29884 37420 29924
rect 37460 29884 37461 29924
rect 37419 29875 37461 29884
rect 1323 29840 1365 29849
rect 1323 29800 1324 29840
rect 1364 29800 1365 29840
rect 1323 29791 1365 29800
rect 1699 29840 1757 29841
rect 1699 29800 1708 29840
rect 1748 29800 1757 29840
rect 1699 29799 1757 29800
rect 2563 29840 2621 29841
rect 2563 29800 2572 29840
rect 2612 29800 2621 29840
rect 2563 29799 2621 29800
rect 4203 29840 4245 29849
rect 4203 29800 4204 29840
rect 4244 29800 4245 29840
rect 4203 29791 4245 29800
rect 4299 29840 4341 29849
rect 4299 29800 4300 29840
rect 4340 29800 4341 29840
rect 4299 29791 4341 29800
rect 4395 29840 4437 29849
rect 4395 29800 4396 29840
rect 4436 29800 4437 29840
rect 4395 29791 4437 29800
rect 4579 29840 4637 29841
rect 4579 29800 4588 29840
rect 4628 29800 4637 29840
rect 4579 29799 4637 29800
rect 4683 29840 4725 29849
rect 4683 29800 4684 29840
rect 4724 29800 4725 29840
rect 4683 29791 4725 29800
rect 4875 29840 4917 29849
rect 4875 29800 4876 29840
rect 4916 29800 4917 29840
rect 4875 29791 4917 29800
rect 5067 29840 5109 29849
rect 5067 29800 5068 29840
rect 5108 29800 5109 29840
rect 5067 29791 5109 29800
rect 5163 29840 5205 29849
rect 5163 29800 5164 29840
rect 5204 29800 5205 29840
rect 5163 29791 5205 29800
rect 5259 29840 5301 29849
rect 5259 29800 5260 29840
rect 5300 29800 5301 29840
rect 5259 29791 5301 29800
rect 5355 29840 5397 29849
rect 5355 29800 5356 29840
rect 5396 29800 5397 29840
rect 5355 29791 5397 29800
rect 6307 29840 6365 29841
rect 6307 29800 6316 29840
rect 6356 29800 6365 29840
rect 6307 29799 6365 29800
rect 7171 29840 7229 29841
rect 7171 29800 7180 29840
rect 7220 29800 7229 29840
rect 7171 29799 7229 29800
rect 7459 29840 7517 29841
rect 7459 29800 7468 29840
rect 7508 29800 7517 29840
rect 7459 29799 7517 29800
rect 8043 29840 8085 29849
rect 8043 29800 8044 29840
rect 8084 29800 8085 29840
rect 8043 29791 8085 29800
rect 8139 29840 8181 29849
rect 8139 29800 8140 29840
rect 8180 29800 8181 29840
rect 8139 29791 8181 29800
rect 8235 29840 8277 29849
rect 8235 29800 8236 29840
rect 8276 29800 8277 29840
rect 8235 29791 8277 29800
rect 8331 29840 8373 29849
rect 8331 29800 8332 29840
rect 8372 29800 8373 29840
rect 8331 29791 8373 29800
rect 8523 29840 8565 29849
rect 8523 29800 8524 29840
rect 8564 29800 8565 29840
rect 8523 29791 8565 29800
rect 8715 29840 8757 29849
rect 8715 29800 8716 29840
rect 8756 29800 8757 29840
rect 8715 29791 8757 29800
rect 8803 29840 8861 29841
rect 8803 29800 8812 29840
rect 8852 29800 8861 29840
rect 8803 29799 8861 29800
rect 9667 29840 9725 29841
rect 9667 29800 9676 29840
rect 9716 29800 9725 29840
rect 9667 29799 9725 29800
rect 10915 29840 10973 29841
rect 10915 29800 10924 29840
rect 10964 29800 10973 29840
rect 10915 29799 10973 29800
rect 11875 29840 11933 29841
rect 11875 29800 11884 29840
rect 11924 29800 11933 29840
rect 11875 29799 11933 29800
rect 12163 29840 12221 29841
rect 12163 29800 12172 29840
rect 12212 29800 12221 29840
rect 12163 29799 12221 29800
rect 13035 29840 13077 29849
rect 13035 29800 13036 29840
rect 13076 29800 13077 29840
rect 13035 29791 13077 29800
rect 14563 29840 14621 29841
rect 14563 29800 14572 29840
rect 14612 29800 14621 29840
rect 14563 29799 14621 29800
rect 15427 29840 15485 29841
rect 15427 29800 15436 29840
rect 15476 29800 15485 29840
rect 15427 29799 15485 29800
rect 15819 29840 15861 29849
rect 15819 29800 15820 29840
rect 15860 29800 15861 29840
rect 15819 29791 15861 29800
rect 16875 29840 16917 29849
rect 16875 29800 16876 29840
rect 16916 29800 16917 29840
rect 16875 29791 16917 29800
rect 17251 29840 17309 29841
rect 17251 29800 17260 29840
rect 17300 29800 17309 29840
rect 17251 29799 17309 29800
rect 18499 29840 18557 29841
rect 18499 29800 18508 29840
rect 18548 29800 18557 29840
rect 18499 29799 18557 29800
rect 19363 29840 19421 29841
rect 19363 29800 19372 29840
rect 19412 29800 19421 29840
rect 19363 29799 19421 29800
rect 21763 29840 21821 29841
rect 21763 29800 21772 29840
rect 21812 29800 21821 29840
rect 21763 29799 21821 29800
rect 21955 29840 22013 29841
rect 21955 29800 21964 29840
rect 22004 29800 22013 29840
rect 21955 29799 22013 29800
rect 22059 29840 22101 29849
rect 22059 29800 22060 29840
rect 22100 29800 22101 29840
rect 22059 29791 22101 29800
rect 22251 29840 22293 29849
rect 22251 29800 22252 29840
rect 22292 29800 22293 29840
rect 22251 29791 22293 29800
rect 22915 29840 22973 29841
rect 22915 29800 22924 29840
rect 22964 29800 22973 29840
rect 22915 29799 22973 29800
rect 23779 29840 23837 29841
rect 23779 29800 23788 29840
rect 23828 29800 23837 29840
rect 23779 29799 23837 29800
rect 25227 29840 25269 29849
rect 25227 29800 25228 29840
rect 25268 29800 25269 29840
rect 25227 29791 25269 29800
rect 25419 29840 25461 29849
rect 25419 29800 25420 29840
rect 25460 29800 25461 29840
rect 25419 29791 25461 29800
rect 25507 29840 25565 29841
rect 25507 29800 25516 29840
rect 25556 29800 25565 29840
rect 25507 29799 25565 29800
rect 25699 29840 25757 29841
rect 25699 29800 25708 29840
rect 25748 29800 25757 29840
rect 25699 29799 25757 29800
rect 26659 29840 26717 29841
rect 26659 29800 26668 29840
rect 26708 29800 26717 29840
rect 26659 29799 26717 29800
rect 27043 29840 27101 29841
rect 27043 29800 27052 29840
rect 27092 29800 27101 29840
rect 27043 29799 27101 29800
rect 27339 29840 27381 29849
rect 27339 29800 27340 29840
rect 27380 29800 27381 29840
rect 27339 29791 27381 29800
rect 27435 29840 27477 29849
rect 27435 29800 27436 29840
rect 27476 29800 27477 29840
rect 27435 29791 27477 29800
rect 29827 29840 29885 29841
rect 29827 29800 29836 29840
rect 29876 29800 29885 29840
rect 29827 29799 29885 29800
rect 30691 29840 30749 29841
rect 30691 29800 30700 29840
rect 30740 29800 30749 29840
rect 30691 29799 30749 29800
rect 32707 29840 32765 29841
rect 32707 29800 32716 29840
rect 32756 29800 32765 29840
rect 32707 29799 32765 29800
rect 32907 29840 32949 29849
rect 32907 29800 32908 29840
rect 32948 29800 32949 29840
rect 32907 29791 32949 29800
rect 33003 29840 33045 29849
rect 33003 29800 33004 29840
rect 33044 29800 33045 29840
rect 33003 29791 33045 29800
rect 33099 29840 33141 29849
rect 33099 29800 33100 29840
rect 33140 29800 33141 29840
rect 33099 29791 33141 29800
rect 33195 29840 33237 29849
rect 33195 29800 33196 29840
rect 33236 29800 33237 29840
rect 33195 29791 33237 29800
rect 33963 29840 34005 29849
rect 33963 29800 33964 29840
rect 34004 29800 34005 29840
rect 33963 29791 34005 29800
rect 34627 29840 34685 29841
rect 34627 29800 34636 29840
rect 34676 29800 34685 29840
rect 34627 29799 34685 29800
rect 35019 29840 35061 29849
rect 35019 29800 35020 29840
rect 35060 29800 35061 29840
rect 35019 29791 35061 29800
rect 35211 29840 35253 29849
rect 35211 29800 35212 29840
rect 35252 29800 35253 29840
rect 35211 29791 35253 29800
rect 35299 29840 35357 29841
rect 35299 29800 35308 29840
rect 35348 29800 35357 29840
rect 35299 29799 35357 29800
rect 35691 29840 35733 29849
rect 35691 29800 35692 29840
rect 35732 29800 35733 29840
rect 35691 29791 35733 29800
rect 35875 29840 35933 29841
rect 35875 29800 35884 29840
rect 35924 29800 35933 29840
rect 35875 29799 35933 29800
rect 36739 29840 36797 29841
rect 36739 29800 36748 29840
rect 36788 29800 36797 29840
rect 36739 29799 36797 29800
rect 36939 29840 36981 29849
rect 36939 29800 36940 29840
rect 36980 29800 36981 29840
rect 36939 29791 36981 29800
rect 37131 29840 37173 29849
rect 37131 29800 37132 29840
rect 37172 29800 37173 29840
rect 38563 29840 38621 29841
rect 37131 29791 37173 29800
rect 37219 29825 37277 29826
rect 37219 29785 37228 29825
rect 37268 29785 37277 29825
rect 38563 29800 38572 29840
rect 38612 29800 38621 29840
rect 38563 29799 38621 29800
rect 39427 29840 39485 29841
rect 39427 29800 39436 29840
rect 39476 29800 39485 29840
rect 39427 29799 39485 29800
rect 39819 29840 39861 29849
rect 39819 29800 39820 29840
rect 39860 29800 39861 29840
rect 39819 29791 39861 29800
rect 40675 29840 40733 29841
rect 40675 29800 40684 29840
rect 40724 29800 40733 29840
rect 40675 29799 40733 29800
rect 40779 29840 40821 29849
rect 40779 29800 40780 29840
rect 40820 29800 40821 29840
rect 40779 29791 40821 29800
rect 40971 29840 41013 29849
rect 40971 29800 40972 29840
rect 41012 29800 41013 29840
rect 40971 29791 41013 29800
rect 41163 29840 41205 29849
rect 41163 29800 41164 29840
rect 41204 29800 41205 29840
rect 41163 29791 41205 29800
rect 41259 29840 41301 29849
rect 41259 29800 41260 29840
rect 41300 29800 41301 29840
rect 41259 29791 41301 29800
rect 41355 29840 41397 29849
rect 41355 29800 41356 29840
rect 41396 29800 41397 29840
rect 41355 29791 41397 29800
rect 41451 29840 41493 29849
rect 41451 29800 41452 29840
rect 41492 29800 41493 29840
rect 41451 29791 41493 29800
rect 42307 29840 42365 29841
rect 42307 29800 42316 29840
rect 42356 29800 42365 29840
rect 42307 29799 42365 29800
rect 42603 29840 42645 29849
rect 42603 29800 42604 29840
rect 42644 29800 42645 29840
rect 42603 29791 42645 29800
rect 42699 29840 42741 29849
rect 42699 29800 42700 29840
rect 42740 29800 42741 29840
rect 42699 29791 42741 29800
rect 42795 29840 42837 29849
rect 42795 29800 42796 29840
rect 42836 29800 42837 29840
rect 42795 29791 42837 29800
rect 43171 29840 43229 29841
rect 43171 29800 43180 29840
rect 43220 29800 43229 29840
rect 43171 29799 43229 29800
rect 44419 29840 44477 29841
rect 44419 29800 44428 29840
rect 44468 29800 44477 29840
rect 44419 29799 44477 29800
rect 45283 29840 45341 29841
rect 45283 29800 45292 29840
rect 45332 29800 45341 29840
rect 45283 29799 45341 29800
rect 47875 29840 47933 29841
rect 47875 29800 47884 29840
rect 47924 29800 47933 29840
rect 47875 29799 47933 29800
rect 37219 29784 37277 29785
rect 8619 29756 8661 29765
rect 8619 29716 8620 29756
rect 8660 29716 8661 29756
rect 8619 29707 8661 29716
rect 17931 29756 17973 29765
rect 17931 29716 17932 29756
rect 17972 29716 17973 29756
rect 17931 29707 17973 29716
rect 18123 29756 18165 29765
rect 18123 29716 18124 29756
rect 18164 29716 18165 29756
rect 18123 29707 18165 29716
rect 22539 29756 22581 29765
rect 22539 29716 22540 29756
rect 22580 29716 22581 29756
rect 22539 29707 22581 29716
rect 25323 29756 25365 29765
rect 25323 29716 25324 29756
rect 25364 29716 25365 29756
rect 25323 29707 25365 29716
rect 29451 29756 29493 29765
rect 29451 29716 29452 29756
rect 29492 29716 29493 29756
rect 29451 29707 29493 29716
rect 35787 29756 35829 29765
rect 35787 29716 35788 29756
rect 35828 29716 35829 29756
rect 35787 29707 35829 29716
rect 37035 29756 37077 29765
rect 37035 29716 37036 29756
rect 37076 29716 37077 29756
rect 37035 29707 37077 29716
rect 43851 29756 43893 29765
rect 43851 29716 43852 29756
rect 43892 29716 43893 29756
rect 43851 29707 43893 29716
rect 44043 29756 44085 29765
rect 44043 29716 44044 29756
rect 44084 29716 44085 29756
rect 44043 29707 44085 29716
rect 4099 29672 4157 29673
rect 4099 29632 4108 29672
rect 4148 29632 4157 29672
rect 4099 29631 4157 29632
rect 5635 29672 5693 29673
rect 5635 29632 5644 29672
rect 5684 29632 5693 29672
rect 5635 29631 5693 29632
rect 6499 29672 6557 29673
rect 6499 29632 6508 29672
rect 6548 29632 6557 29672
rect 6499 29631 6557 29632
rect 7371 29672 7413 29681
rect 7371 29632 7372 29672
rect 7412 29632 7413 29672
rect 7371 29623 7413 29632
rect 8995 29672 9053 29673
rect 8995 29632 9004 29672
rect 9044 29632 9053 29672
rect 8995 29631 9053 29632
rect 20515 29672 20573 29673
rect 20515 29632 20524 29672
rect 20564 29632 20573 29672
rect 20515 29631 20573 29632
rect 21675 29672 21717 29681
rect 21675 29632 21676 29672
rect 21716 29632 21717 29672
rect 21675 29623 21717 29632
rect 24931 29672 24989 29673
rect 24931 29632 24940 29672
rect 24980 29632 24989 29672
rect 24931 29631 24989 29632
rect 26371 29672 26429 29673
rect 26371 29632 26380 29672
rect 26420 29632 26429 29672
rect 26371 29631 26429 29632
rect 31843 29672 31901 29673
rect 31843 29632 31852 29672
rect 31892 29632 31901 29672
rect 31843 29631 31901 29632
rect 32035 29672 32093 29673
rect 32035 29632 32044 29672
rect 32084 29632 32093 29672
rect 32035 29631 32093 29632
rect 35107 29672 35165 29673
rect 35107 29632 35116 29672
rect 35156 29632 35165 29672
rect 35107 29631 35165 29632
rect 40867 29672 40925 29673
rect 40867 29632 40876 29672
rect 40916 29632 40925 29672
rect 40867 29631 40925 29632
rect 42499 29672 42557 29673
rect 42499 29632 42508 29672
rect 42548 29632 42557 29672
rect 42499 29631 42557 29632
rect 46435 29672 46493 29673
rect 46435 29632 46444 29672
rect 46484 29632 46493 29672
rect 46435 29631 46493 29632
rect 47787 29672 47829 29681
rect 47787 29632 47788 29672
rect 47828 29632 47829 29672
rect 47787 29623 47829 29632
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 3715 29336 3773 29337
rect 3715 29296 3724 29336
rect 3764 29296 3773 29336
rect 3715 29295 3773 29296
rect 7947 29336 7989 29345
rect 7947 29296 7948 29336
rect 7988 29296 7989 29336
rect 7947 29287 7989 29296
rect 11779 29336 11837 29337
rect 11779 29296 11788 29336
rect 11828 29296 11837 29336
rect 11779 29295 11837 29296
rect 16675 29336 16733 29337
rect 16675 29296 16684 29336
rect 16724 29296 16733 29336
rect 16675 29295 16733 29296
rect 18691 29336 18749 29337
rect 18691 29296 18700 29336
rect 18740 29296 18749 29336
rect 18691 29295 18749 29296
rect 23107 29336 23165 29337
rect 23107 29296 23116 29336
rect 23156 29296 23165 29336
rect 23107 29295 23165 29296
rect 26571 29336 26613 29345
rect 26571 29296 26572 29336
rect 26612 29296 26613 29336
rect 26571 29287 26613 29296
rect 34243 29336 34301 29337
rect 34243 29296 34252 29336
rect 34292 29296 34301 29336
rect 34243 29295 34301 29296
rect 43747 29336 43805 29337
rect 43747 29296 43756 29336
rect 43796 29296 43805 29336
rect 43747 29295 43805 29296
rect 48451 29336 48509 29337
rect 48451 29296 48460 29336
rect 48500 29296 48509 29336
rect 48451 29295 48509 29296
rect 1323 29252 1365 29261
rect 1323 29212 1324 29252
rect 1364 29212 1365 29252
rect 1323 29203 1365 29212
rect 3915 29252 3957 29261
rect 3915 29212 3916 29252
rect 3956 29212 3957 29252
rect 3915 29203 3957 29212
rect 4875 29252 4917 29261
rect 4875 29212 4876 29252
rect 4916 29212 4917 29252
rect 4875 29203 4917 29212
rect 8715 29252 8757 29261
rect 8715 29212 8716 29252
rect 8756 29212 8757 29252
rect 8715 29203 8757 29212
rect 16971 29252 17013 29261
rect 16971 29212 16972 29252
rect 17012 29212 17013 29252
rect 16971 29203 17013 29212
rect 23499 29252 23541 29261
rect 23499 29212 23500 29252
rect 23540 29212 23541 29252
rect 23499 29203 23541 29212
rect 25899 29252 25941 29261
rect 25899 29212 25900 29252
rect 25940 29212 25941 29252
rect 25899 29203 25941 29212
rect 26859 29252 26901 29261
rect 26859 29212 26860 29252
rect 26900 29212 26901 29252
rect 26859 29203 26901 29212
rect 30987 29252 31029 29261
rect 30987 29212 30988 29252
rect 31028 29212 31029 29252
rect 30987 29203 31029 29212
rect 31851 29252 31893 29261
rect 31851 29212 31852 29252
rect 31892 29212 31893 29252
rect 31851 29203 31893 29212
rect 40395 29252 40437 29261
rect 40395 29212 40396 29252
rect 40436 29212 40437 29252
rect 40395 29203 40437 29212
rect 1699 29168 1757 29169
rect 1699 29128 1708 29168
rect 1748 29128 1757 29168
rect 1699 29127 1757 29128
rect 2563 29168 2621 29169
rect 2563 29128 2572 29168
rect 2612 29128 2621 29168
rect 2563 29127 2621 29128
rect 4579 29168 4637 29169
rect 4579 29128 4588 29168
rect 4628 29128 4637 29168
rect 4579 29127 4637 29128
rect 5251 29168 5309 29169
rect 5251 29128 5260 29168
rect 5300 29128 5309 29168
rect 5251 29127 5309 29128
rect 6115 29168 6173 29169
rect 6115 29128 6124 29168
rect 6164 29128 6173 29168
rect 6115 29127 6173 29128
rect 8419 29168 8477 29169
rect 8419 29128 8428 29168
rect 8468 29128 8477 29168
rect 8419 29127 8477 29128
rect 9091 29168 9149 29169
rect 9091 29128 9100 29168
rect 9140 29128 9149 29168
rect 9091 29127 9149 29128
rect 9955 29168 10013 29169
rect 9955 29128 9964 29168
rect 10004 29128 10013 29168
rect 9955 29127 10013 29128
rect 12451 29168 12509 29169
rect 12451 29128 12460 29168
rect 12500 29128 12509 29168
rect 12451 29127 12509 29128
rect 13515 29168 13557 29177
rect 13515 29128 13516 29168
rect 13556 29128 13557 29168
rect 13515 29119 13557 29128
rect 13699 29168 13757 29169
rect 13699 29128 13708 29168
rect 13748 29128 13757 29168
rect 13699 29127 13757 29128
rect 14563 29168 14621 29169
rect 14563 29128 14572 29168
rect 14612 29128 14621 29168
rect 14563 29127 14621 29128
rect 14851 29168 14909 29169
rect 14851 29128 14860 29168
rect 14900 29128 14909 29168
rect 14851 29127 14909 29128
rect 16107 29168 16149 29177
rect 16107 29128 16108 29168
rect 16148 29128 16149 29168
rect 16107 29119 16149 29128
rect 16483 29168 16541 29169
rect 16483 29128 16492 29168
rect 16532 29128 16541 29168
rect 16483 29127 16541 29128
rect 16587 29168 16629 29177
rect 16587 29128 16588 29168
rect 16628 29128 16629 29168
rect 16587 29119 16629 29128
rect 16779 29168 16821 29177
rect 16779 29128 16780 29168
rect 16820 29128 16821 29168
rect 16779 29119 16821 29128
rect 17635 29168 17693 29169
rect 17635 29128 17644 29168
rect 17684 29128 17693 29168
rect 17635 29127 17693 29128
rect 17827 29168 17885 29169
rect 17827 29128 17836 29168
rect 17876 29128 17885 29168
rect 17827 29127 17885 29128
rect 19363 29168 19421 29169
rect 19363 29128 19372 29168
rect 19412 29128 19421 29168
rect 19363 29127 19421 29128
rect 19563 29168 19605 29177
rect 19563 29128 19564 29168
rect 19604 29128 19605 29168
rect 19563 29119 19605 29128
rect 19755 29168 19797 29177
rect 19755 29128 19756 29168
rect 19796 29128 19797 29168
rect 19755 29119 19797 29128
rect 19843 29168 19901 29169
rect 19843 29128 19852 29168
rect 19892 29128 19901 29168
rect 19843 29127 19901 29128
rect 20619 29168 20661 29177
rect 20619 29128 20620 29168
rect 20660 29128 20661 29168
rect 20619 29119 20661 29128
rect 21475 29168 21533 29169
rect 21475 29128 21484 29168
rect 21524 29128 21533 29168
rect 21475 29127 21533 29128
rect 22539 29168 22581 29177
rect 22539 29128 22540 29168
rect 22580 29128 22581 29168
rect 22539 29119 22581 29128
rect 22635 29168 22677 29177
rect 22635 29128 22636 29168
rect 22676 29128 22677 29168
rect 22635 29119 22677 29128
rect 22731 29168 22773 29177
rect 22731 29128 22732 29168
rect 22772 29128 22773 29168
rect 22731 29119 22773 29128
rect 22827 29168 22869 29177
rect 22827 29128 22828 29168
rect 22868 29128 22869 29168
rect 22827 29119 22869 29128
rect 23019 29168 23061 29177
rect 23019 29128 23020 29168
rect 23060 29128 23061 29168
rect 23019 29119 23061 29128
rect 23211 29168 23253 29177
rect 23211 29128 23212 29168
rect 23252 29128 23253 29168
rect 23211 29119 23253 29128
rect 23299 29168 23357 29169
rect 23299 29128 23308 29168
rect 23348 29128 23357 29168
rect 23299 29127 23357 29128
rect 24163 29168 24221 29169
rect 24163 29128 24172 29168
rect 24212 29128 24221 29168
rect 24163 29127 24221 29128
rect 24939 29168 24981 29177
rect 24939 29128 24940 29168
rect 24980 29128 24981 29168
rect 24939 29119 24981 29128
rect 25035 29168 25077 29177
rect 25035 29128 25036 29168
rect 25076 29128 25077 29168
rect 25035 29119 25077 29128
rect 25131 29168 25173 29177
rect 25131 29128 25132 29168
rect 25172 29128 25173 29168
rect 25131 29119 25173 29128
rect 25227 29168 25269 29177
rect 25227 29128 25228 29168
rect 25268 29128 25269 29168
rect 25227 29119 25269 29128
rect 25507 29168 25565 29169
rect 25507 29128 25516 29168
rect 25556 29128 25565 29168
rect 25507 29127 25565 29128
rect 25803 29168 25845 29177
rect 25803 29128 25804 29168
rect 25844 29128 25845 29168
rect 25803 29119 25845 29128
rect 26659 29168 26717 29169
rect 26659 29128 26668 29168
rect 26708 29128 26717 29168
rect 26659 29127 26717 29128
rect 27523 29168 27581 29169
rect 27523 29128 27532 29168
rect 27572 29128 27581 29168
rect 27523 29127 27581 29128
rect 27715 29168 27773 29169
rect 27715 29128 27724 29168
rect 27764 29128 27773 29168
rect 27715 29127 27773 29128
rect 28107 29168 28149 29177
rect 28107 29128 28108 29168
rect 28148 29128 28149 29168
rect 28107 29119 28149 29128
rect 28203 29168 28245 29177
rect 28203 29128 28204 29168
rect 28244 29128 28245 29168
rect 28203 29119 28245 29128
rect 28299 29168 28341 29177
rect 28299 29128 28300 29168
rect 28340 29128 28341 29168
rect 28299 29119 28341 29128
rect 28395 29168 28437 29177
rect 28395 29128 28396 29168
rect 28436 29128 28437 29168
rect 28395 29119 28437 29128
rect 29251 29168 29309 29169
rect 29251 29128 29260 29168
rect 29300 29128 29309 29168
rect 29251 29127 29309 29128
rect 29443 29168 29501 29169
rect 29443 29128 29452 29168
rect 29492 29128 29501 29168
rect 29443 29127 29501 29128
rect 30403 29168 30461 29169
rect 30403 29128 30412 29168
rect 30452 29128 30461 29168
rect 30403 29127 30461 29128
rect 31083 29168 31125 29177
rect 31083 29128 31084 29168
rect 31124 29128 31125 29168
rect 31083 29119 31125 29128
rect 31363 29168 31421 29169
rect 31363 29128 31372 29168
rect 31412 29128 31421 29168
rect 31363 29127 31421 29128
rect 32227 29168 32285 29169
rect 32227 29128 32236 29168
rect 32276 29128 32285 29168
rect 32227 29127 32285 29128
rect 33091 29168 33149 29169
rect 33091 29128 33100 29168
rect 33140 29128 33149 29168
rect 33091 29127 33149 29128
rect 34435 29168 34493 29169
rect 34435 29128 34444 29168
rect 34484 29128 34493 29168
rect 34435 29127 34493 29128
rect 35683 29168 35741 29169
rect 35683 29128 35692 29168
rect 35732 29128 35741 29168
rect 35683 29127 35741 29128
rect 36547 29168 36605 29169
rect 36547 29128 36556 29168
rect 36596 29128 36605 29168
rect 36547 29127 36605 29128
rect 36939 29168 36981 29177
rect 36939 29128 36940 29168
rect 36980 29128 36981 29168
rect 36939 29119 36981 29128
rect 37227 29168 37269 29177
rect 37227 29128 37228 29168
rect 37268 29128 37269 29168
rect 37227 29119 37269 29128
rect 37323 29168 37365 29177
rect 37323 29128 37324 29168
rect 37364 29128 37365 29168
rect 37323 29119 37365 29128
rect 37419 29168 37461 29177
rect 37419 29128 37420 29168
rect 37460 29128 37461 29168
rect 37419 29119 37461 29128
rect 37515 29168 37557 29177
rect 37515 29128 37516 29168
rect 37556 29128 37557 29168
rect 37515 29119 37557 29128
rect 39523 29168 39581 29169
rect 39523 29128 39532 29168
rect 39572 29128 39581 29168
rect 39523 29127 39581 29128
rect 40771 29168 40829 29169
rect 40771 29128 40780 29168
rect 40820 29128 40829 29168
rect 40771 29127 40829 29128
rect 41635 29168 41693 29169
rect 41635 29128 41644 29168
rect 41684 29128 41693 29168
rect 41635 29127 41693 29128
rect 43075 29168 43133 29169
rect 43075 29128 43084 29168
rect 43124 29128 43133 29168
rect 43075 29127 43133 29128
rect 44043 29168 44085 29177
rect 44043 29128 44044 29168
rect 44084 29128 44085 29168
rect 44043 29119 44085 29128
rect 44139 29168 44181 29177
rect 44139 29128 44140 29168
rect 44180 29128 44181 29168
rect 44139 29119 44181 29128
rect 44235 29168 44277 29177
rect 44235 29128 44236 29168
rect 44276 29128 44277 29168
rect 44235 29119 44277 29128
rect 44331 29168 44373 29177
rect 44331 29128 44332 29168
rect 44372 29128 44373 29168
rect 44331 29119 44373 29128
rect 45475 29168 45533 29169
rect 45475 29128 45484 29168
rect 45524 29128 45533 29168
rect 45475 29127 45533 29128
rect 45867 29168 45909 29177
rect 45867 29128 45868 29168
rect 45908 29128 45909 29168
rect 45867 29119 45909 29128
rect 46243 29168 46301 29169
rect 46243 29128 46252 29168
rect 46292 29128 46301 29168
rect 46243 29127 46301 29128
rect 47107 29168 47165 29169
rect 47107 29128 47116 29168
rect 47156 29128 47165 29168
rect 47107 29127 47165 29128
rect 49123 29168 49181 29169
rect 49123 29128 49132 29168
rect 49172 29128 49181 29168
rect 49123 29127 49181 29128
rect 7275 29084 7317 29093
rect 7275 29044 7276 29084
rect 7316 29044 7317 29084
rect 7275 29035 7317 29044
rect 27819 29084 27861 29093
rect 27819 29044 27820 29084
rect 27860 29044 27861 29084
rect 27819 29035 27861 29044
rect 29163 29084 29205 29093
rect 29163 29044 29164 29084
rect 29204 29044 29205 29084
rect 29163 29035 29205 29044
rect 48267 29084 48309 29093
rect 48267 29044 48268 29084
rect 48308 29044 48309 29084
rect 48267 29035 48309 29044
rect 1131 29000 1173 29009
rect 1131 28960 1132 29000
rect 1172 28960 1173 29000
rect 1131 28951 1173 28960
rect 15915 29000 15957 29009
rect 15915 28960 15916 29000
rect 15956 28960 15957 29000
rect 15915 28951 15957 28960
rect 24747 29000 24789 29009
rect 24747 28960 24748 29000
rect 24788 28960 24789 29000
rect 24747 28951 24789 28960
rect 30691 29000 30749 29001
rect 30691 28960 30700 29000
rect 30740 28960 30749 29000
rect 30691 28959 30749 28960
rect 38091 29000 38133 29009
rect 38091 28960 38092 29000
rect 38132 28960 38133 29000
rect 38091 28951 38133 28960
rect 40195 29000 40253 29001
rect 40195 28960 40204 29000
rect 40244 28960 40253 29000
rect 40195 28959 40253 28960
rect 42787 29000 42845 29001
rect 42787 28960 42796 29000
rect 42836 28960 42845 29000
rect 42787 28959 42845 28960
rect 45195 29000 45237 29009
rect 45195 28960 45196 29000
rect 45236 28960 45237 29000
rect 45195 28951 45237 28960
rect 11107 28916 11165 28917
rect 11107 28876 11116 28916
rect 11156 28876 11165 28916
rect 11107 28875 11165 28876
rect 13611 28916 13653 28925
rect 13611 28876 13612 28916
rect 13652 28876 13653 28916
rect 13611 28867 13653 28876
rect 14475 28916 14517 28925
rect 14475 28876 14476 28916
rect 14516 28876 14517 28916
rect 14475 28867 14517 28876
rect 14763 28916 14805 28925
rect 14763 28876 14764 28916
rect 14804 28876 14805 28916
rect 14763 28867 14805 28876
rect 18499 28916 18557 28917
rect 18499 28876 18508 28916
rect 18548 28876 18557 28916
rect 18499 28875 18557 28876
rect 19563 28916 19605 28925
rect 19563 28876 19564 28916
rect 19604 28876 19605 28916
rect 19563 28867 19605 28876
rect 20811 28916 20853 28925
rect 20811 28876 20812 28916
rect 20852 28876 20853 28916
rect 20811 28867 20853 28876
rect 26179 28916 26237 28917
rect 26179 28876 26188 28916
rect 26228 28876 26237 28916
rect 26179 28875 26237 28876
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 2571 28580 2613 28589
rect 2571 28540 2572 28580
rect 2612 28540 2613 28580
rect 2571 28531 2613 28540
rect 3531 28580 3573 28589
rect 3531 28540 3532 28580
rect 3572 28540 3573 28580
rect 3531 28531 3573 28540
rect 6123 28580 6165 28589
rect 6123 28540 6124 28580
rect 6164 28540 6165 28580
rect 6123 28531 6165 28540
rect 15243 28580 15285 28589
rect 15243 28540 15244 28580
rect 15284 28540 15285 28580
rect 15243 28531 15285 28540
rect 18403 28580 18461 28581
rect 18403 28540 18412 28580
rect 18452 28540 18461 28580
rect 18403 28539 18461 28540
rect 18603 28580 18645 28589
rect 18603 28540 18604 28580
rect 18644 28540 18645 28580
rect 18603 28531 18645 28540
rect 22243 28580 22301 28581
rect 22243 28540 22252 28580
rect 22292 28540 22301 28580
rect 22243 28539 22301 28540
rect 26851 28580 26909 28581
rect 26851 28540 26860 28580
rect 26900 28540 26909 28580
rect 26851 28539 26909 28540
rect 30595 28580 30653 28581
rect 30595 28540 30604 28580
rect 30644 28540 30653 28580
rect 30595 28539 30653 28540
rect 32523 28580 32565 28589
rect 32523 28540 32524 28580
rect 32564 28540 32565 28580
rect 32523 28531 32565 28540
rect 35115 28580 35157 28589
rect 35115 28540 35116 28580
rect 35156 28540 35157 28580
rect 35115 28531 35157 28540
rect 37035 28580 37077 28589
rect 37035 28540 37036 28580
rect 37076 28540 37077 28580
rect 37035 28531 37077 28540
rect 40779 28580 40821 28589
rect 40779 28540 40780 28580
rect 40820 28540 40821 28580
rect 40779 28531 40821 28540
rect 43179 28580 43221 28589
rect 43179 28540 43180 28580
rect 43220 28540 43221 28580
rect 43179 28531 43221 28540
rect 1707 28496 1749 28505
rect 1707 28456 1708 28496
rect 1748 28456 1749 28496
rect 1707 28447 1749 28456
rect 13611 28496 13653 28505
rect 13611 28456 13612 28496
rect 13652 28456 13653 28496
rect 13611 28447 13653 28456
rect 23499 28496 23541 28505
rect 23499 28456 23500 28496
rect 23540 28456 23541 28496
rect 23499 28447 23541 28456
rect 32907 28496 32949 28505
rect 32907 28456 32908 28496
rect 32948 28456 32949 28496
rect 32907 28447 32949 28456
rect 33387 28496 33429 28505
rect 33387 28456 33388 28496
rect 33428 28456 33429 28496
rect 33387 28447 33429 28456
rect 37707 28496 37749 28505
rect 37707 28456 37708 28496
rect 37748 28456 37749 28496
rect 37707 28447 37749 28456
rect 41827 28496 41885 28497
rect 41827 28456 41836 28496
rect 41876 28456 41885 28496
rect 41827 28455 41885 28456
rect 45579 28496 45621 28505
rect 45579 28456 45580 28496
rect 45620 28456 45621 28496
rect 45579 28447 45621 28456
rect 48747 28496 48789 28505
rect 48747 28456 48748 28496
rect 48788 28456 48789 28496
rect 48747 28447 48789 28456
rect 49227 28496 49269 28505
rect 49227 28456 49228 28496
rect 49268 28456 49269 28496
rect 49227 28447 49269 28456
rect 7851 28412 7893 28421
rect 7851 28372 7852 28412
rect 7892 28372 7893 28412
rect 7851 28363 7893 28372
rect 30219 28412 30261 28421
rect 30219 28372 30220 28412
rect 30260 28372 30261 28412
rect 30219 28363 30261 28372
rect 44139 28373 44181 28382
rect 2659 28328 2717 28329
rect 2659 28288 2668 28328
rect 2708 28288 2717 28328
rect 2659 28287 2717 28288
rect 2851 28328 2909 28329
rect 2851 28288 2860 28328
rect 2900 28288 2909 28328
rect 2851 28287 2909 28288
rect 3811 28328 3869 28329
rect 3811 28288 3820 28328
rect 3860 28288 3869 28328
rect 3811 28287 3869 28288
rect 4771 28328 4829 28329
rect 4771 28288 4780 28328
rect 4820 28288 4829 28328
rect 4771 28287 4829 28288
rect 4971 28328 5013 28337
rect 4971 28288 4972 28328
rect 5012 28288 5013 28328
rect 4971 28279 5013 28288
rect 5067 28328 5109 28337
rect 5067 28288 5068 28328
rect 5108 28288 5109 28328
rect 5067 28279 5109 28288
rect 5163 28328 5205 28337
rect 5163 28288 5164 28328
rect 5204 28288 5205 28328
rect 5163 28279 5205 28288
rect 5443 28328 5501 28329
rect 5443 28288 5452 28328
rect 5492 28288 5501 28328
rect 5443 28287 5501 28288
rect 5827 28328 5885 28329
rect 5827 28288 5836 28328
rect 5876 28288 5885 28328
rect 5827 28287 5885 28288
rect 6123 28328 6165 28337
rect 6123 28288 6124 28328
rect 6164 28288 6165 28328
rect 6123 28279 6165 28288
rect 6315 28328 6357 28337
rect 6315 28288 6316 28328
rect 6356 28288 6357 28328
rect 6315 28279 6357 28288
rect 6403 28328 6461 28329
rect 6403 28288 6412 28328
rect 6452 28288 6461 28328
rect 6403 28287 6461 28288
rect 7555 28328 7613 28329
rect 7555 28288 7564 28328
rect 7604 28288 7613 28328
rect 7555 28287 7613 28288
rect 8515 28328 8573 28329
rect 8515 28288 8524 28328
rect 8564 28288 8573 28328
rect 8515 28287 8573 28288
rect 8707 28328 8765 28329
rect 8707 28288 8716 28328
rect 8756 28288 8765 28328
rect 8707 28287 8765 28288
rect 10339 28328 10397 28329
rect 10339 28288 10348 28328
rect 10388 28288 10397 28328
rect 10339 28287 10397 28288
rect 11683 28328 11741 28329
rect 11683 28288 11692 28328
rect 11732 28288 11741 28328
rect 11683 28287 11741 28288
rect 12547 28328 12605 28329
rect 12547 28288 12556 28328
rect 12596 28288 12605 28328
rect 12547 28287 12605 28288
rect 14187 28328 14229 28337
rect 14187 28288 14188 28328
rect 14228 28288 14229 28328
rect 14187 28279 14229 28288
rect 15715 28328 15773 28329
rect 15715 28288 15724 28328
rect 15764 28288 15773 28328
rect 15715 28287 15773 28288
rect 16387 28328 16445 28329
rect 16387 28288 16396 28328
rect 16436 28288 16445 28328
rect 16387 28287 16445 28288
rect 17251 28328 17309 28329
rect 17251 28288 17260 28328
rect 17300 28288 17309 28328
rect 17251 28287 17309 28288
rect 18691 28328 18749 28329
rect 18691 28288 18700 28328
rect 18740 28288 18749 28328
rect 18691 28287 18749 28288
rect 18979 28328 19037 28329
rect 18979 28288 18988 28328
rect 19028 28288 19037 28328
rect 18979 28287 19037 28288
rect 20227 28328 20285 28329
rect 20227 28288 20236 28328
rect 20276 28288 20285 28328
rect 20227 28287 20285 28288
rect 21091 28328 21149 28329
rect 21091 28288 21100 28328
rect 21140 28288 21149 28328
rect 21091 28287 21149 28288
rect 24835 28328 24893 28329
rect 24835 28288 24844 28328
rect 24884 28288 24893 28328
rect 24835 28287 24893 28288
rect 25699 28328 25757 28329
rect 25699 28288 25708 28328
rect 25748 28288 25757 28328
rect 25699 28287 25757 28288
rect 27331 28328 27389 28329
rect 27331 28288 27340 28328
rect 27380 28288 27389 28328
rect 27331 28287 27389 28288
rect 27435 28328 27477 28337
rect 27435 28288 27436 28328
rect 27476 28288 27477 28328
rect 27435 28279 27477 28288
rect 27627 28328 27669 28337
rect 27627 28288 27628 28328
rect 27668 28288 27669 28328
rect 27627 28279 27669 28288
rect 28195 28328 28253 28329
rect 28195 28288 28204 28328
rect 28244 28288 28253 28328
rect 28195 28287 28253 28288
rect 29059 28328 29117 28329
rect 29059 28288 29068 28328
rect 29108 28288 29117 28328
rect 29059 28287 29117 28288
rect 31267 28328 31325 28329
rect 31267 28288 31276 28328
rect 31316 28288 31325 28328
rect 31267 28287 31325 28288
rect 31459 28328 31517 28329
rect 31459 28288 31468 28328
rect 31508 28288 31517 28328
rect 31459 28287 31517 28288
rect 31563 28328 31605 28337
rect 31563 28288 31564 28328
rect 31604 28288 31605 28328
rect 31563 28279 31605 28288
rect 31755 28328 31797 28337
rect 31755 28288 31756 28328
rect 31796 28288 31797 28328
rect 31755 28279 31797 28288
rect 31947 28328 31989 28337
rect 31947 28288 31948 28328
rect 31988 28288 31989 28328
rect 31947 28279 31989 28288
rect 32043 28328 32085 28337
rect 32043 28288 32044 28328
rect 32084 28288 32085 28328
rect 32043 28279 32085 28288
rect 32139 28328 32181 28337
rect 32139 28288 32140 28328
rect 32180 28288 32181 28328
rect 32139 28279 32181 28288
rect 32235 28328 32277 28337
rect 32235 28288 32236 28328
rect 32276 28288 32277 28328
rect 32235 28279 32277 28288
rect 32419 28328 32477 28329
rect 32419 28288 32428 28328
rect 32468 28288 32477 28328
rect 33195 28328 33237 28337
rect 32419 28287 32477 28288
rect 33091 28313 33149 28314
rect 33091 28273 33100 28313
rect 33140 28273 33149 28313
rect 33195 28288 33196 28328
rect 33236 28288 33237 28328
rect 33195 28279 33237 28288
rect 33387 28328 33429 28337
rect 33387 28288 33388 28328
rect 33428 28288 33429 28328
rect 33387 28279 33429 28288
rect 33571 28328 33629 28329
rect 33571 28288 33580 28328
rect 33620 28288 33629 28328
rect 33571 28287 33629 28288
rect 34435 28328 34493 28329
rect 34435 28288 34444 28328
rect 34484 28288 34493 28328
rect 34435 28287 34493 28288
rect 35395 28328 35453 28329
rect 35395 28288 35404 28328
rect 35444 28288 35453 28328
rect 35395 28287 35453 28288
rect 35683 28328 35741 28329
rect 35683 28288 35692 28328
rect 35732 28288 35741 28328
rect 35683 28287 35741 28288
rect 35875 28328 35933 28329
rect 35875 28288 35884 28328
rect 35924 28288 35933 28328
rect 35875 28287 35933 28288
rect 36835 28328 36893 28329
rect 36835 28288 36844 28328
rect 36884 28288 36893 28328
rect 36835 28287 36893 28288
rect 37123 28328 37181 28329
rect 37123 28288 37132 28328
rect 37172 28288 37181 28328
rect 37123 28287 37181 28288
rect 38371 28328 38429 28329
rect 38371 28288 38380 28328
rect 38420 28288 38429 28328
rect 38371 28287 38429 28288
rect 40291 28328 40349 28329
rect 40291 28288 40300 28328
rect 40340 28288 40349 28328
rect 40291 28287 40349 28288
rect 40483 28328 40541 28329
rect 40483 28288 40492 28328
rect 40532 28288 40541 28328
rect 40483 28287 40541 28288
rect 40587 28328 40629 28337
rect 40587 28288 40588 28328
rect 40628 28288 40629 28328
rect 40587 28279 40629 28288
rect 40779 28328 40821 28337
rect 40779 28288 40780 28328
rect 40820 28288 40821 28328
rect 40779 28279 40821 28288
rect 40963 28328 41021 28329
rect 40963 28288 40972 28328
rect 41012 28288 41021 28328
rect 40963 28287 41021 28288
rect 42123 28328 42165 28337
rect 42123 28288 42124 28328
rect 42164 28288 42165 28328
rect 42123 28279 42165 28288
rect 42219 28328 42261 28337
rect 42219 28288 42220 28328
rect 42260 28288 42261 28328
rect 42219 28279 42261 28288
rect 42499 28328 42557 28329
rect 42499 28288 42508 28328
rect 42548 28288 42557 28328
rect 42499 28287 42557 28288
rect 42883 28328 42941 28329
rect 42883 28288 42892 28328
rect 42932 28288 42941 28328
rect 42883 28287 42941 28288
rect 42987 28328 43029 28337
rect 42987 28288 42988 28328
rect 43028 28288 43029 28328
rect 42987 28279 43029 28288
rect 43179 28328 43221 28337
rect 43179 28288 43180 28328
rect 43220 28288 43221 28328
rect 43179 28279 43221 28288
rect 43363 28328 43421 28329
rect 43363 28288 43372 28328
rect 43412 28288 43421 28328
rect 43363 28287 43421 28288
rect 43467 28328 43509 28337
rect 43467 28288 43468 28328
rect 43508 28288 43509 28328
rect 43467 28279 43509 28288
rect 43659 28328 43701 28337
rect 43659 28288 43660 28328
rect 43700 28288 43701 28328
rect 43659 28279 43701 28288
rect 43851 28328 43893 28337
rect 43851 28288 43852 28328
rect 43892 28288 43893 28328
rect 43851 28279 43893 28288
rect 43947 28328 43989 28337
rect 43947 28288 43948 28328
rect 43988 28288 43989 28328
rect 43947 28279 43989 28288
rect 44043 28328 44085 28337
rect 44043 28288 44044 28328
rect 44084 28288 44085 28328
rect 44139 28333 44140 28373
rect 44180 28333 44181 28373
rect 44139 28324 44181 28333
rect 44323 28328 44381 28329
rect 44043 28279 44085 28288
rect 44323 28288 44332 28328
rect 44372 28288 44381 28328
rect 44323 28287 44381 28288
rect 45195 28328 45237 28337
rect 45195 28288 45196 28328
rect 45236 28288 45237 28328
rect 45195 28279 45237 28288
rect 46147 28328 46205 28329
rect 46147 28288 46156 28328
rect 46196 28288 46205 28328
rect 46147 28287 46205 28288
rect 46443 28328 46485 28337
rect 46443 28288 46444 28328
rect 46484 28288 46485 28328
rect 46443 28279 46485 28288
rect 47107 28328 47165 28329
rect 47107 28288 47116 28328
rect 47156 28288 47165 28328
rect 47107 28287 47165 28288
rect 47403 28328 47445 28337
rect 47403 28288 47404 28328
rect 47444 28288 47445 28328
rect 47403 28279 47445 28288
rect 47499 28328 47541 28337
rect 47499 28288 47500 28328
rect 47540 28288 47541 28328
rect 47499 28279 47541 28288
rect 47595 28328 47637 28337
rect 47595 28288 47596 28328
rect 47636 28288 47637 28328
rect 47595 28279 47637 28288
rect 47691 28328 47733 28337
rect 47691 28288 47692 28328
rect 47732 28288 47733 28328
rect 47691 28279 47733 28288
rect 48547 28328 48605 28329
rect 48547 28288 48556 28328
rect 48596 28288 48605 28328
rect 48547 28287 48605 28288
rect 48747 28328 48789 28337
rect 48747 28288 48748 28328
rect 48788 28288 48789 28328
rect 48747 28279 48789 28288
rect 48939 28328 48981 28337
rect 48939 28288 48940 28328
rect 48980 28288 48981 28328
rect 48939 28279 48981 28288
rect 49027 28328 49085 28329
rect 49027 28288 49036 28328
rect 49076 28288 49085 28328
rect 49027 28287 49085 28288
rect 50563 28328 50621 28329
rect 50563 28288 50572 28328
rect 50612 28288 50621 28328
rect 50563 28287 50621 28288
rect 33091 28272 33149 28273
rect 6691 28244 6749 28245
rect 6691 28204 6700 28244
rect 6740 28204 6749 28244
rect 6691 28203 6749 28204
rect 12939 28244 12981 28253
rect 12939 28204 12940 28244
rect 12980 28204 12981 28244
rect 12939 28195 12981 28204
rect 16011 28244 16053 28253
rect 16011 28204 16012 28244
rect 16052 28204 16053 28244
rect 16011 28195 16053 28204
rect 19659 28244 19701 28253
rect 19659 28204 19660 28244
rect 19700 28204 19701 28244
rect 19659 28195 19701 28204
rect 19851 28244 19893 28253
rect 19851 28204 19852 28244
rect 19892 28204 19893 28244
rect 19851 28195 19893 28204
rect 24459 28244 24501 28253
rect 24459 28204 24460 28244
rect 24500 28204 24501 28244
rect 24459 28195 24501 28204
rect 27819 28244 27861 28253
rect 27819 28204 27820 28244
rect 27860 28204 27861 28244
rect 27819 28195 27861 28204
rect 39235 28244 39293 28245
rect 39235 28204 39244 28244
rect 39284 28204 39293 28244
rect 39235 28203 39293 28204
rect 43563 28244 43605 28253
rect 43563 28204 43564 28244
rect 43604 28204 43605 28244
rect 43563 28195 43605 28204
rect 4099 28160 4157 28161
rect 4099 28120 4108 28160
rect 4148 28120 4157 28160
rect 4099 28119 4157 28120
rect 5251 28160 5309 28161
rect 5251 28120 5260 28160
rect 5300 28120 5309 28160
rect 5251 28119 5309 28120
rect 5547 28160 5589 28169
rect 5547 28120 5548 28160
rect 5588 28120 5589 28160
rect 5547 28111 5589 28120
rect 5739 28160 5781 28169
rect 5739 28120 5740 28160
rect 5780 28120 5781 28160
rect 5739 28111 5781 28120
rect 9379 28160 9437 28161
rect 9379 28120 9388 28160
rect 9428 28120 9437 28160
rect 9379 28119 9437 28120
rect 9667 28160 9725 28161
rect 9667 28120 9676 28160
rect 9716 28120 9725 28160
rect 9667 28119 9725 28120
rect 10531 28160 10589 28161
rect 10531 28120 10540 28160
rect 10580 28120 10589 28160
rect 10531 28119 10589 28120
rect 27523 28160 27581 28161
rect 27523 28120 27532 28160
rect 27572 28120 27581 28160
rect 27523 28119 27581 28120
rect 31651 28160 31709 28161
rect 31651 28120 31660 28160
rect 31700 28120 31709 28160
rect 31651 28119 31709 28120
rect 34243 28160 34301 28161
rect 34243 28120 34252 28160
rect 34292 28120 34301 28160
rect 34243 28119 34301 28120
rect 36163 28160 36221 28161
rect 36163 28120 36172 28160
rect 36212 28120 36221 28160
rect 36163 28119 36221 28120
rect 39619 28160 39677 28161
rect 39619 28120 39628 28160
rect 39668 28120 39677 28160
rect 39619 28119 39677 28120
rect 41635 28160 41693 28161
rect 41635 28120 41644 28160
rect 41684 28120 41693 28160
rect 41635 28119 41693 28120
rect 46059 28160 46101 28169
rect 46059 28120 46060 28160
rect 46100 28120 46101 28160
rect 46059 28111 46101 28120
rect 47875 28160 47933 28161
rect 47875 28120 47884 28160
rect 47924 28120 47933 28160
rect 47875 28119 47933 28120
rect 49891 28160 49949 28161
rect 49891 28120 49900 28160
rect 49940 28120 49949 28160
rect 49891 28119 49949 28120
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 23595 27824 23637 27833
rect 23595 27784 23596 27824
rect 23636 27784 23637 27824
rect 23595 27775 23637 27784
rect 33667 27824 33725 27825
rect 33667 27784 33676 27824
rect 33716 27784 33725 27824
rect 33667 27783 33725 27784
rect 5251 27740 5309 27741
rect 5251 27700 5260 27740
rect 5300 27700 5309 27740
rect 5251 27699 5309 27700
rect 9675 27740 9717 27749
rect 9675 27700 9676 27740
rect 9716 27700 9717 27740
rect 9675 27691 9717 27700
rect 11595 27740 11637 27749
rect 11595 27700 11596 27740
rect 11636 27700 11637 27740
rect 11595 27691 11637 27700
rect 15339 27740 15381 27749
rect 15339 27700 15340 27740
rect 15380 27700 15381 27740
rect 15339 27691 15381 27700
rect 17451 27740 17493 27749
rect 17451 27700 17452 27740
rect 17492 27700 17493 27740
rect 17451 27691 17493 27700
rect 20715 27740 20757 27749
rect 20715 27700 20716 27740
rect 20756 27700 20757 27740
rect 20715 27691 20757 27700
rect 25995 27740 26037 27749
rect 25995 27700 25996 27740
rect 26036 27700 26037 27740
rect 25995 27691 26037 27700
rect 29835 27740 29877 27749
rect 29835 27700 29836 27740
rect 29876 27700 29877 27740
rect 29835 27691 29877 27700
rect 31275 27740 31317 27749
rect 31275 27700 31276 27740
rect 31316 27700 31317 27740
rect 31275 27691 31317 27700
rect 34155 27740 34197 27749
rect 34155 27700 34156 27740
rect 34196 27700 34197 27740
rect 34155 27691 34197 27700
rect 39531 27740 39573 27749
rect 39531 27700 39532 27740
rect 39572 27700 39573 27740
rect 39531 27691 39573 27700
rect 42219 27740 42261 27749
rect 42219 27700 42220 27740
rect 42260 27700 42261 27740
rect 42219 27691 42261 27700
rect 47883 27740 47925 27749
rect 47883 27700 47884 27740
rect 47924 27700 47925 27740
rect 47883 27691 47925 27700
rect 1227 27656 1269 27665
rect 1227 27616 1228 27656
rect 1268 27616 1269 27656
rect 1227 27607 1269 27616
rect 1603 27656 1661 27657
rect 1603 27616 1612 27656
rect 1652 27616 1661 27656
rect 1603 27615 1661 27616
rect 2467 27656 2525 27657
rect 2467 27616 2476 27656
rect 2516 27616 2525 27656
rect 2467 27615 2525 27616
rect 3811 27656 3869 27657
rect 3811 27616 3820 27656
rect 3860 27616 3869 27656
rect 3811 27615 3869 27616
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4107 27656 4149 27665
rect 4107 27616 4108 27656
rect 4148 27616 4149 27656
rect 4107 27607 4149 27616
rect 4491 27656 4533 27665
rect 4491 27616 4492 27656
rect 4532 27616 4533 27656
rect 4491 27607 4533 27616
rect 5635 27656 5693 27657
rect 5635 27616 5644 27656
rect 5684 27616 5693 27656
rect 5635 27615 5693 27616
rect 5931 27656 5973 27665
rect 5931 27616 5932 27656
rect 5972 27616 5973 27656
rect 5931 27607 5973 27616
rect 6027 27656 6069 27665
rect 6027 27616 6028 27656
rect 6068 27616 6069 27656
rect 6027 27607 6069 27616
rect 6595 27656 6653 27657
rect 6595 27616 6604 27656
rect 6644 27616 6653 27656
rect 6595 27615 6653 27616
rect 6795 27656 6837 27665
rect 6795 27616 6796 27656
rect 6836 27616 6837 27656
rect 6795 27607 6837 27616
rect 6891 27656 6933 27665
rect 6891 27616 6892 27656
rect 6932 27616 6933 27656
rect 6891 27607 6933 27616
rect 6987 27656 7029 27665
rect 6987 27616 6988 27656
rect 7028 27616 7029 27656
rect 6987 27607 7029 27616
rect 7083 27656 7125 27665
rect 7083 27616 7084 27656
rect 7124 27616 7125 27656
rect 7083 27607 7125 27616
rect 8419 27656 8477 27657
rect 8419 27616 8428 27656
rect 8468 27616 8477 27656
rect 8419 27615 8477 27616
rect 9283 27656 9341 27657
rect 9283 27616 9292 27656
rect 9332 27616 9341 27656
rect 9283 27615 9341 27616
rect 10915 27656 10973 27657
rect 10915 27616 10924 27656
rect 10964 27616 10973 27656
rect 10915 27615 10973 27616
rect 11203 27656 11261 27657
rect 11203 27616 11212 27656
rect 11252 27616 11261 27656
rect 11203 27615 11261 27616
rect 11499 27656 11541 27665
rect 11499 27616 11500 27656
rect 11540 27616 11541 27656
rect 11499 27607 11541 27616
rect 12067 27656 12125 27657
rect 12067 27616 12076 27656
rect 12116 27616 12125 27656
rect 12067 27615 12125 27616
rect 13027 27656 13085 27657
rect 13027 27616 13036 27656
rect 13076 27616 13085 27656
rect 13027 27615 13085 27616
rect 13315 27656 13373 27657
rect 13315 27616 13324 27656
rect 13364 27616 13373 27656
rect 13315 27615 13373 27616
rect 14187 27656 14229 27665
rect 14187 27616 14188 27656
rect 14228 27616 14229 27656
rect 14187 27607 14229 27616
rect 14571 27656 14613 27665
rect 14571 27616 14572 27656
rect 14612 27616 14613 27656
rect 14571 27607 14613 27616
rect 14763 27656 14805 27665
rect 14763 27616 14764 27656
rect 14804 27616 14805 27656
rect 14763 27607 14805 27616
rect 14851 27656 14909 27657
rect 14851 27616 14860 27656
rect 14900 27616 14909 27656
rect 14851 27615 14909 27616
rect 15435 27656 15477 27665
rect 15435 27616 15436 27656
rect 15476 27616 15477 27656
rect 15435 27607 15477 27616
rect 15715 27656 15773 27657
rect 15715 27616 15724 27656
rect 15764 27616 15773 27656
rect 15715 27615 15773 27616
rect 17355 27656 17397 27665
rect 17355 27616 17356 27656
rect 17396 27616 17397 27656
rect 17355 27607 17397 27616
rect 17547 27656 17589 27665
rect 17547 27616 17548 27656
rect 17588 27616 17589 27656
rect 17547 27607 17589 27616
rect 17635 27656 17693 27657
rect 17635 27616 17644 27656
rect 17684 27616 17693 27656
rect 17635 27615 17693 27616
rect 18123 27656 18165 27665
rect 18123 27616 18124 27656
rect 18164 27616 18165 27656
rect 18123 27607 18165 27616
rect 18219 27656 18261 27665
rect 18219 27616 18220 27656
rect 18260 27616 18261 27656
rect 18219 27607 18261 27616
rect 18499 27656 18557 27657
rect 18499 27616 18508 27656
rect 18548 27616 18557 27656
rect 18499 27615 18557 27616
rect 18795 27656 18837 27665
rect 18795 27616 18796 27656
rect 18836 27616 18837 27656
rect 18795 27607 18837 27616
rect 18891 27656 18933 27665
rect 18891 27616 18892 27656
rect 18932 27616 18933 27656
rect 18891 27607 18933 27616
rect 18987 27656 19029 27665
rect 18987 27616 18988 27656
rect 19028 27616 19029 27656
rect 18987 27607 19029 27616
rect 19083 27656 19125 27665
rect 19083 27616 19084 27656
rect 19124 27616 19125 27656
rect 19083 27607 19125 27616
rect 19555 27656 19613 27657
rect 19555 27616 19564 27656
rect 19604 27616 19613 27656
rect 19555 27615 19613 27616
rect 20515 27656 20573 27657
rect 20515 27616 20524 27656
rect 20564 27616 20573 27656
rect 20515 27615 20573 27616
rect 20803 27656 20861 27657
rect 20803 27616 20812 27656
rect 20852 27616 20861 27656
rect 20803 27615 20861 27616
rect 21003 27656 21045 27665
rect 21003 27616 21004 27656
rect 21044 27616 21045 27656
rect 21003 27607 21045 27616
rect 21667 27656 21725 27657
rect 21667 27616 21676 27656
rect 21716 27616 21725 27656
rect 21667 27615 21725 27616
rect 21859 27656 21917 27657
rect 21859 27616 21868 27656
rect 21908 27616 21917 27656
rect 21859 27615 21917 27616
rect 22819 27656 22877 27657
rect 22819 27616 22828 27656
rect 22868 27616 22877 27656
rect 22819 27615 22877 27616
rect 23979 27656 24021 27665
rect 23979 27616 23980 27656
rect 24020 27616 24021 27656
rect 23979 27607 24021 27616
rect 24747 27656 24789 27665
rect 24747 27616 24748 27656
rect 24788 27616 24789 27656
rect 24747 27607 24789 27616
rect 24835 27656 24893 27657
rect 24835 27616 24844 27656
rect 24884 27616 24893 27656
rect 24835 27615 24893 27616
rect 25035 27656 25077 27665
rect 25035 27616 25036 27656
rect 25076 27616 25077 27656
rect 25035 27607 25077 27616
rect 25227 27656 25269 27665
rect 25227 27616 25228 27656
rect 25268 27616 25269 27656
rect 25227 27607 25269 27616
rect 25315 27656 25373 27657
rect 25315 27616 25324 27656
rect 25364 27616 25373 27656
rect 25315 27615 25373 27616
rect 25603 27656 25661 27657
rect 25603 27616 25612 27656
rect 25652 27616 25661 27656
rect 25603 27615 25661 27616
rect 25899 27656 25941 27665
rect 25899 27616 25900 27656
rect 25940 27616 25941 27656
rect 25899 27607 25941 27616
rect 27811 27656 27869 27657
rect 27811 27616 27820 27656
rect 27860 27616 27869 27656
rect 27811 27615 27869 27616
rect 27915 27656 27957 27665
rect 27915 27616 27916 27656
rect 27956 27616 27957 27656
rect 27915 27607 27957 27616
rect 28107 27656 28149 27665
rect 28107 27616 28108 27656
rect 28148 27616 28149 27656
rect 28107 27607 28149 27616
rect 29731 27656 29789 27657
rect 29731 27616 29740 27656
rect 29780 27616 29789 27656
rect 29731 27615 29789 27616
rect 30027 27656 30069 27665
rect 30027 27616 30028 27656
rect 30068 27616 30069 27656
rect 30027 27607 30069 27616
rect 30123 27656 30165 27665
rect 30123 27616 30124 27656
rect 30164 27616 30165 27656
rect 30123 27607 30165 27616
rect 30219 27656 30261 27665
rect 30219 27616 30220 27656
rect 30260 27616 30261 27656
rect 30219 27607 30261 27616
rect 30315 27656 30357 27665
rect 30315 27616 30316 27656
rect 30356 27616 30357 27656
rect 30315 27607 30357 27616
rect 30507 27656 30549 27665
rect 30507 27616 30508 27656
rect 30548 27616 30549 27656
rect 30507 27607 30549 27616
rect 30699 27656 30741 27665
rect 30699 27616 30700 27656
rect 30740 27616 30741 27656
rect 30699 27607 30741 27616
rect 30787 27656 30845 27657
rect 30787 27616 30796 27656
rect 30836 27616 30845 27656
rect 30787 27615 30845 27616
rect 31371 27656 31413 27665
rect 31371 27616 31372 27656
rect 31412 27616 31413 27656
rect 31371 27607 31413 27616
rect 31651 27656 31709 27657
rect 31651 27616 31660 27656
rect 31700 27616 31709 27656
rect 31651 27615 31709 27616
rect 32611 27656 32669 27657
rect 32611 27616 32620 27656
rect 32660 27616 32669 27656
rect 32611 27615 32669 27616
rect 33379 27656 33437 27657
rect 33379 27616 33388 27656
rect 33428 27616 33437 27656
rect 33379 27615 33437 27616
rect 33771 27656 33813 27665
rect 33771 27616 33772 27656
rect 33812 27616 33813 27656
rect 33771 27607 33813 27616
rect 33867 27656 33909 27665
rect 33867 27616 33868 27656
rect 33908 27616 33909 27656
rect 33867 27607 33909 27616
rect 33963 27656 34005 27665
rect 33963 27616 33964 27656
rect 34004 27616 34005 27656
rect 33963 27607 34005 27616
rect 34531 27656 34589 27657
rect 34531 27616 34540 27656
rect 34580 27616 34589 27656
rect 34531 27615 34589 27616
rect 35395 27656 35453 27657
rect 35395 27616 35404 27656
rect 35444 27616 35453 27656
rect 35395 27615 35453 27616
rect 36939 27656 36981 27665
rect 36939 27616 36940 27656
rect 36980 27616 36981 27656
rect 36939 27607 36981 27616
rect 37315 27656 37373 27657
rect 37315 27616 37324 27656
rect 37364 27616 37373 27656
rect 37315 27615 37373 27616
rect 38179 27656 38237 27657
rect 38179 27616 38188 27656
rect 38228 27616 38237 27656
rect 38179 27615 38237 27616
rect 39907 27656 39965 27657
rect 39907 27616 39916 27656
rect 39956 27616 39965 27656
rect 39907 27615 39965 27616
rect 40771 27656 40829 27657
rect 40771 27616 40780 27656
rect 40820 27616 40829 27656
rect 40771 27615 40829 27616
rect 42115 27656 42173 27657
rect 42115 27616 42124 27656
rect 42164 27616 42173 27656
rect 42115 27615 42173 27616
rect 43755 27656 43797 27665
rect 43755 27616 43756 27656
rect 43796 27616 43797 27656
rect 43755 27607 43797 27616
rect 44139 27656 44181 27665
rect 44139 27616 44140 27656
rect 44180 27616 44181 27656
rect 44139 27607 44181 27616
rect 44515 27656 44573 27657
rect 44515 27616 44524 27656
rect 44564 27616 44573 27656
rect 44515 27615 44573 27616
rect 45379 27656 45437 27657
rect 45379 27616 45388 27656
rect 45428 27616 45437 27656
rect 45379 27615 45437 27616
rect 46819 27656 46877 27657
rect 46819 27616 46828 27656
rect 46868 27616 46877 27656
rect 46819 27615 46877 27616
rect 47683 27656 47741 27657
rect 47683 27616 47692 27656
rect 47732 27616 47741 27656
rect 47683 27615 47741 27616
rect 48259 27656 48317 27657
rect 48259 27616 48268 27656
rect 48308 27616 48317 27656
rect 48259 27615 48317 27616
rect 49123 27656 49181 27657
rect 49123 27616 49132 27656
rect 49172 27616 49181 27656
rect 49123 27615 49181 27616
rect 51139 27656 51197 27657
rect 51139 27616 51148 27656
rect 51188 27616 51197 27656
rect 51139 27615 51197 27616
rect 3627 27572 3669 27581
rect 3627 27532 3628 27572
rect 3668 27532 3669 27572
rect 3627 27523 3669 27532
rect 28675 27572 28733 27573
rect 28675 27532 28684 27572
rect 28724 27532 28733 27572
rect 28675 27531 28733 27532
rect 39339 27572 39381 27581
rect 39339 27532 39340 27572
rect 39380 27532 39381 27572
rect 39339 27523 39381 27532
rect 50283 27572 50325 27581
rect 50283 27532 50284 27572
rect 50324 27532 50325 27572
rect 50283 27523 50325 27532
rect 4107 27488 4149 27497
rect 4107 27448 4108 27488
rect 4148 27448 4149 27488
rect 4107 27439 4149 27448
rect 10059 27488 10101 27497
rect 10059 27448 10060 27488
rect 10100 27448 10101 27488
rect 10059 27439 10101 27448
rect 16491 27488 16533 27497
rect 16491 27448 16492 27488
rect 16532 27448 16533 27488
rect 16491 27439 16533 27448
rect 23787 27488 23829 27497
rect 23787 27448 23788 27488
rect 23828 27448 23829 27488
rect 23787 27439 23829 27448
rect 25035 27488 25077 27497
rect 25035 27448 25036 27488
rect 25076 27448 25077 27488
rect 25035 27439 25077 27448
rect 28875 27488 28917 27497
rect 28875 27448 28876 27488
rect 28916 27448 28917 27488
rect 28875 27439 28917 27448
rect 32811 27488 32853 27497
rect 32811 27448 32812 27488
rect 32852 27448 32853 27488
rect 32811 27439 32853 27448
rect 36547 27488 36605 27489
rect 36547 27448 36556 27488
rect 36596 27448 36605 27488
rect 36547 27447 36605 27448
rect 41923 27488 41981 27489
rect 41923 27448 41932 27488
rect 41972 27448 41981 27488
rect 41923 27447 41981 27448
rect 4683 27404 4725 27413
rect 4683 27364 4684 27404
rect 4724 27364 4725 27404
rect 4683 27355 4725 27364
rect 6307 27404 6365 27405
rect 6307 27364 6316 27404
rect 6356 27364 6365 27404
rect 6307 27363 6365 27364
rect 6507 27404 6549 27413
rect 6507 27364 6508 27404
rect 6548 27364 6549 27404
rect 6507 27355 6549 27364
rect 7267 27404 7325 27405
rect 7267 27364 7276 27404
rect 7316 27364 7325 27404
rect 7267 27363 7325 27364
rect 10243 27404 10301 27405
rect 10243 27364 10252 27404
rect 10292 27364 10301 27404
rect 10243 27363 10301 27364
rect 11875 27404 11933 27405
rect 11875 27364 11884 27404
rect 11924 27364 11933 27404
rect 11875 27363 11933 27364
rect 12363 27404 12405 27413
rect 12363 27364 12364 27404
rect 12404 27364 12405 27404
rect 12363 27355 12405 27364
rect 14571 27404 14613 27413
rect 14571 27364 14572 27404
rect 14612 27364 14613 27404
rect 14571 27355 14613 27364
rect 15043 27404 15101 27405
rect 15043 27364 15052 27404
rect 15092 27364 15101 27404
rect 15043 27363 15101 27364
rect 17827 27404 17885 27405
rect 17827 27364 17836 27404
rect 17876 27364 17885 27404
rect 17827 27363 17885 27364
rect 19851 27404 19893 27413
rect 19851 27364 19852 27404
rect 19892 27364 19893 27404
rect 19851 27355 19893 27364
rect 26275 27404 26333 27405
rect 26275 27364 26284 27404
rect 26324 27364 26333 27404
rect 26275 27363 26333 27364
rect 28107 27404 28149 27413
rect 28107 27364 28108 27404
rect 28148 27364 28149 27404
rect 28107 27355 28149 27364
rect 28491 27404 28533 27413
rect 28491 27364 28492 27404
rect 28532 27364 28533 27404
rect 28491 27355 28533 27364
rect 30507 27404 30549 27413
rect 30507 27364 30508 27404
rect 30548 27364 30549 27404
rect 30507 27355 30549 27364
rect 30979 27404 31037 27405
rect 30979 27364 30988 27404
rect 31028 27364 31037 27404
rect 30979 27363 31037 27364
rect 31939 27404 31997 27405
rect 31939 27364 31948 27404
rect 31988 27364 31997 27404
rect 31939 27363 31997 27364
rect 33291 27404 33333 27413
rect 33291 27364 33292 27404
rect 33332 27364 33333 27404
rect 33291 27355 33333 27364
rect 43563 27404 43605 27413
rect 43563 27364 43564 27404
rect 43604 27364 43605 27404
rect 43563 27355 43605 27364
rect 46531 27404 46589 27405
rect 46531 27364 46540 27404
rect 46580 27364 46589 27404
rect 46531 27363 46589 27364
rect 46731 27404 46773 27413
rect 46731 27364 46732 27404
rect 46772 27364 46773 27404
rect 46731 27355 46773 27364
rect 47011 27404 47069 27405
rect 47011 27364 47020 27404
rect 47060 27364 47069 27404
rect 47011 27363 47069 27364
rect 50467 27404 50525 27405
rect 50467 27364 50476 27404
rect 50516 27364 50525 27404
rect 50467 27363 50525 27364
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 2763 27068 2805 27077
rect 2763 27028 2764 27068
rect 2804 27028 2805 27068
rect 2763 27019 2805 27028
rect 4867 27068 4925 27069
rect 4867 27028 4876 27068
rect 4916 27028 4925 27068
rect 4867 27027 4925 27028
rect 8427 27068 8469 27077
rect 8427 27028 8428 27068
rect 8468 27028 8469 27068
rect 8427 27019 8469 27028
rect 9291 27068 9333 27077
rect 9291 27028 9292 27068
rect 9332 27028 9333 27068
rect 9291 27019 9333 27028
rect 12459 27068 12501 27077
rect 12459 27028 12460 27068
rect 12500 27028 12501 27068
rect 12459 27019 12501 27028
rect 17739 27068 17781 27077
rect 17739 27028 17740 27068
rect 17780 27028 17781 27068
rect 17739 27019 17781 27028
rect 20515 27068 20573 27069
rect 20515 27028 20524 27068
rect 20564 27028 20573 27068
rect 20515 27027 20573 27028
rect 24075 27068 24117 27077
rect 24075 27028 24076 27068
rect 24116 27028 24117 27068
rect 24075 27019 24117 27028
rect 30987 27068 31029 27077
rect 30987 27028 30988 27068
rect 31028 27028 31029 27068
rect 30987 27019 31029 27028
rect 34243 27068 34301 27069
rect 34243 27028 34252 27068
rect 34292 27028 34301 27068
rect 34243 27027 34301 27028
rect 37707 27068 37749 27077
rect 37707 27028 37708 27068
rect 37748 27028 37749 27068
rect 37707 27019 37749 27028
rect 39435 27068 39477 27077
rect 39435 27028 39436 27068
rect 39476 27028 39477 27068
rect 39435 27019 39477 27028
rect 40491 27068 40533 27077
rect 40491 27028 40492 27068
rect 40532 27028 40533 27068
rect 40491 27019 40533 27028
rect 42987 27068 43029 27077
rect 42987 27028 42988 27068
rect 43028 27028 43029 27068
rect 42987 27019 43029 27028
rect 45099 27068 45141 27077
rect 45099 27028 45100 27068
rect 45140 27028 45141 27068
rect 45099 27019 45141 27028
rect 45579 27068 45621 27077
rect 45579 27028 45580 27068
rect 45620 27028 45621 27068
rect 45579 27019 45621 27028
rect 46539 27068 46581 27077
rect 46539 27028 46540 27068
rect 46580 27028 46581 27068
rect 46539 27019 46581 27028
rect 51715 27068 51773 27069
rect 51715 27028 51724 27068
rect 51764 27028 51773 27068
rect 51715 27027 51773 27028
rect 2187 26984 2229 26993
rect 2187 26944 2188 26984
rect 2228 26944 2229 26984
rect 2187 26935 2229 26944
rect 9099 26984 9141 26993
rect 9099 26944 9100 26984
rect 9140 26944 9141 26984
rect 9099 26935 9141 26944
rect 11491 26984 11549 26985
rect 11491 26944 11500 26984
rect 11540 26944 11549 26984
rect 11491 26943 11549 26944
rect 13227 26984 13269 26993
rect 13227 26944 13228 26984
rect 13268 26944 13269 26984
rect 13227 26935 13269 26944
rect 23403 26984 23445 26993
rect 23403 26944 23404 26984
rect 23444 26944 23445 26984
rect 23403 26935 23445 26944
rect 38467 26984 38525 26985
rect 38467 26944 38476 26984
rect 38516 26944 38525 26984
rect 38467 26943 38525 26944
rect 40011 26984 40053 26993
rect 40011 26944 40012 26984
rect 40052 26944 40053 26984
rect 40011 26935 40053 26944
rect 27435 26900 27477 26909
rect 27435 26860 27436 26900
rect 27476 26860 27477 26900
rect 27435 26851 27477 26860
rect 30115 26900 30173 26901
rect 30115 26860 30124 26900
rect 30164 26860 30173 26900
rect 30115 26859 30173 26860
rect 13960 26831 14002 26840
rect 2851 26816 2909 26817
rect 2851 26776 2860 26816
rect 2900 26776 2909 26816
rect 2851 26775 2909 26776
rect 3139 26816 3197 26817
rect 3139 26776 3148 26816
rect 3188 26776 3197 26816
rect 3139 26775 3197 26776
rect 3331 26816 3389 26817
rect 3331 26776 3340 26816
rect 3380 26776 3389 26816
rect 3331 26775 3389 26776
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 3915 26816 3957 26825
rect 3915 26776 3916 26816
rect 3956 26776 3957 26816
rect 3915 26767 3957 26776
rect 4011 26816 4053 26825
rect 4011 26776 4012 26816
rect 4052 26776 4053 26816
rect 4011 26767 4053 26776
rect 4107 26816 4149 26825
rect 4107 26776 4108 26816
rect 4148 26776 4149 26816
rect 4107 26767 4149 26776
rect 4395 26816 4437 26825
rect 4395 26776 4396 26816
rect 4436 26776 4437 26816
rect 4395 26767 4437 26776
rect 4491 26816 4533 26825
rect 4491 26776 4492 26816
rect 4532 26776 4533 26816
rect 4491 26767 4533 26776
rect 4587 26816 4629 26825
rect 4587 26776 4588 26816
rect 4628 26776 4629 26816
rect 4587 26767 4629 26776
rect 4683 26816 4725 26825
rect 4683 26776 4684 26816
rect 4724 26776 4725 26816
rect 4683 26767 4725 26776
rect 5539 26816 5597 26817
rect 5539 26776 5548 26816
rect 5588 26776 5597 26816
rect 5539 26775 5597 26776
rect 5739 26816 5781 26825
rect 5739 26776 5740 26816
rect 5780 26776 5781 26816
rect 5739 26767 5781 26776
rect 5931 26816 5973 26825
rect 5931 26776 5932 26816
rect 5972 26776 5973 26816
rect 5931 26767 5973 26776
rect 6019 26816 6077 26817
rect 6019 26776 6028 26816
rect 6068 26776 6077 26816
rect 6019 26775 6077 26776
rect 6219 26816 6261 26825
rect 6219 26776 6220 26816
rect 6260 26776 6261 26816
rect 6219 26767 6261 26776
rect 6403 26816 6461 26817
rect 6403 26776 6412 26816
rect 6452 26776 6461 26816
rect 6403 26775 6461 26776
rect 7555 26816 7613 26817
rect 7555 26776 7564 26816
rect 7604 26776 7613 26816
rect 7555 26775 7613 26776
rect 7843 26816 7901 26817
rect 7843 26776 7852 26816
rect 7892 26776 7901 26816
rect 7843 26775 7901 26776
rect 7947 26816 7989 26825
rect 7947 26776 7948 26816
rect 7988 26776 7989 26816
rect 7947 26767 7989 26776
rect 8139 26816 8181 26825
rect 8139 26776 8140 26816
rect 8180 26776 8181 26816
rect 8139 26767 8181 26776
rect 8331 26816 8373 26825
rect 8331 26776 8332 26816
rect 8372 26776 8373 26816
rect 8331 26767 8373 26776
rect 8515 26816 8573 26817
rect 8515 26776 8524 26816
rect 8564 26776 8573 26816
rect 8515 26775 8573 26776
rect 9291 26816 9333 26825
rect 9291 26776 9292 26816
rect 9332 26776 9333 26816
rect 9291 26767 9333 26776
rect 9483 26816 9525 26825
rect 9483 26776 9484 26816
rect 9524 26776 9525 26816
rect 9483 26767 9525 26776
rect 9571 26816 9629 26817
rect 9571 26776 9580 26816
rect 9620 26776 9629 26816
rect 9571 26775 9629 26776
rect 9771 26816 9813 26825
rect 9771 26776 9772 26816
rect 9812 26776 9813 26816
rect 9771 26767 9813 26776
rect 9867 26816 9909 26825
rect 9867 26776 9868 26816
rect 9908 26776 9909 26816
rect 9867 26767 9909 26776
rect 9963 26816 10005 26825
rect 9963 26776 9964 26816
rect 10004 26776 10005 26816
rect 9963 26767 10005 26776
rect 10251 26816 10293 26825
rect 10251 26776 10252 26816
rect 10292 26776 10293 26816
rect 10251 26767 10293 26776
rect 10347 26816 10389 26825
rect 10347 26776 10348 26816
rect 10388 26776 10389 26816
rect 10347 26767 10389 26776
rect 10443 26816 10485 26825
rect 10443 26776 10444 26816
rect 10484 26776 10485 26816
rect 10443 26767 10485 26776
rect 10539 26816 10581 26825
rect 10539 26776 10540 26816
rect 10580 26776 10581 26816
rect 10539 26767 10581 26776
rect 10819 26816 10877 26817
rect 10819 26776 10828 26816
rect 10868 26776 10877 26816
rect 10819 26775 10877 26776
rect 11115 26816 11157 26825
rect 11115 26776 11116 26816
rect 11156 26776 11157 26816
rect 11115 26767 11157 26776
rect 11683 26816 11741 26817
rect 11683 26776 11692 26816
rect 11732 26776 11741 26816
rect 11683 26775 11741 26776
rect 12459 26816 12501 26825
rect 12459 26776 12460 26816
rect 12500 26776 12501 26816
rect 12459 26767 12501 26776
rect 12651 26816 12693 26825
rect 12651 26776 12652 26816
rect 12692 26776 12693 26816
rect 12651 26767 12693 26776
rect 12739 26816 12797 26817
rect 12739 26776 12748 26816
rect 12788 26776 12797 26816
rect 12739 26775 12797 26776
rect 12931 26816 12989 26817
rect 12931 26776 12940 26816
rect 12980 26776 12989 26816
rect 12931 26775 12989 26776
rect 13035 26816 13077 26825
rect 13035 26776 13036 26816
rect 13076 26776 13077 26816
rect 13035 26767 13077 26776
rect 13227 26816 13269 26825
rect 13227 26776 13228 26816
rect 13268 26776 13269 26816
rect 13227 26767 13269 26776
rect 13411 26816 13469 26817
rect 13411 26776 13420 26816
rect 13460 26776 13469 26816
rect 13411 26775 13469 26776
rect 13507 26816 13565 26817
rect 13507 26776 13516 26816
rect 13556 26776 13565 26816
rect 13507 26775 13565 26776
rect 13707 26816 13749 26825
rect 13707 26776 13708 26816
rect 13748 26776 13749 26816
rect 13707 26767 13749 26776
rect 13803 26816 13845 26825
rect 13803 26776 13804 26816
rect 13844 26776 13845 26816
rect 13960 26791 13961 26831
rect 14001 26791 14002 26831
rect 13960 26782 14002 26791
rect 14179 26816 14237 26817
rect 13803 26767 13845 26776
rect 14179 26776 14188 26816
rect 14228 26776 14237 26816
rect 14179 26775 14237 26776
rect 14275 26816 14333 26817
rect 14275 26776 14284 26816
rect 14324 26776 14333 26816
rect 14275 26775 14333 26776
rect 14475 26816 14517 26825
rect 14475 26776 14476 26816
rect 14516 26776 14517 26816
rect 14475 26767 14517 26776
rect 14571 26816 14613 26825
rect 14571 26776 14572 26816
rect 14612 26776 14613 26816
rect 14571 26767 14613 26776
rect 14718 26816 14776 26817
rect 14718 26776 14727 26816
rect 14767 26776 14776 26816
rect 14718 26775 14776 26776
rect 14955 26816 14997 26825
rect 14955 26776 14956 26816
rect 14996 26776 14997 26816
rect 14955 26767 14997 26776
rect 15139 26816 15197 26817
rect 15139 26776 15148 26816
rect 15188 26776 15197 26816
rect 15139 26775 15197 26776
rect 15331 26816 15389 26817
rect 15331 26776 15340 26816
rect 15380 26776 15389 26816
rect 15331 26775 15389 26776
rect 15435 26816 15477 26825
rect 15435 26776 15436 26816
rect 15476 26776 15477 26816
rect 15435 26767 15477 26776
rect 15627 26816 15669 26825
rect 15627 26776 15628 26816
rect 15668 26776 15669 26816
rect 15627 26767 15669 26776
rect 16003 26816 16061 26817
rect 16003 26776 16012 26816
rect 16052 26776 16061 26816
rect 16003 26775 16061 26776
rect 16107 26816 16149 26825
rect 16107 26776 16108 26816
rect 16148 26776 16149 26816
rect 16107 26767 16149 26776
rect 16299 26816 16341 26825
rect 16299 26776 16300 26816
rect 16340 26776 16341 26816
rect 16299 26767 16341 26776
rect 16579 26816 16637 26817
rect 16579 26776 16588 26816
rect 16628 26776 16637 26816
rect 16579 26775 16637 26776
rect 16771 26816 16829 26817
rect 16771 26776 16780 26816
rect 16820 26776 16829 26816
rect 16771 26775 16829 26776
rect 16963 26816 17021 26817
rect 16963 26776 16972 26816
rect 17012 26776 17021 26816
rect 16963 26775 17021 26776
rect 17163 26816 17205 26825
rect 17163 26776 17164 26816
rect 17204 26776 17205 26816
rect 17163 26767 17205 26776
rect 17827 26816 17885 26817
rect 17827 26776 17836 26816
rect 17876 26776 17885 26816
rect 17827 26775 17885 26776
rect 18123 26816 18165 26825
rect 18123 26776 18124 26816
rect 18164 26776 18165 26816
rect 18123 26767 18165 26776
rect 18219 26816 18261 26825
rect 18219 26776 18220 26816
rect 18260 26776 18261 26816
rect 18219 26767 18261 26776
rect 18315 26816 18357 26825
rect 18315 26776 18316 26816
rect 18356 26776 18357 26816
rect 18315 26767 18357 26776
rect 18603 26816 18645 26825
rect 18603 26776 18604 26816
rect 18644 26776 18645 26816
rect 18603 26767 18645 26776
rect 18699 26816 18741 26825
rect 18699 26776 18700 26816
rect 18740 26776 18741 26816
rect 18699 26767 18741 26776
rect 18795 26816 18837 26825
rect 18795 26776 18796 26816
rect 18836 26776 18837 26816
rect 18795 26767 18837 26776
rect 19083 26816 19125 26825
rect 19083 26776 19084 26816
rect 19124 26776 19125 26816
rect 19083 26767 19125 26776
rect 19275 26816 19317 26825
rect 19275 26776 19276 26816
rect 19316 26776 19317 26816
rect 19275 26767 19317 26776
rect 19363 26816 19421 26817
rect 19363 26776 19372 26816
rect 19412 26776 19421 26816
rect 19363 26775 19421 26776
rect 19563 26816 19605 26825
rect 19563 26776 19564 26816
rect 19604 26776 19605 26816
rect 19563 26767 19605 26776
rect 20227 26816 20285 26817
rect 20227 26776 20236 26816
rect 20276 26776 20285 26816
rect 20227 26775 20285 26776
rect 21667 26816 21725 26817
rect 21667 26776 21676 26816
rect 21716 26776 21725 26816
rect 21667 26775 21725 26776
rect 22531 26816 22589 26817
rect 22531 26776 22540 26816
rect 22580 26776 22589 26816
rect 22531 26775 22589 26776
rect 24459 26816 24501 26825
rect 24459 26776 24460 26816
rect 24500 26776 24501 26816
rect 24459 26767 24501 26776
rect 24939 26816 24981 26825
rect 24939 26776 24940 26816
rect 24980 26776 24981 26816
rect 24939 26767 24981 26776
rect 25035 26816 25077 26825
rect 25035 26776 25036 26816
rect 25076 26776 25077 26816
rect 25035 26767 25077 26776
rect 25131 26816 25173 26825
rect 25131 26776 25132 26816
rect 25172 26776 25173 26816
rect 25131 26767 25173 26776
rect 25419 26816 25461 26825
rect 25419 26776 25420 26816
rect 25460 26776 25461 26816
rect 25419 26767 25461 26776
rect 25611 26816 25653 26825
rect 25611 26776 25612 26816
rect 25652 26776 25653 26816
rect 25611 26767 25653 26776
rect 25699 26816 25757 26817
rect 25699 26776 25708 26816
rect 25748 26776 25757 26816
rect 25699 26775 25757 26776
rect 26563 26816 26621 26817
rect 26563 26776 26572 26816
rect 26612 26776 26621 26816
rect 26563 26775 26621 26776
rect 26955 26816 26997 26825
rect 26955 26776 26956 26816
rect 26996 26776 26997 26816
rect 26955 26767 26997 26776
rect 27051 26816 27093 26825
rect 27051 26776 27052 26816
rect 27092 26776 27093 26816
rect 27051 26767 27093 26776
rect 27531 26816 27573 26825
rect 28491 26821 28533 26830
rect 27531 26776 27532 26816
rect 27572 26776 27573 26816
rect 27531 26767 27573 26776
rect 28003 26816 28061 26817
rect 28003 26776 28012 26816
rect 28052 26776 28061 26816
rect 28003 26775 28061 26776
rect 28491 26781 28492 26821
rect 28532 26781 28533 26821
rect 28491 26772 28533 26781
rect 28875 26816 28917 26825
rect 28875 26776 28876 26816
rect 28916 26776 28917 26816
rect 28875 26767 28917 26776
rect 29067 26816 29109 26825
rect 29067 26776 29068 26816
rect 29108 26776 29109 26816
rect 29067 26767 29109 26776
rect 29155 26816 29213 26817
rect 29155 26776 29164 26816
rect 29204 26776 29213 26816
rect 29155 26775 29213 26776
rect 29547 26816 29589 26825
rect 29547 26776 29548 26816
rect 29588 26776 29589 26816
rect 29547 26767 29589 26776
rect 29643 26816 29685 26825
rect 29643 26776 29644 26816
rect 29684 26776 29685 26816
rect 29643 26767 29685 26776
rect 30507 26816 30549 26825
rect 30507 26776 30508 26816
rect 30548 26776 30549 26816
rect 30507 26767 30549 26776
rect 30603 26816 30645 26825
rect 30603 26776 30604 26816
rect 30644 26776 30645 26816
rect 30603 26767 30645 26776
rect 30699 26816 30741 26825
rect 30699 26776 30700 26816
rect 30740 26776 30741 26816
rect 30699 26767 30741 26776
rect 30987 26816 31029 26825
rect 30987 26776 30988 26816
rect 31028 26776 31029 26816
rect 30987 26767 31029 26776
rect 31179 26816 31221 26825
rect 31179 26776 31180 26816
rect 31220 26776 31221 26816
rect 31179 26767 31221 26776
rect 31267 26816 31325 26817
rect 31267 26776 31276 26816
rect 31316 26776 31325 26816
rect 31267 26775 31325 26776
rect 31851 26816 31893 26825
rect 31851 26776 31852 26816
rect 31892 26776 31893 26816
rect 31851 26767 31893 26776
rect 32227 26816 32285 26817
rect 32227 26776 32236 26816
rect 32276 26776 32285 26816
rect 32227 26775 32285 26776
rect 33091 26816 33149 26817
rect 33091 26776 33100 26816
rect 33140 26776 33149 26816
rect 33091 26775 33149 26776
rect 34627 26816 34685 26817
rect 34627 26776 34636 26816
rect 34676 26776 34685 26816
rect 34627 26775 34685 26776
rect 34731 26816 34773 26825
rect 34731 26776 34732 26816
rect 34772 26776 34773 26816
rect 34731 26767 34773 26776
rect 34923 26816 34965 26825
rect 34923 26776 34924 26816
rect 34964 26776 34965 26816
rect 34923 26767 34965 26776
rect 35395 26816 35453 26817
rect 35395 26776 35404 26816
rect 35444 26776 35453 26816
rect 35395 26775 35453 26776
rect 35587 26816 35645 26817
rect 35587 26776 35596 26816
rect 35636 26776 35645 26816
rect 35587 26775 35645 26776
rect 35787 26816 35829 26825
rect 35787 26776 35788 26816
rect 35828 26776 35829 26816
rect 35787 26767 35829 26776
rect 38179 26816 38237 26817
rect 38179 26776 38188 26816
rect 38228 26776 38237 26816
rect 38179 26775 38237 26776
rect 38763 26816 38805 26825
rect 38763 26776 38764 26816
rect 38804 26776 38805 26816
rect 38763 26767 38805 26776
rect 38859 26816 38901 26825
rect 38859 26776 38860 26816
rect 38900 26776 38901 26816
rect 38859 26767 38901 26776
rect 39139 26816 39197 26817
rect 39139 26776 39148 26816
rect 39188 26776 39197 26816
rect 39139 26775 39197 26776
rect 39435 26816 39477 26825
rect 39435 26776 39436 26816
rect 39476 26776 39477 26816
rect 39435 26767 39477 26776
rect 39627 26816 39669 26825
rect 39627 26776 39628 26816
rect 39668 26776 39669 26816
rect 39627 26767 39669 26776
rect 39715 26816 39773 26817
rect 39715 26776 39724 26816
rect 39764 26776 39773 26816
rect 39715 26775 39773 26776
rect 40387 26816 40445 26817
rect 40387 26776 40396 26816
rect 40436 26776 40445 26816
rect 40387 26775 40445 26776
rect 41059 26816 41117 26817
rect 41059 26776 41068 26816
rect 41108 26776 41117 26816
rect 41059 26775 41117 26776
rect 42019 26816 42077 26817
rect 42019 26776 42028 26816
rect 42068 26776 42077 26816
rect 42019 26775 42077 26776
rect 42691 26816 42749 26817
rect 42691 26776 42700 26816
rect 42740 26776 42749 26816
rect 42691 26775 42749 26776
rect 42795 26816 42837 26825
rect 42795 26776 42796 26816
rect 42836 26776 42837 26816
rect 42795 26767 42837 26776
rect 42987 26816 43029 26825
rect 42987 26776 42988 26816
rect 43028 26776 43029 26816
rect 42987 26767 43029 26776
rect 43179 26816 43221 26825
rect 43179 26776 43180 26816
rect 43220 26776 43221 26816
rect 43179 26767 43221 26776
rect 43275 26816 43317 26825
rect 43275 26776 43276 26816
rect 43316 26776 43317 26816
rect 43275 26767 43317 26776
rect 43371 26816 43413 26825
rect 43371 26776 43372 26816
rect 43412 26776 43413 26816
rect 43371 26767 43413 26776
rect 43467 26816 43509 26825
rect 43467 26776 43468 26816
rect 43508 26776 43509 26816
rect 43467 26767 43509 26776
rect 43651 26816 43709 26817
rect 43651 26776 43660 26816
rect 43700 26776 43709 26816
rect 43651 26775 43709 26776
rect 43755 26816 43797 26825
rect 43755 26776 43756 26816
rect 43796 26776 43797 26816
rect 43755 26767 43797 26776
rect 43947 26816 43989 26825
rect 43947 26776 43948 26816
rect 43988 26776 43989 26816
rect 43947 26767 43989 26776
rect 44803 26816 44861 26817
rect 44803 26776 44812 26816
rect 44852 26776 44861 26816
rect 44803 26775 44861 26776
rect 44995 26816 45053 26817
rect 44995 26776 45004 26816
rect 45044 26776 45053 26816
rect 44995 26775 45053 26776
rect 45283 26816 45341 26817
rect 45283 26776 45292 26816
rect 45332 26776 45341 26816
rect 45283 26775 45341 26776
rect 45387 26816 45429 26825
rect 45387 26776 45388 26816
rect 45428 26776 45429 26816
rect 45387 26767 45429 26776
rect 45579 26816 45621 26825
rect 45579 26776 45580 26816
rect 45620 26776 45621 26816
rect 45579 26767 45621 26776
rect 45859 26816 45917 26817
rect 45859 26776 45868 26816
rect 45908 26776 45917 26816
rect 45859 26775 45917 26776
rect 47875 26816 47933 26817
rect 47875 26776 47884 26816
rect 47924 26776 47933 26816
rect 47875 26775 47933 26776
rect 48163 26816 48221 26817
rect 48163 26776 48172 26816
rect 48212 26776 48221 26816
rect 48163 26775 48221 26776
rect 49699 26816 49757 26817
rect 49699 26776 49708 26816
rect 49748 26776 49757 26816
rect 49699 26775 49757 26776
rect 50563 26816 50621 26817
rect 50563 26776 50572 26816
rect 50612 26776 50621 26816
rect 50563 26775 50621 26776
rect 3819 26732 3861 26741
rect 3819 26692 3820 26732
rect 3860 26692 3861 26732
rect 3819 26683 3861 26692
rect 5835 26732 5877 26741
rect 5835 26692 5836 26732
rect 5876 26692 5877 26732
rect 5835 26683 5877 26692
rect 6315 26732 6357 26741
rect 6315 26692 6316 26732
rect 6356 26692 6357 26732
rect 6315 26683 6357 26692
rect 6691 26732 6749 26733
rect 6691 26692 6700 26732
rect 6740 26692 6749 26732
rect 6691 26691 6749 26692
rect 8043 26732 8085 26741
rect 8043 26692 8044 26732
rect 8084 26692 8085 26732
rect 8043 26683 8085 26692
rect 11211 26732 11253 26741
rect 11211 26692 11212 26732
rect 11252 26692 11253 26732
rect 11211 26683 11253 26692
rect 11787 26732 11829 26741
rect 11787 26692 11788 26732
rect 11828 26692 11829 26732
rect 11787 26683 11829 26692
rect 15051 26732 15093 26741
rect 15051 26692 15052 26732
rect 15092 26692 15093 26732
rect 15051 26683 15093 26692
rect 15531 26732 15573 26741
rect 15531 26692 15532 26732
rect 15572 26692 15573 26732
rect 15531 26683 15573 26692
rect 17067 26732 17109 26741
rect 17067 26692 17068 26732
rect 17108 26692 17109 26732
rect 17067 26683 17109 26692
rect 22923 26732 22965 26741
rect 22923 26692 22924 26732
rect 22964 26692 22965 26732
rect 22923 26683 22965 26692
rect 28971 26732 29013 26741
rect 28971 26692 28972 26732
rect 29012 26692 29013 26732
rect 28971 26683 29013 26692
rect 35691 26732 35733 26741
rect 35691 26692 35692 26732
rect 35732 26692 35733 26732
rect 35691 26683 35733 26692
rect 49027 26732 49085 26733
rect 49027 26692 49036 26732
rect 49076 26692 49085 26732
rect 49027 26691 49085 26692
rect 49323 26732 49365 26741
rect 49323 26692 49324 26732
rect 49364 26692 49365 26732
rect 49323 26683 49365 26692
rect 3051 26648 3093 26657
rect 3051 26608 3052 26648
rect 3092 26608 3093 26648
rect 3051 26599 3093 26608
rect 3523 26648 3581 26649
rect 3523 26608 3532 26648
rect 3572 26608 3581 26648
rect 3523 26607 3581 26608
rect 7083 26648 7125 26657
rect 7083 26608 7084 26648
rect 7124 26608 7125 26648
rect 7083 26599 7125 26608
rect 10051 26648 10109 26649
rect 10051 26608 10060 26648
rect 10100 26608 10109 26648
rect 10051 26607 10109 26608
rect 13795 26648 13853 26649
rect 13795 26608 13804 26648
rect 13844 26608 13853 26648
rect 13795 26607 13853 26608
rect 14371 26648 14429 26649
rect 14371 26608 14380 26648
rect 14420 26608 14429 26648
rect 14371 26607 14429 26608
rect 16195 26648 16253 26649
rect 16195 26608 16204 26648
rect 16244 26608 16253 26648
rect 16195 26607 16253 26608
rect 18019 26648 18077 26649
rect 18019 26608 18028 26648
rect 18068 26608 18077 26648
rect 18019 26607 18077 26608
rect 18883 26648 18941 26649
rect 18883 26608 18892 26648
rect 18932 26608 18941 26648
rect 18883 26607 18941 26608
rect 19171 26648 19229 26649
rect 19171 26608 19180 26648
rect 19220 26608 19229 26648
rect 19171 26607 19229 26608
rect 24835 26648 24893 26649
rect 24835 26608 24844 26648
rect 24884 26608 24893 26648
rect 24835 26607 24893 26608
rect 25507 26648 25565 26649
rect 25507 26608 25516 26648
rect 25556 26608 25565 26648
rect 25507 26607 25565 26608
rect 25891 26648 25949 26649
rect 25891 26608 25900 26648
rect 25940 26608 25949 26648
rect 25891 26607 25949 26608
rect 28683 26648 28725 26657
rect 28683 26608 28684 26648
rect 28724 26608 28725 26648
rect 28683 26599 28725 26608
rect 29347 26648 29405 26649
rect 29347 26608 29356 26648
rect 29396 26608 29405 26648
rect 29347 26607 29405 26608
rect 29931 26648 29973 26657
rect 29931 26608 29932 26648
rect 29972 26608 29973 26648
rect 29931 26599 29973 26608
rect 30787 26648 30845 26649
rect 30787 26608 30796 26648
rect 30836 26608 30845 26648
rect 30787 26607 30845 26608
rect 34819 26648 34877 26649
rect 34819 26608 34828 26648
rect 34868 26608 34877 26648
rect 34819 26607 34877 26608
rect 35307 26648 35349 26657
rect 35307 26608 35308 26648
rect 35348 26608 35349 26648
rect 35307 26599 35349 26608
rect 43843 26648 43901 26649
rect 43843 26608 43852 26648
rect 43892 26608 43901 26648
rect 43843 26607 43901 26608
rect 44131 26648 44189 26649
rect 44131 26608 44140 26648
rect 44180 26608 44189 26648
rect 44131 26607 44189 26608
rect 47203 26648 47261 26649
rect 47203 26608 47212 26648
rect 47252 26608 47261 26648
rect 47203 26607 47261 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 30795 26370 30837 26379
rect 30795 26330 30796 26370
rect 30836 26330 30837 26370
rect 30795 26321 30837 26330
rect 11203 26312 11261 26313
rect 11203 26272 11212 26312
rect 11252 26272 11261 26312
rect 11203 26271 11261 26272
rect 11395 26312 11453 26313
rect 11395 26272 11404 26312
rect 11444 26272 11453 26312
rect 11395 26271 11453 26272
rect 14755 26312 14813 26313
rect 14755 26272 14764 26312
rect 14804 26272 14813 26312
rect 14755 26271 14813 26272
rect 21091 26312 21149 26313
rect 21091 26272 21100 26312
rect 21140 26272 21149 26312
rect 21091 26271 21149 26272
rect 25987 26312 26045 26313
rect 25987 26272 25996 26312
rect 26036 26272 26045 26312
rect 25987 26271 26045 26272
rect 29155 26312 29213 26313
rect 29155 26272 29164 26312
rect 29204 26272 29213 26312
rect 29155 26271 29213 26272
rect 35491 26312 35549 26313
rect 35491 26272 35500 26312
rect 35540 26272 35549 26312
rect 35491 26271 35549 26272
rect 36555 26312 36597 26321
rect 36555 26272 36556 26312
rect 36596 26272 36597 26312
rect 36555 26263 36597 26272
rect 38371 26312 38429 26313
rect 38371 26272 38380 26312
rect 38420 26272 38429 26312
rect 38371 26271 38429 26272
rect 39043 26312 39101 26313
rect 39043 26272 39052 26312
rect 39092 26272 39101 26312
rect 39043 26271 39101 26272
rect 42795 26312 42837 26321
rect 42795 26272 42796 26312
rect 42836 26272 42837 26312
rect 42795 26263 42837 26272
rect 47395 26312 47453 26313
rect 47395 26272 47404 26312
rect 47444 26272 47453 26312
rect 47395 26271 47453 26272
rect 48931 26312 48989 26313
rect 48931 26272 48940 26312
rect 48980 26272 48989 26312
rect 48931 26271 48989 26272
rect 51235 26312 51293 26313
rect 51235 26272 51244 26312
rect 51284 26272 51293 26312
rect 51235 26271 51293 26272
rect 1707 26228 1749 26237
rect 1707 26188 1708 26228
rect 1748 26188 1749 26228
rect 1707 26179 1749 26188
rect 8811 26228 8853 26237
rect 8811 26188 8812 26228
rect 8852 26188 8853 26228
rect 8811 26179 8853 26188
rect 17643 26228 17685 26237
rect 17643 26188 17644 26228
rect 17684 26188 17685 26228
rect 17643 26179 17685 26188
rect 20139 26228 20181 26237
rect 20139 26188 20140 26228
rect 20180 26188 20181 26228
rect 20139 26179 20181 26188
rect 37323 26228 37365 26237
rect 37323 26188 37324 26228
rect 37364 26188 37365 26228
rect 37323 26179 37365 26188
rect 37803 26228 37845 26237
rect 37803 26188 37804 26228
rect 37844 26188 37845 26228
rect 37803 26179 37845 26188
rect 41931 26228 41973 26237
rect 41931 26188 41932 26228
rect 41972 26188 41973 26228
rect 41931 26179 41973 26188
rect 44235 26228 44277 26237
rect 44235 26188 44236 26228
rect 44276 26188 44277 26228
rect 44235 26179 44277 26188
rect 45003 26228 45045 26237
rect 45003 26188 45004 26228
rect 45044 26188 45045 26228
rect 45003 26179 45045 26188
rect 2083 26144 2141 26145
rect 2083 26104 2092 26144
rect 2132 26104 2141 26144
rect 2083 26103 2141 26104
rect 2947 26144 3005 26145
rect 2947 26104 2956 26144
rect 2996 26104 3005 26144
rect 2947 26103 3005 26104
rect 4387 26144 4445 26145
rect 4387 26104 4396 26144
rect 4436 26104 4445 26144
rect 4387 26103 4445 26104
rect 4683 26144 4725 26153
rect 4683 26104 4684 26144
rect 4724 26104 4725 26144
rect 4683 26095 4725 26104
rect 5347 26144 5405 26145
rect 5347 26104 5356 26144
rect 5396 26104 5405 26144
rect 5347 26103 5405 26104
rect 5827 26144 5885 26145
rect 5827 26104 5836 26144
rect 5876 26104 5885 26144
rect 5827 26103 5885 26104
rect 6123 26144 6165 26153
rect 6123 26104 6124 26144
rect 6164 26104 6165 26144
rect 6123 26095 6165 26104
rect 6219 26144 6261 26153
rect 6219 26104 6220 26144
rect 6260 26104 6261 26144
rect 6219 26095 6261 26104
rect 6883 26144 6941 26145
rect 6883 26104 6892 26144
rect 6932 26104 6941 26144
rect 6883 26103 6941 26104
rect 7755 26144 7797 26153
rect 7755 26104 7756 26144
rect 7796 26104 7797 26144
rect 7755 26095 7797 26104
rect 7947 26144 7989 26153
rect 7947 26104 7948 26144
rect 7988 26104 7989 26144
rect 7947 26095 7989 26104
rect 8035 26144 8093 26145
rect 8035 26104 8044 26144
rect 8084 26104 8093 26144
rect 8035 26103 8093 26104
rect 9187 26144 9245 26145
rect 9187 26104 9196 26144
rect 9236 26104 9245 26144
rect 9187 26103 9245 26104
rect 10051 26144 10109 26145
rect 10051 26104 10060 26144
rect 10100 26104 10109 26144
rect 10051 26103 10109 26104
rect 12067 26144 12125 26145
rect 12067 26104 12076 26144
rect 12116 26104 12125 26144
rect 12067 26103 12125 26104
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13803 26144 13845 26153
rect 13803 26104 13804 26144
rect 13844 26104 13845 26144
rect 13803 26095 13845 26104
rect 13891 26144 13949 26145
rect 13891 26104 13900 26144
rect 13940 26104 13949 26144
rect 13891 26103 13949 26104
rect 14083 26144 14141 26145
rect 14083 26104 14092 26144
rect 14132 26104 14141 26144
rect 14083 26103 14141 26104
rect 14187 26144 14229 26153
rect 14187 26104 14188 26144
rect 14228 26104 14229 26144
rect 14187 26095 14229 26104
rect 14379 26144 14421 26153
rect 14379 26104 14380 26144
rect 14420 26104 14421 26144
rect 14379 26095 14421 26104
rect 14563 26144 14621 26145
rect 14563 26104 14572 26144
rect 14612 26104 14621 26144
rect 14563 26103 14621 26104
rect 14667 26144 14709 26153
rect 14667 26104 14668 26144
rect 14708 26104 14709 26144
rect 14667 26095 14709 26104
rect 14859 26144 14901 26153
rect 14859 26104 14860 26144
rect 14900 26104 14901 26144
rect 14859 26095 14901 26104
rect 15243 26144 15285 26153
rect 15243 26104 15244 26144
rect 15284 26104 15285 26144
rect 15243 26095 15285 26104
rect 15339 26144 15381 26153
rect 15339 26104 15340 26144
rect 15380 26104 15381 26144
rect 15339 26095 15381 26104
rect 15427 26144 15485 26145
rect 15427 26104 15436 26144
rect 15476 26104 15485 26144
rect 15427 26103 15485 26104
rect 15715 26144 15773 26145
rect 15715 26104 15724 26144
rect 15764 26104 15773 26144
rect 15715 26103 15773 26104
rect 15811 26144 15869 26145
rect 15811 26104 15820 26144
rect 15860 26104 15869 26144
rect 15811 26103 15869 26104
rect 16011 26144 16053 26153
rect 16011 26104 16012 26144
rect 16052 26104 16053 26144
rect 16011 26095 16053 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16107 26095 16149 26104
rect 16200 26144 16258 26145
rect 16200 26104 16209 26144
rect 16249 26104 16258 26144
rect 16200 26103 16258 26104
rect 16587 26144 16629 26153
rect 16587 26104 16588 26144
rect 16628 26104 16629 26144
rect 16587 26095 16629 26104
rect 16683 26144 16725 26153
rect 16683 26104 16684 26144
rect 16724 26104 16725 26144
rect 16683 26095 16725 26104
rect 16779 26144 16821 26153
rect 16779 26104 16780 26144
rect 16820 26104 16821 26144
rect 16779 26095 16821 26104
rect 16875 26144 16917 26153
rect 16875 26104 16876 26144
rect 16916 26104 16917 26144
rect 16875 26095 16917 26104
rect 17067 26144 17109 26153
rect 17067 26104 17068 26144
rect 17108 26104 17109 26144
rect 17067 26095 17109 26104
rect 17163 26144 17205 26153
rect 17163 26104 17164 26144
rect 17204 26104 17205 26144
rect 17163 26095 17205 26104
rect 17259 26144 17301 26153
rect 17259 26104 17260 26144
rect 17300 26104 17301 26144
rect 17259 26095 17301 26104
rect 17355 26144 17397 26153
rect 17355 26104 17356 26144
rect 17396 26104 17397 26144
rect 17355 26095 17397 26104
rect 17547 26144 17589 26153
rect 17547 26104 17548 26144
rect 17588 26104 17589 26144
rect 17547 26095 17589 26104
rect 17739 26144 17781 26153
rect 17739 26104 17740 26144
rect 17780 26104 17781 26144
rect 17739 26095 17781 26104
rect 17827 26144 17885 26145
rect 17827 26104 17836 26144
rect 17876 26104 17885 26144
rect 17827 26103 17885 26104
rect 18691 26144 18749 26145
rect 18691 26104 18700 26144
rect 18740 26104 18749 26144
rect 18691 26103 18749 26104
rect 19075 26144 19133 26145
rect 19075 26104 19084 26144
rect 19124 26104 19133 26144
rect 19075 26103 19133 26104
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19467 26144 19509 26153
rect 19467 26104 19468 26144
rect 19508 26104 19509 26144
rect 19467 26095 19509 26104
rect 19939 26144 19997 26145
rect 19939 26104 19948 26144
rect 19988 26104 19997 26144
rect 19939 26103 19997 26104
rect 20043 26144 20085 26153
rect 20043 26104 20044 26144
rect 20084 26104 20085 26144
rect 20043 26095 20085 26104
rect 20235 26144 20277 26153
rect 20235 26104 20236 26144
rect 20276 26104 20277 26144
rect 20235 26095 20277 26104
rect 20419 26144 20477 26145
rect 20419 26104 20428 26144
rect 20468 26104 20477 26144
rect 20419 26103 20477 26104
rect 21955 26144 22013 26145
rect 21955 26104 21964 26144
rect 22004 26104 22013 26144
rect 21955 26103 22013 26104
rect 22155 26144 22197 26153
rect 22155 26104 22156 26144
rect 22196 26104 22197 26144
rect 22155 26095 22197 26104
rect 23595 26144 23637 26153
rect 23595 26104 23596 26144
rect 23636 26104 23637 26144
rect 23595 26095 23637 26104
rect 23971 26144 24029 26145
rect 23971 26104 23980 26144
rect 24020 26104 24029 26144
rect 23971 26103 24029 26104
rect 24835 26144 24893 26145
rect 24835 26104 24844 26144
rect 24884 26104 24893 26144
rect 24835 26103 24893 26104
rect 26379 26144 26421 26153
rect 26379 26104 26380 26144
rect 26420 26104 26421 26144
rect 26379 26095 26421 26104
rect 26475 26144 26517 26153
rect 26475 26104 26476 26144
rect 26516 26104 26517 26144
rect 26475 26095 26517 26104
rect 26571 26144 26613 26153
rect 26571 26104 26572 26144
rect 26612 26104 26613 26144
rect 26571 26095 26613 26104
rect 26667 26144 26709 26153
rect 26667 26104 26668 26144
rect 26708 26104 26709 26144
rect 26667 26095 26709 26104
rect 26947 26144 27005 26145
rect 26947 26104 26956 26144
rect 26996 26104 27005 26144
rect 26947 26103 27005 26104
rect 27907 26144 27965 26145
rect 27907 26104 27916 26144
rect 27956 26104 27965 26144
rect 27907 26103 27965 26104
rect 28483 26144 28541 26145
rect 28483 26104 28492 26144
rect 28532 26104 28541 26144
rect 28483 26103 28541 26104
rect 28587 26139 28629 26148
rect 28587 26099 28588 26139
rect 28628 26099 28629 26139
rect 28675 26144 28733 26145
rect 28675 26104 28684 26144
rect 28724 26104 28733 26144
rect 28675 26103 28733 26104
rect 29067 26144 29109 26153
rect 29067 26104 29068 26144
rect 29108 26104 29109 26144
rect 28587 26090 28629 26099
rect 29067 26095 29109 26104
rect 29259 26144 29301 26153
rect 29259 26104 29260 26144
rect 29300 26104 29301 26144
rect 29259 26095 29301 26104
rect 29347 26144 29405 26145
rect 29347 26104 29356 26144
rect 29396 26104 29405 26144
rect 29347 26103 29405 26104
rect 29643 26144 29685 26153
rect 29643 26104 29644 26144
rect 29684 26104 29685 26144
rect 29643 26095 29685 26104
rect 29835 26144 29877 26153
rect 29835 26104 29836 26144
rect 29876 26104 29877 26144
rect 29835 26095 29877 26104
rect 29923 26144 29981 26145
rect 29923 26104 29932 26144
rect 29972 26104 29981 26144
rect 29923 26103 29981 26104
rect 30603 26144 30645 26153
rect 30603 26104 30604 26144
rect 30644 26104 30645 26144
rect 30603 26095 30645 26104
rect 30691 26144 30749 26145
rect 30691 26104 30700 26144
rect 30740 26104 30749 26144
rect 31563 26144 31605 26153
rect 30691 26103 30749 26104
rect 31371 26133 31413 26142
rect 31371 26093 31372 26133
rect 31412 26093 31413 26133
rect 31563 26104 31564 26144
rect 31604 26104 31605 26144
rect 31563 26095 31605 26104
rect 31651 26144 31709 26145
rect 31651 26104 31660 26144
rect 31700 26104 31709 26144
rect 31651 26103 31709 26104
rect 31843 26144 31901 26145
rect 31843 26104 31852 26144
rect 31892 26104 31901 26144
rect 31843 26103 31901 26104
rect 32803 26144 32861 26145
rect 32803 26104 32812 26144
rect 32852 26104 32861 26144
rect 32803 26103 32861 26104
rect 33091 26144 33149 26145
rect 33091 26104 33100 26144
rect 33140 26104 33149 26144
rect 33091 26103 33149 26104
rect 33963 26144 34005 26153
rect 33963 26104 33964 26144
rect 34004 26104 34005 26144
rect 33963 26095 34005 26104
rect 35011 26144 35069 26145
rect 35011 26104 35020 26144
rect 35060 26104 35069 26144
rect 35011 26103 35069 26104
rect 35211 26144 35253 26153
rect 35211 26104 35212 26144
rect 35252 26104 35253 26144
rect 35211 26095 35253 26104
rect 35307 26144 35349 26153
rect 35307 26104 35308 26144
rect 35348 26104 35349 26144
rect 35307 26095 35349 26104
rect 35403 26144 35445 26153
rect 35403 26104 35404 26144
rect 35444 26104 35445 26144
rect 35403 26095 35445 26104
rect 36171 26144 36213 26153
rect 36171 26104 36172 26144
rect 36212 26104 36213 26144
rect 36171 26095 36213 26104
rect 37027 26144 37085 26145
rect 37027 26104 37036 26144
rect 37076 26104 37085 26144
rect 37027 26103 37085 26104
rect 37219 26144 37277 26145
rect 37219 26104 37228 26144
rect 37268 26104 37277 26144
rect 37219 26103 37277 26104
rect 37419 26144 37461 26153
rect 37419 26104 37420 26144
rect 37460 26104 37461 26144
rect 37419 26095 37461 26104
rect 37899 26144 37941 26153
rect 37899 26104 37900 26144
rect 37940 26104 37941 26144
rect 37899 26095 37941 26104
rect 37995 26144 38037 26153
rect 37995 26104 37996 26144
rect 38036 26104 38037 26144
rect 37995 26095 38037 26104
rect 38091 26144 38133 26153
rect 38091 26104 38092 26144
rect 38132 26104 38133 26144
rect 38091 26095 38133 26104
rect 38283 26144 38325 26153
rect 38283 26104 38284 26144
rect 38324 26104 38325 26144
rect 38283 26095 38325 26104
rect 38475 26144 38517 26153
rect 38475 26104 38476 26144
rect 38516 26104 38517 26144
rect 38475 26095 38517 26104
rect 38563 26144 38621 26145
rect 38563 26104 38572 26144
rect 38612 26104 38621 26144
rect 38563 26103 38621 26104
rect 38763 26144 38805 26153
rect 38763 26104 38764 26144
rect 38804 26104 38805 26144
rect 38763 26095 38805 26104
rect 38859 26144 38901 26153
rect 38859 26104 38860 26144
rect 38900 26104 38901 26144
rect 38859 26095 38901 26104
rect 38955 26144 38997 26153
rect 38955 26104 38956 26144
rect 38996 26104 38997 26144
rect 38955 26095 38997 26104
rect 40483 26144 40541 26145
rect 40483 26104 40492 26144
rect 40532 26104 40541 26144
rect 40483 26103 40541 26104
rect 40587 26144 40629 26153
rect 40587 26104 40588 26144
rect 40628 26104 40629 26144
rect 40587 26095 40629 26104
rect 40779 26144 40821 26153
rect 40779 26104 40780 26144
rect 40820 26104 40821 26144
rect 40779 26095 40821 26104
rect 41163 26144 41205 26153
rect 41163 26104 41164 26144
rect 41204 26104 41205 26144
rect 41163 26095 41205 26104
rect 41259 26144 41301 26153
rect 41259 26104 41260 26144
rect 41300 26104 41301 26144
rect 41259 26095 41301 26104
rect 41355 26144 41397 26153
rect 41355 26104 41356 26144
rect 41396 26104 41397 26144
rect 41355 26095 41397 26104
rect 41451 26144 41493 26153
rect 41451 26104 41452 26144
rect 41492 26104 41493 26144
rect 41451 26095 41493 26104
rect 42027 26144 42069 26153
rect 42027 26104 42028 26144
rect 42068 26104 42069 26144
rect 42027 26095 42069 26104
rect 42307 26144 42365 26145
rect 42307 26104 42316 26144
rect 42356 26104 42365 26144
rect 42307 26103 42365 26104
rect 42883 26144 42941 26145
rect 42883 26104 42892 26144
rect 42932 26104 42941 26144
rect 42883 26103 42941 26104
rect 43083 26144 43125 26153
rect 43083 26104 43084 26144
rect 43124 26104 43125 26144
rect 43083 26095 43125 26104
rect 43747 26144 43805 26145
rect 43747 26104 43756 26144
rect 43796 26104 43805 26144
rect 43747 26103 43805 26104
rect 44331 26144 44373 26153
rect 44331 26104 44332 26144
rect 44372 26104 44373 26144
rect 44331 26095 44373 26104
rect 44611 26144 44669 26145
rect 44611 26104 44620 26144
rect 44660 26104 44669 26144
rect 44611 26103 44669 26104
rect 45379 26144 45437 26145
rect 45379 26104 45388 26144
rect 45428 26104 45437 26144
rect 45379 26103 45437 26104
rect 46243 26144 46301 26145
rect 46243 26104 46252 26144
rect 46292 26104 46301 26144
rect 46243 26103 46301 26104
rect 47779 26144 47837 26145
rect 47779 26104 47788 26144
rect 47828 26104 47837 26144
rect 48075 26144 48117 26153
rect 47779 26103 47837 26104
rect 47875 26130 47933 26131
rect 31371 26084 31413 26093
rect 47875 26090 47884 26130
rect 47924 26090 47933 26130
rect 48075 26104 48076 26144
rect 48116 26104 48117 26144
rect 48075 26095 48117 26104
rect 48259 26144 48317 26145
rect 48259 26104 48268 26144
rect 48308 26104 48317 26144
rect 48259 26103 48317 26104
rect 49123 26144 49181 26145
rect 49123 26104 49132 26144
rect 49172 26104 49181 26144
rect 49123 26103 49181 26104
rect 50755 26144 50813 26145
rect 50755 26104 50764 26144
rect 50804 26104 50813 26144
rect 50755 26103 50813 26104
rect 50955 26144 50997 26153
rect 50955 26104 50956 26144
rect 50996 26104 50997 26144
rect 50955 26095 50997 26104
rect 51051 26144 51093 26153
rect 51051 26104 51052 26144
rect 51092 26104 51093 26144
rect 51051 26095 51093 26104
rect 51147 26144 51189 26153
rect 51147 26104 51148 26144
rect 51188 26104 51189 26144
rect 51147 26095 51189 26104
rect 47875 26089 47933 26090
rect 4107 26060 4149 26069
rect 4107 26020 4108 26060
rect 4148 26020 4149 26060
rect 4107 26011 4149 26020
rect 1515 25976 1557 25985
rect 1515 25936 1516 25976
rect 1556 25936 1557 25976
rect 1515 25927 1557 25936
rect 6499 25976 6557 25977
rect 6499 25936 6508 25976
rect 6548 25936 6557 25976
rect 6499 25935 6557 25936
rect 7755 25976 7797 25985
rect 7755 25936 7756 25976
rect 7796 25936 7797 25976
rect 7755 25927 7797 25936
rect 8427 25976 8469 25985
rect 8427 25936 8428 25976
rect 8468 25936 8469 25976
rect 8427 25927 8469 25936
rect 12459 25976 12501 25985
rect 12459 25936 12460 25976
rect 12500 25936 12501 25976
rect 12459 25927 12501 25936
rect 19747 25976 19805 25977
rect 19747 25936 19756 25976
rect 19796 25936 19805 25976
rect 19747 25935 19805 25936
rect 21483 25976 21525 25985
rect 21483 25936 21484 25976
rect 21524 25936 21525 25976
rect 21483 25927 21525 25936
rect 31371 25976 31413 25985
rect 31371 25936 31372 25976
rect 31412 25936 31413 25976
rect 31371 25927 31413 25936
rect 40299 25976 40341 25985
rect 40299 25936 40300 25976
rect 40340 25936 40341 25976
rect 40299 25927 40341 25936
rect 41635 25976 41693 25977
rect 41635 25936 41644 25976
rect 41684 25936 41693 25976
rect 41635 25935 41693 25936
rect 43939 25976 43997 25977
rect 43939 25936 43948 25976
rect 43988 25936 43997 25976
rect 43939 25935 43997 25936
rect 48075 25976 48117 25985
rect 48075 25936 48076 25976
rect 48116 25936 48117 25976
rect 48075 25927 48117 25936
rect 51435 25976 51477 25985
rect 51435 25936 51436 25976
rect 51476 25936 51477 25976
rect 51435 25927 51477 25936
rect 4491 25892 4533 25901
rect 4491 25852 4492 25892
rect 4532 25852 4533 25892
rect 4491 25843 4533 25852
rect 7555 25892 7613 25893
rect 7555 25852 7564 25892
rect 7604 25852 7613 25892
rect 7555 25851 7613 25852
rect 13611 25892 13653 25901
rect 13611 25852 13612 25892
rect 13652 25852 13653 25892
rect 13611 25843 13653 25852
rect 14379 25892 14421 25901
rect 14379 25852 14380 25892
rect 14420 25852 14421 25892
rect 14379 25843 14421 25852
rect 15723 25892 15765 25901
rect 15723 25852 15724 25892
rect 15764 25852 15765 25892
rect 15723 25843 15765 25852
rect 18019 25892 18077 25893
rect 18019 25852 18028 25892
rect 18068 25852 18077 25892
rect 18019 25851 18077 25852
rect 22059 25892 22101 25901
rect 22059 25852 22060 25892
rect 22100 25852 22101 25892
rect 22059 25843 22101 25852
rect 27243 25892 27285 25901
rect 27243 25852 27244 25892
rect 27284 25852 27285 25892
rect 27243 25843 27285 25852
rect 28203 25892 28245 25901
rect 28203 25852 28204 25892
rect 28244 25852 28245 25892
rect 28203 25843 28245 25852
rect 29643 25892 29685 25901
rect 29643 25852 29644 25892
rect 29684 25852 29685 25892
rect 29643 25843 29685 25852
rect 30315 25892 30357 25901
rect 30315 25852 30316 25892
rect 30356 25852 30357 25892
rect 30315 25843 30357 25852
rect 34339 25892 34397 25893
rect 34339 25852 34348 25892
rect 34388 25852 34397 25892
rect 34339 25851 34397 25852
rect 40779 25892 40821 25901
rect 40779 25852 40780 25892
rect 40820 25852 40821 25892
rect 40779 25843 40821 25852
rect 49795 25892 49853 25893
rect 49795 25852 49804 25892
rect 49844 25852 49853 25892
rect 49795 25851 49853 25852
rect 50083 25892 50141 25893
rect 50083 25852 50092 25892
rect 50132 25852 50141 25892
rect 50083 25851 50141 25852
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 3427 25556 3485 25557
rect 3427 25516 3436 25556
rect 3476 25516 3485 25556
rect 3427 25515 3485 25516
rect 6315 25556 6357 25565
rect 6315 25516 6316 25556
rect 6356 25516 6357 25556
rect 6315 25507 6357 25516
rect 13707 25556 13749 25565
rect 13707 25516 13708 25556
rect 13748 25516 13749 25556
rect 13707 25507 13749 25516
rect 15243 25556 15285 25565
rect 15243 25516 15244 25556
rect 15284 25516 15285 25556
rect 15243 25507 15285 25516
rect 17835 25556 17877 25565
rect 17835 25516 17836 25556
rect 17876 25516 17877 25556
rect 17835 25507 17877 25516
rect 20419 25556 20477 25557
rect 20419 25516 20428 25556
rect 20468 25516 20477 25556
rect 20419 25515 20477 25516
rect 20619 25556 20661 25565
rect 20619 25516 20620 25556
rect 20660 25516 20661 25556
rect 20619 25507 20661 25516
rect 27915 25556 27957 25565
rect 27915 25516 27916 25556
rect 27956 25516 27957 25556
rect 27915 25507 27957 25516
rect 32043 25556 32085 25565
rect 32043 25516 32044 25556
rect 32084 25516 32085 25556
rect 32043 25507 32085 25516
rect 36171 25556 36213 25565
rect 36171 25516 36172 25556
rect 36212 25516 36213 25556
rect 36171 25507 36213 25516
rect 39339 25556 39381 25565
rect 39339 25516 39340 25556
rect 39380 25516 39381 25556
rect 39339 25507 39381 25516
rect 42691 25556 42749 25557
rect 42691 25516 42700 25556
rect 42740 25516 42749 25556
rect 42691 25515 42749 25516
rect 43755 25556 43797 25565
rect 43755 25516 43756 25556
rect 43796 25516 43797 25556
rect 43755 25507 43797 25516
rect 11883 25472 11925 25481
rect 11883 25432 11884 25472
rect 11924 25432 11925 25472
rect 11883 25423 11925 25432
rect 16395 25472 16437 25481
rect 16395 25432 16396 25472
rect 16436 25432 16437 25472
rect 16395 25423 16437 25432
rect 22635 25472 22677 25481
rect 22635 25432 22636 25472
rect 22676 25432 22677 25472
rect 22635 25423 22677 25432
rect 30507 25472 30549 25481
rect 30507 25432 30508 25472
rect 30548 25432 30549 25472
rect 30507 25423 30549 25432
rect 45099 25472 45141 25481
rect 45099 25432 45100 25472
rect 45140 25432 45141 25472
rect 45099 25423 45141 25432
rect 9291 25388 9333 25397
rect 9291 25348 9292 25388
rect 9332 25348 9333 25388
rect 9291 25339 9333 25348
rect 12651 25388 12693 25397
rect 12651 25348 12652 25388
rect 12692 25348 12693 25388
rect 26851 25388 26909 25389
rect 26851 25348 26860 25388
rect 26900 25348 26909 25388
rect 12651 25339 12693 25348
rect 22251 25339 22293 25348
rect 12739 25327 12797 25328
rect 1411 25304 1469 25305
rect 1411 25264 1420 25304
rect 1460 25264 1469 25304
rect 1411 25263 1469 25264
rect 2275 25304 2333 25305
rect 2275 25264 2284 25304
rect 2324 25264 2333 25304
rect 2275 25263 2333 25264
rect 4291 25304 4349 25305
rect 4291 25264 4300 25304
rect 4340 25264 4349 25304
rect 4291 25263 4349 25264
rect 4579 25304 4637 25305
rect 4579 25264 4588 25304
rect 4628 25264 4637 25304
rect 4579 25263 4637 25264
rect 5451 25304 5493 25313
rect 5451 25264 5452 25304
rect 5492 25264 5493 25304
rect 5451 25255 5493 25264
rect 5923 25304 5981 25305
rect 5923 25264 5932 25304
rect 5972 25264 5981 25304
rect 5923 25263 5981 25264
rect 6027 25304 6069 25313
rect 6027 25264 6028 25304
rect 6068 25264 6069 25304
rect 6027 25255 6069 25264
rect 7843 25304 7901 25305
rect 7843 25264 7852 25304
rect 7892 25264 7901 25304
rect 7843 25263 7901 25264
rect 8707 25304 8765 25305
rect 8707 25264 8716 25304
rect 8756 25264 8765 25304
rect 8707 25263 8765 25264
rect 9099 25304 9141 25313
rect 9099 25264 9100 25304
rect 9140 25264 9141 25304
rect 9099 25255 9141 25264
rect 9379 25304 9437 25305
rect 9379 25264 9388 25304
rect 9428 25264 9437 25304
rect 9379 25263 9437 25264
rect 9667 25304 9725 25305
rect 9667 25264 9676 25304
rect 9716 25264 9725 25304
rect 9667 25263 9725 25264
rect 9963 25304 10005 25313
rect 9963 25264 9964 25304
rect 10004 25264 10005 25304
rect 9963 25255 10005 25264
rect 10059 25304 10101 25313
rect 10059 25264 10060 25304
rect 10100 25264 10101 25304
rect 10059 25255 10101 25264
rect 10155 25304 10197 25313
rect 10155 25264 10156 25304
rect 10196 25264 10197 25304
rect 10155 25255 10197 25264
rect 10539 25304 10581 25313
rect 10539 25264 10540 25304
rect 10580 25264 10581 25304
rect 10539 25255 10581 25264
rect 10635 25304 10677 25313
rect 10635 25264 10636 25304
rect 10676 25264 10677 25304
rect 10635 25255 10677 25264
rect 10731 25304 10773 25313
rect 10731 25264 10732 25304
rect 10772 25264 10773 25304
rect 10731 25255 10773 25264
rect 10827 25304 10869 25313
rect 10827 25264 10828 25304
rect 10868 25264 10869 25304
rect 10827 25255 10869 25264
rect 11011 25304 11069 25305
rect 11011 25264 11020 25304
rect 11060 25264 11069 25304
rect 11011 25263 11069 25264
rect 11883 25304 11925 25313
rect 11883 25264 11884 25304
rect 11924 25264 11925 25304
rect 11883 25255 11925 25264
rect 12075 25304 12117 25313
rect 12075 25264 12076 25304
rect 12116 25264 12117 25304
rect 12075 25255 12117 25264
rect 12163 25304 12221 25305
rect 12163 25264 12172 25304
rect 12212 25264 12221 25304
rect 12163 25263 12221 25264
rect 12555 25304 12597 25313
rect 12555 25264 12556 25304
rect 12596 25264 12597 25304
rect 12739 25287 12748 25327
rect 12788 25287 12797 25327
rect 12739 25286 12797 25287
rect 13214 25304 13272 25305
rect 12555 25255 12597 25264
rect 13214 25264 13223 25304
rect 13263 25264 13272 25304
rect 13214 25263 13272 25264
rect 13323 25304 13365 25313
rect 13323 25264 13324 25304
rect 13364 25264 13365 25304
rect 13323 25255 13365 25264
rect 13419 25304 13461 25313
rect 13419 25264 13420 25304
rect 13460 25264 13461 25304
rect 13419 25255 13461 25264
rect 13603 25304 13661 25305
rect 13603 25264 13612 25304
rect 13652 25264 13661 25304
rect 13603 25263 13661 25264
rect 13699 25304 13757 25305
rect 13699 25264 13708 25304
rect 13748 25264 13757 25304
rect 13699 25263 13757 25264
rect 13891 25304 13949 25305
rect 13891 25264 13900 25304
rect 13940 25264 13949 25304
rect 13891 25263 13949 25264
rect 14947 25304 15005 25305
rect 14947 25264 14956 25304
rect 14996 25264 15005 25304
rect 14947 25263 15005 25264
rect 15051 25304 15093 25313
rect 15051 25264 15052 25304
rect 15092 25264 15093 25304
rect 15051 25255 15093 25264
rect 15243 25304 15285 25313
rect 15243 25264 15244 25304
rect 15284 25264 15285 25304
rect 15243 25255 15285 25264
rect 16099 25304 16157 25305
rect 16099 25264 16108 25304
rect 16148 25264 16157 25304
rect 16099 25263 16157 25264
rect 16203 25304 16245 25313
rect 16203 25264 16204 25304
rect 16244 25264 16245 25304
rect 16203 25255 16245 25264
rect 16395 25304 16437 25313
rect 16395 25264 16396 25304
rect 16436 25264 16437 25304
rect 16395 25255 16437 25264
rect 17539 25304 17597 25305
rect 17539 25264 17548 25304
rect 17588 25264 17597 25304
rect 17539 25263 17597 25264
rect 17643 25304 17685 25313
rect 17643 25264 17644 25304
rect 17684 25264 17685 25304
rect 17643 25255 17685 25264
rect 17835 25304 17877 25313
rect 17835 25264 17836 25304
rect 17876 25264 17877 25304
rect 17835 25255 17877 25264
rect 18027 25304 18069 25313
rect 18027 25264 18028 25304
rect 18068 25264 18069 25304
rect 18027 25255 18069 25264
rect 18403 25304 18461 25305
rect 18403 25264 18412 25304
rect 18452 25264 18461 25304
rect 18403 25263 18461 25264
rect 19267 25304 19325 25305
rect 19267 25264 19276 25304
rect 19316 25264 19325 25304
rect 19267 25263 19325 25264
rect 20707 25304 20765 25305
rect 20707 25264 20716 25304
rect 20756 25264 20765 25304
rect 20707 25263 20765 25264
rect 20907 25304 20949 25313
rect 20907 25264 20908 25304
rect 20948 25264 20949 25304
rect 20907 25255 20949 25264
rect 21571 25304 21629 25305
rect 21571 25264 21580 25304
rect 21620 25264 21629 25304
rect 21571 25263 21629 25264
rect 22147 25304 22205 25305
rect 22147 25264 22156 25304
rect 22196 25264 22205 25304
rect 22251 25299 22252 25339
rect 22292 25299 22293 25339
rect 26571 25339 26613 25348
rect 26851 25347 26909 25348
rect 37611 25388 37653 25397
rect 37611 25348 37612 25388
rect 37652 25348 37653 25388
rect 37611 25339 37653 25348
rect 37707 25388 37749 25397
rect 37707 25348 37708 25388
rect 37748 25348 37749 25388
rect 37707 25339 37749 25348
rect 46923 25388 46965 25397
rect 46923 25348 46924 25388
rect 46964 25348 46965 25388
rect 46923 25339 46965 25348
rect 47019 25388 47061 25397
rect 47019 25348 47020 25388
rect 47060 25348 47061 25388
rect 47019 25339 47061 25348
rect 49419 25388 49461 25397
rect 49419 25348 49420 25388
rect 49460 25348 49461 25388
rect 49419 25339 49461 25348
rect 23595 25309 23637 25318
rect 22251 25290 22293 25299
rect 22339 25304 22397 25305
rect 22147 25263 22205 25264
rect 22339 25264 22348 25304
rect 22388 25264 22397 25304
rect 22339 25263 22397 25264
rect 22723 25304 22781 25305
rect 22723 25264 22732 25304
rect 22772 25264 22781 25304
rect 22723 25263 22781 25264
rect 23491 25304 23549 25305
rect 23491 25264 23500 25304
rect 23540 25264 23549 25304
rect 23491 25263 23549 25264
rect 23595 25269 23596 25309
rect 23636 25269 23637 25309
rect 23595 25260 23637 25269
rect 23683 25304 23741 25305
rect 23683 25264 23692 25304
rect 23732 25264 23741 25304
rect 23683 25263 23741 25264
rect 24651 25304 24693 25313
rect 24651 25264 24652 25304
rect 24692 25264 24693 25304
rect 24651 25255 24693 25264
rect 24843 25304 24885 25313
rect 24843 25264 24844 25304
rect 24884 25264 24885 25304
rect 24843 25255 24885 25264
rect 24931 25304 24989 25305
rect 24931 25264 24940 25304
rect 24980 25264 24989 25304
rect 24931 25263 24989 25264
rect 26467 25304 26525 25305
rect 26467 25264 26476 25304
rect 26516 25264 26525 25304
rect 26571 25299 26572 25339
rect 26612 25299 26613 25339
rect 36651 25318 36693 25327
rect 26571 25290 26613 25299
rect 26659 25304 26717 25305
rect 26467 25263 26525 25264
rect 26659 25264 26668 25304
rect 26708 25264 26717 25304
rect 26659 25263 26717 25264
rect 27235 25304 27293 25305
rect 27235 25264 27244 25304
rect 27284 25264 27293 25304
rect 27235 25263 27293 25264
rect 28195 25304 28253 25305
rect 28195 25264 28204 25304
rect 28244 25264 28253 25304
rect 28195 25263 28253 25264
rect 28867 25304 28925 25305
rect 28867 25264 28876 25304
rect 28916 25264 28925 25304
rect 28867 25263 28925 25264
rect 29827 25304 29885 25305
rect 29827 25264 29836 25304
rect 29876 25264 29885 25304
rect 29827 25263 29885 25264
rect 30315 25304 30357 25313
rect 30315 25264 30316 25304
rect 30356 25264 30357 25304
rect 30315 25255 30357 25264
rect 32619 25304 32661 25313
rect 32619 25264 32620 25304
rect 32660 25264 32661 25304
rect 32619 25255 32661 25264
rect 33003 25304 33045 25313
rect 33003 25264 33004 25304
rect 33044 25264 33045 25304
rect 33003 25255 33045 25264
rect 33379 25304 33437 25305
rect 33379 25264 33388 25304
rect 33428 25264 33437 25304
rect 33379 25263 33437 25264
rect 34243 25304 34301 25305
rect 34243 25264 34252 25304
rect 34292 25264 34301 25304
rect 34243 25263 34301 25264
rect 35595 25304 35637 25313
rect 35595 25264 35596 25304
rect 35636 25264 35637 25304
rect 35595 25255 35637 25264
rect 35691 25304 35733 25313
rect 35691 25264 35692 25304
rect 35732 25264 35733 25304
rect 35691 25255 35733 25264
rect 35787 25304 35829 25313
rect 35787 25264 35788 25304
rect 35828 25264 35829 25304
rect 35787 25255 35829 25264
rect 35883 25304 35925 25313
rect 35883 25264 35884 25304
rect 35924 25264 35925 25304
rect 35883 25255 35925 25264
rect 36259 25304 36317 25305
rect 36259 25264 36268 25304
rect 36308 25264 36317 25304
rect 36651 25278 36652 25318
rect 36692 25278 36693 25318
rect 45963 25318 46005 25327
rect 36651 25269 36693 25278
rect 37123 25304 37181 25305
rect 36259 25263 36317 25264
rect 37123 25264 37132 25304
rect 37172 25264 37181 25304
rect 37123 25263 37181 25264
rect 38091 25304 38133 25313
rect 38091 25264 38092 25304
rect 38132 25264 38133 25304
rect 38091 25255 38133 25264
rect 38187 25304 38229 25313
rect 38187 25264 38188 25304
rect 38228 25264 38229 25304
rect 38187 25255 38229 25264
rect 39147 25304 39189 25313
rect 39147 25264 39148 25304
rect 39188 25264 39189 25304
rect 39147 25255 39189 25264
rect 40299 25304 40341 25313
rect 40299 25264 40300 25304
rect 40340 25264 40341 25304
rect 40299 25255 40341 25264
rect 40675 25304 40733 25305
rect 40675 25264 40684 25304
rect 40724 25264 40733 25304
rect 40675 25263 40733 25264
rect 41539 25304 41597 25305
rect 41539 25264 41548 25304
rect 41588 25264 41597 25304
rect 41539 25263 41597 25264
rect 42883 25304 42941 25305
rect 42883 25264 42892 25304
rect 42932 25264 42941 25304
rect 42883 25263 42941 25264
rect 43843 25304 43901 25305
rect 43843 25264 43852 25304
rect 43892 25264 43901 25304
rect 43843 25263 43901 25264
rect 44523 25304 44565 25313
rect 44523 25264 44524 25304
rect 44564 25264 44565 25304
rect 44523 25255 44565 25264
rect 44619 25304 44661 25313
rect 44619 25264 44620 25304
rect 44660 25264 44661 25304
rect 44619 25255 44661 25264
rect 44715 25304 44757 25313
rect 44715 25264 44716 25304
rect 44756 25264 44757 25304
rect 44715 25255 44757 25264
rect 44811 25304 44853 25313
rect 44811 25264 44812 25304
rect 44852 25264 44853 25304
rect 44811 25255 44853 25264
rect 45571 25304 45629 25305
rect 45571 25264 45580 25304
rect 45620 25264 45629 25304
rect 45963 25278 45964 25318
rect 46004 25278 46005 25318
rect 45963 25269 46005 25278
rect 46435 25304 46493 25305
rect 45571 25263 45629 25264
rect 46435 25264 46444 25304
rect 46484 25264 46493 25304
rect 46435 25263 46493 25264
rect 47403 25304 47445 25313
rect 47403 25264 47404 25304
rect 47444 25264 47445 25304
rect 47403 25255 47445 25264
rect 47499 25304 47541 25313
rect 47499 25264 47500 25304
rect 47540 25264 47541 25304
rect 47499 25255 47541 25264
rect 47787 25304 47829 25313
rect 47787 25264 47788 25304
rect 47828 25264 47829 25304
rect 47787 25255 47829 25264
rect 47875 25304 47933 25305
rect 47875 25264 47884 25304
rect 47924 25264 47933 25304
rect 47875 25263 47933 25264
rect 48075 25304 48117 25313
rect 48075 25264 48076 25304
rect 48116 25264 48117 25304
rect 48075 25255 48117 25264
rect 48171 25304 48213 25313
rect 48171 25264 48172 25304
rect 48212 25264 48213 25304
rect 48171 25255 48213 25264
rect 48267 25304 48309 25313
rect 48267 25264 48268 25304
rect 48308 25264 48309 25304
rect 48267 25255 48309 25264
rect 48547 25304 48605 25305
rect 48547 25264 48556 25304
rect 48596 25264 48605 25304
rect 48547 25263 48605 25264
rect 50563 25304 50621 25305
rect 50563 25264 50572 25304
rect 50612 25264 50621 25304
rect 50563 25263 50621 25264
rect 51427 25304 51485 25305
rect 51427 25264 51436 25304
rect 51476 25264 51485 25304
rect 51427 25263 51485 25264
rect 51819 25304 51861 25313
rect 51819 25264 51820 25304
rect 51860 25264 51861 25304
rect 51819 25255 51861 25264
rect 1035 25220 1077 25229
rect 1035 25180 1036 25220
rect 1076 25180 1077 25220
rect 1035 25171 1077 25180
rect 3627 25220 3669 25229
rect 3627 25180 3628 25220
rect 3668 25180 3669 25220
rect 3627 25171 3669 25180
rect 24747 25220 24789 25229
rect 24747 25180 24748 25220
rect 24788 25180 24789 25220
rect 24747 25171 24789 25180
rect 26187 25220 26229 25229
rect 26187 25180 26188 25220
rect 26228 25180 26229 25220
rect 26187 25171 26229 25180
rect 36459 25220 36501 25229
rect 36459 25180 36460 25220
rect 36500 25180 36501 25220
rect 36459 25171 36501 25180
rect 43563 25220 43605 25229
rect 43563 25180 43564 25220
rect 43604 25180 43605 25220
rect 43563 25171 43605 25180
rect 45771 25220 45813 25229
rect 45771 25180 45772 25220
rect 45812 25180 45813 25220
rect 45771 25171 45813 25180
rect 6691 25136 6749 25137
rect 6691 25096 6700 25136
rect 6740 25096 6749 25136
rect 6691 25095 6749 25096
rect 9579 25136 9621 25145
rect 9579 25096 9580 25136
rect 9620 25096 9621 25136
rect 9579 25087 9621 25096
rect 9859 25136 9917 25137
rect 9859 25096 9868 25136
rect 9908 25096 9917 25136
rect 9859 25095 9917 25096
rect 11683 25136 11741 25137
rect 11683 25096 11692 25136
rect 11732 25096 11741 25136
rect 11683 25095 11741 25096
rect 14563 25136 14621 25137
rect 14563 25096 14572 25136
rect 14612 25096 14621 25136
rect 14563 25095 14621 25096
rect 21867 25136 21909 25145
rect 21867 25096 21868 25136
rect 21908 25096 21909 25136
rect 21867 25087 21909 25096
rect 23211 25136 23253 25145
rect 23211 25096 23212 25136
rect 23252 25096 23253 25136
rect 23211 25087 23253 25096
rect 35395 25136 35453 25137
rect 35395 25096 35404 25136
rect 35444 25096 35453 25136
rect 35395 25095 35453 25096
rect 45483 25136 45525 25145
rect 45483 25096 45484 25136
rect 45524 25096 45525 25136
rect 45483 25087 45525 25096
rect 48355 25136 48413 25137
rect 48355 25096 48364 25136
rect 48404 25096 48413 25136
rect 48355 25095 48413 25096
rect 49219 25136 49277 25137
rect 49219 25096 49228 25136
rect 49268 25096 49277 25136
rect 49219 25095 49277 25096
rect 5835 25078 5877 25087
rect 5835 25038 5836 25078
rect 5876 25038 5877 25078
rect 5835 25029 5877 25038
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 843 24800 885 24809
rect 843 24760 844 24800
rect 884 24760 885 24800
rect 843 24751 885 24760
rect 1987 24800 2045 24801
rect 1987 24760 1996 24800
rect 2036 24760 2045 24800
rect 1987 24759 2045 24760
rect 4195 24800 4253 24801
rect 4195 24760 4204 24800
rect 4244 24760 4253 24800
rect 4195 24759 4253 24760
rect 6691 24800 6749 24801
rect 6691 24760 6700 24800
rect 6740 24760 6749 24800
rect 6691 24759 6749 24760
rect 9667 24800 9725 24801
rect 9667 24760 9676 24800
rect 9716 24760 9725 24800
rect 9667 24759 9725 24760
rect 10819 24800 10877 24801
rect 10819 24760 10828 24800
rect 10868 24760 10877 24800
rect 10819 24759 10877 24760
rect 17067 24800 17109 24809
rect 17067 24760 17068 24800
rect 17108 24760 17109 24800
rect 17067 24751 17109 24760
rect 24075 24800 24117 24809
rect 24075 24760 24076 24800
rect 24116 24760 24117 24800
rect 24075 24751 24117 24760
rect 25323 24800 25365 24809
rect 25323 24760 25324 24800
rect 25364 24760 25365 24800
rect 25323 24751 25365 24760
rect 26379 24800 26421 24809
rect 26379 24760 26380 24800
rect 26420 24760 26421 24800
rect 26379 24751 26421 24760
rect 27043 24800 27101 24801
rect 27043 24760 27052 24800
rect 27092 24760 27101 24800
rect 27043 24759 27101 24760
rect 31275 24800 31317 24809
rect 31275 24760 31276 24800
rect 31316 24760 31317 24800
rect 31275 24751 31317 24760
rect 35395 24800 35453 24801
rect 35395 24760 35404 24800
rect 35444 24760 35453 24800
rect 35395 24759 35453 24760
rect 41635 24800 41693 24801
rect 41635 24760 41644 24800
rect 41684 24760 41693 24800
rect 41635 24759 41693 24760
rect 41923 24800 41981 24801
rect 41923 24760 41932 24800
rect 41972 24760 41981 24800
rect 41923 24759 41981 24760
rect 46243 24800 46301 24801
rect 46243 24760 46252 24800
rect 46292 24760 46301 24800
rect 46243 24759 46301 24760
rect 47011 24800 47069 24801
rect 47011 24760 47020 24800
rect 47060 24760 47069 24800
rect 47011 24759 47069 24760
rect 48643 24800 48701 24801
rect 48643 24760 48652 24800
rect 48692 24760 48701 24800
rect 48643 24759 48701 24760
rect 49035 24800 49077 24809
rect 49035 24760 49036 24800
rect 49076 24760 49077 24800
rect 49035 24751 49077 24760
rect 4395 24716 4437 24725
rect 4395 24676 4396 24716
rect 4436 24676 4437 24716
rect 4395 24667 4437 24676
rect 6123 24716 6165 24725
rect 6123 24676 6124 24716
rect 6164 24676 6165 24716
rect 6123 24667 6165 24676
rect 10347 24716 10389 24725
rect 10347 24676 10348 24716
rect 10388 24676 10389 24716
rect 10347 24667 10389 24676
rect 13227 24716 13269 24725
rect 13227 24676 13228 24716
rect 13268 24676 13269 24716
rect 13227 24667 13269 24676
rect 27435 24716 27477 24725
rect 27435 24676 27436 24716
rect 27476 24676 27477 24716
rect 27435 24667 27477 24676
rect 33003 24716 33045 24725
rect 33003 24676 33004 24716
rect 33044 24676 33045 24716
rect 33003 24667 33045 24676
rect 38859 24716 38901 24725
rect 38859 24676 38860 24716
rect 38900 24676 38901 24716
rect 38859 24667 38901 24676
rect 44331 24716 44373 24725
rect 44331 24676 44332 24716
rect 44372 24676 44373 24716
rect 44331 24667 44373 24676
rect 49323 24716 49365 24725
rect 49323 24676 49324 24716
rect 49364 24676 49365 24716
rect 49323 24667 49365 24676
rect 30123 24645 30165 24654
rect 931 24632 989 24633
rect 931 24592 940 24632
rect 980 24592 989 24632
rect 931 24591 989 24592
rect 1899 24632 1941 24641
rect 1899 24592 1900 24632
rect 1940 24592 1941 24632
rect 1899 24583 1941 24592
rect 2091 24632 2133 24641
rect 2091 24592 2092 24632
rect 2132 24592 2133 24632
rect 2091 24583 2133 24592
rect 2179 24632 2237 24633
rect 2179 24592 2188 24632
rect 2228 24592 2237 24632
rect 2179 24591 2237 24592
rect 2379 24632 2421 24641
rect 2379 24592 2380 24632
rect 2420 24592 2421 24632
rect 2379 24583 2421 24592
rect 2475 24632 2517 24641
rect 2475 24592 2476 24632
rect 2516 24592 2517 24632
rect 2475 24583 2517 24592
rect 2571 24632 2613 24641
rect 2571 24592 2572 24632
rect 2612 24592 2613 24632
rect 2571 24583 2613 24592
rect 2667 24632 2709 24641
rect 2667 24592 2668 24632
rect 2708 24592 2709 24632
rect 2667 24583 2709 24592
rect 3523 24632 3581 24633
rect 3523 24592 3532 24632
rect 3572 24592 3581 24632
rect 3523 24591 3581 24592
rect 3915 24632 3957 24641
rect 3915 24592 3916 24632
rect 3956 24592 3957 24632
rect 3915 24583 3957 24592
rect 4011 24632 4053 24641
rect 4011 24592 4012 24632
rect 4052 24592 4053 24632
rect 4011 24583 4053 24592
rect 4107 24632 4149 24641
rect 4107 24592 4108 24632
rect 4148 24592 4149 24632
rect 4107 24583 4149 24592
rect 5059 24632 5117 24633
rect 5059 24592 5068 24632
rect 5108 24592 5117 24632
rect 5059 24591 5117 24592
rect 5451 24632 5493 24641
rect 5451 24592 5452 24632
rect 5492 24592 5493 24632
rect 5451 24583 5493 24592
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5547 24583 5589 24592
rect 5643 24632 5685 24641
rect 5643 24592 5644 24632
rect 5684 24592 5685 24632
rect 5643 24583 5685 24592
rect 5739 24632 5781 24641
rect 5739 24592 5740 24632
rect 5780 24592 5781 24632
rect 5739 24583 5781 24592
rect 5923 24632 5981 24633
rect 5923 24592 5932 24632
rect 5972 24592 5981 24632
rect 5923 24591 5981 24592
rect 6027 24632 6069 24641
rect 6027 24592 6028 24632
rect 6068 24592 6069 24632
rect 6027 24583 6069 24592
rect 6219 24632 6261 24641
rect 6219 24592 6220 24632
rect 6260 24592 6261 24632
rect 6219 24583 6261 24592
rect 6411 24632 6453 24641
rect 6411 24592 6412 24632
rect 6452 24592 6453 24632
rect 6411 24583 6453 24592
rect 6507 24632 6549 24641
rect 6507 24592 6508 24632
rect 6548 24592 6549 24632
rect 6507 24583 6549 24592
rect 6603 24632 6645 24641
rect 6603 24592 6604 24632
rect 6644 24592 6645 24632
rect 6603 24583 6645 24592
rect 7555 24632 7613 24633
rect 7555 24592 7564 24632
rect 7604 24592 7613 24632
rect 7555 24591 7613 24592
rect 7755 24632 7797 24641
rect 7755 24592 7756 24632
rect 7796 24592 7797 24632
rect 7755 24583 7797 24592
rect 7947 24632 7989 24641
rect 7947 24592 7948 24632
rect 7988 24592 7989 24632
rect 7947 24583 7989 24592
rect 8619 24632 8661 24641
rect 8619 24592 8620 24632
rect 8660 24592 8661 24632
rect 8619 24583 8661 24592
rect 8803 24632 8861 24633
rect 8803 24592 8812 24632
rect 8852 24592 8861 24632
rect 8803 24591 8861 24592
rect 8995 24632 9053 24633
rect 8995 24592 9004 24632
rect 9044 24592 9053 24632
rect 8995 24591 9053 24592
rect 9955 24632 10013 24633
rect 9955 24592 9964 24632
rect 10004 24592 10013 24632
rect 9955 24591 10013 24592
rect 10251 24632 10293 24641
rect 10251 24592 10252 24632
rect 10292 24592 10293 24632
rect 10251 24583 10293 24592
rect 11971 24632 12029 24633
rect 11971 24592 11980 24632
rect 12020 24592 12029 24632
rect 11971 24591 12029 24592
rect 12835 24632 12893 24633
rect 12835 24592 12844 24632
rect 12884 24592 12893 24632
rect 12835 24591 12893 24592
rect 13507 24632 13565 24633
rect 13507 24592 13516 24632
rect 13556 24592 13565 24632
rect 13507 24591 13565 24592
rect 13803 24632 13845 24641
rect 13803 24592 13804 24632
rect 13844 24592 13845 24632
rect 13803 24583 13845 24592
rect 13899 24632 13941 24641
rect 13899 24592 13900 24632
rect 13940 24592 13941 24632
rect 13899 24583 13941 24592
rect 14467 24632 14525 24633
rect 14467 24592 14476 24632
rect 14516 24592 14525 24632
rect 14467 24591 14525 24592
rect 15427 24632 15485 24633
rect 15427 24592 15436 24632
rect 15476 24592 15485 24632
rect 15427 24591 15485 24592
rect 15531 24632 15573 24641
rect 15531 24592 15532 24632
rect 15572 24592 15573 24632
rect 15531 24583 15573 24592
rect 15723 24632 15765 24641
rect 15723 24592 15724 24632
rect 15764 24592 15765 24632
rect 15723 24583 15765 24592
rect 15915 24632 15957 24641
rect 15915 24592 15916 24632
rect 15956 24592 15957 24632
rect 15915 24583 15957 24592
rect 16011 24632 16053 24641
rect 16011 24592 16012 24632
rect 16052 24592 16053 24632
rect 16011 24583 16053 24592
rect 16107 24632 16149 24641
rect 16107 24592 16108 24632
rect 16148 24592 16149 24632
rect 16107 24583 16149 24592
rect 16203 24632 16245 24641
rect 16203 24592 16204 24632
rect 16244 24592 16245 24632
rect 16203 24583 16245 24592
rect 16963 24632 17021 24633
rect 16963 24592 16972 24632
rect 17012 24592 17021 24632
rect 16963 24591 17021 24592
rect 17259 24632 17301 24641
rect 17259 24592 17260 24632
rect 17300 24592 17301 24632
rect 17259 24583 17301 24592
rect 17923 24632 17981 24633
rect 17923 24592 17932 24632
rect 17972 24592 17981 24632
rect 17923 24591 17981 24592
rect 18123 24632 18165 24641
rect 18123 24592 18124 24632
rect 18164 24592 18165 24632
rect 18123 24583 18165 24592
rect 18219 24632 18261 24641
rect 18219 24592 18220 24632
rect 18260 24592 18261 24632
rect 18219 24583 18261 24592
rect 18315 24632 18357 24641
rect 18315 24592 18316 24632
rect 18356 24592 18357 24632
rect 18315 24583 18357 24592
rect 18411 24632 18453 24641
rect 18411 24592 18412 24632
rect 18452 24592 18453 24632
rect 18411 24583 18453 24592
rect 18691 24632 18749 24633
rect 18691 24592 18700 24632
rect 18740 24592 18749 24632
rect 18691 24591 18749 24592
rect 20907 24632 20949 24641
rect 20907 24592 20908 24632
rect 20948 24592 20949 24632
rect 20907 24583 20949 24592
rect 21003 24632 21045 24641
rect 21003 24592 21004 24632
rect 21044 24592 21045 24632
rect 21003 24583 21045 24592
rect 21099 24632 21141 24641
rect 21099 24592 21100 24632
rect 21140 24592 21141 24632
rect 21099 24583 21141 24592
rect 21195 24632 21237 24641
rect 21195 24592 21196 24632
rect 21236 24592 21237 24632
rect 21195 24583 21237 24592
rect 21763 24632 21821 24633
rect 21763 24592 21772 24632
rect 21812 24592 21821 24632
rect 21763 24591 21821 24592
rect 21867 24627 21909 24636
rect 21867 24587 21868 24627
rect 21908 24587 21909 24627
rect 21955 24632 22013 24633
rect 21955 24592 21964 24632
rect 22004 24592 22013 24632
rect 21955 24591 22013 24592
rect 22243 24632 22301 24633
rect 22243 24592 22252 24632
rect 22292 24592 22301 24632
rect 22243 24591 22301 24592
rect 24547 24632 24605 24633
rect 24547 24592 24556 24632
rect 24596 24592 24605 24632
rect 24547 24591 24605 24592
rect 25707 24632 25749 24641
rect 25707 24592 25708 24632
rect 25748 24592 25749 24632
rect 21867 24578 21909 24587
rect 25707 24583 25749 24592
rect 26083 24632 26141 24633
rect 26083 24592 26092 24632
rect 26132 24592 26141 24632
rect 26083 24591 26141 24592
rect 26187 24632 26229 24641
rect 26187 24592 26188 24632
rect 26228 24592 26229 24632
rect 26187 24583 26229 24592
rect 26467 24632 26525 24633
rect 26467 24592 26476 24632
rect 26516 24592 26525 24632
rect 26467 24591 26525 24592
rect 26955 24632 26997 24641
rect 26955 24592 26956 24632
rect 26996 24592 26997 24632
rect 26955 24583 26997 24592
rect 27147 24632 27189 24641
rect 27147 24592 27148 24632
rect 27188 24592 27189 24632
rect 27147 24583 27189 24592
rect 27235 24632 27293 24633
rect 27235 24592 27244 24632
rect 27284 24592 27293 24632
rect 27235 24591 27293 24592
rect 28099 24632 28157 24633
rect 28099 24592 28108 24632
rect 28148 24592 28157 24632
rect 28099 24591 28157 24592
rect 29251 24632 29309 24633
rect 29251 24592 29260 24632
rect 29300 24592 29309 24632
rect 29251 24591 29309 24592
rect 29635 24632 29693 24633
rect 29635 24592 29644 24632
rect 29684 24592 29693 24632
rect 29635 24591 29693 24592
rect 29835 24632 29877 24641
rect 29835 24592 29836 24632
rect 29876 24592 29877 24632
rect 29835 24583 29877 24592
rect 30019 24632 30077 24633
rect 30019 24592 30028 24632
rect 30068 24592 30077 24632
rect 30123 24605 30124 24645
rect 30164 24605 30165 24645
rect 30123 24596 30165 24605
rect 30315 24632 30357 24641
rect 30019 24591 30077 24592
rect 30315 24592 30316 24632
rect 30356 24592 30357 24632
rect 30315 24583 30357 24592
rect 30787 24632 30845 24633
rect 30787 24592 30796 24632
rect 30836 24592 30845 24632
rect 30787 24591 30845 24592
rect 31659 24632 31701 24641
rect 31659 24592 31660 24632
rect 31700 24592 31701 24632
rect 31659 24583 31701 24592
rect 32131 24632 32189 24633
rect 32131 24592 32140 24632
rect 32180 24592 32189 24632
rect 32131 24591 32189 24592
rect 32907 24632 32949 24641
rect 32907 24592 32908 24632
rect 32948 24592 32949 24632
rect 32907 24583 32949 24592
rect 33091 24632 33149 24633
rect 33091 24592 33100 24632
rect 33140 24592 33149 24632
rect 33091 24591 33149 24592
rect 33291 24632 33333 24641
rect 33291 24592 33292 24632
rect 33332 24592 33333 24632
rect 33291 24583 33333 24592
rect 33955 24632 34013 24633
rect 33955 24592 33964 24632
rect 34004 24592 34013 24632
rect 33955 24591 34013 24592
rect 34243 24632 34301 24633
rect 34243 24592 34252 24632
rect 34292 24592 34301 24632
rect 34243 24591 34301 24592
rect 35203 24632 35261 24633
rect 35203 24592 35212 24632
rect 35252 24592 35261 24632
rect 35203 24591 35261 24592
rect 36067 24632 36125 24633
rect 36067 24592 36076 24632
rect 36116 24592 36125 24632
rect 36067 24591 36125 24592
rect 37699 24632 37757 24633
rect 37699 24592 37708 24632
rect 37748 24592 37757 24632
rect 37699 24591 37757 24592
rect 38571 24632 38613 24641
rect 38571 24592 38572 24632
rect 38612 24592 38613 24632
rect 38571 24583 38613 24592
rect 39051 24627 39093 24636
rect 39051 24587 39052 24627
rect 39092 24587 39093 24627
rect 39523 24632 39581 24633
rect 39523 24592 39532 24632
rect 39572 24592 39581 24632
rect 39523 24591 39581 24592
rect 40107 24632 40149 24641
rect 40107 24592 40108 24632
rect 40148 24592 40149 24632
rect 39051 24578 39093 24587
rect 40107 24583 40149 24592
rect 40491 24632 40533 24641
rect 40491 24592 40492 24632
rect 40532 24592 40533 24632
rect 40491 24583 40533 24592
rect 40587 24632 40629 24641
rect 40587 24592 40588 24632
rect 40628 24592 40629 24632
rect 40587 24583 40629 24592
rect 40971 24632 41013 24641
rect 40971 24592 40972 24632
rect 41012 24592 41013 24632
rect 40971 24583 41013 24592
rect 41067 24632 41109 24641
rect 41067 24592 41068 24632
rect 41108 24592 41109 24632
rect 41067 24583 41109 24592
rect 41163 24632 41205 24641
rect 41163 24592 41164 24632
rect 41204 24592 41205 24632
rect 41163 24583 41205 24592
rect 41259 24632 41301 24641
rect 41259 24592 41260 24632
rect 41300 24592 41301 24632
rect 41259 24583 41301 24592
rect 41443 24632 41501 24633
rect 41443 24592 41452 24632
rect 41492 24592 41501 24632
rect 41443 24591 41501 24592
rect 41547 24632 41589 24641
rect 41547 24592 41548 24632
rect 41588 24592 41589 24632
rect 41547 24583 41589 24592
rect 41739 24632 41781 24641
rect 41739 24592 41740 24632
rect 41780 24592 41781 24632
rect 41739 24583 41781 24592
rect 43075 24632 43133 24633
rect 43075 24592 43084 24632
rect 43124 24592 43133 24632
rect 43075 24591 43133 24592
rect 43939 24632 43997 24633
rect 43939 24592 43948 24632
rect 43988 24592 43997 24632
rect 43939 24591 43997 24592
rect 44707 24632 44765 24633
rect 44707 24592 44716 24632
rect 44756 24592 44765 24632
rect 44707 24591 44765 24592
rect 45667 24632 45725 24633
rect 45667 24592 45676 24632
rect 45716 24592 45725 24632
rect 45667 24591 45725 24592
rect 46347 24632 46389 24641
rect 46347 24592 46348 24632
rect 46388 24592 46389 24632
rect 46347 24583 46389 24592
rect 46443 24632 46485 24641
rect 46443 24592 46444 24632
rect 46484 24592 46485 24632
rect 46443 24583 46485 24592
rect 46539 24632 46581 24641
rect 46539 24592 46540 24632
rect 46580 24592 46581 24632
rect 46539 24583 46581 24592
rect 46731 24632 46773 24641
rect 46731 24592 46732 24632
rect 46772 24592 46773 24632
rect 46731 24583 46773 24592
rect 46827 24632 46869 24641
rect 46827 24592 46828 24632
rect 46868 24592 46869 24632
rect 46827 24583 46869 24592
rect 46923 24632 46965 24641
rect 46923 24592 46924 24632
rect 46964 24592 46965 24632
rect 46923 24583 46965 24592
rect 47203 24632 47261 24633
rect 47203 24592 47212 24632
rect 47252 24592 47261 24632
rect 47203 24591 47261 24592
rect 47307 24632 47349 24641
rect 47307 24592 47308 24632
rect 47348 24592 47349 24632
rect 47307 24583 47349 24592
rect 47499 24632 47541 24641
rect 47499 24592 47500 24632
rect 47540 24592 47541 24632
rect 47499 24583 47541 24592
rect 47683 24632 47741 24633
rect 47683 24592 47692 24632
rect 47732 24592 47741 24632
rect 47683 24591 47741 24592
rect 48555 24632 48597 24641
rect 48555 24592 48556 24632
rect 48596 24592 48597 24632
rect 48555 24583 48597 24592
rect 48747 24632 48789 24641
rect 48747 24592 48748 24632
rect 48788 24592 48789 24632
rect 48747 24583 48789 24592
rect 48835 24632 48893 24633
rect 48835 24592 48844 24632
rect 48884 24592 48893 24632
rect 48835 24591 48893 24592
rect 49123 24632 49181 24633
rect 49123 24592 49132 24632
rect 49172 24592 49181 24632
rect 49123 24591 49181 24592
rect 49699 24632 49757 24633
rect 49699 24592 49708 24632
rect 49748 24592 49757 24632
rect 49699 24591 49757 24592
rect 50563 24632 50621 24633
rect 50563 24592 50572 24632
rect 50612 24592 50621 24632
rect 50563 24591 50621 24592
rect 7851 24548 7893 24557
rect 7851 24508 7852 24548
rect 7892 24508 7893 24548
rect 7851 24499 7893 24508
rect 23115 24548 23157 24557
rect 23115 24508 23116 24548
rect 23156 24508 23157 24548
rect 23115 24499 23157 24508
rect 40011 24548 40053 24557
rect 40011 24508 40012 24548
rect 40052 24508 40053 24548
rect 40011 24499 40053 24508
rect 1323 24464 1365 24473
rect 1323 24424 1324 24464
rect 1364 24424 1365 24464
rect 1323 24415 1365 24424
rect 1707 24464 1749 24473
rect 1707 24424 1708 24464
rect 1748 24424 1749 24464
rect 1707 24415 1749 24424
rect 8139 24464 8181 24473
rect 8139 24424 8140 24464
rect 8180 24424 8181 24464
rect 8139 24415 8181 24424
rect 8715 24464 8757 24473
rect 8715 24424 8716 24464
rect 8756 24424 8757 24464
rect 8715 24415 8757 24424
rect 10627 24464 10685 24465
rect 10627 24424 10636 24464
rect 10676 24424 10685 24464
rect 10627 24423 10685 24424
rect 14179 24464 14237 24465
rect 14179 24424 14188 24464
rect 14228 24424 14237 24464
rect 14179 24423 14237 24424
rect 14763 24464 14805 24473
rect 14763 24424 14764 24464
rect 14804 24424 14805 24464
rect 14763 24415 14805 24424
rect 15723 24464 15765 24473
rect 15723 24424 15724 24464
rect 15764 24424 15765 24464
rect 15723 24415 15765 24424
rect 18891 24464 18933 24473
rect 18891 24424 18892 24464
rect 18932 24424 18933 24464
rect 18891 24415 18933 24424
rect 19275 24464 19317 24473
rect 19275 24424 19276 24464
rect 19316 24424 19317 24464
rect 19275 24415 19317 24424
rect 30315 24464 30357 24473
rect 30315 24424 30316 24464
rect 30356 24424 30357 24464
rect 30315 24415 30357 24424
rect 32715 24464 32757 24473
rect 32715 24424 32716 24464
rect 32756 24424 32757 24464
rect 32715 24415 32757 24424
rect 47499 24464 47541 24473
rect 47499 24424 47500 24464
rect 47540 24424 47541 24464
rect 47499 24415 47541 24424
rect 2851 24380 2909 24381
rect 2851 24340 2860 24380
rect 2900 24340 2909 24380
rect 2851 24339 2909 24340
rect 6883 24380 6941 24381
rect 6883 24340 6892 24380
rect 6932 24340 6941 24380
rect 6883 24339 6941 24340
rect 14379 24380 14421 24389
rect 14379 24340 14380 24380
rect 14420 24340 14421 24380
rect 14379 24331 14421 24340
rect 18603 24380 18645 24389
rect 18603 24340 18604 24380
rect 18644 24340 18645 24380
rect 18603 24331 18645 24340
rect 21483 24380 21525 24389
rect 21483 24340 21484 24380
rect 21524 24340 21525 24380
rect 21483 24331 21525 24340
rect 28587 24380 28629 24389
rect 28587 24340 28588 24380
rect 28628 24340 28629 24380
rect 28587 24331 28629 24340
rect 29739 24380 29781 24389
rect 29739 24340 29740 24380
rect 29780 24340 29781 24380
rect 29739 24331 29781 24340
rect 32043 24380 32085 24389
rect 32043 24340 32044 24380
rect 32084 24340 32085 24380
rect 32043 24331 32085 24340
rect 35395 24380 35453 24381
rect 35395 24340 35404 24380
rect 35444 24340 35453 24380
rect 35395 24339 35453 24340
rect 48355 24380 48413 24381
rect 48355 24340 48364 24380
rect 48404 24340 48413 24380
rect 48355 24339 48413 24340
rect 51715 24380 51773 24381
rect 51715 24340 51724 24380
rect 51764 24340 51773 24380
rect 51715 24339 51773 24340
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 17739 24044 17781 24053
rect 17739 24004 17740 24044
rect 17780 24004 17781 24044
rect 17739 23995 17781 24004
rect 40011 24044 40053 24053
rect 40011 24004 40012 24044
rect 40052 24004 40053 24044
rect 40011 23995 40053 24004
rect 40779 24044 40821 24053
rect 40779 24004 40780 24044
rect 40820 24004 40821 24044
rect 40779 23995 40821 24004
rect 46251 24044 46293 24053
rect 46251 24004 46252 24044
rect 46292 24004 46293 24044
rect 46251 23995 46293 24004
rect 46731 24044 46773 24053
rect 46731 24004 46732 24044
rect 46772 24004 46773 24044
rect 46731 23995 46773 24004
rect 4011 23960 4053 23969
rect 4011 23920 4012 23960
rect 4052 23920 4053 23960
rect 4011 23911 4053 23920
rect 6123 23960 6165 23969
rect 6123 23920 6124 23960
rect 6164 23920 6165 23960
rect 6123 23911 6165 23920
rect 9283 23960 9341 23961
rect 9283 23920 9292 23960
rect 9332 23920 9341 23960
rect 9283 23919 9341 23920
rect 9675 23960 9717 23969
rect 9675 23920 9676 23960
rect 9716 23920 9717 23960
rect 9675 23911 9717 23920
rect 14091 23960 14133 23969
rect 14091 23920 14092 23960
rect 14132 23920 14133 23960
rect 14091 23911 14133 23920
rect 16675 23960 16733 23961
rect 16675 23920 16684 23960
rect 16724 23920 16733 23960
rect 16675 23919 16733 23920
rect 21387 23960 21429 23969
rect 21387 23920 21388 23960
rect 21428 23920 21429 23960
rect 21387 23911 21429 23920
rect 25131 23960 25173 23969
rect 25131 23920 25132 23960
rect 25172 23920 25173 23960
rect 25131 23911 25173 23920
rect 26763 23960 26805 23969
rect 26763 23920 26764 23960
rect 26804 23920 26805 23960
rect 26763 23911 26805 23920
rect 30795 23960 30837 23969
rect 30795 23920 30796 23960
rect 30836 23920 30837 23960
rect 30795 23911 30837 23920
rect 31275 23960 31317 23969
rect 31275 23920 31276 23960
rect 31316 23920 31317 23960
rect 31275 23911 31317 23920
rect 40491 23960 40533 23969
rect 40491 23920 40492 23960
rect 40532 23920 40533 23960
rect 40491 23911 40533 23920
rect 43659 23960 43701 23969
rect 43659 23920 43660 23960
rect 43700 23920 43701 23960
rect 43659 23911 43701 23920
rect 44907 23960 44949 23969
rect 44907 23920 44908 23960
rect 44948 23920 44949 23960
rect 44907 23911 44949 23920
rect 49611 23960 49653 23969
rect 49611 23920 49612 23960
rect 49652 23920 49653 23960
rect 49611 23911 49653 23920
rect 50859 23960 50901 23969
rect 50859 23920 50860 23960
rect 50900 23920 50901 23960
rect 50859 23911 50901 23920
rect 3531 23876 3573 23885
rect 3531 23836 3532 23876
rect 3572 23836 3573 23876
rect 3531 23827 3573 23836
rect 10443 23876 10485 23885
rect 10443 23836 10444 23876
rect 10484 23836 10485 23876
rect 10443 23827 10485 23836
rect 23787 23876 23829 23885
rect 23787 23836 23788 23876
rect 23828 23836 23829 23876
rect 23787 23827 23829 23836
rect 32995 23876 33053 23877
rect 32995 23836 33004 23876
rect 33044 23836 33053 23876
rect 37803 23876 37845 23885
rect 32995 23835 33053 23836
rect 36699 23834 36741 23843
rect 17739 23803 17781 23812
rect 1507 23792 1565 23793
rect 1507 23752 1516 23792
rect 1556 23752 1565 23792
rect 1507 23751 1565 23752
rect 2371 23792 2429 23793
rect 2371 23752 2380 23792
rect 2420 23752 2429 23792
rect 2371 23751 2429 23752
rect 3723 23792 3765 23801
rect 3723 23752 3724 23792
rect 3764 23752 3765 23792
rect 3723 23743 3765 23752
rect 3811 23792 3869 23793
rect 3811 23752 3820 23792
rect 3860 23752 3869 23792
rect 3811 23751 3869 23752
rect 4011 23792 4053 23801
rect 4011 23752 4012 23792
rect 4052 23752 4053 23792
rect 4011 23743 4053 23752
rect 4203 23792 4245 23801
rect 4203 23752 4204 23792
rect 4244 23752 4245 23792
rect 4203 23743 4245 23752
rect 4291 23792 4349 23793
rect 4291 23752 4300 23792
rect 4340 23752 4349 23792
rect 4291 23751 4349 23752
rect 4587 23792 4629 23801
rect 4587 23752 4588 23792
rect 4628 23752 4629 23792
rect 4587 23743 4629 23752
rect 4779 23792 4821 23801
rect 4779 23752 4780 23792
rect 4820 23752 4821 23792
rect 4779 23743 4821 23752
rect 4867 23792 4925 23793
rect 4867 23752 4876 23792
rect 4916 23752 4925 23792
rect 4867 23751 4925 23752
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 5259 23792 5301 23801
rect 5259 23752 5260 23792
rect 5300 23752 5301 23792
rect 5259 23743 5301 23752
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 5451 23792 5493 23801
rect 5451 23752 5452 23792
rect 5492 23752 5493 23792
rect 5451 23743 5493 23752
rect 6595 23792 6653 23793
rect 6595 23752 6604 23792
rect 6644 23752 6653 23792
rect 6595 23751 6653 23752
rect 6891 23792 6933 23801
rect 6891 23752 6892 23792
rect 6932 23752 6933 23792
rect 6891 23743 6933 23752
rect 7267 23792 7325 23793
rect 7267 23752 7276 23792
rect 7316 23752 7325 23792
rect 7267 23751 7325 23752
rect 8131 23792 8189 23793
rect 8131 23752 8140 23792
rect 8180 23752 8189 23792
rect 8131 23751 8189 23752
rect 9963 23792 10005 23801
rect 9963 23752 9964 23792
rect 10004 23752 10005 23792
rect 9963 23743 10005 23752
rect 10059 23792 10101 23801
rect 10059 23752 10060 23792
rect 10100 23752 10101 23792
rect 10059 23743 10101 23752
rect 10155 23792 10197 23801
rect 10155 23752 10156 23792
rect 10196 23752 10197 23792
rect 10155 23743 10197 23752
rect 11211 23792 11253 23801
rect 11211 23752 11212 23792
rect 11252 23752 11253 23792
rect 11211 23743 11253 23752
rect 12747 23792 12789 23801
rect 12747 23752 12748 23792
rect 12788 23752 12789 23792
rect 12747 23743 12789 23752
rect 13795 23792 13853 23793
rect 13795 23752 13804 23792
rect 13844 23752 13853 23792
rect 13795 23751 13853 23752
rect 13899 23792 13941 23801
rect 13899 23752 13900 23792
rect 13940 23752 13941 23792
rect 13899 23743 13941 23752
rect 14091 23792 14133 23801
rect 14091 23752 14092 23792
rect 14132 23752 14133 23792
rect 14091 23743 14133 23752
rect 14283 23792 14325 23801
rect 14283 23752 14284 23792
rect 14324 23752 14325 23792
rect 14283 23743 14325 23752
rect 14659 23792 14717 23793
rect 14659 23752 14668 23792
rect 14708 23752 14717 23792
rect 14659 23751 14717 23752
rect 15523 23792 15581 23793
rect 15523 23752 15532 23792
rect 15572 23752 15581 23792
rect 15523 23751 15581 23752
rect 16971 23792 17013 23801
rect 16971 23752 16972 23792
rect 17012 23752 17013 23792
rect 16971 23743 17013 23752
rect 17067 23792 17109 23801
rect 17067 23752 17068 23792
rect 17108 23752 17109 23792
rect 17067 23743 17109 23752
rect 17443 23792 17501 23793
rect 17443 23752 17452 23792
rect 17492 23752 17501 23792
rect 17443 23751 17501 23752
rect 17547 23792 17589 23801
rect 17547 23752 17548 23792
rect 17588 23752 17589 23792
rect 17739 23763 17740 23803
rect 17780 23763 17781 23803
rect 17739 23754 17781 23763
rect 17923 23792 17981 23793
rect 17547 23743 17589 23752
rect 17923 23752 17932 23792
rect 17972 23752 17981 23792
rect 17923 23751 17981 23752
rect 19459 23792 19517 23793
rect 19459 23752 19468 23792
rect 19508 23752 19517 23792
rect 19459 23751 19517 23752
rect 20707 23792 20765 23793
rect 20707 23752 20716 23792
rect 20756 23752 20765 23792
rect 20707 23751 20765 23752
rect 21579 23792 21621 23801
rect 21579 23752 21580 23792
rect 21620 23752 21621 23792
rect 21579 23743 21621 23752
rect 23019 23792 23061 23801
rect 23019 23752 23020 23792
rect 23060 23752 23061 23792
rect 23019 23743 23061 23752
rect 24363 23792 24405 23801
rect 24363 23752 24364 23792
rect 24404 23752 24405 23792
rect 24363 23743 24405 23752
rect 24459 23792 24501 23801
rect 24459 23752 24460 23792
rect 24500 23752 24501 23792
rect 24459 23743 24501 23752
rect 24643 23792 24701 23793
rect 24643 23752 24652 23792
rect 24692 23752 24701 23792
rect 24643 23751 24701 23752
rect 25603 23792 25661 23793
rect 25603 23752 25612 23792
rect 25652 23752 25661 23792
rect 25603 23751 25661 23752
rect 25899 23792 25941 23801
rect 25899 23752 25900 23792
rect 25940 23752 25941 23792
rect 25899 23743 25941 23752
rect 26563 23792 26621 23793
rect 26563 23752 26572 23792
rect 26612 23752 26621 23792
rect 26563 23751 26621 23752
rect 28195 23792 28253 23793
rect 28195 23752 28204 23792
rect 28244 23752 28253 23792
rect 28195 23751 28253 23752
rect 29443 23792 29501 23793
rect 29443 23752 29452 23792
rect 29492 23752 29501 23792
rect 29443 23751 29501 23752
rect 29739 23792 29781 23801
rect 29739 23752 29740 23792
rect 29780 23752 29781 23792
rect 29739 23743 29781 23752
rect 30403 23792 30461 23793
rect 30403 23752 30412 23792
rect 30452 23752 30461 23792
rect 30403 23751 30461 23752
rect 30979 23792 31037 23793
rect 30979 23752 30988 23792
rect 31028 23752 31037 23792
rect 30979 23751 31037 23752
rect 31083 23792 31125 23801
rect 31083 23752 31084 23792
rect 31124 23752 31125 23792
rect 31083 23743 31125 23752
rect 31275 23792 31317 23801
rect 31275 23752 31276 23792
rect 31316 23752 31317 23792
rect 31275 23743 31317 23752
rect 32131 23792 32189 23793
rect 32131 23752 32140 23792
rect 32180 23752 32189 23792
rect 32131 23751 32189 23752
rect 32331 23792 32373 23801
rect 32331 23752 32332 23792
rect 32372 23752 32373 23792
rect 32331 23743 32373 23752
rect 32427 23792 32469 23801
rect 32427 23752 32428 23792
rect 32468 23752 32469 23792
rect 32427 23743 32469 23752
rect 32523 23792 32565 23801
rect 32523 23752 32524 23792
rect 32564 23752 32565 23792
rect 32523 23743 32565 23752
rect 32619 23792 32661 23801
rect 32619 23752 32620 23792
rect 32660 23752 32661 23792
rect 32619 23743 32661 23752
rect 33387 23792 33429 23801
rect 33387 23752 33388 23792
rect 33428 23752 33429 23792
rect 33387 23743 33429 23752
rect 33483 23792 33525 23801
rect 33483 23752 33484 23792
rect 33524 23752 33525 23792
rect 33483 23743 33525 23752
rect 33579 23792 33621 23801
rect 33579 23752 33580 23792
rect 33620 23752 33621 23792
rect 33579 23743 33621 23752
rect 33675 23792 33717 23801
rect 33675 23752 33676 23792
rect 33716 23752 33717 23792
rect 33675 23743 33717 23752
rect 33867 23792 33909 23801
rect 33867 23752 33868 23792
rect 33908 23752 33909 23792
rect 33867 23743 33909 23752
rect 33963 23792 34005 23801
rect 33963 23752 33964 23792
rect 34004 23752 34005 23792
rect 33963 23743 34005 23752
rect 34059 23792 34101 23801
rect 34059 23752 34060 23792
rect 34100 23752 34101 23792
rect 34059 23743 34101 23752
rect 34155 23792 34197 23801
rect 34155 23752 34156 23792
rect 34196 23752 34197 23792
rect 34155 23743 34197 23752
rect 34339 23792 34397 23793
rect 34339 23752 34348 23792
rect 34388 23752 34397 23792
rect 34339 23751 34397 23752
rect 34443 23792 34485 23801
rect 34443 23752 34444 23792
rect 34484 23752 34485 23792
rect 34443 23743 34485 23752
rect 34635 23792 34677 23801
rect 36699 23794 36700 23834
rect 36740 23794 36741 23834
rect 37803 23836 37804 23876
rect 37844 23836 37845 23876
rect 37803 23827 37845 23836
rect 46531 23876 46589 23877
rect 46531 23836 46540 23876
rect 46580 23836 46589 23876
rect 46531 23835 46589 23836
rect 47883 23876 47925 23885
rect 47883 23836 47884 23876
rect 47924 23836 47925 23876
rect 47883 23827 47925 23836
rect 34635 23752 34636 23792
rect 34676 23752 34677 23792
rect 34635 23743 34677 23752
rect 35491 23792 35549 23793
rect 35491 23752 35500 23792
rect 35540 23752 35549 23792
rect 35491 23751 35549 23752
rect 36355 23792 36413 23793
rect 36355 23752 36364 23792
rect 36404 23752 36413 23792
rect 36699 23785 36741 23794
rect 37219 23792 37277 23793
rect 36355 23751 36413 23752
rect 37219 23752 37228 23792
rect 37268 23752 37277 23792
rect 37219 23751 37277 23752
rect 37707 23792 37749 23801
rect 37707 23752 37708 23792
rect 37748 23752 37749 23792
rect 37707 23743 37749 23752
rect 38187 23792 38229 23801
rect 38187 23752 38188 23792
rect 38228 23752 38229 23792
rect 38187 23743 38229 23752
rect 38283 23792 38325 23801
rect 38283 23752 38284 23792
rect 38324 23752 38325 23792
rect 38283 23743 38325 23752
rect 39235 23792 39293 23793
rect 39235 23752 39244 23792
rect 39284 23752 39293 23792
rect 39235 23751 39293 23752
rect 40099 23792 40157 23793
rect 40099 23752 40108 23792
rect 40148 23752 40157 23792
rect 40099 23751 40157 23752
rect 40867 23792 40925 23793
rect 40867 23752 40876 23792
rect 40916 23752 40925 23792
rect 40867 23751 40925 23752
rect 41731 23792 41789 23793
rect 41731 23752 41740 23792
rect 41780 23752 41789 23792
rect 41731 23751 41789 23752
rect 41931 23792 41973 23801
rect 41931 23752 41932 23792
rect 41972 23752 41973 23792
rect 41931 23743 41973 23752
rect 42027 23792 42069 23801
rect 42027 23752 42028 23792
rect 42068 23752 42069 23792
rect 42027 23743 42069 23752
rect 42123 23792 42165 23801
rect 42123 23752 42124 23792
rect 42164 23752 42165 23792
rect 42123 23743 42165 23752
rect 43267 23792 43325 23793
rect 43267 23752 43276 23792
rect 43316 23752 43325 23792
rect 43267 23751 43325 23752
rect 45771 23792 45813 23801
rect 45771 23752 45772 23792
rect 45812 23752 45813 23792
rect 45771 23743 45813 23752
rect 45867 23792 45909 23801
rect 45867 23752 45868 23792
rect 45908 23752 45909 23792
rect 45867 23743 45909 23752
rect 45963 23792 46005 23801
rect 45963 23752 45964 23792
rect 46004 23752 46005 23792
rect 45963 23743 46005 23752
rect 46155 23792 46197 23801
rect 46155 23752 46156 23792
rect 46196 23752 46197 23792
rect 46155 23743 46197 23752
rect 46339 23792 46397 23793
rect 46339 23752 46348 23792
rect 46388 23752 46397 23792
rect 46339 23751 46397 23752
rect 47587 23792 47645 23793
rect 47587 23752 47596 23792
rect 47636 23752 47645 23792
rect 47587 23751 47645 23752
rect 48739 23792 48797 23793
rect 48739 23752 48748 23792
rect 48788 23752 48797 23792
rect 48739 23751 48797 23752
rect 49123 23792 49181 23793
rect 49123 23752 49132 23792
rect 49172 23752 49181 23792
rect 49123 23751 49181 23752
rect 49803 23792 49845 23801
rect 49803 23752 49804 23792
rect 49844 23752 49845 23792
rect 49803 23743 49845 23752
rect 50467 23792 50525 23793
rect 50467 23752 50476 23792
rect 50516 23752 50525 23792
rect 50467 23751 50525 23752
rect 1131 23708 1173 23717
rect 1131 23668 1132 23708
rect 1172 23668 1173 23708
rect 1131 23659 1173 23668
rect 4683 23708 4725 23717
rect 4683 23668 4684 23708
rect 4724 23668 4725 23708
rect 4683 23659 4725 23668
rect 11971 23708 12029 23709
rect 11971 23668 11980 23708
rect 12020 23668 12029 23708
rect 11971 23667 12029 23668
rect 27331 23708 27389 23709
rect 27331 23668 27340 23708
rect 27380 23668 27389 23708
rect 27331 23667 27389 23668
rect 34539 23708 34581 23717
rect 34539 23668 34540 23708
rect 34580 23668 34581 23708
rect 34539 23659 34581 23668
rect 36555 23708 36597 23717
rect 36555 23668 36556 23708
rect 36596 23668 36597 23708
rect 36555 23659 36597 23668
rect 42603 23708 42645 23717
rect 42603 23668 42604 23708
rect 42644 23668 42645 23708
rect 42603 23659 42645 23668
rect 9859 23624 9917 23625
rect 9859 23584 9868 23624
rect 9908 23584 9917 23624
rect 9859 23583 9917 23584
rect 17251 23624 17309 23625
rect 17251 23584 17260 23624
rect 17300 23584 17309 23624
rect 17251 23583 17309 23584
rect 18595 23624 18653 23625
rect 18595 23584 18604 23624
rect 18644 23584 18653 23624
rect 18595 23583 18653 23584
rect 18787 23624 18845 23625
rect 18787 23584 18796 23624
rect 18836 23584 18845 23624
rect 18787 23583 18845 23584
rect 23403 23624 23445 23633
rect 23403 23584 23404 23624
rect 23444 23584 23445 23624
rect 23403 23575 23445 23584
rect 24163 23624 24221 23625
rect 24163 23584 24172 23624
rect 24212 23584 24221 23624
rect 24163 23583 24221 23584
rect 28971 23624 29013 23633
rect 28971 23584 28972 23624
rect 29012 23584 29013 23624
rect 28971 23575 29013 23584
rect 31459 23624 31517 23625
rect 31459 23584 31468 23624
rect 31508 23584 31517 23624
rect 31459 23583 31517 23584
rect 33195 23624 33237 23633
rect 33195 23584 33196 23624
rect 33236 23584 33237 23624
rect 33195 23575 33237 23584
rect 34819 23624 34877 23625
rect 34819 23584 34828 23624
rect 34868 23584 34877 23624
rect 34819 23583 34877 23584
rect 35683 23624 35741 23625
rect 35683 23584 35692 23624
rect 35732 23584 35741 23624
rect 35683 23583 35741 23584
rect 38563 23624 38621 23625
rect 38563 23584 38572 23624
rect 38612 23584 38621 23624
rect 38563 23583 38621 23584
rect 41059 23624 41117 23625
rect 41059 23584 41068 23624
rect 41108 23584 41117 23624
rect 41059 23583 41117 23584
rect 42211 23624 42269 23625
rect 42211 23584 42220 23624
rect 42260 23584 42269 23624
rect 42211 23583 42269 23584
rect 45667 23624 45725 23625
rect 45667 23584 45676 23624
rect 45716 23584 45725 23624
rect 45667 23583 45725 23584
rect 46915 23624 46973 23625
rect 46915 23584 46924 23624
rect 46964 23584 46973 23624
rect 46915 23583 46973 23584
rect 49035 23624 49077 23633
rect 49035 23584 49036 23624
rect 49076 23584 49077 23624
rect 49035 23575 49077 23584
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 3811 23288 3869 23289
rect 3811 23248 3820 23288
rect 3860 23248 3869 23288
rect 3811 23247 3869 23248
rect 5635 23288 5693 23289
rect 5635 23248 5644 23288
rect 5684 23248 5693 23288
rect 5635 23247 5693 23248
rect 5931 23288 5973 23297
rect 5931 23248 5932 23288
rect 5972 23248 5973 23288
rect 5931 23239 5973 23248
rect 18019 23288 18077 23289
rect 18019 23248 18028 23288
rect 18068 23248 18077 23288
rect 18019 23247 18077 23248
rect 20803 23288 20861 23289
rect 20803 23248 20812 23288
rect 20852 23248 20861 23288
rect 20803 23247 20861 23248
rect 22155 23288 22197 23297
rect 22155 23248 22156 23288
rect 22196 23248 22197 23288
rect 22155 23239 22197 23248
rect 33475 23288 33533 23289
rect 33475 23248 33484 23288
rect 33524 23248 33533 23288
rect 33475 23247 33533 23248
rect 33667 23288 33725 23289
rect 33667 23248 33676 23288
rect 33716 23248 33725 23288
rect 33667 23247 33725 23248
rect 37315 23288 37373 23289
rect 37315 23248 37324 23288
rect 37364 23248 37373 23288
rect 37315 23247 37373 23248
rect 38667 23288 38709 23297
rect 38667 23248 38668 23288
rect 38708 23248 38709 23288
rect 38667 23239 38709 23248
rect 39531 23288 39573 23297
rect 39531 23248 39532 23288
rect 39572 23248 39573 23288
rect 39531 23239 39573 23248
rect 43363 23288 43421 23289
rect 43363 23248 43372 23288
rect 43412 23248 43421 23288
rect 43363 23247 43421 23248
rect 46819 23288 46877 23289
rect 46819 23248 46828 23288
rect 46868 23248 46877 23288
rect 46819 23247 46877 23248
rect 50179 23288 50237 23289
rect 50179 23248 50188 23288
rect 50228 23248 50237 23288
rect 50179 23247 50237 23248
rect 1419 23204 1461 23213
rect 1419 23164 1420 23204
rect 1460 23164 1461 23204
rect 1419 23155 1461 23164
rect 12835 23204 12893 23205
rect 12835 23164 12844 23204
rect 12884 23164 12893 23204
rect 12835 23163 12893 23164
rect 16491 23204 16533 23213
rect 16491 23164 16492 23204
rect 16532 23164 16533 23204
rect 16491 23155 16533 23164
rect 18411 23204 18453 23213
rect 18411 23164 18412 23204
rect 18452 23164 18453 23204
rect 18411 23155 18453 23164
rect 28867 23204 28925 23205
rect 28867 23164 28876 23204
rect 28916 23164 28925 23204
rect 28867 23163 28925 23164
rect 31083 23204 31125 23213
rect 31083 23164 31084 23204
rect 31124 23164 31125 23204
rect 31083 23155 31125 23164
rect 34923 23204 34965 23213
rect 34923 23164 34924 23204
rect 34964 23164 34965 23204
rect 34923 23155 34965 23164
rect 40683 23204 40725 23213
rect 40683 23164 40684 23204
rect 40724 23164 40725 23204
rect 40683 23155 40725 23164
rect 47787 23204 47829 23213
rect 47787 23164 47788 23204
rect 47828 23164 47829 23204
rect 47787 23155 47829 23164
rect 17547 23141 17589 23150
rect 1795 23120 1853 23121
rect 1795 23080 1804 23120
rect 1844 23080 1853 23120
rect 1795 23079 1853 23080
rect 2659 23120 2717 23121
rect 2659 23080 2668 23120
rect 2708 23080 2717 23120
rect 2659 23079 2717 23080
rect 4099 23120 4157 23121
rect 4099 23080 4108 23120
rect 4148 23080 4157 23120
rect 4099 23079 4157 23080
rect 4963 23120 5021 23121
rect 4963 23080 4972 23120
rect 5012 23080 5021 23120
rect 4963 23079 5021 23080
rect 5835 23120 5877 23129
rect 5835 23080 5836 23120
rect 5876 23080 5877 23120
rect 5835 23071 5877 23080
rect 6123 23120 6165 23129
rect 6123 23080 6124 23120
rect 6164 23080 6165 23120
rect 6123 23071 6165 23080
rect 7171 23120 7229 23121
rect 7171 23080 7180 23120
rect 7220 23080 7229 23120
rect 7171 23079 7229 23080
rect 8035 23120 8093 23121
rect 8035 23080 8044 23120
rect 8084 23080 8093 23120
rect 8035 23079 8093 23080
rect 8707 23120 8765 23121
rect 8707 23080 8716 23120
rect 8756 23080 8765 23120
rect 8707 23079 8765 23080
rect 8811 23120 8853 23129
rect 8811 23080 8812 23120
rect 8852 23080 8853 23120
rect 8811 23071 8853 23080
rect 9003 23120 9045 23129
rect 9003 23080 9004 23120
rect 9044 23080 9045 23120
rect 9003 23071 9045 23080
rect 9859 23120 9917 23121
rect 9859 23080 9868 23120
rect 9908 23080 9917 23120
rect 9859 23079 9917 23080
rect 10723 23120 10781 23121
rect 10723 23080 10732 23120
rect 10772 23080 10781 23120
rect 10723 23079 10781 23080
rect 11587 23120 11645 23121
rect 11587 23080 11596 23120
rect 11636 23080 11645 23120
rect 11587 23079 11645 23080
rect 11875 23120 11933 23121
rect 11875 23080 11884 23120
rect 11924 23080 11933 23120
rect 11875 23079 11933 23080
rect 13699 23120 13757 23121
rect 13699 23080 13708 23120
rect 13748 23080 13757 23120
rect 13699 23079 13757 23080
rect 14475 23120 14517 23129
rect 14475 23080 14476 23120
rect 14516 23080 14517 23120
rect 14475 23071 14517 23080
rect 15139 23120 15197 23121
rect 15139 23080 15148 23120
rect 15188 23080 15197 23120
rect 15139 23079 15197 23080
rect 15435 23120 15477 23129
rect 15435 23080 15436 23120
rect 15476 23080 15477 23120
rect 15435 23071 15477 23080
rect 15531 23120 15573 23129
rect 15531 23080 15532 23120
rect 15572 23080 15573 23120
rect 15531 23071 15573 23080
rect 15627 23120 15669 23129
rect 15627 23080 15628 23120
rect 15668 23080 15669 23120
rect 15627 23071 15669 23080
rect 15723 23120 15765 23129
rect 15723 23080 15724 23120
rect 15764 23080 15765 23120
rect 15723 23071 15765 23080
rect 16395 23120 16437 23129
rect 16395 23080 16396 23120
rect 16436 23080 16437 23120
rect 16395 23071 16437 23080
rect 16579 23120 16637 23121
rect 16579 23080 16588 23120
rect 16628 23080 16637 23120
rect 16579 23079 16637 23080
rect 16771 23120 16829 23121
rect 16771 23080 16780 23120
rect 16820 23080 16829 23120
rect 16771 23079 16829 23080
rect 16875 23120 16917 23129
rect 16875 23080 16876 23120
rect 16916 23080 16917 23120
rect 16875 23071 16917 23080
rect 17067 23120 17109 23129
rect 17067 23080 17068 23120
rect 17108 23080 17109 23120
rect 17067 23071 17109 23080
rect 17451 23120 17493 23129
rect 17451 23080 17452 23120
rect 17492 23080 17493 23120
rect 17547 23101 17548 23141
rect 17588 23101 17589 23141
rect 17547 23092 17589 23101
rect 17643 23120 17685 23129
rect 17451 23071 17493 23080
rect 17643 23080 17644 23120
rect 17684 23080 17685 23120
rect 17643 23071 17685 23080
rect 17739 23120 17781 23129
rect 17739 23080 17740 23120
rect 17780 23080 17781 23120
rect 17739 23071 17781 23080
rect 17931 23120 17973 23129
rect 17931 23080 17932 23120
rect 17972 23080 17973 23120
rect 17931 23071 17973 23080
rect 18123 23120 18165 23129
rect 18123 23080 18124 23120
rect 18164 23080 18165 23120
rect 18123 23071 18165 23080
rect 18211 23120 18269 23121
rect 18211 23080 18220 23120
rect 18260 23080 18269 23120
rect 18211 23079 18269 23080
rect 18787 23120 18845 23121
rect 18787 23080 18796 23120
rect 18836 23080 18845 23120
rect 18787 23079 18845 23080
rect 19651 23120 19709 23121
rect 19651 23080 19660 23120
rect 19700 23080 19709 23120
rect 19651 23079 19709 23080
rect 22539 23120 22581 23129
rect 22539 23080 22540 23120
rect 22580 23080 22581 23120
rect 22539 23071 22581 23080
rect 22923 23120 22965 23129
rect 22923 23080 22924 23120
rect 22964 23080 22965 23120
rect 22923 23071 22965 23080
rect 23299 23120 23357 23121
rect 23299 23080 23308 23120
rect 23348 23080 23357 23120
rect 23299 23079 23357 23080
rect 24163 23120 24221 23121
rect 24163 23080 24172 23120
rect 24212 23080 24221 23120
rect 24163 23079 24221 23080
rect 25411 23120 25469 23121
rect 25411 23080 25420 23120
rect 25460 23080 25469 23120
rect 25411 23079 25469 23080
rect 25803 23120 25845 23129
rect 25803 23080 25804 23120
rect 25844 23080 25845 23120
rect 25803 23071 25845 23080
rect 26179 23120 26237 23121
rect 26179 23080 26188 23120
rect 26228 23080 26237 23120
rect 26179 23079 26237 23080
rect 27043 23120 27101 23121
rect 27043 23080 27052 23120
rect 27092 23080 27101 23120
rect 27043 23079 27101 23080
rect 28203 23120 28245 23129
rect 28203 23080 28204 23120
rect 28244 23080 28245 23120
rect 28203 23071 28245 23080
rect 29643 23120 29685 23129
rect 29643 23080 29644 23120
rect 29684 23080 29685 23120
rect 29643 23071 29685 23080
rect 30315 23120 30357 23129
rect 30315 23080 30316 23120
rect 30356 23080 30357 23120
rect 30315 23071 30357 23080
rect 30411 23120 30453 23129
rect 30411 23080 30412 23120
rect 30452 23080 30453 23120
rect 30411 23071 30453 23080
rect 30691 23120 30749 23121
rect 30691 23080 30700 23120
rect 30740 23080 30749 23120
rect 30691 23079 30749 23080
rect 31459 23120 31517 23121
rect 31459 23080 31468 23120
rect 31508 23080 31517 23120
rect 31459 23079 31517 23080
rect 32323 23120 32381 23121
rect 32323 23080 32332 23120
rect 32372 23080 32381 23120
rect 32323 23079 32381 23080
rect 34339 23120 34397 23121
rect 34339 23080 34348 23120
rect 34388 23080 34397 23120
rect 34339 23079 34397 23080
rect 35299 23120 35357 23121
rect 35299 23080 35308 23120
rect 35348 23080 35357 23120
rect 35299 23079 35357 23080
rect 36163 23120 36221 23121
rect 36163 23080 36172 23120
rect 36212 23080 36221 23120
rect 36163 23079 36221 23080
rect 38563 23120 38621 23121
rect 38563 23080 38572 23120
rect 38612 23080 38621 23120
rect 38563 23079 38621 23080
rect 38955 23120 38997 23129
rect 38955 23080 38956 23120
rect 38996 23080 38997 23120
rect 38955 23071 38997 23080
rect 39051 23120 39093 23129
rect 39051 23080 39052 23120
rect 39092 23080 39093 23120
rect 39051 23071 39093 23080
rect 39147 23120 39189 23129
rect 39147 23080 39148 23120
rect 39188 23080 39189 23120
rect 39147 23071 39189 23080
rect 39243 23120 39285 23129
rect 39243 23080 39244 23120
rect 39284 23080 39285 23120
rect 39243 23071 39285 23080
rect 39427 23120 39485 23121
rect 39427 23080 39436 23120
rect 39476 23080 39485 23120
rect 39427 23079 39485 23080
rect 39723 23120 39765 23129
rect 39723 23080 39724 23120
rect 39764 23080 39765 23120
rect 39723 23071 39765 23080
rect 40387 23120 40445 23121
rect 40387 23080 40396 23120
rect 40436 23080 40445 23120
rect 40387 23079 40445 23080
rect 41059 23120 41117 23121
rect 41059 23080 41068 23120
rect 41108 23080 41117 23120
rect 41059 23079 41117 23080
rect 41923 23120 41981 23121
rect 41923 23080 41932 23120
rect 41972 23080 41981 23120
rect 41923 23079 41981 23080
rect 43467 23120 43509 23129
rect 43467 23080 43468 23120
rect 43508 23080 43509 23120
rect 43467 23071 43509 23080
rect 43563 23120 43605 23129
rect 43563 23080 43564 23120
rect 43604 23080 43605 23120
rect 43563 23071 43605 23080
rect 43659 23120 43701 23129
rect 43659 23080 43660 23120
rect 43700 23080 43701 23120
rect 43659 23071 43701 23080
rect 43939 23120 43997 23121
rect 43939 23080 43948 23120
rect 43988 23080 43997 23120
rect 43939 23079 43997 23080
rect 44227 23120 44285 23121
rect 44227 23080 44236 23120
rect 44276 23080 44285 23120
rect 44227 23079 44285 23080
rect 44427 23120 44469 23129
rect 44427 23080 44428 23120
rect 44468 23080 44469 23120
rect 44427 23071 44469 23080
rect 44803 23120 44861 23121
rect 44803 23080 44812 23120
rect 44852 23080 44861 23120
rect 44803 23079 44861 23080
rect 45667 23120 45725 23121
rect 45667 23080 45676 23120
rect 45716 23080 45725 23120
rect 45667 23079 45725 23080
rect 47211 23120 47253 23129
rect 47211 23080 47212 23120
rect 47252 23080 47253 23120
rect 47211 23071 47253 23080
rect 47307 23120 47349 23129
rect 47307 23080 47308 23120
rect 47348 23080 47349 23120
rect 47307 23071 47349 23080
rect 47403 23120 47445 23129
rect 47403 23080 47404 23120
rect 47444 23080 47445 23120
rect 47403 23071 47445 23080
rect 47499 23120 47541 23129
rect 47499 23080 47500 23120
rect 47540 23080 47541 23120
rect 47499 23071 47541 23080
rect 48163 23120 48221 23121
rect 48163 23080 48172 23120
rect 48212 23080 48221 23120
rect 48163 23079 48221 23080
rect 49027 23120 49085 23121
rect 49027 23080 49036 23120
rect 49076 23080 49085 23120
rect 49027 23079 49085 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 16099 23036 16157 23037
rect 16099 22996 16108 23036
rect 16148 22996 16157 23036
rect 16099 22995 16157 22996
rect 9003 22952 9045 22961
rect 9003 22912 9004 22952
rect 9044 22912 9045 22952
rect 9003 22903 9045 22912
rect 14283 22952 14325 22961
rect 14283 22912 14284 22952
rect 14324 22912 14325 22952
rect 14283 22903 14325 22912
rect 15915 22952 15957 22961
rect 15915 22912 15916 22952
rect 15956 22912 15957 22952
rect 15915 22903 15957 22912
rect 30019 22952 30077 22953
rect 30019 22912 30028 22952
rect 30068 22912 30077 22952
rect 30019 22911 30077 22912
rect 34731 22952 34773 22961
rect 34731 22912 34732 22952
rect 34772 22912 34773 22952
rect 34731 22903 34773 22912
rect 37803 22952 37845 22961
rect 37803 22912 37804 22952
rect 37844 22912 37845 22952
rect 37803 22903 37845 22912
rect 43075 22952 43133 22953
rect 43075 22912 43084 22952
rect 43124 22912 43133 22952
rect 43075 22911 43133 22912
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 4771 22868 4829 22869
rect 4771 22828 4780 22868
rect 4820 22828 4829 22868
rect 4771 22827 4829 22828
rect 5635 22868 5693 22869
rect 5635 22828 5644 22868
rect 5684 22828 5693 22868
rect 5635 22827 5693 22828
rect 6499 22868 6557 22869
rect 6499 22828 6508 22868
rect 6548 22828 6557 22868
rect 6499 22827 6557 22828
rect 7363 22868 7421 22869
rect 7363 22828 7372 22868
rect 7412 22828 7421 22868
rect 7363 22827 7421 22828
rect 9187 22868 9245 22869
rect 9187 22828 9196 22868
rect 9236 22828 9245 22868
rect 9187 22827 9245 22828
rect 10051 22868 10109 22869
rect 10051 22828 10060 22868
rect 10100 22828 10109 22868
rect 10051 22827 10109 22828
rect 10915 22868 10973 22869
rect 10915 22828 10924 22868
rect 10964 22828 10973 22868
rect 10915 22827 10973 22828
rect 12547 22868 12605 22869
rect 12547 22828 12556 22868
rect 12596 22828 12605 22868
rect 12547 22827 12605 22828
rect 17067 22868 17109 22877
rect 17067 22828 17068 22868
rect 17108 22828 17109 22868
rect 17067 22819 17109 22828
rect 43851 22868 43893 22877
rect 43851 22828 43852 22868
rect 43892 22828 43893 22868
rect 43851 22819 43893 22828
rect 44139 22868 44181 22877
rect 44139 22828 44140 22868
rect 44180 22828 44181 22868
rect 44139 22819 44181 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 4099 22532 4157 22533
rect 4099 22492 4108 22532
rect 4148 22492 4157 22532
rect 4099 22491 4157 22492
rect 6411 22532 6453 22541
rect 6411 22492 6412 22532
rect 6452 22492 6453 22532
rect 6411 22483 6453 22492
rect 8515 22532 8573 22533
rect 8515 22492 8524 22532
rect 8564 22492 8573 22532
rect 8515 22491 8573 22492
rect 11971 22532 12029 22533
rect 11971 22492 11980 22532
rect 12020 22492 12029 22532
rect 11971 22491 12029 22492
rect 14179 22532 14237 22533
rect 14179 22492 14188 22532
rect 14228 22492 14237 22532
rect 14179 22491 14237 22492
rect 14859 22532 14901 22541
rect 14859 22492 14860 22532
rect 14900 22492 14901 22532
rect 14859 22483 14901 22492
rect 16299 22532 16341 22541
rect 16299 22492 16300 22532
rect 16340 22492 16341 22532
rect 16299 22483 16341 22492
rect 22339 22532 22397 22533
rect 22339 22492 22348 22532
rect 22388 22492 22397 22532
rect 22339 22491 22397 22492
rect 29155 22532 29213 22533
rect 29155 22492 29164 22532
rect 29204 22492 29213 22532
rect 29155 22491 29213 22492
rect 34251 22532 34293 22541
rect 34251 22492 34252 22532
rect 34292 22492 34293 22532
rect 34251 22483 34293 22492
rect 39715 22532 39773 22533
rect 39715 22492 39724 22532
rect 39764 22492 39773 22532
rect 39715 22491 39773 22492
rect 41451 22532 41493 22541
rect 41451 22492 41452 22532
rect 41492 22492 41493 22532
rect 41451 22483 41493 22492
rect 43083 22532 43125 22541
rect 43083 22492 43084 22532
rect 43124 22492 43125 22532
rect 43083 22483 43125 22492
rect 48355 22532 48413 22533
rect 48355 22492 48364 22532
rect 48404 22492 48413 22532
rect 48355 22491 48413 22492
rect 1515 22448 1557 22457
rect 1515 22408 1516 22448
rect 1556 22408 1557 22448
rect 1515 22399 1557 22408
rect 5931 22448 5973 22457
rect 5931 22408 5932 22448
rect 5972 22408 5973 22448
rect 5931 22399 5973 22408
rect 12931 22448 12989 22449
rect 12931 22408 12940 22448
rect 12980 22408 12989 22448
rect 12931 22407 12989 22408
rect 19755 22448 19797 22457
rect 19755 22408 19756 22448
rect 19796 22408 19797 22448
rect 19755 22399 19797 22408
rect 23403 22448 23445 22457
rect 23403 22408 23404 22448
rect 23444 22408 23445 22448
rect 23403 22399 23445 22408
rect 27243 22448 27285 22457
rect 27243 22408 27244 22448
rect 27284 22408 27285 22448
rect 27243 22399 27285 22408
rect 47595 22448 47637 22457
rect 47595 22408 47596 22448
rect 47636 22408 47637 22448
rect 47595 22399 47637 22408
rect 51619 22448 51677 22449
rect 51619 22408 51628 22448
rect 51668 22408 51677 22448
rect 51619 22407 51677 22408
rect 34443 22364 34485 22373
rect 34443 22324 34444 22364
rect 34484 22324 34485 22364
rect 34443 22315 34485 22324
rect 40387 22364 40445 22365
rect 40387 22324 40396 22364
rect 40436 22324 40445 22364
rect 40387 22323 40445 22324
rect 2083 22280 2141 22281
rect 2083 22240 2092 22280
rect 2132 22240 2141 22280
rect 2083 22239 2141 22240
rect 2947 22280 3005 22281
rect 2947 22240 2956 22280
rect 2996 22240 3005 22280
rect 2947 22239 3005 22240
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4395 22280 4437 22289
rect 4395 22240 4396 22280
rect 4436 22240 4437 22280
rect 4395 22231 4437 22240
rect 4491 22280 4533 22289
rect 4491 22240 4492 22280
rect 4532 22240 4533 22280
rect 4491 22231 4533 22240
rect 4587 22280 4629 22289
rect 4587 22240 4588 22280
rect 4628 22240 4629 22280
rect 4587 22231 4629 22240
rect 4779 22280 4821 22289
rect 4779 22240 4780 22280
rect 4820 22240 4821 22280
rect 4779 22231 4821 22240
rect 4971 22280 5013 22289
rect 4971 22240 4972 22280
rect 5012 22240 5013 22280
rect 4971 22231 5013 22240
rect 5059 22280 5117 22281
rect 5059 22240 5068 22280
rect 5108 22240 5117 22280
rect 5059 22239 5117 22240
rect 5539 22280 5597 22281
rect 5539 22240 5548 22280
rect 5588 22240 5597 22280
rect 5539 22239 5597 22240
rect 6115 22280 6173 22281
rect 6115 22240 6124 22280
rect 6164 22240 6173 22280
rect 6115 22239 6173 22240
rect 6219 22280 6261 22289
rect 6219 22240 6220 22280
rect 6260 22240 6261 22280
rect 6219 22231 6261 22240
rect 6411 22280 6453 22289
rect 6411 22240 6412 22280
rect 6452 22240 6453 22280
rect 6411 22231 6453 22240
rect 7267 22280 7325 22281
rect 7267 22240 7276 22280
rect 7316 22240 7325 22280
rect 7267 22239 7325 22240
rect 7467 22280 7509 22289
rect 7467 22240 7468 22280
rect 7508 22240 7509 22280
rect 7467 22231 7509 22240
rect 7555 22280 7613 22281
rect 7555 22240 7564 22280
rect 7604 22240 7613 22280
rect 7555 22239 7613 22240
rect 7843 22280 7901 22281
rect 7843 22240 7852 22280
rect 7892 22240 7901 22280
rect 7843 22239 7901 22240
rect 8139 22280 8181 22289
rect 8139 22240 8140 22280
rect 8180 22240 8181 22280
rect 8139 22231 8181 22240
rect 9283 22280 9341 22281
rect 9283 22240 9292 22280
rect 9332 22240 9341 22280
rect 9283 22239 9341 22240
rect 9579 22280 9621 22289
rect 9579 22240 9580 22280
rect 9620 22240 9621 22280
rect 9579 22231 9621 22240
rect 9955 22280 10013 22281
rect 9955 22240 9964 22280
rect 10004 22240 10013 22280
rect 9955 22239 10013 22240
rect 10819 22280 10877 22281
rect 10819 22240 10828 22280
rect 10868 22240 10877 22280
rect 10819 22239 10877 22240
rect 12259 22280 12317 22281
rect 12259 22240 12268 22280
rect 12308 22240 12317 22280
rect 12259 22239 12317 22240
rect 12555 22280 12597 22289
rect 12555 22240 12556 22280
rect 12596 22240 12597 22280
rect 12555 22231 12597 22240
rect 12651 22280 12693 22289
rect 12651 22240 12652 22280
rect 12692 22240 12693 22280
rect 12651 22231 12693 22240
rect 13507 22280 13565 22281
rect 13507 22240 13516 22280
rect 13556 22240 13565 22280
rect 13507 22239 13565 22240
rect 13803 22280 13845 22289
rect 13803 22240 13804 22280
rect 13844 22240 13845 22280
rect 13803 22231 13845 22240
rect 14563 22280 14621 22281
rect 14563 22240 14572 22280
rect 14612 22240 14621 22280
rect 14563 22239 14621 22240
rect 14667 22280 14709 22289
rect 14667 22240 14668 22280
rect 14708 22240 14709 22280
rect 14667 22231 14709 22240
rect 14859 22280 14901 22289
rect 14859 22240 14860 22280
rect 14900 22240 14901 22280
rect 14859 22231 14901 22240
rect 15139 22280 15197 22281
rect 15139 22240 15148 22280
rect 15188 22240 15197 22280
rect 15139 22239 15197 22240
rect 16099 22280 16157 22281
rect 16099 22240 16108 22280
rect 16148 22240 16157 22280
rect 16099 22239 16157 22240
rect 16387 22280 16445 22281
rect 16387 22240 16396 22280
rect 16436 22240 16445 22280
rect 16387 22239 16445 22240
rect 16587 22280 16629 22289
rect 16587 22240 16588 22280
rect 16628 22240 16629 22280
rect 16587 22231 16629 22240
rect 17251 22280 17309 22281
rect 17251 22240 17260 22280
rect 17300 22240 17309 22280
rect 17251 22239 17309 22240
rect 17451 22280 17493 22289
rect 17451 22240 17452 22280
rect 17492 22240 17493 22280
rect 17451 22231 17493 22240
rect 17547 22280 17589 22289
rect 17547 22240 17548 22280
rect 17588 22240 17589 22280
rect 17547 22231 17589 22240
rect 17643 22280 17685 22289
rect 17643 22240 17644 22280
rect 17684 22240 17685 22280
rect 17643 22231 17685 22240
rect 17739 22280 17781 22289
rect 17739 22240 17740 22280
rect 17780 22240 17781 22280
rect 17739 22231 17781 22240
rect 18211 22280 18269 22281
rect 18211 22240 18220 22280
rect 18260 22240 18269 22280
rect 18211 22239 18269 22240
rect 20323 22280 20381 22281
rect 20323 22240 20332 22280
rect 20372 22240 20381 22280
rect 20323 22239 20381 22240
rect 21187 22280 21245 22281
rect 21187 22240 21196 22280
rect 21236 22240 21245 22280
rect 21187 22239 21245 22240
rect 23203 22280 23261 22281
rect 23203 22240 23212 22280
rect 23252 22240 23261 22280
rect 23203 22239 23261 22240
rect 24355 22280 24413 22281
rect 24355 22240 24364 22280
rect 24404 22240 24413 22280
rect 24355 22239 24413 22240
rect 30307 22280 30365 22281
rect 30307 22240 30316 22280
rect 30356 22240 30365 22280
rect 30307 22239 30365 22240
rect 31171 22280 31229 22281
rect 31171 22240 31180 22280
rect 31220 22240 31229 22280
rect 31171 22239 31229 22240
rect 32419 22280 32477 22281
rect 32419 22240 32428 22280
rect 32468 22240 32477 22280
rect 32419 22239 32477 22240
rect 32619 22280 32661 22289
rect 32619 22240 32620 22280
rect 32660 22240 32661 22280
rect 32619 22231 32661 22240
rect 32811 22280 32853 22289
rect 32811 22240 32812 22280
rect 32852 22240 32853 22280
rect 32811 22231 32853 22240
rect 32899 22280 32957 22281
rect 32899 22240 32908 22280
rect 32948 22240 32957 22280
rect 32899 22239 32957 22240
rect 33763 22280 33821 22281
rect 33763 22240 33772 22280
rect 33812 22240 33821 22280
rect 33763 22239 33821 22240
rect 34147 22280 34205 22281
rect 34147 22240 34156 22280
rect 34196 22240 34205 22280
rect 34147 22239 34205 22240
rect 34531 22280 34589 22281
rect 34531 22240 34540 22280
rect 34580 22240 34589 22280
rect 34531 22239 34589 22240
rect 34819 22280 34877 22281
rect 34819 22240 34828 22280
rect 34868 22240 34877 22280
rect 34819 22239 34877 22240
rect 35691 22280 35733 22289
rect 35691 22240 35692 22280
rect 35732 22240 35733 22280
rect 35691 22231 35733 22240
rect 37699 22280 37757 22281
rect 37699 22240 37708 22280
rect 37748 22240 37757 22280
rect 37699 22239 37757 22240
rect 38563 22280 38621 22281
rect 38563 22240 38572 22280
rect 38612 22240 38621 22280
rect 38563 22239 38621 22240
rect 40195 22280 40253 22281
rect 40195 22240 40204 22280
rect 40244 22240 40253 22280
rect 40195 22239 40253 22240
rect 40779 22280 40821 22289
rect 40779 22240 40780 22280
rect 40820 22240 40821 22280
rect 40779 22231 40821 22240
rect 40875 22280 40917 22289
rect 40875 22240 40876 22280
rect 40916 22240 40917 22280
rect 40875 22231 40917 22240
rect 40963 22280 41021 22281
rect 40963 22240 40972 22280
rect 41012 22240 41021 22280
rect 40963 22239 41021 22240
rect 41155 22280 41213 22281
rect 41155 22240 41164 22280
rect 41204 22240 41213 22280
rect 41155 22239 41213 22240
rect 41259 22280 41301 22289
rect 41259 22240 41260 22280
rect 41300 22240 41301 22280
rect 41259 22231 41301 22240
rect 41451 22280 41493 22289
rect 41451 22240 41452 22280
rect 41492 22240 41493 22280
rect 41451 22231 41493 22240
rect 41643 22280 41685 22289
rect 41643 22240 41644 22280
rect 41684 22240 41685 22280
rect 41643 22231 41685 22240
rect 41739 22280 41781 22289
rect 41739 22240 41740 22280
rect 41780 22240 41781 22280
rect 41739 22231 41781 22240
rect 41835 22280 41877 22289
rect 41835 22240 41836 22280
rect 41876 22240 41877 22280
rect 41835 22231 41877 22240
rect 41931 22280 41973 22289
rect 41931 22240 41932 22280
rect 41972 22240 41973 22280
rect 41931 22231 41973 22240
rect 42787 22280 42845 22281
rect 42787 22240 42796 22280
rect 42836 22240 42845 22280
rect 42787 22239 42845 22240
rect 42987 22280 43029 22289
rect 42987 22240 42988 22280
rect 43028 22240 43029 22280
rect 42987 22231 43029 22240
rect 43171 22280 43229 22281
rect 43171 22240 43180 22280
rect 43220 22240 43229 22280
rect 43171 22239 43229 22240
rect 43363 22280 43421 22281
rect 43363 22240 43372 22280
rect 43412 22240 43421 22280
rect 43363 22239 43421 22240
rect 43467 22280 43509 22289
rect 43467 22240 43468 22280
rect 43508 22240 43509 22280
rect 43467 22231 43509 22240
rect 43659 22280 43701 22289
rect 43659 22240 43660 22280
rect 43700 22240 43701 22280
rect 43659 22231 43701 22240
rect 43851 22280 43893 22289
rect 43851 22240 43852 22280
rect 43892 22240 43893 22280
rect 43851 22231 43893 22240
rect 43947 22280 43989 22289
rect 43947 22240 43948 22280
rect 43988 22240 43989 22280
rect 43947 22231 43989 22240
rect 44043 22280 44085 22289
rect 44043 22240 44044 22280
rect 44084 22240 44085 22280
rect 44043 22231 44085 22240
rect 44139 22280 44181 22289
rect 44139 22240 44140 22280
rect 44180 22240 44181 22280
rect 44139 22231 44181 22240
rect 44331 22280 44373 22289
rect 44331 22240 44332 22280
rect 44372 22240 44373 22280
rect 44331 22231 44373 22240
rect 44427 22280 44469 22289
rect 44427 22240 44428 22280
rect 44468 22240 44469 22280
rect 44427 22231 44469 22240
rect 44523 22280 44565 22289
rect 44523 22240 44524 22280
rect 44564 22240 44565 22280
rect 44523 22231 44565 22240
rect 44803 22280 44861 22281
rect 44803 22240 44812 22280
rect 44852 22240 44861 22280
rect 44803 22239 44861 22240
rect 44995 22280 45053 22281
rect 44995 22240 45004 22280
rect 45044 22240 45053 22280
rect 44995 22239 45053 22240
rect 45379 22280 45437 22281
rect 45379 22240 45388 22280
rect 45428 22240 45437 22280
rect 45379 22239 45437 22240
rect 45579 22280 45621 22289
rect 45579 22240 45580 22280
rect 45620 22240 45621 22280
rect 45579 22231 45621 22240
rect 45771 22280 45813 22289
rect 45771 22240 45772 22280
rect 45812 22240 45813 22280
rect 45771 22231 45813 22240
rect 45859 22280 45917 22281
rect 45859 22240 45868 22280
rect 45908 22240 45917 22280
rect 45859 22239 45917 22240
rect 46059 22280 46101 22289
rect 46059 22240 46060 22280
rect 46100 22240 46101 22280
rect 46059 22231 46101 22240
rect 46155 22280 46197 22289
rect 46155 22240 46156 22280
rect 46196 22240 46197 22280
rect 46155 22231 46197 22240
rect 46251 22280 46293 22289
rect 46251 22240 46252 22280
rect 46292 22240 46293 22280
rect 46251 22231 46293 22240
rect 46347 22280 46389 22289
rect 46347 22240 46348 22280
rect 46388 22240 46389 22280
rect 46347 22231 46389 22240
rect 47203 22280 47261 22281
rect 47203 22240 47212 22280
rect 47252 22240 47261 22280
rect 47203 22239 47261 22240
rect 47779 22280 47837 22281
rect 47779 22240 47788 22280
rect 47828 22240 47837 22280
rect 47779 22239 47837 22240
rect 47883 22280 47925 22289
rect 47883 22240 47884 22280
rect 47924 22240 47925 22280
rect 47883 22231 47925 22240
rect 48075 22280 48117 22289
rect 48075 22240 48076 22280
rect 48116 22240 48117 22280
rect 48075 22231 48117 22240
rect 49027 22280 49085 22281
rect 49027 22240 49036 22280
rect 49076 22240 49085 22280
rect 49027 22239 49085 22240
rect 49603 22280 49661 22281
rect 49603 22240 49612 22280
rect 49652 22240 49661 22280
rect 49603 22239 49661 22240
rect 50467 22280 50525 22281
rect 50467 22240 50476 22280
rect 50516 22240 50525 22280
rect 50467 22239 50525 22240
rect 1707 22196 1749 22205
rect 1707 22156 1708 22196
rect 1748 22156 1749 22196
rect 1707 22147 1749 22156
rect 4875 22196 4917 22205
rect 4875 22156 4876 22196
rect 4916 22156 4917 22196
rect 4875 22147 4917 22156
rect 8235 22196 8277 22205
rect 8235 22156 8236 22196
rect 8276 22156 8277 22196
rect 8235 22147 8277 22156
rect 13899 22196 13941 22205
rect 13899 22156 13900 22196
rect 13940 22156 13941 22196
rect 13899 22147 13941 22156
rect 19947 22196 19989 22205
rect 19947 22156 19948 22196
rect 19988 22156 19989 22196
rect 19947 22147 19989 22156
rect 31563 22196 31605 22205
rect 31563 22156 31564 22196
rect 31604 22156 31605 22196
rect 31563 22147 31605 22156
rect 31755 22196 31797 22205
rect 31755 22156 31756 22196
rect 31796 22156 31797 22196
rect 31755 22147 31797 22156
rect 32715 22196 32757 22205
rect 32715 22156 32716 22196
rect 32756 22156 32757 22196
rect 32715 22147 32757 22156
rect 37323 22196 37365 22205
rect 37323 22156 37324 22196
rect 37364 22156 37365 22196
rect 37323 22147 37365 22156
rect 40107 22196 40149 22205
rect 40107 22156 40108 22196
rect 40148 22156 40149 22196
rect 40107 22147 40149 22156
rect 45675 22196 45717 22205
rect 45675 22156 45676 22196
rect 45716 22156 45717 22196
rect 45675 22147 45717 22156
rect 46539 22196 46581 22205
rect 46539 22156 46540 22196
rect 46580 22156 46581 22196
rect 46539 22147 46581 22156
rect 47979 22196 48021 22205
rect 47979 22156 47980 22196
rect 48020 22156 48021 22196
rect 47979 22147 48021 22156
rect 49227 22196 49269 22205
rect 49227 22156 49228 22196
rect 49268 22156 49269 22196
rect 49227 22147 49269 22156
rect 643 22112 701 22113
rect 643 22072 652 22112
rect 692 22072 701 22112
rect 643 22071 701 22072
rect 5451 22112 5493 22121
rect 5451 22072 5452 22112
rect 5492 22072 5493 22112
rect 5451 22063 5493 22072
rect 6595 22112 6653 22113
rect 6595 22072 6604 22112
rect 6644 22072 6653 22112
rect 6595 22071 6653 22072
rect 9387 22112 9429 22121
rect 9387 22072 9388 22112
rect 9428 22072 9429 22112
rect 9387 22063 9429 22072
rect 18699 22112 18741 22121
rect 18699 22072 18700 22112
rect 18740 22072 18741 22112
rect 18699 22063 18741 22072
rect 22531 22112 22589 22113
rect 22531 22072 22540 22112
rect 22580 22072 22589 22112
rect 22531 22071 22589 22072
rect 24163 22112 24221 22113
rect 24163 22072 24172 22112
rect 24212 22072 24221 22112
rect 24163 22071 24221 22072
rect 24451 22112 24509 22113
rect 24451 22072 24460 22112
rect 24500 22072 24509 22112
rect 24451 22071 24509 22072
rect 33091 22112 33149 22113
rect 33091 22072 33100 22112
rect 33140 22072 33149 22112
rect 33091 22071 33149 22072
rect 42115 22112 42173 22113
rect 42115 22072 42124 22112
rect 42164 22072 42173 22112
rect 42115 22071 42173 22072
rect 43555 22112 43613 22113
rect 43555 22072 43564 22112
rect 43604 22072 43613 22112
rect 43555 22071 43613 22072
rect 44611 22112 44669 22113
rect 44611 22072 44620 22112
rect 44660 22072 44669 22112
rect 44611 22071 44669 22072
rect 45291 22112 45333 22121
rect 45291 22072 45292 22112
rect 45332 22072 45333 22112
rect 45291 22063 45333 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 4483 21776 4541 21777
rect 4483 21736 4492 21776
rect 4532 21736 4541 21776
rect 4483 21735 4541 21736
rect 5539 21776 5597 21777
rect 5539 21736 5548 21776
rect 5588 21736 5597 21776
rect 5539 21735 5597 21736
rect 16387 21776 16445 21777
rect 16387 21736 16396 21776
rect 16436 21736 16445 21776
rect 16387 21735 16445 21736
rect 18979 21776 19037 21777
rect 18979 21736 18988 21776
rect 19028 21736 19037 21776
rect 18979 21735 19037 21736
rect 19459 21776 19517 21777
rect 19459 21736 19468 21776
rect 19508 21736 19517 21776
rect 19459 21735 19517 21736
rect 22635 21776 22677 21785
rect 22635 21736 22636 21776
rect 22676 21736 22677 21776
rect 22635 21727 22677 21736
rect 25891 21776 25949 21777
rect 25891 21736 25900 21776
rect 25940 21736 25949 21776
rect 25891 21735 25949 21736
rect 26475 21776 26517 21785
rect 26475 21736 26476 21776
rect 26516 21736 26517 21776
rect 26475 21727 26517 21736
rect 29155 21776 29213 21777
rect 29155 21736 29164 21776
rect 29204 21736 29213 21776
rect 29155 21735 29213 21736
rect 32611 21776 32669 21777
rect 32611 21736 32620 21776
rect 32660 21736 32669 21776
rect 32611 21735 32669 21736
rect 35203 21776 35261 21777
rect 35203 21736 35212 21776
rect 35252 21736 35261 21776
rect 35203 21735 35261 21736
rect 39331 21776 39389 21777
rect 39331 21736 39340 21776
rect 39380 21736 39389 21776
rect 39331 21735 39389 21736
rect 41251 21776 41309 21777
rect 41251 21736 41260 21776
rect 41300 21736 41309 21776
rect 41251 21735 41309 21736
rect 42603 21776 42645 21785
rect 42603 21736 42604 21776
rect 42644 21736 42645 21776
rect 42603 21727 42645 21736
rect 45195 21776 45237 21785
rect 45195 21736 45196 21776
rect 45236 21736 45237 21776
rect 45195 21727 45237 21736
rect 46155 21776 46197 21785
rect 46155 21736 46156 21776
rect 46196 21736 46197 21776
rect 46155 21727 46197 21736
rect 6123 21692 6165 21701
rect 6123 21652 6124 21692
rect 6164 21652 6165 21692
rect 6123 21643 6165 21652
rect 13995 21692 14037 21701
rect 13995 21652 13996 21692
rect 14036 21652 14037 21692
rect 13995 21643 14037 21652
rect 16587 21692 16629 21701
rect 16587 21652 16588 21692
rect 16628 21652 16629 21692
rect 16587 21643 16629 21652
rect 26763 21692 26805 21701
rect 26763 21652 26764 21692
rect 26804 21652 26805 21692
rect 26763 21643 26805 21652
rect 32811 21692 32853 21701
rect 32811 21652 32812 21692
rect 32852 21652 32853 21692
rect 32811 21643 32853 21652
rect 38379 21692 38421 21701
rect 38379 21652 38380 21692
rect 38420 21652 38421 21692
rect 38379 21643 38421 21652
rect 47595 21692 47637 21701
rect 47595 21652 47596 21692
rect 47636 21652 47637 21692
rect 47595 21643 47637 21652
rect 2091 21608 2133 21617
rect 2091 21568 2092 21608
rect 2132 21568 2133 21608
rect 2091 21559 2133 21568
rect 2467 21608 2525 21609
rect 2467 21568 2476 21608
rect 2516 21568 2525 21608
rect 2467 21567 2525 21568
rect 3331 21608 3389 21609
rect 3331 21568 3340 21608
rect 3380 21568 3389 21608
rect 3331 21567 3389 21568
rect 4867 21608 4925 21609
rect 4867 21568 4876 21608
rect 4916 21568 4925 21608
rect 4867 21567 4925 21568
rect 5067 21608 5109 21617
rect 5067 21568 5068 21608
rect 5108 21568 5109 21608
rect 5067 21559 5109 21568
rect 5259 21608 5301 21617
rect 5259 21568 5260 21608
rect 5300 21568 5301 21608
rect 5259 21559 5301 21568
rect 5347 21608 5405 21609
rect 5347 21568 5356 21608
rect 5396 21568 5405 21608
rect 5347 21567 5405 21568
rect 5643 21608 5685 21617
rect 5643 21568 5644 21608
rect 5684 21568 5685 21608
rect 5643 21559 5685 21568
rect 5739 21608 5781 21617
rect 5739 21568 5740 21608
rect 5780 21568 5781 21608
rect 5739 21559 5781 21568
rect 5835 21608 5877 21617
rect 5835 21568 5836 21608
rect 5876 21568 5877 21608
rect 5835 21559 5877 21568
rect 6499 21608 6557 21609
rect 6499 21568 6508 21608
rect 6548 21568 6557 21608
rect 6499 21567 6557 21568
rect 7363 21608 7421 21609
rect 7363 21568 7372 21608
rect 7412 21568 7421 21608
rect 7363 21567 7421 21568
rect 9579 21608 9621 21617
rect 9579 21568 9580 21608
rect 9620 21568 9621 21608
rect 9579 21559 9621 21568
rect 9675 21608 9717 21617
rect 9675 21568 9676 21608
rect 9716 21568 9717 21608
rect 9675 21559 9717 21568
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 9867 21608 9909 21617
rect 9867 21568 9868 21608
rect 9908 21568 9909 21608
rect 9867 21559 9909 21568
rect 10147 21608 10205 21609
rect 10147 21568 10156 21608
rect 10196 21568 10205 21608
rect 10147 21567 10205 21568
rect 11307 21608 11349 21617
rect 11307 21568 11308 21608
rect 11348 21568 11349 21608
rect 11307 21559 11349 21568
rect 11403 21608 11445 21617
rect 11403 21568 11404 21608
rect 11444 21568 11445 21608
rect 11403 21559 11445 21568
rect 11499 21608 11541 21617
rect 11499 21568 11500 21608
rect 11540 21568 11541 21608
rect 11499 21559 11541 21568
rect 11595 21608 11637 21617
rect 11595 21568 11596 21608
rect 11636 21568 11637 21608
rect 11595 21559 11637 21568
rect 11779 21608 11837 21609
rect 11779 21568 11788 21608
rect 11828 21568 11837 21608
rect 11779 21567 11837 21568
rect 13027 21608 13085 21609
rect 13027 21568 13036 21608
rect 13076 21568 13085 21608
rect 13027 21567 13085 21568
rect 14371 21608 14429 21609
rect 14371 21568 14380 21608
rect 14420 21568 14429 21608
rect 14371 21567 14429 21568
rect 15235 21608 15293 21609
rect 15235 21568 15244 21608
rect 15284 21568 15293 21608
rect 15235 21567 15293 21568
rect 16963 21608 17021 21609
rect 16963 21568 16972 21608
rect 17012 21568 17021 21608
rect 16963 21567 17021 21568
rect 17827 21608 17885 21609
rect 17827 21568 17836 21608
rect 17876 21568 17885 21608
rect 17827 21567 17885 21568
rect 20995 21608 21053 21609
rect 20995 21568 21004 21608
rect 21044 21568 21053 21608
rect 20995 21567 21053 21568
rect 21195 21608 21237 21617
rect 21195 21568 21196 21608
rect 21236 21568 21237 21608
rect 21195 21559 21237 21568
rect 21291 21608 21333 21617
rect 21291 21568 21292 21608
rect 21332 21568 21333 21608
rect 21291 21559 21333 21568
rect 21387 21608 21429 21617
rect 21387 21568 21388 21608
rect 21428 21568 21429 21608
rect 21387 21559 21429 21568
rect 21483 21608 21525 21617
rect 21483 21568 21484 21608
rect 21524 21568 21525 21608
rect 21483 21559 21525 21568
rect 22539 21608 22581 21617
rect 22539 21568 22540 21608
rect 22580 21568 22581 21608
rect 22539 21559 22581 21568
rect 22731 21608 22773 21617
rect 22731 21568 22732 21608
rect 22772 21568 22773 21608
rect 22731 21559 22773 21568
rect 22923 21608 22965 21617
rect 22923 21568 22924 21608
rect 22964 21568 22965 21608
rect 22923 21559 22965 21568
rect 23587 21608 23645 21609
rect 23587 21568 23596 21608
rect 23636 21568 23645 21608
rect 23587 21567 23645 21568
rect 23787 21608 23829 21617
rect 23787 21568 23788 21608
rect 23828 21568 23829 21608
rect 23787 21559 23829 21568
rect 23979 21608 24021 21617
rect 23979 21568 23980 21608
rect 24020 21568 24021 21608
rect 23979 21559 24021 21568
rect 24843 21608 24885 21617
rect 24843 21568 24844 21608
rect 24884 21568 24885 21608
rect 24843 21559 24885 21568
rect 24939 21608 24981 21617
rect 24939 21568 24940 21608
rect 24980 21568 24981 21608
rect 24939 21559 24981 21568
rect 25035 21608 25077 21617
rect 25035 21568 25036 21608
rect 25076 21568 25077 21608
rect 25035 21559 25077 21568
rect 25131 21608 25173 21617
rect 25131 21568 25132 21608
rect 25172 21568 25173 21608
rect 25131 21559 25173 21568
rect 25323 21608 25365 21617
rect 25323 21568 25324 21608
rect 25364 21568 25365 21608
rect 25323 21559 25365 21568
rect 25419 21608 25461 21617
rect 25419 21568 25420 21608
rect 25460 21568 25461 21608
rect 25419 21559 25461 21568
rect 25515 21608 25557 21617
rect 25515 21568 25516 21608
rect 25556 21568 25557 21608
rect 25515 21559 25557 21568
rect 25611 21608 25653 21617
rect 25611 21568 25612 21608
rect 25652 21568 25653 21608
rect 25611 21559 25653 21568
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 25803 21559 25845 21568
rect 25995 21608 26037 21617
rect 25995 21568 25996 21608
rect 26036 21568 26037 21608
rect 25995 21559 26037 21568
rect 26083 21608 26141 21609
rect 26083 21568 26092 21608
rect 26132 21568 26141 21608
rect 26083 21567 26141 21568
rect 26379 21608 26421 21617
rect 26379 21568 26380 21608
rect 26420 21568 26421 21608
rect 26379 21559 26421 21568
rect 26571 21608 26613 21617
rect 26571 21568 26572 21608
rect 26612 21568 26613 21608
rect 26571 21559 26613 21568
rect 27139 21608 27197 21609
rect 27139 21568 27148 21608
rect 27188 21568 27197 21608
rect 27139 21567 27197 21568
rect 28003 21608 28061 21609
rect 28003 21568 28012 21608
rect 28052 21568 28061 21608
rect 28003 21567 28061 21568
rect 30979 21608 31037 21609
rect 30979 21568 30988 21608
rect 31028 21568 31037 21608
rect 30979 21567 31037 21568
rect 31083 21608 31125 21617
rect 31083 21568 31084 21608
rect 31124 21568 31125 21608
rect 31083 21559 31125 21568
rect 31275 21608 31317 21617
rect 31275 21568 31276 21608
rect 31316 21568 31317 21608
rect 31275 21559 31317 21568
rect 31467 21608 31509 21617
rect 31467 21568 31468 21608
rect 31508 21568 31509 21608
rect 31467 21559 31509 21568
rect 31563 21608 31605 21617
rect 31563 21568 31564 21608
rect 31604 21568 31605 21608
rect 31563 21559 31605 21568
rect 31659 21608 31701 21617
rect 31659 21568 31660 21608
rect 31700 21568 31701 21608
rect 31659 21559 31701 21568
rect 31755 21608 31797 21617
rect 31755 21568 31756 21608
rect 31796 21568 31797 21608
rect 31755 21559 31797 21568
rect 32331 21608 32373 21617
rect 32331 21568 32332 21608
rect 32372 21568 32373 21608
rect 32331 21559 32373 21568
rect 32427 21608 32469 21617
rect 32427 21568 32428 21608
rect 32468 21568 32469 21608
rect 32427 21559 32469 21568
rect 32523 21608 32565 21617
rect 32523 21568 32524 21608
rect 32564 21568 32565 21608
rect 32523 21559 32565 21568
rect 33187 21608 33245 21609
rect 33187 21568 33196 21608
rect 33236 21568 33245 21608
rect 33187 21567 33245 21568
rect 34051 21608 34109 21609
rect 34051 21568 34060 21608
rect 34100 21568 34109 21608
rect 34051 21567 34109 21568
rect 35587 21608 35645 21609
rect 35587 21568 35596 21608
rect 35636 21568 35645 21608
rect 35587 21567 35645 21568
rect 37411 21608 37469 21609
rect 37411 21568 37420 21608
rect 37460 21568 37469 21608
rect 37411 21567 37469 21568
rect 37899 21608 37941 21617
rect 37899 21568 37900 21608
rect 37940 21568 37941 21608
rect 37899 21559 37941 21568
rect 37995 21608 38037 21617
rect 37995 21568 37996 21608
rect 38036 21568 38037 21608
rect 37995 21559 38037 21568
rect 38091 21608 38133 21617
rect 38091 21568 38092 21608
rect 38132 21568 38133 21608
rect 38091 21559 38133 21568
rect 38187 21608 38229 21617
rect 38187 21568 38188 21608
rect 38228 21568 38229 21608
rect 38187 21559 38229 21568
rect 39043 21608 39101 21609
rect 39043 21568 39052 21608
rect 39092 21568 39101 21608
rect 39043 21567 39101 21568
rect 39243 21608 39285 21617
rect 39243 21568 39244 21608
rect 39284 21568 39285 21608
rect 39243 21559 39285 21568
rect 39435 21608 39477 21617
rect 39435 21568 39436 21608
rect 39476 21568 39477 21608
rect 39435 21559 39477 21568
rect 39523 21608 39581 21609
rect 39523 21568 39532 21608
rect 39572 21568 39581 21608
rect 39523 21567 39581 21568
rect 40299 21608 40341 21617
rect 40299 21568 40300 21608
rect 40340 21568 40341 21608
rect 40299 21559 40341 21568
rect 40395 21608 40437 21617
rect 40395 21568 40396 21608
rect 40436 21568 40437 21608
rect 40395 21559 40437 21568
rect 40491 21608 40533 21617
rect 40491 21568 40492 21608
rect 40532 21568 40533 21608
rect 40491 21559 40533 21568
rect 40587 21608 40629 21617
rect 40587 21568 40588 21608
rect 40628 21568 40629 21608
rect 40587 21559 40629 21568
rect 40779 21608 40821 21617
rect 40779 21568 40780 21608
rect 40820 21568 40821 21608
rect 40779 21559 40821 21568
rect 40971 21608 41013 21617
rect 40971 21568 40972 21608
rect 41012 21568 41013 21608
rect 40971 21559 41013 21568
rect 41059 21608 41117 21609
rect 41059 21568 41068 21608
rect 41108 21568 41117 21608
rect 41059 21567 41117 21568
rect 41923 21608 41981 21609
rect 41923 21568 41932 21608
rect 41972 21568 41981 21608
rect 41923 21567 41981 21568
rect 42115 21608 42173 21609
rect 42115 21568 42124 21608
rect 42164 21568 42173 21608
rect 42115 21567 42173 21568
rect 43075 21608 43133 21609
rect 43075 21568 43084 21608
rect 43124 21568 43133 21608
rect 43075 21567 43133 21568
rect 43371 21608 43413 21617
rect 43371 21568 43372 21608
rect 43412 21568 43413 21608
rect 43371 21559 43413 21568
rect 44035 21608 44093 21609
rect 44035 21568 44044 21608
rect 44084 21568 44093 21608
rect 44035 21567 44093 21568
rect 44227 21608 44285 21609
rect 44227 21568 44236 21608
rect 44276 21568 44285 21608
rect 44227 21567 44285 21568
rect 44331 21608 44373 21617
rect 44331 21568 44332 21608
rect 44372 21568 44373 21608
rect 44331 21559 44373 21568
rect 44523 21608 44565 21617
rect 44523 21568 44524 21608
rect 44564 21568 44565 21608
rect 44523 21559 44565 21568
rect 45579 21608 45621 21617
rect 45579 21568 45580 21608
rect 45620 21568 45621 21608
rect 45579 21559 45621 21568
rect 47019 21608 47061 21617
rect 47019 21568 47020 21608
rect 47060 21568 47061 21608
rect 47019 21559 47061 21568
rect 47115 21608 47157 21617
rect 47115 21568 47116 21608
rect 47156 21568 47157 21608
rect 47115 21559 47157 21568
rect 47211 21608 47253 21617
rect 47211 21568 47212 21608
rect 47252 21568 47253 21608
rect 47211 21559 47253 21568
rect 47307 21608 47349 21617
rect 47307 21568 47308 21608
rect 47348 21568 47349 21608
rect 47307 21559 47349 21568
rect 47499 21608 47541 21617
rect 47499 21568 47500 21608
rect 47540 21568 47541 21608
rect 47499 21559 47541 21568
rect 47691 21608 47733 21617
rect 47691 21568 47692 21608
rect 47732 21568 47733 21608
rect 47691 21559 47733 21568
rect 47779 21608 47837 21609
rect 47779 21568 47788 21608
rect 47828 21568 47837 21608
rect 47779 21567 47837 21568
rect 47971 21608 48029 21609
rect 47971 21568 47980 21608
rect 48020 21568 48029 21608
rect 47971 21567 48029 21568
rect 20131 21549 20189 21550
rect 8523 21524 8565 21533
rect 8523 21484 8524 21524
rect 8564 21484 8565 21524
rect 20131 21509 20140 21549
rect 20180 21509 20189 21549
rect 20131 21508 20189 21509
rect 21859 21524 21917 21525
rect 8523 21475 8565 21484
rect 21859 21484 21868 21524
rect 21908 21484 21917 21524
rect 21859 21483 21917 21484
rect 23883 21524 23925 21533
rect 23883 21484 23884 21524
rect 23924 21484 23925 21524
rect 23883 21475 23925 21484
rect 36459 21524 36501 21533
rect 36459 21484 36460 21524
rect 36500 21484 36501 21524
rect 36459 21475 36501 21484
rect 46339 21524 46397 21525
rect 46339 21484 46348 21524
rect 46388 21484 46397 21524
rect 46339 21483 46397 21484
rect 48651 21524 48693 21533
rect 48651 21484 48652 21524
rect 48692 21484 48693 21524
rect 48651 21475 48693 21484
rect 1899 21440 1941 21449
rect 1899 21400 1900 21440
rect 1940 21400 1941 21440
rect 1899 21391 1941 21400
rect 5067 21440 5109 21449
rect 5067 21400 5068 21440
rect 5108 21400 5109 21440
rect 5067 21391 5109 21400
rect 12651 21440 12693 21449
rect 12651 21400 12652 21440
rect 12692 21400 12693 21440
rect 12651 21391 12693 21400
rect 20323 21440 20381 21441
rect 20323 21400 20332 21440
rect 20372 21400 20381 21440
rect 20323 21399 20381 21400
rect 21675 21440 21717 21449
rect 21675 21400 21676 21440
rect 21716 21400 21717 21440
rect 21675 21391 21717 21400
rect 29835 21440 29877 21449
rect 29835 21400 29836 21440
rect 29876 21400 29877 21440
rect 29835 21391 29877 21400
rect 31275 21440 31317 21449
rect 31275 21400 31276 21440
rect 31316 21400 31317 21440
rect 31275 21391 31317 21400
rect 32139 21440 32181 21449
rect 32139 21400 32140 21440
rect 32180 21400 32181 21440
rect 32139 21391 32181 21400
rect 36739 21440 36797 21441
rect 36739 21400 36748 21440
rect 36788 21400 36797 21440
rect 36739 21399 36797 21400
rect 40107 21440 40149 21449
rect 40107 21400 40108 21440
rect 40148 21400 40149 21440
rect 40107 21391 40149 21400
rect 44523 21440 44565 21449
rect 44523 21400 44524 21440
rect 44564 21400 44565 21440
rect 44523 21391 44565 21400
rect 46731 21440 46773 21449
rect 46731 21400 46732 21440
rect 46772 21400 46773 21440
rect 46731 21391 46773 21400
rect 49035 21440 49077 21449
rect 49035 21400 49036 21440
rect 49076 21400 49077 21440
rect 49035 21391 49077 21400
rect 49707 21440 49749 21449
rect 49707 21400 49708 21440
rect 49748 21400 49749 21440
rect 49707 21391 49749 21400
rect 4779 21356 4821 21365
rect 4779 21316 4780 21356
rect 4820 21316 4821 21356
rect 4779 21307 4821 21316
rect 10443 21356 10485 21365
rect 10443 21316 10444 21356
rect 10484 21316 10485 21356
rect 10443 21307 10485 21316
rect 12451 21356 12509 21357
rect 12451 21316 12460 21356
rect 12500 21316 12509 21356
rect 12451 21315 12509 21316
rect 13131 21356 13173 21365
rect 13131 21316 13132 21356
rect 13172 21316 13173 21356
rect 13131 21307 13173 21316
rect 40779 21356 40821 21365
rect 40779 21316 40780 21356
rect 40820 21316 40821 21356
rect 40779 21307 40821 21316
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 4395 21020 4437 21029
rect 4395 20980 4396 21020
rect 4436 20980 4437 21020
rect 4395 20971 4437 20980
rect 6027 21020 6069 21029
rect 6027 20980 6028 21020
rect 6068 20980 6069 21020
rect 6027 20971 6069 20980
rect 14083 21020 14141 21021
rect 14083 20980 14092 21020
rect 14132 20980 14141 21020
rect 14083 20979 14141 20980
rect 14667 21020 14709 21029
rect 14667 20980 14668 21020
rect 14708 20980 14709 21020
rect 14667 20971 14709 20980
rect 15627 21020 15669 21029
rect 15627 20980 15628 21020
rect 15668 20980 15669 21020
rect 15627 20971 15669 20980
rect 25507 21020 25565 21021
rect 25507 20980 25516 21020
rect 25556 20980 25565 21020
rect 25507 20979 25565 20980
rect 32235 21020 32277 21029
rect 32235 20980 32236 21020
rect 32276 20980 32277 21020
rect 32235 20971 32277 20980
rect 33099 21020 33141 21029
rect 33099 20980 33100 21020
rect 33140 20980 33141 21020
rect 33099 20971 33141 20980
rect 42883 21020 42941 21021
rect 42883 20980 42892 21020
rect 42932 20980 42941 21020
rect 42883 20979 42941 20980
rect 44227 21020 44285 21021
rect 44227 20980 44236 21020
rect 44276 20980 44285 21020
rect 44227 20979 44285 20980
rect 10635 20936 10677 20945
rect 10635 20896 10636 20936
rect 10676 20896 10677 20936
rect 10635 20887 10677 20896
rect 16491 20936 16533 20945
rect 16491 20896 16492 20936
rect 16532 20896 16533 20936
rect 16491 20887 16533 20896
rect 17067 20936 17109 20945
rect 17067 20896 17068 20936
rect 17108 20896 17109 20936
rect 23787 20936 23829 20945
rect 17067 20887 17109 20896
rect 23595 20910 23637 20919
rect 23595 20870 23596 20910
rect 23636 20870 23637 20910
rect 23787 20896 23788 20936
rect 23828 20896 23829 20936
rect 23787 20887 23829 20896
rect 30027 20936 30069 20945
rect 30027 20896 30028 20936
rect 30068 20896 30069 20936
rect 30027 20887 30069 20896
rect 23595 20861 23637 20870
rect 6211 20852 6269 20853
rect 6211 20812 6220 20852
rect 6260 20812 6269 20852
rect 6211 20811 6269 20812
rect 19947 20852 19989 20861
rect 19947 20812 19948 20852
rect 19988 20812 19989 20852
rect 19947 20803 19989 20812
rect 30795 20852 30837 20861
rect 30795 20812 30796 20852
rect 30836 20812 30837 20852
rect 30795 20803 30837 20812
rect 39339 20852 39381 20861
rect 39339 20812 39340 20852
rect 39380 20812 39381 20852
rect 39339 20803 39381 20812
rect 21671 20787 21729 20788
rect 21571 20782 21629 20783
rect 4483 20768 4541 20769
rect 4483 20728 4492 20768
rect 4532 20728 4541 20768
rect 4483 20727 4541 20728
rect 4683 20768 4725 20777
rect 4683 20728 4684 20768
rect 4724 20728 4725 20768
rect 4683 20719 4725 20728
rect 4779 20768 4821 20777
rect 4779 20728 4780 20768
rect 4820 20728 4821 20768
rect 4779 20719 4821 20728
rect 4875 20768 4917 20777
rect 4875 20728 4876 20768
rect 4916 20728 4917 20768
rect 4875 20719 4917 20728
rect 4971 20768 5013 20777
rect 4971 20728 4972 20768
rect 5012 20728 5013 20768
rect 4971 20719 5013 20728
rect 5547 20768 5589 20777
rect 5547 20728 5548 20768
rect 5588 20728 5589 20768
rect 5547 20719 5589 20728
rect 5739 20768 5781 20777
rect 5739 20728 5740 20768
rect 5780 20728 5781 20768
rect 5739 20719 5781 20728
rect 6411 20768 6453 20777
rect 6411 20728 6412 20768
rect 6452 20728 6453 20768
rect 6411 20719 6453 20728
rect 6507 20768 6549 20777
rect 6507 20728 6508 20768
rect 6548 20728 6549 20768
rect 6507 20719 6549 20728
rect 6603 20768 6645 20777
rect 6603 20728 6604 20768
rect 6644 20728 6645 20768
rect 6603 20719 6645 20728
rect 6699 20768 6741 20777
rect 6699 20728 6700 20768
rect 6740 20728 6741 20768
rect 6699 20719 6741 20728
rect 6883 20768 6941 20769
rect 6883 20728 6892 20768
rect 6932 20728 6941 20768
rect 6883 20727 6941 20728
rect 7755 20768 7797 20777
rect 7755 20728 7756 20768
rect 7796 20728 7797 20768
rect 7755 20719 7797 20728
rect 8803 20768 8861 20769
rect 8803 20728 8812 20768
rect 8852 20728 8861 20768
rect 8803 20727 8861 20728
rect 8907 20768 8949 20777
rect 8907 20728 8908 20768
rect 8948 20728 8949 20768
rect 8907 20719 8949 20728
rect 9099 20768 9141 20777
rect 9099 20728 9100 20768
rect 9140 20728 9141 20768
rect 9099 20719 9141 20728
rect 9955 20768 10013 20769
rect 9955 20728 9964 20768
rect 10004 20728 10013 20768
rect 9955 20727 10013 20728
rect 10339 20768 10397 20769
rect 10339 20728 10348 20768
rect 10388 20728 10397 20768
rect 10339 20727 10397 20728
rect 10443 20768 10485 20777
rect 10443 20728 10444 20768
rect 10484 20728 10485 20768
rect 10443 20719 10485 20728
rect 10635 20768 10677 20777
rect 10635 20728 10636 20768
rect 10676 20728 10677 20768
rect 10635 20719 10677 20728
rect 10819 20768 10877 20769
rect 10819 20728 10828 20768
rect 10868 20728 10877 20768
rect 10819 20727 10877 20728
rect 12067 20768 12125 20769
rect 12067 20728 12076 20768
rect 12116 20728 12125 20768
rect 12067 20727 12125 20728
rect 12931 20768 12989 20769
rect 12931 20728 12940 20768
rect 12980 20728 12989 20768
rect 12931 20727 12989 20728
rect 14563 20768 14621 20769
rect 14563 20728 14572 20768
rect 14612 20728 14621 20768
rect 14563 20727 14621 20728
rect 15139 20768 15197 20769
rect 15139 20728 15148 20768
rect 15188 20728 15197 20768
rect 15139 20727 15197 20728
rect 19851 20768 19893 20777
rect 19851 20728 19852 20768
rect 19892 20728 19893 20768
rect 19851 20719 19893 20728
rect 20043 20768 20085 20777
rect 20043 20728 20044 20768
rect 20084 20728 20085 20768
rect 20043 20719 20085 20728
rect 20515 20768 20573 20769
rect 20515 20728 20524 20768
rect 20564 20728 20573 20768
rect 20515 20727 20573 20728
rect 20611 20768 20669 20769
rect 20611 20728 20620 20768
rect 20660 20728 20669 20768
rect 20611 20727 20669 20728
rect 21387 20768 21429 20777
rect 21387 20728 21388 20768
rect 21428 20728 21429 20768
rect 21571 20742 21580 20782
rect 21620 20742 21629 20782
rect 21671 20747 21680 20787
rect 21720 20747 21729 20787
rect 38379 20782 38421 20791
rect 21671 20746 21729 20747
rect 21867 20768 21909 20777
rect 21571 20741 21629 20742
rect 21387 20719 21429 20728
rect 21867 20728 21868 20768
rect 21908 20728 21909 20768
rect 21867 20719 21909 20728
rect 21963 20768 22005 20777
rect 21963 20728 21964 20768
rect 22004 20728 22005 20768
rect 21963 20719 22005 20728
rect 22059 20768 22101 20777
rect 22059 20728 22060 20768
rect 22100 20728 22101 20768
rect 22059 20719 22101 20728
rect 22539 20768 22581 20777
rect 22539 20728 22540 20768
rect 22580 20728 22581 20768
rect 22539 20719 22581 20728
rect 22635 20768 22677 20777
rect 22635 20728 22636 20768
rect 22676 20728 22677 20768
rect 22635 20719 22677 20728
rect 22731 20768 22773 20777
rect 22731 20728 22732 20768
rect 22772 20728 22773 20768
rect 22731 20719 22773 20728
rect 22827 20768 22869 20777
rect 22827 20728 22828 20768
rect 22868 20728 22869 20768
rect 22827 20719 22869 20728
rect 23019 20768 23061 20777
rect 23019 20728 23020 20768
rect 23060 20728 23061 20768
rect 23019 20719 23061 20728
rect 23115 20768 23157 20777
rect 23115 20728 23116 20768
rect 23156 20728 23157 20768
rect 23115 20719 23157 20728
rect 23211 20768 23253 20777
rect 23211 20728 23212 20768
rect 23252 20728 23253 20768
rect 23211 20719 23253 20728
rect 23307 20768 23349 20777
rect 23307 20728 23308 20768
rect 23348 20728 23349 20768
rect 23307 20719 23349 20728
rect 23595 20768 23637 20777
rect 23595 20728 23596 20768
rect 23636 20728 23637 20768
rect 23595 20719 23637 20728
rect 24075 20768 24117 20777
rect 24075 20728 24076 20768
rect 24116 20728 24117 20768
rect 24075 20719 24117 20728
rect 24171 20768 24213 20777
rect 24171 20728 24172 20768
rect 24212 20728 24213 20768
rect 24171 20719 24213 20728
rect 24267 20768 24309 20777
rect 24267 20728 24268 20768
rect 24308 20728 24309 20768
rect 24267 20719 24309 20728
rect 25027 20768 25085 20769
rect 25027 20728 25036 20768
rect 25076 20728 25085 20768
rect 25027 20727 25085 20728
rect 25227 20768 25269 20777
rect 25227 20728 25228 20768
rect 25268 20728 25269 20768
rect 25227 20719 25269 20728
rect 25315 20768 25373 20769
rect 25315 20728 25324 20768
rect 25364 20728 25373 20768
rect 25315 20727 25373 20728
rect 25699 20768 25757 20769
rect 25699 20728 25708 20768
rect 25748 20728 25757 20768
rect 25699 20727 25757 20728
rect 26083 20768 26141 20769
rect 26083 20728 26092 20768
rect 26132 20728 26141 20768
rect 26083 20727 26141 20728
rect 26467 20768 26525 20769
rect 26467 20728 26476 20768
rect 26516 20728 26525 20768
rect 26467 20727 26525 20728
rect 27427 20768 27485 20769
rect 27427 20728 27436 20768
rect 27476 20728 27485 20768
rect 27427 20727 27485 20728
rect 31651 20768 31709 20769
rect 31651 20728 31660 20768
rect 31700 20728 31709 20768
rect 31651 20727 31709 20728
rect 32323 20768 32381 20769
rect 32323 20728 32332 20768
rect 32372 20728 32381 20768
rect 32323 20727 32381 20728
rect 32715 20768 32757 20777
rect 32715 20728 32716 20768
rect 32756 20728 32757 20768
rect 32715 20719 32757 20728
rect 35595 20768 35637 20777
rect 35595 20728 35596 20768
rect 35636 20728 35637 20768
rect 35595 20719 35637 20728
rect 35971 20768 36029 20769
rect 35971 20728 35980 20768
rect 36020 20728 36029 20768
rect 35971 20727 36029 20728
rect 36835 20768 36893 20769
rect 36835 20728 36844 20768
rect 36884 20728 36893 20768
rect 38379 20742 38380 20782
rect 38420 20742 38421 20782
rect 38379 20733 38421 20742
rect 38851 20768 38909 20769
rect 36835 20727 36893 20728
rect 38851 20728 38860 20768
rect 38900 20728 38909 20768
rect 38851 20727 38909 20728
rect 39435 20768 39477 20777
rect 39435 20728 39436 20768
rect 39476 20728 39477 20768
rect 39435 20719 39477 20728
rect 39819 20768 39861 20777
rect 39819 20728 39820 20768
rect 39860 20728 39861 20768
rect 39819 20719 39861 20728
rect 39915 20768 39957 20777
rect 39915 20728 39916 20768
rect 39956 20728 39957 20768
rect 39915 20719 39957 20728
rect 40491 20768 40533 20777
rect 40491 20728 40492 20768
rect 40532 20728 40533 20768
rect 40491 20719 40533 20728
rect 40867 20768 40925 20769
rect 40867 20728 40876 20768
rect 40916 20728 40925 20768
rect 40867 20727 40925 20728
rect 41731 20768 41789 20769
rect 41731 20728 41740 20768
rect 41780 20728 41789 20768
rect 41731 20727 41789 20728
rect 43075 20768 43133 20769
rect 43075 20728 43084 20768
rect 43124 20728 43133 20768
rect 43075 20727 43133 20728
rect 44035 20768 44093 20769
rect 44035 20728 44044 20768
rect 44084 20728 44093 20768
rect 44035 20727 44093 20728
rect 44899 20768 44957 20769
rect 44899 20728 44908 20768
rect 44948 20728 44957 20768
rect 44899 20727 44957 20728
rect 45379 20768 45437 20769
rect 45379 20728 45388 20768
rect 45428 20728 45437 20768
rect 45379 20727 45437 20728
rect 46339 20768 46397 20769
rect 46339 20728 46348 20768
rect 46388 20728 46397 20768
rect 46339 20727 46397 20728
rect 46531 20768 46589 20769
rect 46531 20728 46540 20768
rect 46580 20728 46589 20768
rect 46531 20727 46589 20728
rect 49027 20768 49085 20769
rect 49027 20728 49036 20768
rect 49076 20728 49085 20768
rect 49027 20727 49085 20728
rect 49891 20768 49949 20769
rect 49891 20728 49900 20768
rect 49940 20728 49949 20768
rect 49891 20727 49949 20728
rect 50283 20768 50325 20777
rect 50283 20728 50284 20768
rect 50324 20728 50325 20768
rect 50283 20719 50325 20728
rect 9003 20684 9045 20693
rect 9003 20644 9004 20684
rect 9044 20644 9045 20684
rect 9003 20635 9045 20644
rect 11499 20684 11541 20693
rect 11499 20644 11500 20684
rect 11540 20644 11541 20684
rect 11499 20635 11541 20644
rect 11691 20684 11733 20693
rect 11691 20644 11692 20684
rect 11732 20644 11733 20684
rect 11691 20635 11733 20644
rect 26179 20684 26237 20685
rect 26179 20644 26188 20684
rect 26228 20644 26237 20684
rect 26179 20643 26237 20644
rect 643 20600 701 20601
rect 643 20560 652 20600
rect 692 20560 701 20600
rect 643 20559 701 20560
rect 5643 20600 5685 20609
rect 5643 20560 5644 20600
rect 5684 20560 5685 20600
rect 5643 20551 5685 20560
rect 6027 20600 6069 20609
rect 6027 20560 6028 20600
rect 6068 20560 6069 20600
rect 6027 20551 6069 20560
rect 9283 20600 9341 20601
rect 9283 20560 9292 20600
rect 9332 20560 9341 20600
rect 9283 20559 9341 20560
rect 20811 20600 20853 20609
rect 20811 20560 20812 20600
rect 20852 20560 20853 20600
rect 20811 20551 20853 20560
rect 21475 20600 21533 20601
rect 21475 20560 21484 20600
rect 21524 20560 21533 20600
rect 21475 20559 21533 20560
rect 22147 20600 22205 20601
rect 22147 20560 22156 20600
rect 22196 20560 22205 20600
rect 22147 20559 22205 20560
rect 23971 20600 24029 20601
rect 23971 20560 23980 20600
rect 24020 20560 24029 20600
rect 23971 20559 24029 20560
rect 37987 20600 38045 20601
rect 37987 20560 37996 20600
rect 38036 20560 38045 20600
rect 37987 20559 38045 20560
rect 38187 20600 38229 20609
rect 38187 20560 38188 20600
rect 38228 20560 38229 20600
rect 38187 20551 38229 20560
rect 43747 20600 43805 20601
rect 43747 20560 43756 20600
rect 43796 20560 43805 20600
rect 43747 20559 43805 20560
rect 43947 20600 43989 20609
rect 43947 20560 43948 20600
rect 43988 20560 43989 20600
rect 43947 20551 43989 20560
rect 47203 20600 47261 20601
rect 47203 20560 47212 20600
rect 47252 20560 47261 20600
rect 47203 20559 47261 20560
rect 47875 20600 47933 20601
rect 47875 20560 47884 20600
rect 47924 20560 47933 20600
rect 47875 20559 47933 20560
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 643 20264 701 20265
rect 643 20224 652 20264
rect 692 20224 701 20264
rect 643 20223 701 20224
rect 4099 20264 4157 20265
rect 4099 20224 4108 20264
rect 4148 20224 4157 20264
rect 4099 20223 4157 20224
rect 8035 20264 8093 20265
rect 8035 20224 8044 20264
rect 8084 20224 8093 20264
rect 8035 20223 8093 20224
rect 14083 20264 14141 20265
rect 14083 20224 14092 20264
rect 14132 20224 14141 20264
rect 14083 20223 14141 20224
rect 18987 20264 19029 20273
rect 18987 20224 18988 20264
rect 19028 20224 19029 20264
rect 18987 20215 19029 20224
rect 25027 20264 25085 20265
rect 25027 20224 25036 20264
rect 25076 20224 25085 20264
rect 25027 20223 25085 20224
rect 29059 20264 29117 20265
rect 29059 20224 29068 20264
rect 29108 20224 29117 20264
rect 29059 20223 29117 20224
rect 41923 20264 41981 20265
rect 41923 20224 41932 20264
rect 41972 20224 41981 20264
rect 41923 20223 41981 20224
rect 45187 20264 45245 20265
rect 45187 20224 45196 20264
rect 45236 20224 45245 20264
rect 45187 20223 45245 20224
rect 8811 20180 8853 20189
rect 8811 20140 8812 20180
rect 8852 20140 8853 20180
rect 8811 20131 8853 20140
rect 24459 20180 24501 20189
rect 24459 20140 24460 20180
rect 24500 20140 24501 20180
rect 24459 20131 24501 20140
rect 24739 20180 24797 20181
rect 24739 20140 24748 20180
rect 24788 20140 24797 20180
rect 24739 20139 24797 20140
rect 25507 20180 25565 20181
rect 25507 20140 25516 20180
rect 25556 20140 25565 20180
rect 25507 20139 25565 20140
rect 27811 20180 27869 20181
rect 27811 20140 27820 20180
rect 27860 20140 27869 20180
rect 27811 20139 27869 20140
rect 37803 20180 37845 20189
rect 37803 20140 37804 20180
rect 37844 20140 37845 20180
rect 37803 20131 37845 20140
rect 38379 20180 38421 20189
rect 38379 20140 38380 20180
rect 38420 20140 38421 20180
rect 38379 20131 38421 20140
rect 39243 20180 39285 20189
rect 39243 20140 39244 20180
rect 39284 20140 39285 20180
rect 39243 20131 39285 20140
rect 44619 20180 44661 20189
rect 44619 20140 44620 20180
rect 44660 20140 44661 20180
rect 44619 20131 44661 20140
rect 47595 20180 47637 20189
rect 47595 20140 47596 20180
rect 47636 20140 47637 20180
rect 47595 20131 47637 20140
rect 23875 20117 23933 20118
rect 4003 20096 4061 20097
rect 4003 20056 4012 20096
rect 4052 20056 4061 20096
rect 4003 20055 4061 20056
rect 4875 20096 4917 20105
rect 4875 20056 4876 20096
rect 4916 20056 4917 20096
rect 4875 20047 4917 20056
rect 5067 20096 5109 20105
rect 5067 20056 5068 20096
rect 5108 20056 5109 20096
rect 5067 20047 5109 20056
rect 5643 20096 5685 20105
rect 5643 20056 5644 20096
rect 5684 20056 5685 20096
rect 5643 20047 5685 20056
rect 6019 20096 6077 20097
rect 6019 20056 6028 20096
rect 6068 20056 6077 20096
rect 6019 20055 6077 20056
rect 6883 20096 6941 20097
rect 6883 20056 6892 20096
rect 6932 20056 6941 20096
rect 6883 20055 6941 20056
rect 8515 20096 8573 20097
rect 8515 20056 8524 20096
rect 8564 20056 8573 20096
rect 8515 20055 8573 20056
rect 9187 20096 9245 20097
rect 9187 20056 9196 20096
rect 9236 20056 9245 20096
rect 9187 20055 9245 20056
rect 10051 20096 10109 20097
rect 10051 20056 10060 20096
rect 10100 20056 10109 20096
rect 10051 20055 10109 20056
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 11403 20047 11445 20056
rect 11595 20096 11637 20105
rect 11595 20056 11596 20096
rect 11636 20056 11637 20096
rect 11595 20047 11637 20056
rect 11683 20096 11741 20097
rect 11683 20056 11692 20096
rect 11732 20056 11741 20096
rect 11683 20055 11741 20056
rect 12547 20096 12605 20097
rect 12547 20056 12556 20096
rect 12596 20056 12605 20096
rect 12547 20055 12605 20056
rect 13123 20096 13181 20097
rect 13123 20056 13132 20096
rect 13172 20056 13181 20096
rect 13123 20055 13181 20056
rect 13411 20096 13469 20097
rect 13411 20056 13420 20096
rect 13460 20056 13469 20096
rect 13411 20055 13469 20056
rect 14275 20096 14333 20097
rect 14275 20056 14284 20096
rect 14324 20056 14333 20096
rect 14275 20055 14333 20056
rect 15235 20096 15293 20097
rect 15235 20056 15244 20096
rect 15284 20056 15293 20096
rect 15235 20055 15293 20056
rect 15619 20096 15677 20097
rect 15619 20056 15628 20096
rect 15668 20056 15677 20096
rect 15619 20055 15677 20056
rect 17155 20096 17213 20097
rect 17155 20056 17164 20096
rect 17204 20056 17213 20096
rect 17155 20055 17213 20056
rect 17259 20096 17301 20105
rect 17259 20056 17260 20096
rect 17300 20056 17301 20096
rect 17259 20047 17301 20056
rect 17451 20096 17493 20105
rect 17451 20056 17452 20096
rect 17492 20056 17493 20096
rect 17451 20047 17493 20056
rect 18307 20096 18365 20097
rect 18307 20056 18316 20096
rect 18356 20056 18365 20096
rect 18307 20055 18365 20056
rect 19171 20096 19229 20097
rect 19171 20056 19180 20096
rect 19220 20056 19229 20096
rect 19171 20055 19229 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 20323 20096 20381 20097
rect 20323 20056 20332 20096
rect 20372 20056 20381 20096
rect 20323 20055 20381 20056
rect 21187 20096 21245 20097
rect 21187 20056 21196 20096
rect 21236 20056 21245 20096
rect 21187 20055 21245 20056
rect 21283 20096 21341 20097
rect 21283 20056 21292 20096
rect 21332 20056 21341 20096
rect 21283 20055 21341 20056
rect 21763 20096 21821 20097
rect 21763 20056 21772 20096
rect 21812 20056 21821 20096
rect 21763 20055 21821 20056
rect 21963 20096 22005 20105
rect 21963 20056 21964 20096
rect 22004 20056 22005 20096
rect 21963 20047 22005 20056
rect 22051 20096 22109 20097
rect 22051 20056 22060 20096
rect 22100 20056 22109 20096
rect 22051 20055 22109 20056
rect 22539 20096 22581 20105
rect 22539 20056 22540 20096
rect 22580 20056 22581 20096
rect 22539 20047 22581 20056
rect 22627 20096 22685 20097
rect 22627 20056 22636 20096
rect 22676 20056 22685 20096
rect 22627 20055 22685 20056
rect 23307 20096 23349 20105
rect 23307 20056 23308 20096
rect 23348 20056 23349 20096
rect 23307 20047 23349 20056
rect 23395 20096 23453 20097
rect 23395 20056 23404 20096
rect 23444 20056 23453 20096
rect 23875 20077 23884 20117
rect 23924 20077 23933 20117
rect 23875 20076 23933 20077
rect 24075 20096 24117 20105
rect 23395 20055 23453 20056
rect 24075 20056 24076 20096
rect 24116 20056 24117 20096
rect 24075 20047 24117 20056
rect 24259 20096 24317 20097
rect 24259 20056 24268 20096
rect 24308 20056 24317 20096
rect 24259 20055 24317 20056
rect 24363 20096 24405 20105
rect 24363 20056 24364 20096
rect 24404 20056 24405 20096
rect 24363 20047 24405 20056
rect 24555 20096 24597 20105
rect 24555 20056 24556 20096
rect 24596 20056 24597 20096
rect 24555 20047 24597 20056
rect 24939 20096 24981 20105
rect 24939 20056 24940 20096
rect 24980 20056 24981 20096
rect 24939 20047 24981 20056
rect 25035 20096 25077 20105
rect 25035 20056 25036 20096
rect 25076 20056 25077 20096
rect 25035 20047 25077 20056
rect 25603 20096 25661 20097
rect 25603 20056 25612 20096
rect 25652 20056 25661 20096
rect 25603 20055 25661 20056
rect 25987 20096 26045 20097
rect 25987 20056 25996 20096
rect 26036 20056 26045 20096
rect 25987 20055 26045 20056
rect 26563 20096 26621 20097
rect 26563 20056 26572 20096
rect 26612 20056 26621 20096
rect 26563 20055 26621 20056
rect 27523 20096 27581 20097
rect 27523 20056 27532 20096
rect 27572 20056 27581 20096
rect 27523 20055 27581 20056
rect 28587 20096 28629 20105
rect 28587 20056 28588 20096
rect 28628 20056 28629 20096
rect 28587 20047 28629 20056
rect 29155 20096 29213 20097
rect 29155 20056 29164 20096
rect 29204 20056 29213 20096
rect 29155 20055 29213 20056
rect 29547 20096 29589 20105
rect 29547 20056 29548 20096
rect 29588 20056 29589 20096
rect 29547 20047 29589 20056
rect 29923 20096 29981 20097
rect 29923 20056 29932 20096
rect 29972 20056 29981 20096
rect 29923 20055 29981 20056
rect 30787 20096 30845 20097
rect 30787 20056 30796 20096
rect 30836 20056 30845 20096
rect 30787 20055 30845 20056
rect 32035 20096 32093 20097
rect 32035 20056 32044 20096
rect 32084 20056 32093 20096
rect 32035 20055 32093 20056
rect 36643 20096 36701 20097
rect 36643 20056 36652 20096
rect 36692 20056 36701 20096
rect 36643 20055 36701 20056
rect 37507 20096 37565 20097
rect 37507 20056 37516 20096
rect 37556 20056 37565 20096
rect 37507 20055 37565 20056
rect 37899 20096 37941 20105
rect 37899 20056 37900 20096
rect 37940 20056 37941 20096
rect 37899 20047 37941 20056
rect 37995 20096 38037 20105
rect 37995 20056 37996 20096
rect 38036 20056 38037 20096
rect 37995 20047 38037 20056
rect 38091 20096 38133 20105
rect 38091 20056 38092 20096
rect 38132 20056 38133 20096
rect 38091 20047 38133 20056
rect 38283 20096 38325 20105
rect 38283 20056 38284 20096
rect 38324 20056 38325 20096
rect 38283 20047 38325 20056
rect 38475 20096 38517 20105
rect 38475 20056 38476 20096
rect 38516 20056 38517 20096
rect 38475 20047 38517 20056
rect 38563 20096 38621 20097
rect 38563 20056 38572 20096
rect 38612 20056 38621 20096
rect 38563 20055 38621 20056
rect 38763 20096 38805 20105
rect 38763 20056 38764 20096
rect 38804 20056 38805 20096
rect 38763 20047 38805 20056
rect 38947 20096 39005 20097
rect 38947 20056 38956 20096
rect 38996 20056 39005 20096
rect 38947 20055 39005 20056
rect 39331 20096 39389 20097
rect 39331 20056 39340 20096
rect 39380 20056 39389 20096
rect 39331 20055 39389 20056
rect 39619 20096 39677 20097
rect 39619 20056 39628 20096
rect 39668 20056 39677 20096
rect 39619 20055 39677 20056
rect 40387 20096 40445 20097
rect 40387 20056 40396 20096
rect 40436 20056 40445 20096
rect 40387 20055 40445 20056
rect 41259 20096 41301 20105
rect 41259 20056 41260 20096
rect 41300 20056 41301 20096
rect 41259 20047 41301 20056
rect 41731 20096 41789 20097
rect 41731 20056 41740 20096
rect 41780 20056 41789 20096
rect 41731 20055 41789 20056
rect 41835 20096 41877 20105
rect 41835 20056 41836 20096
rect 41876 20056 41877 20096
rect 41835 20047 41877 20056
rect 42027 20096 42069 20105
rect 42027 20056 42028 20096
rect 42068 20056 42069 20096
rect 42027 20047 42069 20056
rect 43363 20096 43421 20097
rect 43363 20056 43372 20096
rect 43412 20056 43421 20096
rect 43363 20055 43421 20056
rect 44227 20096 44285 20097
rect 44227 20056 44236 20096
rect 44276 20056 44285 20096
rect 44227 20055 44285 20056
rect 46339 20096 46397 20097
rect 46339 20056 46348 20096
rect 46388 20056 46397 20096
rect 46339 20055 46397 20056
rect 47203 20096 47261 20097
rect 47203 20056 47212 20096
rect 47252 20056 47261 20096
rect 47203 20055 47261 20056
rect 11211 20012 11253 20021
rect 11211 19972 11212 20012
rect 11252 19972 11253 20012
rect 11211 19963 11253 19972
rect 13227 20012 13269 20021
rect 13227 19972 13228 20012
rect 13268 19972 13269 20012
rect 13227 19963 13269 19972
rect 18787 20012 18845 20013
rect 18787 19972 18796 20012
rect 18836 19972 18845 20012
rect 18787 19971 18845 19972
rect 19659 20012 19701 20021
rect 19659 19972 19660 20012
rect 19700 19972 19701 20012
rect 19659 19963 19701 19972
rect 20995 20012 21053 20013
rect 20995 19972 21004 20012
rect 21044 19972 21053 20012
rect 20995 19971 21053 19972
rect 22915 20012 22973 20013
rect 22915 19972 22924 20012
rect 22964 19972 22973 20012
rect 22915 19971 22973 19972
rect 23683 20012 23741 20013
rect 23683 19972 23692 20012
rect 23732 19972 23741 20012
rect 23683 19971 23741 19972
rect 36555 20012 36597 20021
rect 36555 19972 36556 20012
rect 36596 19972 36597 20012
rect 36555 19963 36597 19972
rect 38859 20012 38901 20021
rect 38859 19972 38860 20012
rect 38900 19972 38901 20012
rect 38859 19963 38901 19972
rect 42219 20012 42261 20021
rect 42219 19972 42220 20012
rect 42260 19972 42261 20012
rect 42219 19963 42261 19972
rect 2379 19928 2421 19937
rect 2379 19888 2380 19928
rect 2420 19888 2421 19928
rect 2379 19879 2421 19888
rect 5451 19928 5493 19937
rect 5451 19888 5452 19928
rect 5492 19888 5493 19928
rect 5451 19879 5493 19888
rect 12747 19928 12789 19937
rect 12747 19888 12748 19928
rect 12788 19888 12789 19928
rect 12747 19879 12789 19888
rect 16971 19928 17013 19937
rect 16971 19888 16972 19928
rect 17012 19888 17013 19928
rect 16971 19879 17013 19888
rect 33003 19928 33045 19937
rect 33003 19888 33004 19928
rect 33044 19888 33045 19928
rect 33003 19879 33045 19888
rect 33771 19928 33813 19937
rect 33771 19888 33772 19928
rect 33812 19888 33813 19928
rect 33771 19879 33813 19888
rect 36075 19928 36117 19937
rect 36075 19888 36076 19928
rect 36116 19888 36117 19928
rect 36075 19879 36117 19888
rect 3811 19844 3869 19845
rect 3811 19804 3820 19844
rect 3860 19804 3869 19844
rect 3811 19803 3869 19804
rect 4875 19844 4917 19853
rect 4875 19804 4876 19844
rect 4916 19804 4917 19844
rect 4875 19795 4917 19804
rect 8427 19844 8469 19853
rect 8427 19804 8428 19844
rect 8468 19804 8469 19844
rect 8427 19795 8469 19804
rect 11403 19844 11445 19853
rect 11403 19804 11404 19844
rect 11444 19804 11445 19844
rect 11403 19795 11445 19804
rect 11875 19844 11933 19845
rect 11875 19804 11884 19844
rect 11924 19804 11933 19844
rect 11875 19803 11933 19804
rect 16299 19844 16341 19853
rect 16299 19804 16300 19844
rect 16340 19804 16341 19844
rect 16299 19795 16341 19804
rect 17451 19844 17493 19853
rect 17451 19804 17452 19844
rect 17492 19804 17493 19844
rect 17451 19795 17493 19804
rect 17635 19844 17693 19845
rect 17635 19804 17644 19844
rect 17684 19804 17693 19844
rect 17635 19803 17693 19804
rect 19467 19844 19509 19853
rect 19467 19804 19468 19844
rect 19508 19804 19509 19844
rect 19467 19795 19509 19804
rect 21771 19844 21813 19853
rect 21771 19804 21772 19844
rect 21812 19804 21813 19844
rect 21771 19795 21813 19804
rect 23979 19844 24021 19853
rect 23979 19804 23980 19844
rect 24020 19804 24021 19844
rect 23979 19795 24021 19804
rect 26859 19844 26901 19853
rect 26859 19804 26860 19844
rect 26900 19804 26901 19844
rect 26859 19795 26901 19804
rect 28203 19844 28245 19853
rect 28203 19804 28204 19844
rect 28244 19804 28245 19844
rect 28203 19795 28245 19804
rect 29347 19844 29405 19845
rect 29347 19804 29356 19844
rect 29396 19804 29405 19844
rect 29347 19803 29405 19804
rect 36835 19844 36893 19845
rect 36835 19804 36844 19844
rect 36884 19804 36893 19844
rect 36835 19803 36893 19804
rect 39531 19844 39573 19853
rect 39531 19804 39532 19844
rect 39572 19804 39573 19844
rect 39531 19795 39573 19804
rect 40683 19844 40725 19853
rect 40683 19804 40684 19844
rect 40724 19804 40725 19844
rect 40683 19795 40725 19804
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 6507 19508 6549 19517
rect 6507 19468 6508 19508
rect 6548 19468 6549 19508
rect 6507 19459 6549 19468
rect 14275 19508 14333 19509
rect 14275 19468 14284 19508
rect 14324 19468 14333 19508
rect 14275 19467 14333 19468
rect 20907 19508 20949 19517
rect 20907 19468 20908 19508
rect 20948 19468 20949 19508
rect 20907 19459 20949 19468
rect 25707 19508 25749 19517
rect 25707 19468 25708 19508
rect 25748 19468 25749 19508
rect 25707 19459 25749 19468
rect 27147 19508 27189 19517
rect 27147 19468 27148 19508
rect 27188 19468 27189 19508
rect 27147 19459 27189 19468
rect 30315 19508 30357 19517
rect 30315 19468 30316 19508
rect 30356 19468 30357 19508
rect 30315 19459 30357 19468
rect 38187 19508 38229 19517
rect 38187 19468 38188 19508
rect 38228 19468 38229 19508
rect 38187 19459 38229 19468
rect 43171 19508 43229 19509
rect 43171 19468 43180 19508
rect 43220 19468 43229 19508
rect 43171 19467 43229 19468
rect 8523 19424 8565 19433
rect 8523 19384 8524 19424
rect 8564 19384 8565 19424
rect 8523 19375 8565 19384
rect 9291 19424 9333 19433
rect 9291 19384 9292 19424
rect 9332 19384 9333 19424
rect 9291 19375 9333 19384
rect 21483 19424 21525 19433
rect 21483 19384 21484 19424
rect 21524 19384 21525 19424
rect 21483 19375 21525 19384
rect 32331 19424 32373 19433
rect 32331 19384 32332 19424
rect 32372 19384 32373 19424
rect 32331 19375 32373 19384
rect 35211 19424 35253 19433
rect 35211 19384 35212 19424
rect 35252 19384 35253 19424
rect 35211 19375 35253 19384
rect 39147 19424 39189 19433
rect 39147 19384 39148 19424
rect 39188 19384 39189 19424
rect 39147 19375 39189 19384
rect 42891 19424 42933 19433
rect 42891 19384 42892 19424
rect 42932 19384 42933 19424
rect 42891 19375 42933 19384
rect 45099 19424 45141 19433
rect 45099 19384 45100 19424
rect 45140 19384 45141 19424
rect 45099 19375 45141 19384
rect 4299 19340 4341 19349
rect 4299 19300 4300 19340
rect 4340 19300 4341 19340
rect 4299 19291 4341 19300
rect 8707 19340 8765 19341
rect 8707 19300 8716 19340
rect 8756 19300 8765 19340
rect 8707 19299 8765 19300
rect 2275 19256 2333 19257
rect 2275 19216 2284 19256
rect 2324 19216 2333 19256
rect 2275 19215 2333 19216
rect 3139 19256 3197 19257
rect 3139 19216 3148 19256
rect 3188 19216 3197 19256
rect 3139 19215 3197 19216
rect 4675 19256 4733 19257
rect 4675 19216 4684 19256
rect 4724 19216 4733 19256
rect 4675 19215 4733 19216
rect 5547 19256 5589 19265
rect 5547 19216 5548 19256
rect 5588 19216 5589 19256
rect 5547 19207 5589 19216
rect 5739 19256 5781 19265
rect 5739 19216 5740 19256
rect 5780 19216 5781 19256
rect 5739 19207 5781 19216
rect 5827 19256 5885 19257
rect 5827 19216 5836 19256
rect 5876 19216 5885 19256
rect 5827 19215 5885 19216
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6219 19256 6261 19265
rect 6219 19216 6220 19256
rect 6260 19216 6261 19256
rect 6219 19207 6261 19216
rect 6315 19256 6357 19265
rect 6315 19216 6316 19256
rect 6356 19216 6357 19256
rect 6315 19207 6357 19216
rect 6507 19256 6549 19265
rect 6507 19216 6508 19256
rect 6548 19216 6549 19256
rect 6507 19207 6549 19216
rect 6699 19256 6741 19265
rect 6699 19216 6700 19256
rect 6740 19216 6741 19256
rect 6699 19207 6741 19216
rect 6787 19256 6845 19257
rect 6787 19216 6796 19256
rect 6836 19216 6845 19256
rect 6787 19215 6845 19216
rect 6979 19256 7037 19257
rect 6979 19216 6988 19256
rect 7028 19216 7037 19256
rect 6979 19215 7037 19216
rect 7179 19256 7221 19265
rect 7179 19216 7180 19256
rect 7220 19216 7221 19256
rect 7179 19207 7221 19216
rect 7851 19256 7893 19265
rect 7851 19216 7852 19256
rect 7892 19216 7893 19256
rect 7851 19207 7893 19216
rect 8043 19256 8085 19265
rect 8043 19216 8044 19256
rect 8084 19216 8085 19256
rect 8043 19207 8085 19216
rect 10627 19256 10685 19257
rect 10627 19216 10636 19256
rect 10676 19216 10685 19256
rect 10627 19215 10685 19216
rect 11019 19256 11061 19265
rect 11019 19216 11020 19256
rect 11060 19216 11061 19256
rect 11019 19207 11061 19216
rect 11115 19256 11157 19265
rect 11115 19216 11116 19256
rect 11156 19216 11157 19256
rect 11115 19207 11157 19216
rect 11211 19256 11253 19265
rect 11211 19216 11212 19256
rect 11252 19216 11253 19256
rect 11211 19207 11253 19216
rect 11307 19256 11349 19265
rect 11307 19216 11308 19256
rect 11348 19216 11349 19256
rect 11307 19207 11349 19216
rect 11883 19256 11925 19265
rect 11883 19216 11884 19256
rect 11924 19216 11925 19256
rect 11883 19207 11925 19216
rect 12259 19256 12317 19257
rect 12259 19216 12268 19256
rect 12308 19216 12317 19256
rect 12259 19215 12317 19216
rect 13123 19256 13181 19257
rect 13123 19216 13132 19256
rect 13172 19216 13181 19256
rect 13123 19215 13181 19216
rect 14859 19256 14901 19265
rect 14859 19216 14860 19256
rect 14900 19216 14901 19256
rect 14859 19207 14901 19216
rect 16099 19256 16157 19257
rect 16099 19216 16108 19256
rect 16148 19216 16157 19256
rect 16099 19215 16157 19216
rect 17347 19256 17405 19257
rect 17347 19216 17356 19256
rect 17396 19216 17405 19256
rect 17347 19215 17405 19216
rect 18211 19256 18269 19257
rect 18211 19216 18220 19256
rect 18260 19216 18269 19256
rect 18211 19215 18269 19216
rect 19651 19256 19709 19257
rect 19651 19216 19660 19256
rect 19700 19216 19709 19256
rect 19651 19215 19709 19216
rect 20803 19256 20861 19257
rect 20803 19216 20812 19256
rect 20852 19216 20861 19256
rect 20803 19215 20861 19216
rect 21003 19256 21045 19265
rect 21003 19216 21004 19256
rect 21044 19216 21045 19256
rect 21003 19207 21045 19216
rect 22147 19256 22205 19257
rect 22147 19216 22156 19256
rect 22196 19216 22205 19256
rect 22147 19215 22205 19216
rect 22435 19256 22493 19257
rect 22435 19216 22444 19256
rect 22484 19216 22493 19256
rect 22435 19215 22493 19216
rect 22635 19256 22677 19265
rect 22635 19216 22636 19256
rect 22676 19216 22677 19256
rect 22635 19207 22677 19216
rect 22723 19256 22781 19257
rect 22723 19216 22732 19256
rect 22772 19216 22781 19256
rect 22723 19215 22781 19216
rect 23211 19256 23253 19265
rect 23211 19216 23212 19256
rect 23252 19216 23253 19256
rect 23211 19207 23253 19216
rect 23307 19256 23349 19265
rect 23307 19216 23308 19256
rect 23348 19216 23349 19256
rect 23307 19207 23349 19216
rect 23403 19256 23445 19265
rect 23403 19216 23404 19256
rect 23444 19216 23445 19256
rect 23403 19207 23445 19216
rect 23499 19256 23541 19265
rect 23499 19216 23500 19256
rect 23540 19216 23541 19256
rect 23499 19207 23541 19216
rect 23691 19256 23733 19265
rect 23691 19216 23692 19256
rect 23732 19216 23733 19256
rect 23691 19207 23733 19216
rect 23787 19256 23829 19265
rect 23787 19216 23788 19256
rect 23828 19216 23829 19256
rect 23787 19207 23829 19216
rect 23883 19256 23925 19265
rect 23883 19216 23884 19256
rect 23924 19216 23925 19256
rect 23883 19207 23925 19216
rect 23979 19256 24021 19265
rect 23979 19216 23980 19256
rect 24020 19216 24021 19256
rect 23979 19207 24021 19216
rect 25227 19256 25269 19265
rect 25227 19216 25228 19256
rect 25268 19216 25269 19256
rect 25227 19207 25269 19216
rect 25323 19256 25365 19265
rect 25323 19216 25324 19256
rect 25364 19216 25365 19256
rect 25323 19207 25365 19216
rect 25419 19256 25461 19265
rect 25419 19216 25420 19256
rect 25460 19216 25461 19256
rect 25419 19207 25461 19216
rect 25707 19256 25749 19265
rect 25707 19216 25708 19256
rect 25748 19216 25749 19256
rect 25707 19207 25749 19216
rect 25899 19256 25941 19265
rect 25899 19216 25900 19256
rect 25940 19216 25941 19256
rect 25899 19207 25941 19216
rect 25987 19256 26045 19257
rect 25987 19216 25996 19256
rect 26036 19216 26045 19256
rect 25987 19215 26045 19216
rect 26955 19256 26997 19265
rect 26955 19216 26956 19256
rect 26996 19216 26997 19256
rect 26955 19207 26997 19216
rect 28291 19256 28349 19257
rect 28291 19216 28300 19256
rect 28340 19216 28349 19256
rect 28291 19215 28349 19216
rect 28579 19256 28637 19257
rect 28579 19216 28588 19256
rect 28628 19216 28637 19256
rect 28579 19215 28637 19216
rect 28771 19256 28829 19257
rect 28771 19216 28780 19256
rect 28820 19216 28829 19256
rect 28771 19215 28829 19216
rect 29155 19256 29213 19257
rect 29155 19216 29164 19256
rect 29204 19216 29213 19256
rect 29155 19215 29213 19216
rect 29739 19256 29781 19265
rect 29739 19216 29740 19256
rect 29780 19216 29781 19256
rect 29739 19207 29781 19216
rect 29827 19256 29885 19257
rect 29827 19216 29836 19256
rect 29876 19216 29885 19256
rect 29827 19215 29885 19216
rect 30315 19256 30357 19265
rect 30315 19216 30316 19256
rect 30356 19216 30357 19256
rect 30315 19207 30357 19216
rect 30507 19256 30549 19265
rect 30507 19216 30508 19256
rect 30548 19216 30549 19256
rect 30507 19207 30549 19216
rect 32139 19256 32181 19265
rect 32139 19216 32140 19256
rect 32180 19216 32181 19256
rect 32139 19207 32181 19216
rect 32331 19256 32373 19265
rect 32331 19216 32332 19256
rect 32372 19216 32373 19256
rect 32331 19207 32373 19216
rect 32523 19256 32565 19265
rect 32523 19216 32524 19256
rect 32564 19216 32565 19256
rect 32523 19207 32565 19216
rect 32899 19256 32957 19257
rect 32899 19216 32908 19256
rect 32948 19216 32957 19256
rect 32899 19215 32957 19216
rect 33763 19256 33821 19257
rect 33763 19216 33772 19256
rect 33812 19216 33821 19256
rect 33763 19215 33821 19216
rect 34923 19256 34965 19265
rect 34923 19216 34924 19256
rect 34964 19216 34965 19256
rect 34923 19207 34965 19216
rect 35587 19256 35645 19257
rect 35587 19216 35596 19256
rect 35636 19216 35645 19256
rect 35587 19215 35645 19216
rect 36547 19256 36605 19257
rect 36547 19216 36556 19256
rect 36596 19216 36605 19256
rect 36547 19215 36605 19216
rect 36835 19256 36893 19257
rect 36835 19216 36844 19256
rect 36884 19216 36893 19256
rect 36835 19215 36893 19216
rect 37795 19256 37853 19257
rect 37795 19216 37804 19256
rect 37844 19216 37853 19256
rect 37795 19215 37853 19216
rect 38187 19256 38229 19265
rect 38187 19216 38188 19256
rect 38228 19216 38229 19256
rect 38187 19207 38229 19216
rect 38379 19256 38421 19265
rect 38379 19216 38380 19256
rect 38420 19216 38421 19256
rect 38379 19207 38421 19216
rect 38467 19256 38525 19257
rect 38467 19216 38476 19256
rect 38516 19216 38525 19256
rect 38467 19215 38525 19216
rect 38763 19256 38805 19265
rect 38763 19216 38764 19256
rect 38804 19216 38805 19256
rect 38763 19207 38805 19216
rect 38859 19256 38901 19265
rect 38859 19216 38860 19256
rect 38900 19216 38901 19256
rect 38859 19207 38901 19216
rect 38955 19256 38997 19265
rect 38955 19216 38956 19256
rect 38996 19216 38997 19256
rect 38955 19207 38997 19216
rect 39619 19256 39677 19257
rect 39619 19216 39628 19256
rect 39668 19216 39677 19256
rect 39619 19215 39677 19216
rect 39915 19256 39957 19265
rect 39915 19216 39916 19256
rect 39956 19216 39957 19256
rect 39915 19207 39957 19216
rect 40011 19256 40053 19265
rect 40011 19216 40012 19256
rect 40052 19216 40053 19256
rect 40011 19207 40053 19216
rect 40107 19256 40149 19265
rect 40107 19216 40108 19256
rect 40148 19216 40149 19256
rect 40107 19207 40149 19216
rect 41059 19256 41117 19257
rect 41059 19216 41068 19256
rect 41108 19216 41117 19256
rect 41059 19215 41117 19216
rect 42219 19256 42261 19265
rect 42219 19216 42220 19256
rect 42260 19216 42261 19256
rect 42219 19207 42261 19216
rect 42315 19256 42357 19265
rect 42315 19216 42316 19256
rect 42356 19216 42357 19256
rect 42315 19207 42357 19216
rect 42411 19256 42453 19265
rect 42411 19216 42412 19256
rect 42452 19216 42453 19256
rect 42411 19207 42453 19216
rect 42507 19256 42549 19265
rect 42507 19216 42508 19256
rect 42548 19216 42549 19256
rect 42507 19207 42549 19216
rect 43843 19256 43901 19257
rect 43843 19216 43852 19256
rect 43892 19216 43901 19256
rect 43843 19215 43901 19216
rect 44035 19256 44093 19257
rect 44035 19216 44044 19256
rect 44084 19216 44093 19256
rect 44035 19215 44093 19216
rect 1899 19172 1941 19181
rect 1899 19132 1900 19172
rect 1940 19132 1941 19172
rect 1899 19123 1941 19132
rect 7083 19172 7125 19181
rect 7083 19132 7084 19172
rect 7124 19132 7125 19172
rect 7083 19123 7125 19132
rect 16971 19172 17013 19181
rect 16971 19132 16972 19172
rect 17012 19132 17013 19172
rect 16971 19123 17013 19132
rect 20515 19172 20573 19173
rect 20515 19132 20524 19172
rect 20564 19132 20573 19172
rect 20515 19131 20573 19132
rect 40395 19172 40437 19181
rect 40395 19132 40396 19172
rect 40436 19132 40437 19172
rect 40395 19123 40437 19132
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 5347 19088 5405 19089
rect 5347 19048 5356 19088
rect 5396 19048 5405 19088
rect 5347 19047 5405 19048
rect 5635 19088 5693 19089
rect 5635 19048 5644 19088
rect 5684 19048 5693 19088
rect 5635 19047 5693 19048
rect 7947 19088 7989 19097
rect 7947 19048 7948 19088
rect 7988 19048 7989 19088
rect 7947 19039 7989 19048
rect 9955 19088 10013 19089
rect 9955 19048 9964 19088
rect 10004 19048 10013 19088
rect 9955 19047 10013 19048
rect 15243 19088 15285 19097
rect 15243 19048 15244 19088
rect 15284 19048 15285 19088
rect 15243 19039 15285 19048
rect 16771 19088 16829 19089
rect 16771 19048 16780 19088
rect 16820 19048 16829 19088
rect 16771 19047 16829 19048
rect 19363 19088 19421 19089
rect 19363 19048 19372 19088
rect 19412 19048 19421 19088
rect 19363 19047 19421 19048
rect 22443 19088 22485 19097
rect 22443 19048 22444 19088
rect 22484 19048 22485 19088
rect 22443 19039 22485 19048
rect 25507 19088 25565 19089
rect 25507 19048 25516 19088
rect 25556 19048 25565 19088
rect 25507 19047 25565 19048
rect 27339 19088 27381 19097
rect 27339 19048 27340 19088
rect 27380 19048 27381 19088
rect 27339 19039 27381 19048
rect 28107 19088 28149 19097
rect 28107 19048 28108 19088
rect 28148 19048 28149 19088
rect 28107 19039 28149 19048
rect 29259 19088 29301 19097
rect 29259 19048 29260 19088
rect 29300 19048 29301 19088
rect 29259 19039 29301 19048
rect 30123 19088 30165 19097
rect 30123 19048 30124 19088
rect 30164 19048 30165 19088
rect 30123 19039 30165 19048
rect 38659 19088 38717 19089
rect 38659 19048 38668 19088
rect 38708 19048 38717 19088
rect 38659 19047 38717 19048
rect 39723 19088 39765 19097
rect 39723 19048 39724 19088
rect 39764 19048 39765 19088
rect 39723 19039 39765 19048
rect 40195 19088 40253 19089
rect 40195 19048 40204 19088
rect 40244 19048 40253 19088
rect 40195 19047 40253 19048
rect 44707 19088 44765 19089
rect 44707 19048 44716 19088
rect 44756 19048 44765 19088
rect 44707 19047 44765 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 22627 18794 22685 18795
rect 643 18752 701 18753
rect 643 18712 652 18752
rect 692 18712 701 18752
rect 643 18711 701 18712
rect 2859 18752 2901 18761
rect 2859 18712 2860 18752
rect 2900 18712 2901 18752
rect 2859 18703 2901 18712
rect 3235 18752 3293 18753
rect 3235 18712 3244 18752
rect 3284 18712 3293 18752
rect 3235 18711 3293 18712
rect 3523 18752 3581 18753
rect 3523 18712 3532 18752
rect 3572 18712 3581 18752
rect 3523 18711 3581 18712
rect 9291 18752 9333 18761
rect 9291 18712 9292 18752
rect 9332 18712 9333 18752
rect 9291 18703 9333 18712
rect 9955 18752 10013 18753
rect 9955 18712 9964 18752
rect 10004 18712 10013 18752
rect 9955 18711 10013 18712
rect 14755 18752 14813 18753
rect 14755 18712 14764 18752
rect 14804 18712 14813 18752
rect 14755 18711 14813 18712
rect 17347 18752 17405 18753
rect 17347 18712 17356 18752
rect 17396 18712 17405 18752
rect 17347 18711 17405 18712
rect 19083 18752 19125 18761
rect 22627 18754 22636 18794
rect 22676 18754 22685 18794
rect 22627 18753 22685 18754
rect 19083 18712 19084 18752
rect 19124 18712 19125 18752
rect 19083 18703 19125 18712
rect 20899 18752 20957 18753
rect 20899 18712 20908 18752
rect 20948 18712 20957 18752
rect 20899 18711 20957 18712
rect 21379 18752 21437 18753
rect 21379 18712 21388 18752
rect 21428 18712 21437 18752
rect 21379 18711 21437 18712
rect 27907 18752 27965 18753
rect 27907 18712 27916 18752
rect 27956 18712 27965 18752
rect 27907 18711 27965 18712
rect 32899 18752 32957 18753
rect 32899 18712 32908 18752
rect 32948 18712 32957 18752
rect 32899 18711 32957 18712
rect 40483 18752 40541 18753
rect 40483 18712 40492 18752
rect 40532 18712 40541 18752
rect 40483 18711 40541 18712
rect 17163 18668 17205 18677
rect 17163 18628 17164 18668
rect 17204 18628 17205 18668
rect 17163 18619 17205 18628
rect 21091 18668 21149 18669
rect 21091 18628 21100 18668
rect 21140 18628 21149 18668
rect 21091 18627 21149 18628
rect 28195 18668 28253 18669
rect 28195 18628 28204 18668
rect 28244 18628 28253 18668
rect 28195 18627 28253 18628
rect 32139 18668 32181 18677
rect 32139 18628 32140 18668
rect 32180 18628 32181 18668
rect 32139 18619 32181 18628
rect 37899 18668 37941 18677
rect 37899 18628 37900 18668
rect 37940 18628 37941 18668
rect 37899 18619 37941 18628
rect 2763 18584 2805 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 2955 18584 2997 18593
rect 2955 18544 2956 18584
rect 2996 18544 2997 18584
rect 2955 18535 2997 18544
rect 3051 18584 3093 18593
rect 3051 18544 3052 18584
rect 3092 18544 3093 18584
rect 3051 18535 3093 18544
rect 3427 18584 3485 18585
rect 3427 18544 3436 18584
rect 3476 18544 3485 18584
rect 3427 18543 3485 18544
rect 3715 18584 3773 18585
rect 3715 18544 3724 18584
rect 3764 18544 3773 18584
rect 3715 18543 3773 18544
rect 4579 18584 4637 18585
rect 4579 18544 4588 18584
rect 4628 18544 4637 18584
rect 4579 18543 4637 18544
rect 5835 18584 5877 18593
rect 5835 18544 5836 18584
rect 5876 18544 5877 18584
rect 5835 18535 5877 18544
rect 6211 18584 6269 18585
rect 6211 18544 6220 18584
rect 6260 18544 6269 18584
rect 6211 18543 6269 18544
rect 6411 18584 6453 18593
rect 6411 18544 6412 18584
rect 6452 18544 6453 18584
rect 6411 18535 6453 18544
rect 6499 18584 6557 18585
rect 6499 18544 6508 18584
rect 6548 18544 6557 18584
rect 6499 18543 6557 18544
rect 6699 18584 6741 18593
rect 6699 18544 6700 18584
rect 6740 18544 6741 18584
rect 6699 18535 6741 18544
rect 6795 18584 6837 18593
rect 6795 18544 6796 18584
rect 6836 18544 6837 18584
rect 6795 18535 6837 18544
rect 6891 18584 6933 18593
rect 6891 18544 6892 18584
rect 6932 18544 6933 18584
rect 6891 18535 6933 18544
rect 6987 18584 7029 18593
rect 6987 18544 6988 18584
rect 7028 18544 7029 18584
rect 6987 18535 7029 18544
rect 7179 18584 7221 18593
rect 7179 18544 7180 18584
rect 7220 18544 7221 18584
rect 7179 18535 7221 18544
rect 7843 18584 7901 18585
rect 7843 18544 7852 18584
rect 7892 18544 7901 18584
rect 7843 18543 7901 18544
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 8235 18584 8277 18593
rect 8235 18544 8236 18584
rect 8276 18544 8277 18584
rect 8235 18535 8277 18544
rect 8323 18584 8381 18585
rect 8323 18544 8332 18584
rect 8372 18544 8381 18584
rect 8323 18543 8381 18544
rect 8803 18584 8861 18585
rect 8803 18544 8812 18584
rect 8852 18544 8861 18584
rect 8803 18543 8861 18544
rect 10627 18584 10685 18585
rect 10627 18544 10636 18584
rect 10676 18544 10685 18584
rect 10627 18543 10685 18544
rect 15907 18584 15965 18585
rect 15907 18544 15916 18584
rect 15956 18544 15965 18584
rect 15907 18543 15965 18544
rect 16771 18584 16829 18585
rect 16771 18544 16780 18584
rect 16820 18544 16829 18584
rect 16771 18543 16829 18544
rect 18019 18584 18077 18585
rect 18019 18544 18028 18584
rect 18068 18544 18077 18584
rect 18019 18543 18077 18544
rect 18883 18584 18941 18585
rect 18883 18544 18892 18584
rect 18932 18544 18941 18584
rect 18883 18543 18941 18544
rect 19075 18584 19133 18585
rect 19075 18544 19084 18584
rect 19124 18544 19133 18584
rect 19075 18543 19133 18544
rect 19275 18584 19317 18593
rect 19275 18544 19276 18584
rect 19316 18544 19317 18584
rect 19275 18535 19317 18544
rect 19363 18584 19421 18585
rect 19363 18544 19372 18584
rect 19412 18544 19421 18584
rect 19363 18543 19421 18544
rect 19563 18584 19605 18593
rect 19563 18544 19564 18584
rect 19604 18544 19605 18584
rect 19563 18535 19605 18544
rect 19747 18584 19805 18585
rect 19747 18544 19756 18584
rect 19796 18544 19805 18584
rect 19747 18543 19805 18544
rect 20619 18584 20661 18593
rect 20619 18544 20620 18584
rect 20660 18544 20661 18584
rect 20619 18535 20661 18544
rect 20715 18584 20757 18593
rect 20715 18544 20716 18584
rect 20756 18544 20757 18584
rect 20715 18535 20757 18544
rect 21291 18584 21333 18593
rect 21291 18544 21292 18584
rect 21332 18544 21333 18584
rect 21291 18535 21333 18544
rect 21387 18584 21429 18593
rect 21387 18544 21388 18584
rect 21428 18544 21429 18584
rect 21387 18535 21429 18544
rect 22435 18584 22493 18585
rect 22435 18544 22444 18584
rect 22484 18544 22493 18584
rect 22435 18543 22493 18544
rect 22622 18584 22664 18593
rect 22622 18544 22623 18584
rect 22663 18544 22664 18584
rect 22622 18535 22664 18544
rect 24171 18584 24213 18593
rect 24171 18544 24172 18584
rect 24212 18544 24213 18584
rect 24171 18535 24213 18544
rect 24363 18584 24405 18593
rect 24363 18544 24364 18584
rect 24404 18544 24405 18584
rect 24363 18535 24405 18544
rect 24459 18584 24501 18593
rect 24459 18544 24460 18584
rect 24500 18544 24501 18584
rect 24459 18535 24501 18544
rect 24651 18584 24693 18593
rect 24651 18544 24652 18584
rect 24692 18544 24693 18584
rect 24651 18535 24693 18544
rect 24843 18584 24885 18593
rect 24843 18544 24844 18584
rect 24884 18544 24885 18584
rect 24843 18535 24885 18544
rect 26083 18584 26141 18585
rect 26083 18544 26092 18584
rect 26132 18544 26141 18584
rect 26083 18543 26141 18544
rect 28003 18584 28061 18585
rect 28003 18544 28012 18584
rect 28052 18544 28061 18584
rect 28003 18543 28061 18544
rect 28675 18584 28733 18585
rect 28675 18544 28684 18584
rect 28724 18544 28733 18584
rect 28675 18543 28733 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 28779 18535 28821 18544
rect 29355 18584 29397 18593
rect 29355 18544 29356 18584
rect 29396 18544 29397 18584
rect 29355 18535 29397 18544
rect 29547 18584 29589 18593
rect 29547 18544 29548 18584
rect 29588 18544 29589 18584
rect 29547 18535 29589 18544
rect 29635 18584 29693 18585
rect 29635 18544 29644 18584
rect 29684 18544 29693 18584
rect 29635 18543 29693 18544
rect 29835 18584 29877 18593
rect 29835 18544 29836 18584
rect 29876 18544 29877 18584
rect 29835 18535 29877 18544
rect 30019 18584 30077 18585
rect 30019 18544 30028 18584
rect 30068 18544 30077 18584
rect 30019 18543 30077 18544
rect 30315 18584 30357 18593
rect 30315 18544 30316 18584
rect 30356 18544 30357 18584
rect 30315 18535 30357 18544
rect 30507 18584 30549 18593
rect 30507 18544 30508 18584
rect 30548 18544 30549 18584
rect 30507 18535 30549 18544
rect 32523 18584 32565 18593
rect 32523 18544 32524 18584
rect 32564 18544 32565 18584
rect 32523 18535 32565 18544
rect 33003 18584 33045 18593
rect 33003 18544 33004 18584
rect 33044 18544 33045 18584
rect 33003 18535 33045 18544
rect 33099 18584 33141 18593
rect 33099 18544 33100 18584
rect 33140 18544 33141 18584
rect 33099 18535 33141 18544
rect 33195 18584 33237 18593
rect 33195 18544 33196 18584
rect 33236 18544 33237 18584
rect 33195 18535 33237 18544
rect 33667 18584 33725 18585
rect 33667 18544 33676 18584
rect 33716 18544 33725 18584
rect 33667 18543 33725 18544
rect 34347 18584 34389 18593
rect 34347 18544 34348 18584
rect 34388 18544 34389 18584
rect 34347 18535 34389 18544
rect 34539 18584 34581 18593
rect 34539 18544 34540 18584
rect 34580 18544 34581 18584
rect 34539 18535 34581 18544
rect 34915 18584 34973 18585
rect 34915 18544 34924 18584
rect 34964 18544 34973 18584
rect 34915 18543 34973 18544
rect 35779 18584 35837 18585
rect 35779 18544 35788 18584
rect 35828 18544 35837 18584
rect 35779 18543 35837 18544
rect 37027 18584 37085 18585
rect 37027 18544 37036 18584
rect 37076 18544 37085 18584
rect 37027 18543 37085 18544
rect 38275 18584 38333 18585
rect 38275 18544 38284 18584
rect 38324 18544 38333 18584
rect 38275 18543 38333 18544
rect 39139 18584 39197 18585
rect 39139 18544 39148 18584
rect 39188 18544 39197 18584
rect 39139 18543 39197 18544
rect 41635 18584 41693 18585
rect 41635 18544 41644 18584
rect 41684 18544 41693 18584
rect 41635 18543 41693 18544
rect 42499 18584 42557 18585
rect 42499 18544 42508 18584
rect 42548 18544 42557 18584
rect 42499 18543 42557 18544
rect 42891 18584 42933 18593
rect 42891 18544 42892 18584
rect 42932 18544 42933 18584
rect 42891 18535 42933 18544
rect 44227 18584 44285 18585
rect 44227 18544 44236 18584
rect 44276 18544 44285 18584
rect 44227 18543 44285 18544
rect 45475 18584 45533 18585
rect 45475 18544 45484 18584
rect 45524 18544 45533 18584
rect 45475 18543 45533 18544
rect 46339 18584 46397 18585
rect 46339 18544 46348 18584
rect 46388 18544 46397 18584
rect 46339 18543 46397 18544
rect 46731 18584 46773 18593
rect 46731 18544 46732 18584
rect 46772 18544 46773 18584
rect 46731 18535 46773 18544
rect 5643 18500 5685 18509
rect 5643 18460 5644 18500
rect 5684 18460 5685 18500
rect 5643 18451 5685 18460
rect 24747 18500 24789 18509
rect 24747 18460 24748 18500
rect 24788 18460 24789 18500
rect 24747 18451 24789 18460
rect 27523 18500 27581 18501
rect 27523 18460 27532 18500
rect 27572 18460 27581 18500
rect 27523 18459 27581 18460
rect 37411 18500 37469 18501
rect 37411 18460 37420 18500
rect 37460 18460 37469 18500
rect 37411 18459 37469 18460
rect 1707 18416 1749 18425
rect 1707 18376 1708 18416
rect 1748 18376 1749 18416
rect 1707 18367 1749 18376
rect 6403 18416 6461 18417
rect 6403 18376 6412 18416
rect 6452 18376 6461 18416
rect 6403 18375 6461 18376
rect 10827 18416 10869 18425
rect 10827 18376 10828 18416
rect 10868 18376 10869 18416
rect 10827 18367 10869 18376
rect 12555 18416 12597 18425
rect 12555 18376 12556 18416
rect 12596 18376 12597 18416
rect 12555 18367 12597 18376
rect 24451 18416 24509 18417
rect 24451 18376 24460 18416
rect 24500 18376 24509 18416
rect 24451 18375 24509 18376
rect 27723 18416 27765 18425
rect 27723 18376 27724 18416
rect 27764 18376 27765 18416
rect 27723 18367 27765 18376
rect 4387 18332 4445 18333
rect 4387 18292 4396 18332
rect 4436 18292 4445 18332
rect 4387 18291 4445 18292
rect 5251 18332 5309 18333
rect 5251 18292 5260 18332
rect 5300 18292 5309 18332
rect 5251 18291 5309 18292
rect 5835 18332 5877 18341
rect 5835 18292 5836 18332
rect 5876 18292 5877 18332
rect 5835 18283 5877 18292
rect 8043 18332 8085 18341
rect 8043 18292 8044 18332
rect 8084 18292 8085 18332
rect 8043 18283 8085 18292
rect 9291 18332 9333 18341
rect 9291 18292 9292 18332
rect 9332 18292 9333 18332
rect 9291 18283 9333 18292
rect 18211 18332 18269 18333
rect 18211 18292 18220 18332
rect 18260 18292 18269 18332
rect 18211 18291 18269 18292
rect 19659 18332 19701 18341
rect 19659 18292 19660 18332
rect 19700 18292 19701 18332
rect 19659 18283 19701 18292
rect 25611 18332 25653 18341
rect 25611 18292 25612 18332
rect 25652 18292 25653 18332
rect 25611 18283 25653 18292
rect 28491 18332 28533 18341
rect 28491 18292 28492 18332
rect 28532 18292 28533 18332
rect 28491 18283 28533 18292
rect 29355 18332 29397 18341
rect 29355 18292 29356 18332
rect 29396 18292 29397 18332
rect 29355 18283 29397 18292
rect 29931 18332 29973 18341
rect 29931 18292 29932 18332
rect 29972 18292 29973 18332
rect 29931 18283 29973 18292
rect 30315 18332 30357 18341
rect 30315 18292 30316 18332
rect 30356 18292 30357 18332
rect 30315 18283 30357 18292
rect 40291 18332 40349 18333
rect 40291 18292 40300 18332
rect 40340 18292 40349 18332
rect 40291 18291 40349 18292
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 5443 17996 5501 17997
rect 5443 17956 5452 17996
rect 5492 17956 5501 17996
rect 5443 17955 5501 17956
rect 11107 17996 11165 17997
rect 11107 17956 11116 17996
rect 11156 17956 11165 17996
rect 11107 17955 11165 17956
rect 14475 17996 14517 18005
rect 14475 17956 14476 17996
rect 14516 17956 14517 17996
rect 14475 17947 14517 17956
rect 18987 17996 19029 18005
rect 18987 17956 18988 17996
rect 19028 17956 19029 17996
rect 18987 17947 19029 17956
rect 1035 17912 1077 17921
rect 1035 17872 1036 17912
rect 1076 17872 1077 17912
rect 1035 17863 1077 17872
rect 6603 17912 6645 17921
rect 6603 17872 6604 17912
rect 6644 17872 6645 17912
rect 6603 17863 6645 17872
rect 21091 17912 21149 17913
rect 21091 17872 21100 17912
rect 21140 17872 21149 17912
rect 21091 17871 21149 17872
rect 24843 17912 24885 17921
rect 24843 17872 24844 17912
rect 24884 17872 24885 17912
rect 24843 17863 24885 17872
rect 28011 17912 28053 17921
rect 28011 17872 28012 17912
rect 28052 17872 28053 17912
rect 28011 17863 28053 17872
rect 29355 17912 29397 17921
rect 29355 17872 29356 17912
rect 29396 17872 29397 17912
rect 29355 17863 29397 17872
rect 30027 17912 30069 17921
rect 30027 17872 30028 17912
rect 30068 17872 30069 17912
rect 30027 17863 30069 17872
rect 30987 17912 31029 17921
rect 30987 17872 30988 17912
rect 31028 17872 31029 17912
rect 30987 17863 31029 17872
rect 32427 17912 32469 17921
rect 32427 17872 32428 17912
rect 32468 17872 32469 17912
rect 32427 17863 32469 17872
rect 35979 17912 36021 17921
rect 35979 17872 35980 17912
rect 36020 17872 36021 17912
rect 35979 17863 36021 17872
rect 40491 17912 40533 17921
rect 40491 17872 40492 17912
rect 40532 17872 40533 17912
rect 40491 17863 40533 17872
rect 41739 17912 41781 17921
rect 41739 17872 41740 17912
rect 41780 17872 41781 17912
rect 41739 17863 41781 17872
rect 3627 17828 3669 17837
rect 3627 17788 3628 17828
rect 3668 17788 3669 17828
rect 3627 17779 3669 17788
rect 17163 17828 17205 17837
rect 17163 17788 17164 17828
rect 17204 17788 17205 17828
rect 17163 17779 17205 17788
rect 20811 17828 20853 17837
rect 20811 17788 20812 17828
rect 20852 17788 20853 17828
rect 20811 17779 20853 17788
rect 24747 17828 24789 17837
rect 24747 17788 24748 17828
rect 24788 17788 24789 17828
rect 24747 17779 24789 17788
rect 24939 17828 24981 17837
rect 24939 17788 24940 17828
rect 24980 17788 24981 17828
rect 24939 17779 24981 17788
rect 28963 17828 29021 17829
rect 28963 17788 28972 17828
rect 29012 17788 29021 17828
rect 28963 17787 29021 17788
rect 1603 17744 1661 17745
rect 1603 17704 1612 17744
rect 1652 17704 1661 17744
rect 1603 17703 1661 17704
rect 2467 17744 2525 17745
rect 2467 17704 2476 17744
rect 2516 17704 2525 17744
rect 2467 17703 2525 17704
rect 3907 17744 3965 17745
rect 3907 17704 3916 17744
rect 3956 17704 3965 17744
rect 3907 17703 3965 17704
rect 4771 17744 4829 17745
rect 4771 17704 4780 17744
rect 4820 17704 4829 17744
rect 4771 17703 4829 17704
rect 5835 17744 5877 17753
rect 5835 17704 5836 17744
rect 5876 17704 5877 17744
rect 5835 17695 5877 17704
rect 5931 17744 5973 17753
rect 5931 17704 5932 17744
rect 5972 17704 5973 17744
rect 5931 17695 5973 17704
rect 6027 17744 6069 17753
rect 6027 17704 6028 17744
rect 6068 17704 6069 17744
rect 6027 17695 6069 17704
rect 6123 17744 6165 17753
rect 6123 17704 6124 17744
rect 6164 17704 6165 17744
rect 6123 17695 6165 17704
rect 6507 17744 6549 17753
rect 6507 17704 6508 17744
rect 6548 17704 6549 17744
rect 6507 17695 6549 17704
rect 6699 17744 6741 17753
rect 6699 17704 6700 17744
rect 6740 17704 6741 17744
rect 6699 17695 6741 17704
rect 6795 17744 6837 17753
rect 6795 17704 6796 17744
rect 6836 17704 6837 17744
rect 6795 17695 6837 17704
rect 6987 17744 7029 17753
rect 6987 17704 6988 17744
rect 7028 17704 7029 17744
rect 6987 17695 7029 17704
rect 7363 17744 7421 17745
rect 7363 17704 7372 17744
rect 7412 17704 7421 17744
rect 7363 17703 7421 17704
rect 7843 17744 7901 17745
rect 7843 17704 7852 17744
rect 7892 17704 7901 17744
rect 7843 17703 7901 17704
rect 9091 17744 9149 17745
rect 9091 17704 9100 17744
rect 9140 17704 9149 17744
rect 9091 17703 9149 17704
rect 9955 17744 10013 17745
rect 9955 17704 9964 17744
rect 10004 17704 10013 17744
rect 9955 17703 10013 17704
rect 12075 17744 12117 17753
rect 12075 17704 12076 17744
rect 12116 17704 12117 17744
rect 12075 17695 12117 17704
rect 12451 17744 12509 17745
rect 12451 17704 12460 17744
rect 12500 17704 12509 17744
rect 12451 17703 12509 17704
rect 13315 17744 13373 17745
rect 13315 17704 13324 17744
rect 13364 17704 13373 17744
rect 13315 17703 13373 17704
rect 15139 17744 15197 17745
rect 15139 17704 15148 17744
rect 15188 17704 15197 17744
rect 15139 17703 15197 17704
rect 16003 17744 16061 17745
rect 16003 17704 16012 17744
rect 16052 17704 16061 17744
rect 16003 17703 16061 17704
rect 17355 17744 17397 17753
rect 17355 17704 17356 17744
rect 17396 17704 17397 17744
rect 17355 17695 17397 17704
rect 17451 17744 17493 17753
rect 17451 17704 17452 17744
rect 17492 17704 17493 17744
rect 17451 17695 17493 17704
rect 17547 17744 17589 17753
rect 17547 17704 17548 17744
rect 17588 17704 17589 17744
rect 17547 17695 17589 17704
rect 17643 17744 17685 17753
rect 17643 17704 17644 17744
rect 17684 17704 17685 17744
rect 17643 17695 17685 17704
rect 17827 17744 17885 17745
rect 17827 17704 17836 17744
rect 17876 17704 17885 17744
rect 17827 17703 17885 17704
rect 18507 17744 18549 17753
rect 18507 17704 18508 17744
rect 18548 17704 18549 17744
rect 18507 17695 18549 17704
rect 18691 17744 18749 17745
rect 18691 17704 18700 17744
rect 18740 17704 18749 17744
rect 18691 17703 18749 17704
rect 18795 17744 18837 17753
rect 18795 17704 18796 17744
rect 18836 17704 18837 17744
rect 18795 17695 18837 17704
rect 18979 17744 19037 17745
rect 18979 17704 18988 17744
rect 19028 17704 19037 17744
rect 18979 17703 19037 17704
rect 19171 17744 19229 17745
rect 19171 17704 19180 17744
rect 19220 17704 19229 17744
rect 19171 17703 19229 17704
rect 19275 17744 19317 17753
rect 19275 17704 19276 17744
rect 19316 17704 19317 17744
rect 19275 17695 19317 17704
rect 19467 17744 19509 17753
rect 19467 17704 19468 17744
rect 19508 17704 19509 17744
rect 19467 17695 19509 17704
rect 19747 17744 19805 17745
rect 19747 17704 19756 17744
rect 19796 17704 19805 17744
rect 19747 17703 19805 17704
rect 20619 17744 20661 17753
rect 20619 17704 20620 17744
rect 20660 17704 20661 17744
rect 20619 17695 20661 17704
rect 20715 17744 20757 17753
rect 20715 17704 20716 17744
rect 20756 17704 20757 17744
rect 20715 17695 20757 17704
rect 20907 17744 20949 17753
rect 20907 17704 20908 17744
rect 20948 17704 20949 17744
rect 20907 17695 20949 17704
rect 21291 17744 21333 17753
rect 21291 17704 21292 17744
rect 21332 17704 21333 17744
rect 21291 17695 21333 17704
rect 21387 17744 21429 17753
rect 21387 17704 21388 17744
rect 21428 17704 21429 17744
rect 21387 17695 21429 17704
rect 21483 17744 21525 17753
rect 21483 17704 21484 17744
rect 21524 17704 21525 17744
rect 21483 17695 21525 17704
rect 21579 17744 21621 17753
rect 21579 17704 21580 17744
rect 21620 17704 21621 17744
rect 21579 17695 21621 17704
rect 21955 17744 22013 17745
rect 21955 17704 21964 17744
rect 22004 17704 22013 17744
rect 21955 17703 22013 17704
rect 22819 17744 22877 17745
rect 22819 17704 22828 17744
rect 22868 17704 22877 17744
rect 22819 17703 22877 17704
rect 23779 17744 23837 17745
rect 23779 17704 23788 17744
rect 23828 17704 23837 17744
rect 23779 17703 23837 17704
rect 24259 17744 24317 17745
rect 24259 17704 24268 17744
rect 24308 17704 24317 17744
rect 24259 17703 24317 17704
rect 24651 17744 24693 17753
rect 24651 17704 24652 17744
rect 24692 17704 24693 17744
rect 24651 17695 24693 17704
rect 25027 17744 25085 17745
rect 25027 17704 25036 17744
rect 25076 17704 25085 17744
rect 25027 17703 25085 17704
rect 25411 17744 25469 17745
rect 25411 17704 25420 17744
rect 25460 17704 25469 17744
rect 25411 17703 25469 17704
rect 26371 17744 26429 17745
rect 26371 17704 26380 17744
rect 26420 17704 26429 17744
rect 26371 17703 26429 17704
rect 27523 17744 27581 17745
rect 27523 17704 27532 17744
rect 27572 17704 27581 17744
rect 27523 17703 27581 17704
rect 28011 17744 28053 17753
rect 28011 17704 28012 17744
rect 28052 17704 28053 17744
rect 28011 17695 28053 17704
rect 28675 17744 28733 17745
rect 28675 17704 28684 17744
rect 28724 17704 28733 17744
rect 28675 17703 28733 17704
rect 28771 17744 28829 17745
rect 28771 17704 28780 17744
rect 28820 17704 28829 17744
rect 28771 17703 28829 17704
rect 29355 17744 29397 17753
rect 29355 17704 29356 17744
rect 29396 17704 29397 17744
rect 29355 17695 29397 17704
rect 29731 17744 29789 17745
rect 29731 17704 29740 17744
rect 29780 17704 29789 17744
rect 29731 17703 29789 17704
rect 29835 17744 29877 17753
rect 29835 17704 29836 17744
rect 29876 17704 29877 17744
rect 29835 17695 29877 17704
rect 30019 17744 30077 17745
rect 30019 17704 30028 17744
rect 30068 17704 30077 17744
rect 30019 17703 30077 17704
rect 30507 17744 30549 17753
rect 30507 17704 30508 17744
rect 30548 17704 30549 17744
rect 30507 17695 30549 17704
rect 30699 17744 30741 17753
rect 30699 17704 30700 17744
rect 30740 17704 30741 17744
rect 30699 17695 30741 17704
rect 30787 17744 30845 17745
rect 30787 17704 30796 17744
rect 30836 17704 30845 17744
rect 30787 17703 30845 17704
rect 30987 17744 31029 17753
rect 30987 17704 30988 17744
rect 31028 17704 31029 17744
rect 30987 17695 31029 17704
rect 31179 17744 31221 17753
rect 31179 17704 31180 17744
rect 31220 17704 31221 17744
rect 31179 17695 31221 17704
rect 31851 17744 31893 17753
rect 31851 17704 31852 17744
rect 31892 17704 31893 17744
rect 31851 17695 31893 17704
rect 33099 17744 33141 17753
rect 33099 17704 33100 17744
rect 33140 17704 33141 17744
rect 33099 17695 33141 17704
rect 33195 17744 33237 17753
rect 33195 17704 33196 17744
rect 33236 17704 33237 17744
rect 33195 17695 33237 17704
rect 33291 17744 33333 17753
rect 33291 17704 33292 17744
rect 33332 17704 33333 17744
rect 33291 17695 33333 17704
rect 34243 17744 34301 17745
rect 34243 17704 34252 17744
rect 34292 17704 34301 17744
rect 34243 17703 34301 17704
rect 34435 17744 34493 17745
rect 34435 17704 34444 17744
rect 34484 17704 34493 17744
rect 34435 17703 34493 17704
rect 35307 17744 35349 17753
rect 35307 17704 35308 17744
rect 35348 17704 35349 17744
rect 35307 17695 35349 17704
rect 36835 17744 36893 17745
rect 36835 17704 36844 17744
rect 36884 17704 36893 17744
rect 36835 17703 36893 17704
rect 37707 17744 37749 17753
rect 37707 17704 37708 17744
rect 37748 17704 37749 17744
rect 37707 17695 37749 17704
rect 38859 17744 38901 17753
rect 38859 17704 38860 17744
rect 38900 17704 38901 17744
rect 38859 17695 38901 17704
rect 39523 17744 39581 17745
rect 39523 17704 39532 17744
rect 39572 17704 39581 17744
rect 39523 17703 39581 17704
rect 40195 17744 40253 17745
rect 40195 17704 40204 17744
rect 40244 17704 40253 17744
rect 40195 17703 40253 17704
rect 40299 17744 40341 17753
rect 40299 17704 40300 17744
rect 40340 17704 40341 17744
rect 40299 17695 40341 17704
rect 40491 17744 40533 17753
rect 40491 17704 40492 17744
rect 40532 17704 40533 17744
rect 40491 17695 40533 17704
rect 40675 17744 40733 17745
rect 40675 17704 40684 17744
rect 40724 17704 40733 17744
rect 40675 17703 40733 17704
rect 41355 17744 41397 17753
rect 41355 17704 41356 17744
rect 41396 17704 41397 17744
rect 41355 17695 41397 17704
rect 1227 17660 1269 17669
rect 1227 17620 1228 17660
rect 1268 17620 1269 17660
rect 1227 17611 1269 17620
rect 4587 17660 4629 17669
rect 4587 17620 4588 17660
rect 4628 17620 4629 17660
rect 4587 17611 4629 17620
rect 7467 17660 7509 17669
rect 7467 17620 7468 17660
rect 7508 17620 7509 17660
rect 7467 17611 7509 17620
rect 8523 17660 8565 17669
rect 8523 17620 8524 17660
rect 8564 17620 8565 17660
rect 8523 17611 8565 17620
rect 8715 17660 8757 17669
rect 8715 17620 8716 17660
rect 8756 17620 8757 17660
rect 8715 17611 8757 17620
rect 14763 17660 14805 17669
rect 14763 17620 14764 17660
rect 14804 17620 14805 17660
rect 14763 17611 14805 17620
rect 24451 17660 24509 17661
rect 24451 17620 24460 17660
rect 24500 17620 24509 17660
rect 24451 17619 24509 17620
rect 26659 17660 26717 17661
rect 26659 17620 26668 17660
rect 26708 17620 26717 17660
rect 26659 17619 26717 17620
rect 33387 17660 33429 17669
rect 33387 17620 33388 17660
rect 33428 17620 33429 17660
rect 33387 17611 33429 17620
rect 33579 17660 33621 17669
rect 33579 17620 33580 17660
rect 33620 17620 33621 17660
rect 33579 17611 33621 17620
rect 5635 17576 5693 17577
rect 5635 17536 5644 17576
rect 5684 17536 5693 17576
rect 5635 17535 5693 17536
rect 19363 17576 19421 17577
rect 19363 17536 19372 17576
rect 19412 17536 19421 17576
rect 19363 17535 19421 17536
rect 19659 17576 19701 17585
rect 19659 17536 19660 17576
rect 19700 17536 19701 17576
rect 19659 17527 19701 17536
rect 22147 17576 22205 17577
rect 22147 17536 22156 17576
rect 22196 17536 22205 17576
rect 22147 17535 22205 17536
rect 22339 17576 22397 17577
rect 22339 17536 22348 17576
rect 22388 17536 22397 17576
rect 22339 17535 22397 17536
rect 24163 17576 24221 17577
rect 24163 17536 24172 17576
rect 24212 17536 24221 17576
rect 24163 17535 24221 17536
rect 28203 17576 28245 17585
rect 28203 17536 28204 17576
rect 28244 17536 28245 17576
rect 28203 17527 28245 17536
rect 29547 17576 29589 17585
rect 29547 17536 29548 17576
rect 29588 17536 29589 17576
rect 29547 17527 29589 17536
rect 30595 17576 30653 17577
rect 30595 17536 30604 17576
rect 30644 17536 30653 17576
rect 30595 17535 30653 17536
rect 37323 17576 37365 17585
rect 37323 17536 37324 17576
rect 37364 17536 37365 17576
rect 37323 17527 37365 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 6987 17298 7029 17307
rect 6987 17258 6988 17298
rect 7028 17258 7029 17298
rect 6987 17249 7029 17258
rect 643 17240 701 17241
rect 643 17200 652 17240
rect 692 17200 701 17240
rect 643 17199 701 17200
rect 3715 17240 3773 17241
rect 3715 17200 3724 17240
rect 3764 17200 3773 17240
rect 3715 17199 3773 17200
rect 6219 17240 6261 17249
rect 6219 17200 6220 17240
rect 6260 17200 6261 17240
rect 6219 17191 6261 17200
rect 16291 17240 16349 17241
rect 16291 17200 16300 17240
rect 16340 17200 16349 17240
rect 16291 17199 16349 17200
rect 18307 17240 18365 17241
rect 18307 17200 18316 17240
rect 18356 17200 18365 17240
rect 18307 17199 18365 17200
rect 18411 17240 18453 17249
rect 18411 17200 18412 17240
rect 18452 17200 18453 17240
rect 18411 17191 18453 17200
rect 18691 17240 18749 17241
rect 18691 17200 18700 17240
rect 18740 17200 18749 17240
rect 18691 17199 18749 17200
rect 21867 17240 21909 17249
rect 21867 17200 21868 17240
rect 21908 17200 21909 17240
rect 21867 17191 21909 17200
rect 22531 17240 22589 17241
rect 22531 17200 22540 17240
rect 22580 17200 22589 17240
rect 22531 17199 22589 17200
rect 24843 17240 24885 17249
rect 24843 17200 24844 17240
rect 24884 17200 24885 17240
rect 24843 17191 24885 17200
rect 25227 17240 25269 17249
rect 25227 17200 25228 17240
rect 25268 17200 25269 17240
rect 25227 17191 25269 17200
rect 26571 17240 26613 17249
rect 26571 17200 26572 17240
rect 26612 17200 26613 17240
rect 26571 17191 26613 17200
rect 16011 17156 16053 17165
rect 16011 17116 16012 17156
rect 16052 17116 16053 17156
rect 16011 17107 16053 17116
rect 18211 17156 18269 17157
rect 18211 17116 18220 17156
rect 18260 17116 18269 17156
rect 18211 17115 18269 17116
rect 18787 17156 18845 17157
rect 18787 17116 18796 17156
rect 18836 17116 18845 17156
rect 18787 17115 18845 17116
rect 22251 17156 22293 17165
rect 22251 17116 22252 17156
rect 22292 17116 22293 17156
rect 22251 17107 22293 17116
rect 43267 17156 43325 17157
rect 43267 17116 43276 17156
rect 43316 17116 43325 17156
rect 43267 17115 43325 17116
rect 1323 17072 1365 17081
rect 1323 17032 1324 17072
rect 1364 17032 1365 17072
rect 1323 17023 1365 17032
rect 1699 17072 1757 17073
rect 1699 17032 1708 17072
rect 1748 17032 1757 17072
rect 1699 17031 1757 17032
rect 2563 17072 2621 17073
rect 2563 17032 2572 17072
rect 2612 17032 2621 17072
rect 2563 17031 2621 17032
rect 3907 17072 3965 17073
rect 3907 17032 3916 17072
rect 3956 17032 3965 17072
rect 3907 17031 3965 17032
rect 4867 17072 4925 17073
rect 4867 17032 4876 17072
rect 4916 17032 4925 17072
rect 4867 17031 4925 17032
rect 5923 17072 5981 17073
rect 5923 17032 5932 17072
rect 5972 17032 5981 17072
rect 5923 17031 5981 17032
rect 6115 17072 6173 17073
rect 6115 17032 6124 17072
rect 6164 17032 6173 17072
rect 6115 17031 6173 17032
rect 6403 17072 6461 17073
rect 6403 17032 6412 17072
rect 6452 17032 6461 17072
rect 6403 17031 6461 17032
rect 6507 17072 6549 17081
rect 6507 17032 6508 17072
rect 6548 17032 6549 17072
rect 6507 17023 6549 17032
rect 7179 17072 7221 17081
rect 7179 17032 7180 17072
rect 7220 17032 7221 17072
rect 7075 17030 7133 17031
rect 6603 16988 6645 16997
rect 7075 16990 7084 17030
rect 7124 16990 7133 17030
rect 7179 17023 7221 17032
rect 8323 17072 8381 17073
rect 8323 17032 8332 17072
rect 8372 17032 8381 17072
rect 8323 17031 8381 17032
rect 8515 17072 8573 17073
rect 8515 17032 8524 17072
rect 8564 17032 8573 17072
rect 8515 17031 8573 17032
rect 9195 17072 9237 17081
rect 9195 17032 9196 17072
rect 9236 17032 9237 17072
rect 9195 17023 9237 17032
rect 9387 17072 9429 17081
rect 9387 17032 9388 17072
rect 9428 17032 9429 17072
rect 9387 17023 9429 17032
rect 9763 17072 9821 17073
rect 9763 17032 9772 17072
rect 9812 17032 9821 17072
rect 9763 17031 9821 17032
rect 10627 17072 10685 17073
rect 10627 17032 10636 17072
rect 10676 17032 10685 17072
rect 10627 17031 10685 17032
rect 11787 17072 11829 17081
rect 11787 17032 11788 17072
rect 11828 17032 11829 17072
rect 11787 17023 11829 17032
rect 13987 17072 14045 17073
rect 13987 17032 13996 17072
rect 14036 17032 14045 17072
rect 13987 17031 14045 17032
rect 15915 17072 15957 17081
rect 15915 17032 15916 17072
rect 15956 17032 15957 17072
rect 15915 17023 15957 17032
rect 16099 17072 16157 17073
rect 16099 17032 16108 17072
rect 16148 17032 16157 17072
rect 16099 17031 16157 17032
rect 16963 17072 17021 17073
rect 16963 17032 16972 17072
rect 17012 17032 17021 17072
rect 16963 17031 17021 17032
rect 17163 17072 17205 17081
rect 17163 17032 17164 17072
rect 17204 17032 17205 17072
rect 17163 17023 17205 17032
rect 17827 17072 17885 17073
rect 17827 17032 17836 17072
rect 17876 17032 17885 17072
rect 17827 17031 17885 17032
rect 18027 17072 18069 17081
rect 18027 17032 18028 17072
rect 18068 17032 18069 17072
rect 18027 17023 18069 17032
rect 18123 17072 18165 17081
rect 18123 17032 18124 17072
rect 18164 17032 18165 17072
rect 18123 17023 18165 17032
rect 18891 17072 18933 17081
rect 18891 17032 18892 17072
rect 18932 17032 18933 17072
rect 18891 17023 18933 17032
rect 18987 17072 19029 17081
rect 18987 17032 18988 17072
rect 19028 17032 19029 17072
rect 18987 17023 19029 17032
rect 19171 17072 19229 17073
rect 19171 17032 19180 17072
rect 19220 17032 19229 17072
rect 19171 17031 19229 17032
rect 20043 17072 20085 17081
rect 20043 17032 20044 17072
rect 20084 17032 20085 17072
rect 20043 17023 20085 17032
rect 21003 17072 21045 17081
rect 21003 17032 21004 17072
rect 21044 17032 21045 17072
rect 21003 17023 21045 17032
rect 21187 17072 21245 17073
rect 21187 17032 21196 17072
rect 21236 17032 21245 17072
rect 21187 17031 21245 17032
rect 21955 17072 22013 17073
rect 21955 17032 21964 17072
rect 22004 17032 22013 17072
rect 21955 17031 22013 17032
rect 22155 17072 22197 17081
rect 22155 17032 22156 17072
rect 22196 17032 22197 17072
rect 22155 17023 22197 17032
rect 22339 17072 22397 17073
rect 22339 17032 22348 17072
rect 22388 17032 22397 17072
rect 22339 17031 22397 17032
rect 22627 17072 22685 17073
rect 22627 17032 22636 17072
rect 22676 17032 22685 17072
rect 22627 17031 22685 17032
rect 24267 17072 24309 17081
rect 24267 17032 24268 17072
rect 24308 17032 24309 17072
rect 24267 17023 24309 17032
rect 24747 17072 24789 17081
rect 24747 17032 24748 17072
rect 24788 17032 24789 17072
rect 24747 17023 24789 17032
rect 24939 17072 24981 17081
rect 24939 17032 24940 17072
rect 24980 17032 24981 17072
rect 24939 17023 24981 17032
rect 25131 17072 25173 17081
rect 25131 17032 25132 17072
rect 25172 17032 25173 17072
rect 25131 17023 25173 17032
rect 25419 17072 25461 17081
rect 25419 17032 25420 17072
rect 25460 17032 25461 17072
rect 25419 17023 25461 17032
rect 25611 17072 25653 17081
rect 25611 17032 25612 17072
rect 25652 17032 25653 17072
rect 25611 17023 25653 17032
rect 25707 17072 25749 17081
rect 25707 17032 25708 17072
rect 25748 17032 25749 17072
rect 25707 17023 25749 17032
rect 25803 17072 25845 17081
rect 25803 17032 25804 17072
rect 25844 17032 25845 17072
rect 25803 17023 25845 17032
rect 25899 17072 25941 17081
rect 25899 17032 25900 17072
rect 25940 17032 25941 17072
rect 25899 17023 25941 17032
rect 26371 17072 26429 17073
rect 26371 17032 26380 17072
rect 26420 17032 26429 17072
rect 26371 17031 26429 17032
rect 26563 17072 26621 17073
rect 26563 17032 26572 17072
rect 26612 17032 26621 17072
rect 26563 17031 26621 17032
rect 27531 17072 27573 17081
rect 27531 17032 27532 17072
rect 27572 17032 27573 17072
rect 27531 17023 27573 17032
rect 27907 17072 27965 17073
rect 27907 17032 27916 17072
rect 27956 17032 27965 17072
rect 27907 17031 27965 17032
rect 28107 17072 28149 17081
rect 28107 17032 28108 17072
rect 28148 17032 28149 17072
rect 28107 17023 28149 17032
rect 28203 17072 28245 17081
rect 28203 17032 28204 17072
rect 28244 17032 28245 17072
rect 28203 17023 28245 17032
rect 28299 17072 28341 17081
rect 28299 17032 28300 17072
rect 28340 17032 28341 17072
rect 28299 17023 28341 17032
rect 28395 17072 28437 17081
rect 28395 17032 28396 17072
rect 28436 17032 28437 17072
rect 28395 17023 28437 17032
rect 28587 17072 28629 17081
rect 28587 17032 28588 17072
rect 28628 17032 28629 17072
rect 28587 17023 28629 17032
rect 28683 17072 28725 17081
rect 28683 17032 28684 17072
rect 28724 17032 28725 17072
rect 28683 17023 28725 17032
rect 28779 17072 28821 17081
rect 28779 17032 28780 17072
rect 28820 17032 28821 17072
rect 28779 17023 28821 17032
rect 28875 17072 28917 17081
rect 28875 17032 28876 17072
rect 28916 17032 28917 17072
rect 28875 17023 28917 17032
rect 29067 17072 29109 17081
rect 29067 17032 29068 17072
rect 29108 17032 29109 17072
rect 29067 17023 29109 17032
rect 29259 17072 29301 17081
rect 29259 17032 29260 17072
rect 29300 17032 29301 17072
rect 29259 17023 29301 17032
rect 29347 17072 29405 17073
rect 29347 17032 29356 17072
rect 29396 17032 29405 17072
rect 29347 17031 29405 17032
rect 29547 17072 29589 17081
rect 29547 17032 29548 17072
rect 29588 17032 29589 17072
rect 29547 17023 29589 17032
rect 29923 17072 29981 17073
rect 29923 17032 29932 17072
rect 29972 17032 29981 17072
rect 29923 17031 29981 17032
rect 30403 17072 30461 17073
rect 30403 17032 30412 17072
rect 30452 17032 30461 17072
rect 30403 17031 30461 17032
rect 30507 17072 30549 17081
rect 30507 17032 30508 17072
rect 30548 17032 30549 17072
rect 30507 17023 30549 17032
rect 30699 17072 30741 17081
rect 30699 17032 30700 17072
rect 30740 17032 30741 17072
rect 30699 17023 30741 17032
rect 30891 17072 30933 17081
rect 30891 17032 30892 17072
rect 30932 17032 30933 17072
rect 30891 17023 30933 17032
rect 30987 17072 31029 17081
rect 30987 17032 30988 17072
rect 31028 17032 31029 17072
rect 30987 17023 31029 17032
rect 31083 17072 31125 17081
rect 31083 17032 31084 17072
rect 31124 17032 31125 17072
rect 31083 17023 31125 17032
rect 31179 17072 31221 17081
rect 31179 17032 31180 17072
rect 31220 17032 31221 17072
rect 31179 17023 31221 17032
rect 31363 17072 31421 17073
rect 31363 17032 31372 17072
rect 31412 17032 31421 17072
rect 31363 17031 31421 17032
rect 31467 17072 31509 17081
rect 31467 17032 31468 17072
rect 31508 17032 31509 17072
rect 31467 17023 31509 17032
rect 32611 17072 32669 17073
rect 32611 17032 32620 17072
rect 32660 17032 32669 17072
rect 32611 17031 32669 17032
rect 33291 17072 33333 17081
rect 33291 17032 33292 17072
rect 33332 17032 33333 17072
rect 33291 17023 33333 17032
rect 33667 17072 33725 17073
rect 33667 17032 33676 17072
rect 33716 17032 33725 17072
rect 33667 17031 33725 17032
rect 34531 17072 34589 17073
rect 34531 17032 34540 17072
rect 34580 17032 34589 17072
rect 34531 17031 34589 17032
rect 36643 17072 36701 17073
rect 36643 17032 36652 17072
rect 36692 17032 36701 17072
rect 36643 17031 36701 17032
rect 37323 17072 37365 17081
rect 37323 17032 37324 17072
rect 37364 17032 37365 17072
rect 37323 17023 37365 17032
rect 37699 17072 37757 17073
rect 37699 17032 37708 17072
rect 37748 17032 37757 17072
rect 37699 17031 37757 17032
rect 38563 17072 38621 17073
rect 38563 17032 38572 17072
rect 38612 17032 38621 17072
rect 38563 17031 38621 17032
rect 42883 17072 42941 17073
rect 42883 17032 42892 17072
rect 42932 17032 42941 17072
rect 42883 17031 42941 17032
rect 44131 17072 44189 17073
rect 44131 17032 44140 17072
rect 44180 17032 44189 17072
rect 44131 17031 44189 17032
rect 7075 16989 7133 16990
rect 6603 16948 6604 16988
rect 6644 16948 6645 16988
rect 6603 16939 6645 16948
rect 24459 16988 24501 16997
rect 24459 16948 24460 16988
rect 24500 16948 24501 16988
rect 24459 16939 24501 16948
rect 27627 16988 27669 16997
rect 27627 16948 27628 16988
rect 27668 16948 27669 16988
rect 27627 16939 27669 16948
rect 27819 16988 27861 16997
rect 27819 16948 27820 16988
rect 27860 16948 27861 16988
rect 27819 16939 27861 16948
rect 29643 16988 29685 16997
rect 29643 16948 29644 16988
rect 29684 16948 29685 16988
rect 29643 16939 29685 16948
rect 29835 16988 29877 16997
rect 29835 16948 29836 16988
rect 29876 16948 29877 16988
rect 29835 16939 29877 16948
rect 31563 16988 31605 16997
rect 31563 16948 31564 16988
rect 31604 16948 31605 16988
rect 31563 16939 31605 16948
rect 35691 16988 35733 16997
rect 35691 16948 35692 16988
rect 35732 16948 35733 16988
rect 35691 16939 35733 16948
rect 37027 16988 37085 16989
rect 37027 16948 37036 16988
rect 37076 16948 37085 16988
rect 37027 16947 37085 16948
rect 39723 16988 39765 16997
rect 39723 16948 39724 16988
rect 39764 16948 39765 16988
rect 39723 16939 39765 16948
rect 6699 16904 6741 16913
rect 6699 16864 6700 16904
rect 6740 16864 6741 16904
rect 6699 16855 6741 16864
rect 6795 16904 6837 16913
rect 6795 16864 6796 16904
rect 6836 16864 6837 16904
rect 6795 16855 6837 16864
rect 7467 16904 7509 16913
rect 7467 16864 7468 16904
rect 7508 16864 7509 16904
rect 7467 16855 7509 16864
rect 12075 16904 12117 16913
rect 12075 16864 12076 16904
rect 12116 16864 12117 16904
rect 12075 16855 12117 16864
rect 15243 16904 15285 16913
rect 15243 16864 15244 16904
rect 15284 16864 15285 16904
rect 15243 16855 15285 16864
rect 27723 16904 27765 16913
rect 27723 16864 27724 16904
rect 27764 16864 27765 16904
rect 27723 16855 27765 16864
rect 29067 16904 29109 16913
rect 29067 16864 29068 16904
rect 29108 16864 29109 16904
rect 29067 16855 29109 16864
rect 29739 16904 29781 16913
rect 29739 16864 29740 16904
rect 29780 16864 29781 16904
rect 29739 16855 29781 16864
rect 30699 16904 30741 16913
rect 30699 16864 30700 16904
rect 30740 16864 30741 16904
rect 30699 16855 30741 16864
rect 31659 16904 31701 16913
rect 31659 16864 31660 16904
rect 31700 16864 31701 16904
rect 31659 16855 31701 16864
rect 5251 16820 5309 16821
rect 5251 16780 5260 16820
rect 5300 16780 5309 16820
rect 5251 16779 5309 16780
rect 7651 16820 7709 16821
rect 7651 16780 7660 16820
rect 7700 16780 7709 16820
rect 7651 16779 7709 16780
rect 14659 16820 14717 16821
rect 14659 16780 14668 16820
rect 14708 16780 14717 16820
rect 14659 16779 14717 16780
rect 18699 16820 18741 16829
rect 18699 16780 18700 16820
rect 18740 16780 18741 16820
rect 18699 16771 18741 16780
rect 21099 16820 21141 16829
rect 21099 16780 21100 16820
rect 21140 16780 21141 16820
rect 21099 16771 21141 16780
rect 22819 16820 22877 16821
rect 22819 16780 22828 16820
rect 22868 16780 22877 16820
rect 22819 16779 22877 16780
rect 24267 16820 24309 16829
rect 24267 16780 24268 16820
rect 24308 16780 24309 16820
rect 24267 16771 24309 16780
rect 31755 16820 31797 16829
rect 31755 16780 31756 16820
rect 31796 16780 31797 16820
rect 31755 16771 31797 16780
rect 31939 16820 31997 16821
rect 31939 16780 31948 16820
rect 31988 16780 31997 16820
rect 31939 16779 31997 16780
rect 35971 16820 36029 16821
rect 35971 16780 35980 16820
rect 36020 16780 36029 16820
rect 35971 16779 36029 16780
rect 36843 16820 36885 16829
rect 36843 16780 36844 16820
rect 36884 16780 36885 16820
rect 36843 16771 36885 16780
rect 42603 16820 42645 16829
rect 42603 16780 42604 16820
rect 42644 16780 42645 16820
rect 42603 16771 42645 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 8331 16484 8373 16493
rect 8331 16444 8332 16484
rect 8372 16444 8373 16484
rect 8331 16435 8373 16444
rect 29643 16484 29685 16493
rect 29643 16444 29644 16484
rect 29684 16444 29685 16484
rect 29643 16435 29685 16444
rect 36939 16484 36981 16493
rect 36939 16444 36940 16484
rect 36980 16444 36981 16484
rect 36939 16435 36981 16444
rect 939 16400 981 16409
rect 939 16360 940 16400
rect 980 16360 981 16400
rect 939 16351 981 16360
rect 2091 16400 2133 16409
rect 2091 16360 2092 16400
rect 2132 16360 2133 16400
rect 2091 16351 2133 16360
rect 10251 16400 10293 16409
rect 10251 16360 10252 16400
rect 10292 16360 10293 16400
rect 10251 16351 10293 16360
rect 13603 16400 13661 16401
rect 13603 16360 13612 16400
rect 13652 16360 13661 16400
rect 13603 16359 13661 16360
rect 16203 16400 16245 16409
rect 16203 16360 16204 16400
rect 16244 16360 16245 16400
rect 16203 16351 16245 16360
rect 16587 16400 16629 16409
rect 16587 16360 16588 16400
rect 16628 16360 16629 16400
rect 16587 16351 16629 16360
rect 17547 16400 17589 16409
rect 17547 16360 17548 16400
rect 17588 16360 17589 16400
rect 17547 16351 17589 16360
rect 21763 16400 21821 16401
rect 21763 16360 21772 16400
rect 21812 16360 21821 16400
rect 21763 16359 21821 16360
rect 27243 16400 27285 16409
rect 27243 16360 27244 16400
rect 27284 16360 27285 16400
rect 27243 16351 27285 16360
rect 31179 16400 31221 16409
rect 31179 16360 31180 16400
rect 31220 16360 31221 16400
rect 31179 16351 31221 16360
rect 32619 16400 32661 16409
rect 32619 16360 32620 16400
rect 32660 16360 32661 16400
rect 32619 16351 32661 16360
rect 37803 16400 37845 16409
rect 37803 16360 37804 16400
rect 37844 16360 37845 16400
rect 37803 16351 37845 16360
rect 38187 16400 38229 16409
rect 38187 16360 38188 16400
rect 38228 16360 38229 16400
rect 38187 16351 38229 16360
rect 16387 16316 16445 16317
rect 16387 16276 16396 16316
rect 16436 16276 16445 16316
rect 16387 16275 16445 16276
rect 21579 16316 21621 16325
rect 21579 16276 21580 16316
rect 21620 16276 21621 16316
rect 21579 16267 21621 16276
rect 27147 16316 27189 16325
rect 27147 16276 27148 16316
rect 27188 16276 27189 16316
rect 27147 16267 27189 16276
rect 27339 16316 27381 16325
rect 27339 16276 27340 16316
rect 27380 16276 27381 16316
rect 27339 16267 27381 16276
rect 34155 16316 34197 16325
rect 34155 16276 34156 16316
rect 34196 16276 34197 16316
rect 34155 16267 34197 16276
rect 35211 16316 35253 16325
rect 35211 16276 35212 16316
rect 35252 16276 35253 16316
rect 35211 16267 35253 16276
rect 41643 16316 41685 16325
rect 41643 16276 41644 16316
rect 41684 16276 41685 16316
rect 41643 16267 41685 16276
rect 1131 16232 1173 16241
rect 1131 16192 1132 16232
rect 1172 16192 1173 16232
rect 1131 16183 1173 16192
rect 1323 16232 1365 16241
rect 1323 16192 1324 16232
rect 1364 16192 1365 16232
rect 1323 16183 1365 16192
rect 1515 16232 1557 16241
rect 1515 16192 1516 16232
rect 1556 16192 1557 16232
rect 1515 16183 1557 16192
rect 1611 16232 1653 16241
rect 1611 16192 1612 16232
rect 1652 16192 1653 16232
rect 1611 16183 1653 16192
rect 1803 16232 1845 16241
rect 1803 16192 1804 16232
rect 1844 16192 1845 16232
rect 1803 16183 1845 16192
rect 1995 16232 2037 16241
rect 1995 16192 1996 16232
rect 2036 16192 2037 16232
rect 1995 16183 2037 16192
rect 2187 16232 2229 16241
rect 2187 16192 2188 16232
rect 2228 16192 2229 16232
rect 2187 16183 2229 16192
rect 2283 16232 2325 16241
rect 2283 16192 2284 16232
rect 2324 16192 2325 16232
rect 2283 16183 2325 16192
rect 3139 16232 3197 16233
rect 3139 16192 3148 16232
rect 3188 16192 3197 16232
rect 3139 16191 3197 16192
rect 4003 16232 4061 16233
rect 4003 16192 4012 16232
rect 4052 16192 4061 16232
rect 4003 16191 4061 16192
rect 4203 16232 4245 16241
rect 4203 16192 4204 16232
rect 4244 16192 4245 16232
rect 4203 16183 4245 16192
rect 4867 16232 4925 16233
rect 4867 16192 4876 16232
rect 4916 16192 4925 16232
rect 4867 16191 4925 16192
rect 5259 16232 5301 16241
rect 5259 16192 5260 16232
rect 5300 16192 5301 16232
rect 5259 16183 5301 16192
rect 5355 16232 5397 16241
rect 5355 16192 5356 16232
rect 5396 16192 5397 16232
rect 5355 16183 5397 16192
rect 6403 16232 6461 16233
rect 6403 16192 6412 16232
rect 6452 16192 6461 16232
rect 6403 16191 6461 16192
rect 6595 16232 6653 16233
rect 6595 16192 6604 16232
rect 6644 16192 6653 16232
rect 6595 16191 6653 16192
rect 7275 16232 7317 16241
rect 7275 16192 7276 16232
rect 7316 16192 7317 16232
rect 7275 16183 7317 16192
rect 8131 16232 8189 16233
rect 8131 16192 8140 16232
rect 8180 16192 8189 16232
rect 8131 16191 8189 16192
rect 8331 16232 8373 16241
rect 8331 16192 8332 16232
rect 8372 16192 8373 16232
rect 8331 16183 8373 16192
rect 8619 16232 8661 16241
rect 8619 16192 8620 16232
rect 8660 16192 8661 16232
rect 8619 16183 8661 16192
rect 9571 16232 9629 16233
rect 9571 16192 9580 16232
rect 9620 16192 9629 16232
rect 9571 16191 9629 16192
rect 10915 16232 10973 16233
rect 10915 16192 10924 16232
rect 10964 16192 10973 16232
rect 10915 16191 10973 16192
rect 11587 16232 11645 16233
rect 11587 16192 11596 16232
rect 11636 16192 11645 16232
rect 11587 16191 11645 16192
rect 12451 16232 12509 16233
rect 12451 16192 12460 16232
rect 12500 16192 12509 16232
rect 12451 16191 12509 16192
rect 14187 16232 14229 16241
rect 14187 16192 14188 16232
rect 14228 16192 14229 16232
rect 14187 16183 14229 16192
rect 15043 16232 15101 16233
rect 15043 16192 15052 16232
rect 15092 16192 15101 16232
rect 15043 16191 15101 16192
rect 16011 16232 16053 16241
rect 16011 16192 16012 16232
rect 16052 16192 16053 16232
rect 16011 16183 16053 16192
rect 16203 16232 16245 16241
rect 16203 16192 16204 16232
rect 16244 16192 16245 16232
rect 16203 16183 16245 16192
rect 16779 16232 16821 16241
rect 16779 16192 16780 16232
rect 16820 16192 16821 16232
rect 16779 16183 16821 16192
rect 16875 16232 16917 16241
rect 16875 16192 16876 16232
rect 16916 16192 16917 16232
rect 16875 16183 16917 16192
rect 16971 16232 17013 16241
rect 16971 16192 16972 16232
rect 17012 16192 17013 16232
rect 16971 16183 17013 16192
rect 17067 16232 17109 16241
rect 17067 16192 17068 16232
rect 17108 16192 17109 16232
rect 17067 16183 17109 16192
rect 17251 16232 17309 16233
rect 17251 16192 17260 16232
rect 17300 16192 17309 16232
rect 17251 16191 17309 16192
rect 17355 16232 17397 16241
rect 17355 16192 17356 16232
rect 17396 16192 17397 16232
rect 17355 16183 17397 16192
rect 17547 16232 17589 16241
rect 17547 16192 17548 16232
rect 17588 16192 17589 16232
rect 17547 16183 17589 16192
rect 18691 16232 18749 16233
rect 18691 16192 18700 16232
rect 18740 16192 18749 16232
rect 18691 16191 18749 16192
rect 20131 16232 20189 16233
rect 20131 16192 20140 16232
rect 20180 16192 20189 16232
rect 20131 16191 20189 16192
rect 20235 16232 20277 16241
rect 20235 16192 20236 16232
rect 20276 16192 20277 16232
rect 20235 16183 20277 16192
rect 20419 16232 20477 16233
rect 20419 16192 20428 16232
rect 20468 16192 20477 16232
rect 20419 16191 20477 16192
rect 20619 16232 20661 16241
rect 20619 16192 20620 16232
rect 20660 16192 20661 16232
rect 20619 16183 20661 16192
rect 20811 16232 20853 16241
rect 20811 16192 20812 16232
rect 20852 16192 20853 16232
rect 20811 16183 20853 16192
rect 20907 16232 20949 16241
rect 20907 16192 20908 16232
rect 20948 16192 20949 16232
rect 20907 16183 20949 16192
rect 21771 16232 21813 16241
rect 21771 16192 21772 16232
rect 21812 16192 21813 16232
rect 21771 16183 21813 16192
rect 23883 16232 23925 16241
rect 23883 16192 23884 16232
rect 23924 16192 23925 16232
rect 23883 16183 23925 16192
rect 24075 16232 24117 16241
rect 24075 16192 24076 16232
rect 24116 16192 24117 16232
rect 24075 16183 24117 16192
rect 25219 16232 25277 16233
rect 25219 16192 25228 16232
rect 25268 16192 25277 16232
rect 25219 16191 25277 16192
rect 25891 16232 25949 16233
rect 25891 16192 25900 16232
rect 25940 16192 25949 16232
rect 25891 16191 25949 16192
rect 27051 16232 27093 16241
rect 27051 16192 27052 16232
rect 27092 16192 27093 16232
rect 27051 16183 27093 16192
rect 27427 16232 27485 16233
rect 27427 16192 27436 16232
rect 27476 16192 27485 16232
rect 27427 16191 27485 16192
rect 27915 16232 27957 16241
rect 27915 16192 27916 16232
rect 27956 16192 27957 16232
rect 27915 16183 27957 16192
rect 28011 16232 28053 16241
rect 28011 16192 28012 16232
rect 28052 16192 28053 16232
rect 28011 16183 28053 16192
rect 28099 16232 28157 16233
rect 28099 16192 28108 16232
rect 28148 16192 28157 16232
rect 28099 16191 28157 16192
rect 29347 16232 29405 16233
rect 29347 16192 29356 16232
rect 29396 16192 29405 16232
rect 29347 16191 29405 16192
rect 29451 16232 29493 16241
rect 29451 16192 29452 16232
rect 29492 16192 29493 16232
rect 29451 16183 29493 16192
rect 29643 16232 29685 16241
rect 29643 16192 29644 16232
rect 29684 16192 29685 16232
rect 29643 16183 29685 16192
rect 30403 16232 30461 16233
rect 30403 16192 30412 16232
rect 30452 16192 30461 16232
rect 30403 16191 30461 16192
rect 30507 16232 30549 16241
rect 30507 16192 30508 16232
rect 30548 16192 30549 16232
rect 30507 16183 30549 16192
rect 30691 16232 30749 16233
rect 30691 16192 30700 16232
rect 30740 16192 30749 16232
rect 30691 16191 30749 16192
rect 31075 16232 31133 16233
rect 31075 16192 31084 16232
rect 31124 16192 31133 16232
rect 31075 16191 31133 16192
rect 31275 16232 31317 16241
rect 31275 16192 31276 16232
rect 31316 16192 31317 16232
rect 31275 16183 31317 16192
rect 32131 16232 32189 16233
rect 32131 16192 32140 16232
rect 32180 16192 32189 16232
rect 32131 16191 32189 16192
rect 32331 16232 32373 16241
rect 32331 16192 32332 16232
rect 32372 16192 32373 16232
rect 32331 16183 32373 16192
rect 32427 16232 32469 16241
rect 32427 16192 32428 16232
rect 32468 16192 32469 16232
rect 32427 16183 32469 16192
rect 34059 16232 34101 16241
rect 34059 16192 34060 16232
rect 34100 16192 34101 16232
rect 34059 16183 34101 16192
rect 34251 16232 34293 16241
rect 34251 16192 34252 16232
rect 34292 16192 34293 16232
rect 34251 16183 34293 16192
rect 35979 16232 36021 16241
rect 35979 16192 35980 16232
rect 36020 16192 36021 16232
rect 35979 16183 36021 16192
rect 36651 16232 36693 16241
rect 36651 16192 36652 16232
rect 36692 16192 36693 16232
rect 36651 16183 36693 16192
rect 36939 16232 36981 16241
rect 36939 16192 36940 16232
rect 36980 16192 36981 16232
rect 37323 16232 37365 16241
rect 36939 16183 36981 16192
rect 37131 16211 37173 16220
rect 37131 16171 37132 16211
rect 37172 16171 37173 16211
rect 37131 16162 37173 16171
rect 37227 16211 37269 16220
rect 37227 16171 37228 16211
rect 37268 16171 37269 16211
rect 37323 16192 37324 16232
rect 37364 16192 37365 16232
rect 37323 16183 37365 16192
rect 37995 16232 38037 16241
rect 37995 16192 37996 16232
rect 38036 16192 38037 16232
rect 37995 16183 38037 16192
rect 38187 16232 38229 16241
rect 38187 16192 38188 16232
rect 38228 16192 38229 16232
rect 38187 16183 38229 16192
rect 38371 16232 38429 16233
rect 38371 16192 38380 16232
rect 38420 16192 38429 16232
rect 38371 16191 38429 16192
rect 39619 16232 39677 16233
rect 39619 16192 39628 16232
rect 39668 16192 39677 16232
rect 39619 16191 39677 16192
rect 40483 16232 40541 16233
rect 40483 16192 40492 16232
rect 40532 16192 40541 16232
rect 40483 16191 40541 16192
rect 41827 16232 41885 16233
rect 41827 16192 41836 16232
rect 41876 16192 41885 16232
rect 41827 16191 41885 16192
rect 37227 16162 37269 16171
rect 1227 16148 1269 16157
rect 1227 16108 1228 16148
rect 1268 16108 1269 16148
rect 1227 16099 1269 16108
rect 5059 16148 5117 16149
rect 5059 16108 5068 16148
rect 5108 16108 5117 16148
rect 5059 16107 5117 16108
rect 11211 16148 11253 16157
rect 11211 16108 11212 16148
rect 11252 16108 11253 16148
rect 11211 16099 11253 16108
rect 32515 16148 32573 16149
rect 32515 16108 32524 16148
rect 32564 16108 32573 16148
rect 32515 16107 32573 16108
rect 39051 16148 39093 16157
rect 39051 16108 39052 16148
rect 39092 16108 39093 16148
rect 39051 16099 39093 16108
rect 39243 16148 39285 16157
rect 39243 16108 39244 16148
rect 39284 16108 39285 16148
rect 39243 16099 39285 16108
rect 1707 16064 1749 16073
rect 1707 16024 1708 16064
rect 1748 16024 1749 16064
rect 1707 16015 1749 16024
rect 2467 16064 2525 16065
rect 2467 16024 2476 16064
rect 2516 16024 2525 16064
rect 2467 16023 2525 16024
rect 3331 16064 3389 16065
rect 3331 16024 3340 16064
rect 3380 16024 3389 16064
rect 3331 16023 3389 16024
rect 5347 16064 5405 16065
rect 5347 16024 5356 16064
rect 5396 16024 5405 16064
rect 5347 16023 5405 16024
rect 5731 16064 5789 16065
rect 5731 16024 5740 16064
rect 5780 16024 5789 16064
rect 5731 16023 5789 16024
rect 7459 16064 7517 16065
rect 7459 16024 7468 16064
rect 7508 16024 7517 16064
rect 7459 16023 7517 16024
rect 8899 16064 8957 16065
rect 8899 16024 8908 16064
rect 8948 16024 8957 16064
rect 8899 16023 8957 16024
rect 18219 16064 18261 16073
rect 18219 16024 18220 16064
rect 18260 16024 18261 16064
rect 18219 16015 18261 16024
rect 20427 16064 20469 16073
rect 20427 16024 20428 16064
rect 20468 16024 20469 16064
rect 20427 16015 20469 16024
rect 20899 16064 20957 16065
rect 20899 16024 20908 16064
rect 20948 16024 20957 16064
rect 20899 16023 20957 16024
rect 23979 16064 24021 16073
rect 23979 16024 23980 16064
rect 24020 16024 24021 16064
rect 23979 16015 24021 16024
rect 24747 16064 24789 16073
rect 24747 16024 24748 16064
rect 24788 16024 24789 16064
rect 24747 16015 24789 16024
rect 25507 16064 25565 16065
rect 25507 16024 25516 16064
rect 25556 16024 25565 16064
rect 25507 16023 25565 16024
rect 25699 16064 25757 16065
rect 25699 16024 25708 16064
rect 25748 16024 25757 16064
rect 25699 16023 25757 16024
rect 30699 16064 30741 16073
rect 30699 16024 30700 16064
rect 30740 16024 30741 16064
rect 30699 16015 30741 16024
rect 31459 16064 31517 16065
rect 31459 16024 31468 16064
rect 31508 16024 31517 16064
rect 31459 16023 31517 16024
rect 32611 16064 32669 16065
rect 32611 16024 32620 16064
rect 32660 16024 32669 16064
rect 32611 16023 32669 16024
rect 37411 16064 37469 16065
rect 37411 16024 37420 16064
rect 37460 16024 37469 16064
rect 37411 16023 37469 16024
rect 42499 16064 42557 16065
rect 42499 16024 42508 16064
rect 42548 16024 42557 16064
rect 42499 16023 42557 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 739 15728 797 15729
rect 739 15688 748 15728
rect 788 15688 797 15728
rect 739 15687 797 15688
rect 3915 15728 3957 15737
rect 3915 15688 3916 15728
rect 3956 15688 3957 15728
rect 3915 15679 3957 15688
rect 7075 15728 7133 15729
rect 7075 15688 7084 15728
rect 7124 15688 7133 15728
rect 7075 15687 7133 15688
rect 7651 15728 7709 15729
rect 7651 15688 7660 15728
rect 7700 15688 7709 15728
rect 7651 15687 7709 15688
rect 10339 15728 10397 15729
rect 10339 15688 10348 15728
rect 10388 15688 10397 15728
rect 10339 15687 10397 15688
rect 20139 15728 20181 15737
rect 20139 15688 20140 15728
rect 20180 15688 20181 15728
rect 20139 15679 20181 15688
rect 21771 15732 21813 15741
rect 21771 15692 21772 15732
rect 21812 15692 21813 15732
rect 21771 15683 21813 15692
rect 28483 15728 28541 15729
rect 28483 15688 28492 15728
rect 28532 15688 28541 15728
rect 28483 15687 28541 15688
rect 29251 15728 29309 15729
rect 29251 15688 29260 15728
rect 29300 15688 29309 15728
rect 29251 15687 29309 15688
rect 29923 15728 29981 15729
rect 29923 15688 29932 15728
rect 29972 15688 29981 15728
rect 29923 15687 29981 15688
rect 33571 15728 33629 15729
rect 33571 15688 33580 15728
rect 33620 15688 33629 15728
rect 33571 15687 33629 15688
rect 38083 15728 38141 15729
rect 38083 15688 38092 15728
rect 38132 15688 38141 15728
rect 38083 15687 38141 15688
rect 7947 15644 7989 15653
rect 7947 15604 7948 15644
rect 7988 15604 7989 15644
rect 7947 15595 7989 15604
rect 26083 15644 26141 15645
rect 26083 15604 26092 15644
rect 26132 15604 26141 15644
rect 26083 15603 26141 15604
rect 27331 15644 27389 15645
rect 27331 15604 27340 15644
rect 27380 15604 27389 15644
rect 27331 15603 27389 15604
rect 28579 15644 28637 15645
rect 28579 15604 28588 15644
rect 28628 15604 28637 15644
rect 28579 15603 28637 15604
rect 29827 15644 29885 15645
rect 29827 15604 29836 15644
rect 29876 15604 29885 15644
rect 29827 15603 29885 15604
rect 1131 15560 1173 15569
rect 1131 15520 1132 15560
rect 1172 15520 1173 15560
rect 1131 15511 1173 15520
rect 1507 15560 1565 15561
rect 1507 15520 1516 15560
rect 1556 15520 1565 15560
rect 1507 15519 1565 15520
rect 2371 15560 2429 15561
rect 2371 15520 2380 15560
rect 2420 15520 2429 15560
rect 2371 15519 2429 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 4011 15560 4053 15569
rect 4011 15520 4012 15560
rect 4052 15520 4053 15560
rect 4011 15511 4053 15520
rect 4867 15560 4925 15561
rect 4867 15520 4876 15560
rect 4916 15520 4925 15560
rect 4867 15519 4925 15520
rect 5163 15560 5205 15569
rect 5163 15520 5164 15560
rect 5204 15520 5205 15560
rect 5163 15511 5205 15520
rect 5355 15560 5397 15569
rect 5355 15520 5356 15560
rect 5396 15520 5397 15560
rect 5355 15511 5397 15520
rect 5451 15560 5493 15569
rect 5451 15520 5452 15560
rect 5492 15520 5493 15560
rect 5451 15511 5493 15520
rect 5635 15560 5693 15561
rect 5635 15520 5644 15560
rect 5684 15520 5693 15560
rect 5635 15519 5693 15520
rect 6507 15560 6549 15569
rect 6507 15520 6508 15560
rect 6548 15520 6549 15560
rect 6507 15511 6549 15520
rect 6603 15560 6645 15569
rect 6603 15520 6604 15560
rect 6644 15520 6645 15560
rect 6603 15511 6645 15520
rect 6699 15560 6741 15569
rect 6699 15520 6700 15560
rect 6740 15520 6741 15560
rect 6699 15511 6741 15520
rect 6795 15560 6837 15569
rect 6795 15520 6796 15560
rect 6836 15520 6837 15560
rect 6795 15511 6837 15520
rect 6987 15560 7029 15569
rect 6987 15520 6988 15560
rect 7028 15520 7029 15560
rect 6987 15511 7029 15520
rect 7179 15560 7221 15569
rect 7179 15520 7180 15560
rect 7220 15520 7221 15560
rect 7179 15511 7221 15520
rect 7267 15560 7325 15561
rect 7267 15520 7276 15560
rect 7316 15520 7325 15560
rect 7267 15519 7325 15520
rect 7459 15560 7517 15561
rect 7459 15520 7468 15560
rect 7508 15520 7517 15560
rect 7459 15519 7517 15520
rect 7563 15560 7605 15569
rect 7563 15520 7564 15560
rect 7604 15520 7605 15560
rect 7563 15511 7605 15520
rect 7755 15560 7797 15569
rect 7755 15520 7756 15560
rect 7796 15520 7797 15560
rect 7755 15511 7797 15520
rect 8323 15560 8381 15561
rect 8323 15520 8332 15560
rect 8372 15520 8381 15560
rect 8323 15519 8381 15520
rect 9187 15560 9245 15561
rect 9187 15520 9196 15560
rect 9236 15520 9245 15560
rect 9187 15519 9245 15520
rect 11979 15560 12021 15569
rect 11979 15520 11980 15560
rect 12020 15520 12021 15560
rect 11979 15511 12021 15520
rect 12547 15560 12605 15561
rect 12547 15520 12556 15560
rect 12596 15520 12605 15560
rect 12547 15519 12605 15520
rect 14371 15560 14429 15561
rect 14371 15520 14380 15560
rect 14420 15520 14429 15560
rect 14371 15519 14429 15520
rect 15235 15560 15293 15561
rect 15235 15520 15244 15560
rect 15284 15520 15293 15560
rect 15235 15519 15293 15520
rect 15627 15560 15669 15569
rect 15627 15520 15628 15560
rect 15668 15520 15669 15560
rect 15627 15511 15669 15520
rect 15819 15560 15861 15569
rect 15819 15520 15820 15560
rect 15860 15520 15861 15560
rect 15819 15511 15861 15520
rect 16483 15560 16541 15561
rect 16483 15520 16492 15560
rect 16532 15520 16541 15560
rect 16483 15519 16541 15520
rect 17643 15560 17685 15569
rect 17643 15520 17644 15560
rect 17684 15520 17685 15560
rect 17643 15511 17685 15520
rect 18411 15560 18453 15569
rect 18411 15520 18412 15560
rect 18452 15520 18453 15560
rect 18411 15511 18453 15520
rect 18507 15560 18549 15569
rect 18507 15520 18508 15560
rect 18548 15520 18549 15560
rect 18507 15511 18549 15520
rect 18595 15560 18653 15561
rect 18595 15520 18604 15560
rect 18644 15520 18653 15560
rect 18595 15519 18653 15520
rect 18795 15560 18837 15569
rect 18795 15520 18796 15560
rect 18836 15520 18837 15560
rect 18795 15511 18837 15520
rect 18891 15560 18933 15569
rect 18891 15520 18892 15560
rect 18932 15520 18933 15560
rect 18891 15511 18933 15520
rect 18987 15560 19029 15569
rect 18987 15520 18988 15560
rect 19028 15520 19029 15560
rect 18987 15511 19029 15520
rect 19083 15560 19125 15569
rect 19083 15520 19084 15560
rect 19124 15520 19125 15560
rect 19083 15511 19125 15520
rect 19275 15560 19317 15569
rect 19275 15520 19276 15560
rect 19316 15520 19317 15560
rect 19275 15511 19317 15520
rect 19467 15560 19509 15569
rect 19467 15520 19468 15560
rect 19508 15520 19509 15560
rect 19467 15511 19509 15520
rect 19659 15560 19701 15569
rect 19659 15520 19660 15560
rect 19700 15520 19701 15560
rect 19659 15511 19701 15520
rect 19755 15560 19797 15569
rect 19755 15520 19756 15560
rect 19796 15520 19797 15560
rect 19755 15511 19797 15520
rect 19947 15560 19989 15569
rect 19947 15520 19948 15560
rect 19988 15520 19989 15560
rect 19947 15511 19989 15520
rect 20131 15560 20189 15561
rect 20131 15520 20140 15560
rect 20180 15520 20189 15560
rect 20131 15519 20189 15520
rect 20331 15560 20373 15569
rect 20331 15520 20332 15560
rect 20372 15520 20373 15560
rect 20331 15511 20373 15520
rect 20419 15560 20477 15561
rect 20419 15520 20428 15560
rect 20468 15520 20477 15560
rect 20419 15519 20477 15520
rect 20619 15560 20661 15569
rect 20619 15520 20620 15560
rect 20660 15520 20661 15560
rect 20619 15511 20661 15520
rect 20715 15560 20757 15569
rect 20715 15520 20716 15560
rect 20756 15520 20757 15560
rect 20715 15511 20757 15520
rect 20811 15560 20853 15569
rect 20811 15520 20812 15560
rect 20852 15520 20853 15560
rect 20811 15511 20853 15520
rect 20907 15560 20949 15569
rect 20907 15520 20908 15560
rect 20948 15520 20949 15560
rect 20907 15511 20949 15520
rect 21859 15560 21917 15561
rect 21859 15520 21868 15560
rect 21908 15520 21917 15560
rect 21859 15519 21917 15520
rect 21963 15560 22005 15569
rect 21963 15520 21964 15560
rect 22004 15520 22005 15560
rect 21963 15511 22005 15520
rect 25219 15560 25277 15561
rect 25219 15520 25228 15560
rect 25268 15520 25277 15560
rect 25219 15519 25277 15520
rect 26859 15560 26901 15569
rect 26859 15520 26860 15560
rect 26900 15520 26901 15560
rect 26859 15511 26901 15520
rect 27523 15560 27581 15561
rect 27523 15520 27532 15560
rect 27572 15520 27581 15560
rect 27523 15519 27581 15520
rect 27811 15560 27869 15561
rect 27811 15520 27820 15560
rect 27860 15520 27869 15560
rect 27811 15519 27869 15520
rect 28683 15560 28725 15569
rect 28683 15520 28684 15560
rect 28724 15520 28725 15560
rect 28683 15511 28725 15520
rect 28779 15560 28821 15569
rect 28779 15520 28780 15560
rect 28820 15520 28821 15560
rect 28779 15511 28821 15520
rect 28971 15560 29013 15569
rect 28971 15520 28972 15560
rect 29012 15520 29013 15560
rect 28971 15511 29013 15520
rect 29067 15560 29109 15569
rect 29067 15520 29068 15560
rect 29108 15520 29109 15560
rect 29067 15511 29109 15520
rect 29163 15560 29205 15569
rect 29163 15520 29164 15560
rect 29204 15520 29205 15560
rect 29163 15511 29205 15520
rect 29643 15560 29685 15569
rect 29643 15520 29644 15560
rect 29684 15520 29685 15560
rect 29643 15511 29685 15520
rect 29739 15560 29781 15569
rect 29739 15520 29740 15560
rect 29780 15520 29781 15560
rect 29739 15511 29781 15520
rect 30307 15560 30365 15561
rect 30307 15520 30316 15560
rect 30356 15520 30365 15560
rect 30307 15519 30365 15520
rect 31467 15560 31509 15569
rect 31467 15520 31468 15560
rect 31508 15520 31509 15560
rect 31467 15511 31509 15520
rect 31563 15560 31605 15569
rect 31563 15520 31564 15560
rect 31604 15520 31605 15560
rect 31563 15511 31605 15520
rect 31659 15560 31701 15569
rect 31659 15520 31660 15560
rect 31700 15520 31701 15560
rect 31659 15511 31701 15520
rect 31755 15560 31797 15569
rect 31755 15520 31756 15560
rect 31796 15520 31797 15560
rect 31755 15511 31797 15520
rect 32331 15560 32373 15569
rect 32331 15520 32332 15560
rect 32372 15520 32373 15560
rect 32331 15511 32373 15520
rect 32523 15560 32565 15569
rect 32523 15520 32524 15560
rect 32564 15520 32565 15560
rect 32523 15511 32565 15520
rect 32619 15560 32661 15569
rect 32619 15520 32620 15560
rect 32660 15520 32661 15560
rect 32619 15511 32661 15520
rect 33091 15560 33149 15561
rect 33091 15520 33100 15560
rect 33140 15520 33149 15560
rect 33091 15519 33149 15520
rect 33195 15560 33237 15569
rect 33195 15520 33196 15560
rect 33236 15520 33237 15560
rect 33195 15511 33237 15520
rect 33387 15560 33429 15569
rect 33387 15520 33388 15560
rect 33428 15520 33429 15560
rect 33387 15511 33429 15520
rect 33667 15560 33725 15561
rect 33667 15520 33676 15560
rect 33716 15520 33725 15560
rect 33667 15519 33725 15520
rect 34059 15560 34101 15569
rect 34059 15520 34060 15560
rect 34100 15520 34101 15560
rect 34059 15511 34101 15520
rect 34155 15560 34197 15569
rect 34155 15520 34156 15560
rect 34196 15520 34197 15560
rect 34155 15511 34197 15520
rect 34251 15560 34293 15569
rect 34251 15520 34252 15560
rect 34292 15520 34293 15560
rect 34251 15511 34293 15520
rect 34347 15560 34389 15569
rect 34347 15520 34348 15560
rect 34388 15520 34389 15560
rect 34347 15511 34389 15520
rect 34531 15560 34589 15561
rect 34531 15520 34540 15560
rect 34580 15520 34589 15560
rect 34531 15519 34589 15520
rect 35211 15560 35253 15569
rect 35211 15520 35212 15560
rect 35252 15520 35253 15560
rect 35211 15511 35253 15520
rect 35403 15560 35445 15569
rect 35403 15520 35404 15560
rect 35444 15520 35445 15560
rect 35403 15511 35445 15520
rect 35779 15560 35837 15561
rect 35779 15520 35788 15560
rect 35828 15520 35837 15560
rect 35779 15519 35837 15520
rect 36643 15560 36701 15561
rect 36643 15520 36652 15560
rect 36692 15520 36701 15560
rect 36643 15519 36701 15520
rect 38187 15560 38229 15569
rect 38187 15520 38188 15560
rect 38228 15520 38229 15560
rect 38187 15511 38229 15520
rect 38283 15560 38325 15569
rect 38283 15520 38284 15560
rect 38324 15520 38325 15560
rect 38283 15511 38325 15520
rect 38379 15560 38421 15569
rect 38379 15520 38380 15560
rect 38420 15520 38421 15560
rect 38379 15511 38421 15520
rect 40963 15560 41021 15561
rect 40963 15520 40972 15560
rect 41012 15520 41021 15560
rect 40963 15519 41021 15520
rect 41923 15560 41981 15561
rect 41923 15520 41932 15560
rect 41972 15520 41981 15560
rect 41923 15519 41981 15520
rect 43939 15560 43997 15561
rect 43939 15520 43948 15560
rect 43988 15520 43997 15560
rect 43939 15519 43997 15520
rect 5259 15476 5301 15485
rect 5259 15436 5260 15476
rect 5300 15436 5301 15476
rect 5259 15427 5301 15436
rect 11211 15476 11253 15485
rect 11211 15436 11212 15476
rect 11252 15436 11253 15476
rect 11211 15427 11253 15436
rect 23875 15476 23933 15477
rect 23875 15436 23884 15476
rect 23924 15436 23933 15476
rect 23875 15435 23933 15436
rect 24363 15476 24405 15485
rect 24363 15436 24364 15476
rect 24404 15436 24405 15476
rect 24363 15427 24405 15436
rect 19467 15392 19509 15401
rect 19467 15352 19468 15392
rect 19508 15352 19509 15392
rect 19467 15343 19509 15352
rect 19651 15392 19709 15393
rect 19651 15352 19660 15392
rect 19700 15352 19709 15392
rect 19651 15351 19709 15352
rect 28675 15392 28733 15393
rect 28675 15352 28684 15392
rect 28724 15352 28733 15392
rect 28675 15351 28733 15352
rect 29931 15392 29973 15401
rect 29931 15352 29932 15392
rect 29972 15352 29973 15392
rect 29931 15343 29973 15352
rect 32611 15392 32669 15393
rect 32611 15352 32620 15392
rect 32660 15352 32669 15392
rect 32611 15351 32669 15352
rect 39723 15392 39765 15401
rect 39723 15352 39724 15392
rect 39764 15352 39765 15392
rect 39723 15343 39765 15352
rect 3531 15308 3573 15317
rect 3531 15268 3532 15308
rect 3572 15268 3573 15308
rect 3531 15259 3573 15268
rect 4195 15308 4253 15309
rect 4195 15268 4204 15308
rect 4244 15268 4253 15308
rect 4195 15267 4253 15268
rect 6307 15308 6365 15309
rect 6307 15268 6316 15308
rect 6356 15268 6365 15308
rect 6307 15267 6365 15268
rect 12651 15308 12693 15317
rect 12651 15268 12652 15308
rect 12692 15268 12693 15308
rect 12651 15259 12693 15268
rect 13227 15308 13269 15317
rect 13227 15268 13228 15308
rect 13268 15268 13269 15308
rect 13227 15259 13269 15268
rect 17067 15308 17109 15317
rect 17067 15268 17068 15308
rect 17108 15268 17109 15308
rect 17067 15259 17109 15268
rect 22251 15308 22293 15317
rect 22251 15268 22252 15308
rect 22292 15268 22293 15308
rect 22251 15259 22293 15268
rect 23691 15308 23733 15317
rect 23691 15268 23692 15308
rect 23732 15268 23733 15308
rect 23691 15259 23733 15268
rect 26283 15308 26325 15317
rect 26283 15268 26284 15308
rect 26324 15268 26325 15308
rect 26283 15259 26325 15268
rect 30603 15308 30645 15317
rect 30603 15268 30604 15308
rect 30644 15268 30645 15308
rect 30603 15259 30645 15268
rect 33387 15308 33429 15317
rect 33387 15268 33388 15308
rect 33428 15268 33429 15308
rect 33387 15259 33429 15268
rect 33859 15308 33917 15309
rect 33859 15268 33868 15308
rect 33908 15268 33917 15308
rect 33859 15267 33917 15268
rect 37803 15308 37845 15317
rect 37803 15268 37804 15308
rect 37844 15268 37845 15308
rect 37803 15259 37845 15268
rect 44427 15308 44469 15317
rect 44427 15268 44428 15308
rect 44468 15268 44469 15308
rect 44427 15259 44469 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 4771 14972 4829 14973
rect 4771 14932 4780 14972
rect 4820 14932 4829 14972
rect 4771 14931 4829 14932
rect 5635 14972 5693 14973
rect 5635 14932 5644 14972
rect 5684 14932 5693 14972
rect 5635 14931 5693 14932
rect 11107 14972 11165 14973
rect 11107 14932 11116 14972
rect 11156 14932 11165 14972
rect 11107 14931 11165 14932
rect 11979 14972 12021 14981
rect 11979 14932 11980 14972
rect 12020 14932 12021 14972
rect 11979 14923 12021 14932
rect 13803 14972 13845 14981
rect 13803 14932 13804 14972
rect 13844 14932 13845 14972
rect 13803 14923 13845 14932
rect 24835 14972 24893 14973
rect 24835 14932 24844 14972
rect 24884 14932 24893 14972
rect 24835 14931 24893 14932
rect 27243 14972 27285 14981
rect 27243 14932 27244 14972
rect 27284 14932 27285 14972
rect 27243 14923 27285 14932
rect 30891 14972 30933 14981
rect 30891 14932 30892 14972
rect 30932 14932 30933 14972
rect 30891 14923 30933 14932
rect 31467 14972 31509 14981
rect 31467 14932 31468 14972
rect 31508 14932 31509 14972
rect 31467 14923 31509 14932
rect 32427 14972 32469 14981
rect 32427 14932 32428 14972
rect 32468 14932 32469 14972
rect 32427 14923 32469 14932
rect 34443 14972 34485 14981
rect 34443 14932 34444 14972
rect 34484 14932 34485 14972
rect 34443 14923 34485 14932
rect 1707 14888 1749 14897
rect 1707 14848 1708 14888
rect 1748 14848 1749 14888
rect 1707 14839 1749 14848
rect 8235 14888 8277 14897
rect 8235 14848 8236 14888
rect 8276 14848 8277 14888
rect 8235 14839 8277 14848
rect 8523 14888 8565 14897
rect 8523 14848 8524 14888
rect 8564 14848 8565 14888
rect 8523 14839 8565 14848
rect 9867 14888 9909 14897
rect 9867 14848 9868 14888
rect 9908 14848 9909 14888
rect 9867 14839 9909 14848
rect 16683 14888 16725 14897
rect 16683 14848 16684 14888
rect 16724 14848 16725 14888
rect 16683 14839 16725 14848
rect 19083 14888 19125 14897
rect 19083 14848 19084 14888
rect 19124 14848 19125 14888
rect 21003 14888 21045 14897
rect 19083 14839 19125 14848
rect 19179 14846 19221 14855
rect 10051 14804 10109 14805
rect 10051 14764 10060 14804
rect 10100 14764 10109 14804
rect 10051 14763 10109 14764
rect 18987 14804 19029 14813
rect 18987 14764 18988 14804
rect 19028 14764 19029 14804
rect 19179 14806 19180 14846
rect 19220 14806 19221 14846
rect 21003 14848 21004 14888
rect 21044 14848 21045 14888
rect 21003 14839 21045 14848
rect 22251 14888 22293 14897
rect 22251 14848 22252 14888
rect 22292 14848 22293 14888
rect 22251 14839 22293 14848
rect 25123 14888 25181 14889
rect 25123 14848 25132 14888
rect 25172 14848 25181 14888
rect 25123 14847 25181 14848
rect 31083 14888 31125 14897
rect 31083 14848 31084 14888
rect 31124 14848 31125 14888
rect 31083 14839 31125 14848
rect 33291 14888 33333 14897
rect 33291 14848 33292 14888
rect 33332 14848 33333 14888
rect 33291 14839 33333 14848
rect 37899 14888 37941 14897
rect 37899 14848 37900 14888
rect 37940 14848 37941 14888
rect 37899 14839 37941 14848
rect 39051 14888 39093 14897
rect 39051 14848 39052 14888
rect 39092 14848 39093 14888
rect 39051 14839 39093 14848
rect 41355 14888 41397 14897
rect 41355 14848 41356 14888
rect 41396 14848 41397 14888
rect 41355 14839 41397 14848
rect 46915 14888 46973 14889
rect 46915 14848 46924 14888
rect 46964 14848 46973 14888
rect 46915 14847 46973 14848
rect 19179 14797 19221 14806
rect 20907 14804 20949 14813
rect 18987 14755 19029 14764
rect 20907 14764 20908 14804
rect 20948 14764 20949 14804
rect 20907 14755 20949 14764
rect 21099 14804 21141 14813
rect 21099 14764 21100 14804
rect 21140 14764 21141 14804
rect 21099 14755 21141 14764
rect 22155 14804 22197 14813
rect 22155 14764 22156 14804
rect 22196 14764 22197 14804
rect 22155 14755 22197 14764
rect 22347 14804 22389 14813
rect 22347 14764 22348 14804
rect 22388 14764 22389 14804
rect 22347 14755 22389 14764
rect 26859 14804 26901 14813
rect 26859 14764 26860 14804
rect 26900 14764 26901 14804
rect 26859 14755 26901 14764
rect 30691 14804 30749 14805
rect 30691 14764 30700 14804
rect 30740 14764 30749 14804
rect 30691 14763 30749 14764
rect 33195 14804 33237 14813
rect 33195 14764 33196 14804
rect 33236 14764 33237 14804
rect 33195 14755 33237 14764
rect 33387 14804 33429 14813
rect 33387 14764 33388 14804
rect 33428 14764 33429 14804
rect 33387 14755 33429 14764
rect 27331 14743 27389 14744
rect 2379 14720 2421 14729
rect 2379 14680 2380 14720
rect 2420 14680 2421 14720
rect 2379 14671 2421 14680
rect 2755 14720 2813 14721
rect 2755 14680 2764 14720
rect 2804 14680 2813 14720
rect 2755 14679 2813 14680
rect 3619 14720 3677 14721
rect 3619 14680 3628 14720
rect 3668 14680 3677 14720
rect 3619 14679 3677 14680
rect 5163 14720 5205 14729
rect 5163 14680 5164 14720
rect 5204 14680 5205 14720
rect 5163 14671 5205 14680
rect 5259 14720 5301 14729
rect 5259 14680 5260 14720
rect 5300 14680 5301 14720
rect 5259 14671 5301 14680
rect 5355 14720 5397 14729
rect 5355 14680 5356 14720
rect 5396 14680 5397 14720
rect 5355 14671 5397 14680
rect 5451 14720 5493 14729
rect 5451 14680 5452 14720
rect 5492 14680 5493 14720
rect 5451 14671 5493 14680
rect 5835 14720 5877 14729
rect 5835 14680 5836 14720
rect 5876 14680 5877 14720
rect 5835 14671 5877 14680
rect 6211 14720 6269 14721
rect 6211 14680 6220 14720
rect 6260 14680 6269 14720
rect 6211 14679 6269 14680
rect 7075 14720 7133 14721
rect 7075 14680 7084 14720
rect 7124 14680 7133 14720
rect 7075 14679 7133 14680
rect 8907 14720 8949 14729
rect 8907 14680 8908 14720
rect 8948 14680 8949 14720
rect 8907 14671 8949 14680
rect 9099 14720 9141 14729
rect 9099 14680 9100 14720
rect 9140 14680 9141 14720
rect 9099 14671 9141 14680
rect 10435 14720 10493 14721
rect 10435 14680 10444 14720
rect 10484 14680 10493 14720
rect 10435 14679 10493 14680
rect 11299 14720 11357 14721
rect 11299 14680 11308 14720
rect 11348 14680 11357 14720
rect 11299 14679 11357 14680
rect 12259 14720 12317 14721
rect 12259 14680 12268 14720
rect 12308 14680 12317 14720
rect 12843 14720 12885 14729
rect 12259 14679 12317 14680
rect 12651 14699 12693 14708
rect 12651 14659 12652 14699
rect 12692 14659 12693 14699
rect 12651 14650 12693 14659
rect 12747 14699 12789 14708
rect 12747 14659 12748 14699
rect 12788 14659 12789 14699
rect 12843 14680 12844 14720
rect 12884 14680 12885 14720
rect 12843 14671 12885 14680
rect 13227 14720 13269 14729
rect 13227 14680 13228 14720
rect 13268 14680 13269 14720
rect 13227 14671 13269 14680
rect 14947 14720 15005 14721
rect 14947 14680 14956 14720
rect 14996 14680 15005 14720
rect 14947 14679 15005 14680
rect 15235 14720 15293 14721
rect 15235 14680 15244 14720
rect 15284 14680 15293 14720
rect 15235 14679 15293 14680
rect 15339 14720 15381 14729
rect 15339 14680 15340 14720
rect 15380 14680 15381 14720
rect 15339 14671 15381 14680
rect 15531 14720 15573 14729
rect 15531 14680 15532 14720
rect 15572 14680 15573 14720
rect 15531 14671 15573 14680
rect 15715 14720 15773 14721
rect 15715 14680 15724 14720
rect 15764 14680 15773 14720
rect 15715 14679 15773 14680
rect 16195 14720 16253 14721
rect 16195 14680 16204 14720
rect 16244 14680 16253 14720
rect 16195 14679 16253 14680
rect 16299 14720 16341 14729
rect 16299 14680 16300 14720
rect 16340 14680 16341 14720
rect 16299 14671 16341 14680
rect 16491 14720 16533 14729
rect 16491 14680 16492 14720
rect 16532 14680 16533 14720
rect 16491 14671 16533 14680
rect 16683 14720 16725 14729
rect 16683 14680 16684 14720
rect 16724 14680 16725 14720
rect 16683 14671 16725 14680
rect 16963 14720 17021 14721
rect 16963 14680 16972 14720
rect 17012 14680 17021 14720
rect 16963 14679 17021 14680
rect 18123 14720 18165 14729
rect 18123 14680 18124 14720
rect 18164 14680 18165 14720
rect 18123 14671 18165 14680
rect 18499 14720 18557 14721
rect 18499 14680 18508 14720
rect 18548 14680 18557 14720
rect 18499 14679 18557 14680
rect 18883 14720 18941 14721
rect 18883 14680 18892 14720
rect 18932 14680 18941 14720
rect 18883 14679 18941 14680
rect 19275 14720 19317 14729
rect 19275 14680 19276 14720
rect 19316 14680 19317 14720
rect 19275 14671 19317 14680
rect 19755 14720 19797 14729
rect 19755 14680 19756 14720
rect 19796 14680 19797 14720
rect 19755 14671 19797 14680
rect 19851 14720 19893 14729
rect 19851 14680 19852 14720
rect 19892 14680 19893 14720
rect 19851 14671 19893 14680
rect 20043 14720 20085 14729
rect 20043 14680 20044 14720
rect 20084 14680 20085 14720
rect 20043 14671 20085 14680
rect 20331 14720 20373 14729
rect 20331 14680 20332 14720
rect 20372 14680 20373 14720
rect 20331 14671 20373 14680
rect 20427 14720 20469 14729
rect 20427 14680 20428 14720
rect 20468 14680 20469 14720
rect 20427 14671 20469 14680
rect 20523 14720 20565 14729
rect 20523 14680 20524 14720
rect 20564 14680 20565 14720
rect 20523 14671 20565 14680
rect 20619 14720 20661 14729
rect 20619 14680 20620 14720
rect 20660 14680 20661 14720
rect 20619 14671 20661 14680
rect 20803 14720 20861 14721
rect 20803 14680 20812 14720
rect 20852 14680 20861 14720
rect 20803 14679 20861 14680
rect 21195 14720 21237 14729
rect 21195 14680 21196 14720
rect 21236 14680 21237 14720
rect 21195 14671 21237 14680
rect 21379 14720 21437 14721
rect 21379 14680 21388 14720
rect 21428 14680 21437 14720
rect 21379 14679 21437 14680
rect 21483 14720 21525 14729
rect 21483 14680 21484 14720
rect 21524 14680 21525 14720
rect 21483 14671 21525 14680
rect 21579 14720 21621 14729
rect 21579 14680 21580 14720
rect 21620 14680 21621 14720
rect 21579 14671 21621 14680
rect 22051 14720 22109 14721
rect 22051 14680 22060 14720
rect 22100 14680 22109 14720
rect 22051 14679 22109 14680
rect 22443 14720 22485 14729
rect 22443 14680 22444 14720
rect 22484 14680 22485 14720
rect 22443 14671 22485 14680
rect 23595 14720 23637 14729
rect 23595 14680 23596 14720
rect 23636 14680 23637 14720
rect 23595 14671 23637 14680
rect 23691 14720 23733 14729
rect 23691 14680 23692 14720
rect 23732 14680 23733 14720
rect 23691 14671 23733 14680
rect 23787 14720 23829 14729
rect 23787 14680 23788 14720
rect 23828 14680 23829 14720
rect 23787 14671 23829 14680
rect 23979 14720 24021 14729
rect 23979 14680 23980 14720
rect 24020 14680 24021 14720
rect 23979 14671 24021 14680
rect 24075 14720 24117 14729
rect 24075 14680 24076 14720
rect 24116 14680 24117 14720
rect 24075 14671 24117 14680
rect 24163 14720 24221 14721
rect 24163 14680 24172 14720
rect 24212 14680 24221 14720
rect 24163 14679 24221 14680
rect 24355 14720 24413 14721
rect 24355 14680 24364 14720
rect 24404 14680 24413 14720
rect 24355 14679 24413 14680
rect 24555 14720 24597 14729
rect 24555 14680 24556 14720
rect 24596 14680 24597 14720
rect 24555 14671 24597 14680
rect 24643 14720 24701 14721
rect 24643 14680 24652 14720
rect 24692 14680 24701 14720
rect 24643 14679 24701 14680
rect 25419 14720 25461 14729
rect 25419 14680 25420 14720
rect 25460 14680 25461 14720
rect 25419 14671 25461 14680
rect 25515 14720 25557 14729
rect 25515 14680 25516 14720
rect 25556 14680 25557 14720
rect 25515 14671 25557 14680
rect 25795 14720 25853 14721
rect 25795 14680 25804 14720
rect 25844 14680 25853 14720
rect 25795 14679 25853 14680
rect 26179 14720 26237 14721
rect 26179 14680 26188 14720
rect 26228 14680 26237 14720
rect 26179 14679 26237 14680
rect 26763 14720 26805 14729
rect 26763 14680 26764 14720
rect 26804 14680 26805 14720
rect 26763 14671 26805 14680
rect 26947 14720 27005 14721
rect 26947 14680 26956 14720
rect 26996 14680 27005 14720
rect 26947 14679 27005 14680
rect 27147 14720 27189 14729
rect 27147 14680 27148 14720
rect 27188 14680 27189 14720
rect 27331 14703 27340 14743
rect 27380 14703 27389 14743
rect 27331 14702 27389 14703
rect 27531 14720 27573 14729
rect 27147 14671 27189 14680
rect 27531 14680 27532 14720
rect 27572 14680 27573 14720
rect 27531 14671 27573 14680
rect 27715 14720 27773 14721
rect 27715 14680 27724 14720
rect 27764 14680 27773 14720
rect 27715 14679 27773 14680
rect 28107 14720 28149 14729
rect 28107 14680 28108 14720
rect 28148 14680 28149 14720
rect 28107 14671 28149 14680
rect 28195 14720 28253 14721
rect 28195 14680 28204 14720
rect 28244 14680 28253 14720
rect 28195 14679 28253 14680
rect 28675 14720 28733 14721
rect 28675 14680 28684 14720
rect 28724 14680 28733 14720
rect 28675 14679 28733 14680
rect 28779 14720 28821 14729
rect 28779 14680 28780 14720
rect 28820 14680 28821 14720
rect 28779 14671 28821 14680
rect 28971 14720 29013 14729
rect 28971 14680 28972 14720
rect 29012 14680 29013 14720
rect 28971 14671 29013 14680
rect 29163 14720 29205 14729
rect 29163 14680 29164 14720
rect 29204 14680 29205 14720
rect 29163 14671 29205 14680
rect 29259 14720 29301 14729
rect 29259 14680 29260 14720
rect 29300 14680 29301 14720
rect 29259 14671 29301 14680
rect 29355 14720 29397 14729
rect 29355 14680 29356 14720
rect 29396 14680 29397 14720
rect 29355 14671 29397 14680
rect 29451 14720 29493 14729
rect 29451 14680 29452 14720
rect 29492 14680 29493 14720
rect 29451 14671 29493 14680
rect 29635 14720 29693 14721
rect 29635 14680 29644 14720
rect 29684 14680 29693 14720
rect 29635 14679 29693 14680
rect 29739 14720 29781 14729
rect 29739 14680 29740 14720
rect 29780 14680 29781 14720
rect 29739 14671 29781 14680
rect 29931 14720 29973 14729
rect 29931 14680 29932 14720
rect 29972 14680 29973 14720
rect 29931 14671 29973 14680
rect 31083 14720 31125 14729
rect 31083 14680 31084 14720
rect 31124 14680 31125 14720
rect 31083 14671 31125 14680
rect 31275 14720 31317 14729
rect 31275 14680 31276 14720
rect 31316 14680 31317 14720
rect 31275 14671 31317 14680
rect 31467 14720 31509 14729
rect 31467 14680 31468 14720
rect 31508 14680 31509 14720
rect 31747 14720 31805 14721
rect 31467 14671 31509 14680
rect 31659 14678 31701 14687
rect 31747 14680 31756 14720
rect 31796 14680 31805 14720
rect 31747 14679 31805 14680
rect 31947 14720 31989 14729
rect 31947 14680 31948 14720
rect 31988 14680 31989 14720
rect 12747 14650 12789 14659
rect 15435 14636 15477 14645
rect 15435 14596 15436 14636
rect 15476 14596 15477 14636
rect 15435 14587 15477 14596
rect 15819 14636 15861 14645
rect 15819 14596 15820 14636
rect 15860 14596 15861 14636
rect 15819 14587 15861 14596
rect 18603 14636 18645 14645
rect 18603 14596 18604 14636
rect 18644 14596 18645 14636
rect 18603 14587 18645 14596
rect 27627 14636 27669 14645
rect 27627 14596 27628 14636
rect 27668 14596 27669 14636
rect 27627 14587 27669 14596
rect 29835 14636 29877 14645
rect 29835 14596 29836 14636
rect 29876 14596 29877 14636
rect 31659 14638 31660 14678
rect 31700 14638 31701 14678
rect 31947 14671 31989 14680
rect 32043 14720 32085 14729
rect 32043 14680 32044 14720
rect 32084 14680 32085 14720
rect 32043 14671 32085 14680
rect 32139 14720 32181 14729
rect 32139 14680 32140 14720
rect 32180 14680 32181 14720
rect 32139 14671 32181 14680
rect 32235 14720 32277 14729
rect 32235 14680 32236 14720
rect 32276 14680 32277 14720
rect 32235 14671 32277 14680
rect 32715 14720 32757 14729
rect 32715 14680 32716 14720
rect 32756 14680 32757 14720
rect 32715 14671 32757 14680
rect 32803 14720 32861 14721
rect 32803 14680 32812 14720
rect 32852 14680 32861 14720
rect 32803 14679 32861 14680
rect 33099 14720 33141 14729
rect 33099 14680 33100 14720
rect 33140 14680 33141 14720
rect 33099 14671 33141 14680
rect 33475 14720 33533 14721
rect 33475 14680 33484 14720
rect 33524 14680 33533 14720
rect 33475 14679 33533 14680
rect 33675 14720 33717 14729
rect 33675 14680 33676 14720
rect 33716 14680 33717 14720
rect 33675 14671 33717 14680
rect 33771 14720 33813 14729
rect 33771 14680 33772 14720
rect 33812 14680 33813 14720
rect 33771 14671 33813 14680
rect 33867 14720 33909 14729
rect 33867 14680 33868 14720
rect 33908 14680 33909 14720
rect 33867 14671 33909 14680
rect 33963 14720 34005 14729
rect 33963 14680 33964 14720
rect 34004 14680 34005 14720
rect 33963 14671 34005 14680
rect 34147 14720 34205 14721
rect 34147 14680 34156 14720
rect 34196 14680 34205 14720
rect 34147 14679 34205 14680
rect 34251 14720 34293 14729
rect 34251 14680 34252 14720
rect 34292 14680 34293 14720
rect 34251 14671 34293 14680
rect 34443 14720 34485 14729
rect 34443 14680 34444 14720
rect 34484 14680 34485 14720
rect 34443 14671 34485 14680
rect 34635 14720 34677 14729
rect 34635 14680 34636 14720
rect 34676 14680 34677 14720
rect 34635 14671 34677 14680
rect 34731 14720 34773 14729
rect 34731 14680 34732 14720
rect 34772 14680 34773 14720
rect 34731 14671 34773 14680
rect 34819 14720 34877 14721
rect 34819 14680 34828 14720
rect 34868 14680 34877 14720
rect 34819 14679 34877 14680
rect 37603 14720 37661 14721
rect 37603 14680 37612 14720
rect 37652 14680 37661 14720
rect 37603 14679 37661 14680
rect 39715 14720 39773 14721
rect 39715 14680 39724 14720
rect 39764 14680 39773 14720
rect 39715 14679 39773 14680
rect 40963 14720 41021 14721
rect 40963 14680 40972 14720
rect 41012 14680 41021 14720
rect 40963 14679 41021 14680
rect 41067 14720 41109 14729
rect 41067 14680 41068 14720
rect 41108 14680 41109 14720
rect 41067 14671 41109 14680
rect 41739 14720 41781 14729
rect 41739 14680 41740 14720
rect 41780 14680 41781 14720
rect 41739 14671 41781 14680
rect 42115 14720 42173 14721
rect 42115 14680 42124 14720
rect 42164 14680 42173 14720
rect 42115 14679 42173 14680
rect 42979 14720 43037 14721
rect 42979 14680 42988 14720
rect 43028 14680 43037 14720
rect 42979 14679 43037 14680
rect 44139 14720 44181 14729
rect 44139 14680 44140 14720
rect 44180 14680 44181 14720
rect 44139 14671 44181 14680
rect 44515 14720 44573 14721
rect 44515 14680 44524 14720
rect 44564 14680 44573 14720
rect 44515 14679 44573 14680
rect 45667 14720 45725 14721
rect 45667 14680 45676 14720
rect 45716 14680 45725 14720
rect 45667 14679 45725 14680
rect 46539 14720 46581 14729
rect 46539 14680 46540 14720
rect 46580 14680 46581 14720
rect 46539 14671 46581 14680
rect 47587 14720 47645 14721
rect 47587 14680 47596 14720
rect 47636 14680 47645 14720
rect 47587 14679 47645 14680
rect 31659 14629 31701 14638
rect 29835 14587 29877 14596
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 1027 14552 1085 14553
rect 1027 14512 1036 14552
rect 1076 14512 1085 14552
rect 1027 14511 1085 14512
rect 9003 14552 9045 14561
rect 9003 14512 9004 14552
rect 9044 14512 9045 14552
rect 9003 14503 9045 14512
rect 11787 14552 11829 14561
rect 11787 14512 11788 14552
rect 11828 14512 11829 14552
rect 11787 14503 11829 14512
rect 12547 14552 12605 14553
rect 12547 14512 12556 14552
rect 12596 14512 12605 14552
rect 12547 14511 12605 14512
rect 14275 14552 14333 14553
rect 14275 14512 14284 14552
rect 14324 14512 14333 14552
rect 14275 14511 14333 14512
rect 17451 14552 17493 14561
rect 17451 14512 17452 14552
rect 17492 14512 17493 14552
rect 17451 14503 17493 14512
rect 19947 14552 19989 14561
rect 19947 14512 19948 14552
rect 19988 14512 19989 14552
rect 19947 14503 19989 14512
rect 23491 14552 23549 14553
rect 23491 14512 23500 14552
rect 23540 14512 23549 14552
rect 23491 14511 23549 14512
rect 26083 14552 26141 14553
rect 26083 14512 26092 14552
rect 26132 14512 26141 14552
rect 26083 14511 26141 14512
rect 26371 14552 26429 14553
rect 26371 14512 26380 14552
rect 26420 14512 26429 14552
rect 26371 14511 26429 14512
rect 28491 14552 28533 14561
rect 28491 14512 28492 14552
rect 28532 14512 28533 14552
rect 28491 14503 28533 14512
rect 28867 14552 28925 14553
rect 28867 14512 28876 14552
rect 28916 14512 28925 14552
rect 28867 14511 28925 14512
rect 32907 14548 32949 14557
rect 32907 14508 32908 14548
rect 32948 14508 32949 14548
rect 32907 14499 32949 14508
rect 40875 14548 40917 14557
rect 40875 14508 40876 14548
rect 40916 14508 40917 14548
rect 40875 14499 40917 14508
rect 45003 14552 45045 14561
rect 45003 14512 45004 14552
rect 45044 14512 45045 14552
rect 45003 14503 45045 14512
rect 46915 14552 46973 14553
rect 46915 14512 46924 14552
rect 46964 14512 46973 14552
rect 46915 14511 46973 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 643 14216 701 14217
rect 643 14176 652 14216
rect 692 14176 701 14216
rect 643 14175 701 14176
rect 4003 14216 4061 14217
rect 4003 14176 4012 14216
rect 4052 14176 4061 14216
rect 4003 14175 4061 14176
rect 4291 14216 4349 14217
rect 4291 14176 4300 14216
rect 4340 14176 4349 14216
rect 4291 14175 4349 14176
rect 5643 14216 5685 14225
rect 5643 14176 5644 14216
rect 5684 14176 5685 14216
rect 5643 14167 5685 14176
rect 6315 14216 6357 14225
rect 6315 14176 6316 14216
rect 6356 14176 6357 14216
rect 6315 14167 6357 14176
rect 6603 14216 6645 14225
rect 6603 14176 6604 14216
rect 6644 14176 6645 14216
rect 6603 14167 6645 14176
rect 9763 14216 9821 14217
rect 9763 14176 9772 14216
rect 9812 14176 9821 14216
rect 9763 14175 9821 14176
rect 15619 14216 15677 14217
rect 15619 14176 15628 14216
rect 15668 14176 15677 14216
rect 15619 14175 15677 14176
rect 17155 14216 17213 14217
rect 17155 14176 17164 14216
rect 17204 14176 17213 14216
rect 17155 14175 17213 14176
rect 18403 14216 18461 14217
rect 18403 14176 18412 14216
rect 18452 14176 18461 14216
rect 18403 14175 18461 14176
rect 21091 14216 21149 14217
rect 21091 14176 21100 14216
rect 21140 14176 21149 14216
rect 21091 14175 21149 14176
rect 22243 14216 22301 14217
rect 22243 14176 22252 14216
rect 22292 14176 22301 14216
rect 22243 14175 22301 14176
rect 22435 14216 22493 14217
rect 22435 14176 22444 14216
rect 22484 14176 22493 14216
rect 22435 14175 22493 14176
rect 23107 14216 23165 14217
rect 23107 14176 23116 14216
rect 23156 14176 23165 14216
rect 23107 14175 23165 14176
rect 26091 14216 26133 14225
rect 26091 14176 26092 14216
rect 26132 14176 26133 14216
rect 26091 14167 26133 14176
rect 35203 14216 35261 14217
rect 35203 14176 35212 14216
rect 35252 14176 35261 14216
rect 35203 14175 35261 14176
rect 36163 14216 36221 14217
rect 36163 14176 36172 14216
rect 36212 14176 36221 14216
rect 36163 14175 36221 14176
rect 37123 14216 37181 14217
rect 37123 14176 37132 14216
rect 37172 14176 37181 14216
rect 37123 14175 37181 14176
rect 38379 14216 38421 14225
rect 38379 14176 38380 14216
rect 38420 14176 38421 14216
rect 38379 14167 38421 14176
rect 41731 14216 41789 14217
rect 41731 14176 41740 14216
rect 41780 14176 41789 14216
rect 41731 14175 41789 14176
rect 42019 14216 42077 14217
rect 42019 14176 42028 14216
rect 42068 14176 42077 14216
rect 42019 14175 42077 14176
rect 20043 14132 20085 14141
rect 20043 14092 20044 14132
rect 20084 14092 20085 14132
rect 20043 14083 20085 14092
rect 22923 14132 22965 14141
rect 22923 14092 22924 14132
rect 22964 14092 22965 14132
rect 22923 14083 22965 14092
rect 27435 14132 27477 14141
rect 27435 14092 27436 14132
rect 27476 14092 27477 14132
rect 27435 14083 27477 14092
rect 31939 14069 31997 14070
rect 18696 14057 18754 14058
rect 3243 14048 3285 14057
rect 3243 14008 3244 14048
rect 3284 14008 3285 14048
rect 3243 13999 3285 14008
rect 3435 14048 3477 14057
rect 3435 14008 3436 14048
rect 3476 14008 3477 14048
rect 4579 14048 4637 14049
rect 3435 13999 3477 14008
rect 4195 14031 4253 14032
rect 4195 13991 4204 14031
rect 4244 13991 4253 14031
rect 4579 14008 4588 14048
rect 4628 14008 4637 14048
rect 4579 14007 4637 14008
rect 4683 14048 4725 14057
rect 4683 14008 4684 14048
rect 4724 14008 4725 14048
rect 4683 13999 4725 14008
rect 4867 14048 4925 14049
rect 4867 14008 4876 14048
rect 4916 14008 4925 14048
rect 4867 14007 4925 14008
rect 5067 14048 5109 14057
rect 5067 14008 5068 14048
rect 5108 14008 5109 14048
rect 5067 13999 5109 14008
rect 5163 14048 5205 14057
rect 5163 14008 5164 14048
rect 5204 14008 5205 14048
rect 5163 13999 5205 14008
rect 5355 14048 5397 14057
rect 5355 14008 5356 14048
rect 5396 14008 5397 14048
rect 5355 13999 5397 14008
rect 5547 14048 5589 14057
rect 5547 14008 5548 14048
rect 5588 14008 5589 14048
rect 5547 13999 5589 14008
rect 5739 14048 5781 14057
rect 5739 14008 5740 14048
rect 5780 14008 5781 14048
rect 5739 13999 5781 14008
rect 5835 14048 5877 14057
rect 5835 14008 5836 14048
rect 5876 14008 5877 14048
rect 5835 13999 5877 14008
rect 6019 14048 6077 14049
rect 6019 14008 6028 14048
rect 6068 14008 6077 14048
rect 6019 14007 6077 14008
rect 6123 14048 6165 14057
rect 6123 14008 6124 14048
rect 6164 14008 6165 14048
rect 6123 13999 6165 14008
rect 6307 14048 6365 14049
rect 6307 14008 6316 14048
rect 6356 14008 6365 14048
rect 6307 14007 6365 14008
rect 6691 14048 6749 14049
rect 6691 14008 6700 14048
rect 6740 14008 6749 14048
rect 6691 14007 6749 14008
rect 8035 14048 8093 14049
rect 8035 14008 8044 14048
rect 8084 14008 8093 14048
rect 8035 14007 8093 14008
rect 10915 14048 10973 14049
rect 10915 14008 10924 14048
rect 10964 14008 10973 14048
rect 10915 14007 10973 14008
rect 11779 14048 11837 14049
rect 11779 14008 11788 14048
rect 11828 14008 11837 14048
rect 11779 14007 11837 14008
rect 12171 14048 12213 14057
rect 12171 14008 12172 14048
rect 12212 14008 12213 14048
rect 12171 13999 12213 14008
rect 12459 14048 12501 14057
rect 12459 14008 12460 14048
rect 12500 14008 12501 14048
rect 12459 13999 12501 14008
rect 13123 14048 13181 14049
rect 13123 14008 13132 14048
rect 13172 14008 13181 14048
rect 13123 14007 13181 14008
rect 13795 14048 13853 14049
rect 13795 14008 13804 14048
rect 13844 14008 13853 14048
rect 13795 14007 13853 14008
rect 14755 14048 14813 14049
rect 14755 14008 14764 14048
rect 14804 14008 14813 14048
rect 14755 14007 14813 14008
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 15819 14048 15861 14057
rect 15819 14008 15820 14048
rect 15860 14008 15861 14048
rect 15819 13999 15861 14008
rect 15915 14048 15957 14057
rect 15915 14008 15916 14048
rect 15956 14008 15957 14048
rect 15915 13999 15957 14008
rect 17059 14048 17117 14049
rect 17059 14008 17068 14048
rect 17108 14008 17117 14048
rect 17059 14007 17117 14008
rect 17451 14048 17493 14057
rect 17451 14008 17452 14048
rect 17492 14008 17493 14048
rect 17451 13999 17493 14008
rect 18115 14048 18173 14049
rect 18115 14008 18124 14048
rect 18164 14008 18173 14048
rect 18115 14007 18173 14008
rect 18603 14048 18645 14057
rect 18603 14008 18604 14048
rect 18644 14008 18645 14048
rect 18696 14017 18705 14057
rect 18745 14017 18754 14057
rect 18696 14016 18754 14017
rect 18891 14048 18933 14057
rect 18603 13999 18645 14008
rect 18891 14008 18892 14048
rect 18932 14008 18933 14048
rect 18891 13999 18933 14008
rect 18987 14048 19029 14057
rect 18987 14008 18988 14048
rect 19028 14008 19029 14048
rect 18987 13999 19029 14008
rect 19083 14048 19125 14057
rect 19083 14008 19084 14048
rect 19124 14008 19125 14048
rect 19083 13999 19125 14008
rect 19179 14048 19221 14057
rect 19179 14008 19180 14048
rect 19220 14008 19221 14048
rect 19179 13999 19221 14008
rect 19651 14048 19709 14049
rect 19651 14008 19660 14048
rect 19700 14008 19709 14048
rect 19651 14007 19709 14008
rect 19947 14048 19989 14057
rect 19947 14008 19948 14048
rect 19988 14008 19989 14048
rect 19947 13999 19989 14008
rect 20611 14048 20669 14049
rect 20611 14008 20620 14048
rect 20660 14008 20669 14048
rect 20611 14007 20669 14008
rect 20707 14048 20765 14049
rect 20707 14008 20716 14048
rect 20756 14008 20765 14048
rect 20707 14007 20765 14008
rect 20907 14048 20949 14057
rect 20907 14008 20908 14048
rect 20948 14008 20949 14048
rect 20907 13999 20949 14008
rect 21003 14048 21045 14057
rect 21003 14008 21004 14048
rect 21044 14008 21045 14048
rect 21003 13999 21045 14008
rect 21096 14048 21154 14049
rect 21096 14008 21105 14048
rect 21145 14008 21154 14048
rect 21096 14007 21154 14008
rect 21387 14048 21429 14057
rect 21387 14008 21388 14048
rect 21428 14008 21429 14048
rect 21387 13999 21429 14008
rect 21763 14048 21821 14049
rect 21763 14008 21772 14048
rect 21812 14008 21821 14048
rect 21763 14007 21821 14008
rect 21963 14048 22005 14057
rect 21963 14008 21964 14048
rect 22004 14008 22005 14048
rect 21963 13999 22005 14008
rect 22635 14048 22677 14057
rect 22635 14008 22636 14048
rect 22676 14008 22677 14048
rect 22635 13999 22677 14008
rect 24259 14048 24317 14049
rect 24259 14008 24268 14048
rect 24308 14008 24317 14048
rect 24259 14007 24317 14008
rect 26475 14048 26517 14057
rect 26475 14008 26476 14048
rect 26516 14008 26517 14048
rect 26475 13999 26517 14008
rect 27531 14048 27573 14057
rect 27531 14008 27532 14048
rect 27572 14008 27573 14048
rect 27531 13999 27573 14008
rect 27811 14048 27869 14049
rect 27811 14008 27820 14048
rect 27860 14008 27869 14048
rect 27811 14007 27869 14008
rect 28203 14048 28245 14057
rect 28203 14008 28204 14048
rect 28244 14008 28245 14048
rect 28203 13999 28245 14008
rect 28299 14048 28341 14057
rect 28299 14008 28300 14048
rect 28340 14008 28341 14048
rect 28299 13999 28341 14008
rect 28395 14048 28437 14057
rect 28395 14008 28396 14048
rect 28436 14008 28437 14048
rect 28395 13999 28437 14008
rect 28491 14048 28533 14057
rect 28491 14008 28492 14048
rect 28532 14008 28533 14048
rect 28491 13999 28533 14008
rect 30219 14048 30261 14057
rect 30219 14008 30220 14048
rect 30260 14008 30261 14048
rect 30219 13999 30261 14008
rect 30315 14048 30357 14057
rect 30315 14008 30316 14048
rect 30356 14008 30357 14048
rect 30315 13999 30357 14008
rect 30411 14048 30453 14057
rect 30411 14008 30412 14048
rect 30452 14008 30453 14048
rect 30411 13999 30453 14008
rect 30507 14048 30549 14057
rect 30507 14008 30508 14048
rect 30548 14008 30549 14048
rect 30507 13999 30549 14008
rect 31755 14048 31797 14057
rect 31755 14008 31756 14048
rect 31796 14008 31797 14048
rect 31939 14029 31948 14069
rect 31988 14029 31997 14069
rect 31939 14028 31997 14029
rect 32131 14048 32189 14049
rect 31755 13999 31797 14008
rect 32131 14008 32140 14048
rect 32180 14008 32189 14048
rect 32131 14007 32189 14008
rect 32523 14048 32565 14057
rect 32523 14008 32524 14048
rect 32564 14008 32565 14048
rect 32523 13999 32565 14008
rect 32707 14048 32765 14049
rect 32707 14008 32716 14048
rect 32756 14008 32765 14048
rect 32707 14007 32765 14008
rect 33099 14048 33141 14057
rect 33099 14008 33100 14048
rect 33140 14008 33141 14048
rect 33099 13999 33141 14008
rect 33291 14048 33333 14057
rect 33291 14008 33292 14048
rect 33332 14008 33333 14048
rect 33291 13999 33333 14008
rect 33667 14048 33725 14049
rect 33667 14008 33676 14048
rect 33716 14008 33725 14048
rect 33667 14007 33725 14008
rect 33867 14048 33909 14057
rect 33867 14008 33868 14048
rect 33908 14008 33909 14048
rect 33867 13999 33909 14008
rect 34155 14048 34197 14057
rect 34155 14008 34156 14048
rect 34196 14008 34197 14048
rect 34155 13999 34197 14008
rect 34923 14048 34965 14057
rect 34923 14008 34924 14048
rect 34964 14008 34965 14048
rect 34923 13999 34965 14008
rect 35019 14048 35061 14057
rect 35019 14008 35020 14048
rect 35060 14008 35061 14048
rect 35019 13999 35061 14008
rect 35403 14048 35445 14057
rect 35403 14008 35404 14048
rect 35444 14008 35445 14048
rect 35403 13999 35445 14008
rect 35691 14048 35733 14057
rect 35691 14008 35692 14048
rect 35732 14008 35733 14048
rect 35691 13999 35733 14008
rect 35883 14048 35925 14057
rect 35883 14008 35884 14048
rect 35924 14008 35925 14048
rect 35883 13999 35925 14008
rect 35979 14048 36021 14057
rect 35979 14008 35980 14048
rect 36020 14008 36021 14048
rect 35979 13999 36021 14008
rect 36363 14048 36405 14057
rect 36363 14008 36364 14048
rect 36404 14008 36405 14048
rect 36363 13999 36405 14008
rect 36555 14048 36597 14057
rect 36555 14008 36556 14048
rect 36596 14008 36597 14048
rect 36555 13999 36597 14008
rect 36643 14048 36701 14049
rect 36643 14008 36652 14048
rect 36692 14008 36701 14048
rect 36643 14007 36701 14008
rect 36843 14048 36885 14057
rect 36843 14008 36844 14048
rect 36884 14008 36885 14048
rect 36843 13999 36885 14008
rect 36939 14048 36981 14057
rect 36939 14008 36940 14048
rect 36980 14008 36981 14048
rect 36939 13999 36981 14008
rect 37323 14048 37365 14057
rect 37323 14008 37324 14048
rect 37364 14008 37365 14048
rect 37323 13999 37365 14008
rect 37611 14048 37653 14057
rect 37611 14008 37612 14048
rect 37652 14008 37653 14048
rect 37611 13999 37653 14008
rect 37995 14048 38037 14057
rect 37995 14008 37996 14048
rect 38036 14008 38037 14048
rect 37995 13999 38037 14008
rect 38851 14048 38909 14049
rect 38851 14008 38860 14048
rect 38900 14008 38909 14048
rect 38851 14007 38909 14008
rect 40683 14048 40725 14057
rect 40683 14008 40684 14048
rect 40724 14008 40725 14048
rect 40683 13999 40725 14008
rect 41539 14048 41597 14049
rect 41539 14008 41548 14048
rect 41588 14008 41597 14048
rect 41539 14007 41597 14008
rect 41923 14048 41981 14049
rect 41923 14008 41932 14048
rect 41972 14008 41981 14048
rect 41923 14007 41981 14008
rect 42499 14048 42557 14049
rect 42499 14008 42508 14048
rect 42548 14008 42557 14048
rect 42499 14007 42557 14008
rect 43459 14048 43517 14049
rect 43459 14008 43468 14048
rect 43508 14008 43517 14048
rect 43459 14007 43517 14008
rect 44139 14048 44181 14057
rect 44139 14008 44140 14048
rect 44180 14008 44181 14048
rect 44139 13999 44181 14008
rect 44515 14048 44573 14049
rect 44515 14008 44524 14048
rect 44564 14008 44573 14048
rect 44515 14007 44573 14008
rect 45379 14048 45437 14049
rect 45379 14008 45388 14048
rect 45428 14008 45437 14048
rect 45379 14007 45437 14008
rect 46627 14048 46685 14049
rect 46627 14008 46636 14048
rect 46676 14008 46685 14048
rect 46627 14007 46685 14008
rect 4195 13990 4253 13991
rect 17643 13964 17685 13973
rect 17643 13924 17644 13964
rect 17684 13924 17685 13964
rect 17643 13915 17685 13924
rect 21483 13964 21525 13973
rect 21483 13924 21484 13964
rect 21524 13924 21525 13964
rect 21483 13915 21525 13924
rect 21675 13964 21717 13973
rect 21675 13924 21676 13964
rect 21716 13924 21717 13964
rect 21675 13915 21717 13924
rect 32235 13964 32277 13973
rect 32235 13924 32236 13964
rect 32276 13924 32277 13964
rect 32235 13915 32277 13924
rect 32427 13964 32469 13973
rect 32427 13924 32428 13964
rect 32468 13924 32469 13964
rect 32427 13915 32469 13924
rect 32811 13962 32853 13971
rect 32811 13922 32812 13962
rect 32852 13922 32853 13962
rect 32811 13913 32853 13922
rect 33003 13964 33045 13973
rect 33003 13924 33004 13964
rect 33044 13924 33045 13964
rect 33003 13915 33045 13924
rect 33387 13964 33429 13973
rect 33387 13924 33388 13964
rect 33428 13924 33429 13964
rect 33387 13915 33429 13924
rect 33579 13964 33621 13973
rect 33579 13924 33580 13964
rect 33620 13924 33621 13964
rect 33579 13915 33621 13924
rect 34059 13964 34101 13973
rect 34059 13924 34060 13964
rect 34100 13924 34101 13964
rect 34059 13915 34101 13924
rect 3819 13880 3861 13889
rect 3819 13840 3820 13880
rect 3860 13840 3861 13880
rect 3819 13831 3861 13840
rect 4875 13880 4917 13889
rect 4875 13840 4876 13880
rect 4916 13840 4917 13880
rect 4875 13831 4917 13840
rect 5059 13880 5117 13881
rect 5059 13840 5068 13880
rect 5108 13840 5117 13880
rect 5059 13839 5117 13840
rect 7371 13880 7413 13889
rect 7371 13840 7372 13880
rect 7412 13840 7413 13880
rect 7371 13831 7413 13840
rect 8811 13880 8853 13889
rect 8811 13840 8812 13880
rect 8852 13840 8853 13880
rect 8811 13831 8853 13840
rect 14091 13880 14133 13889
rect 14091 13840 14092 13880
rect 14132 13840 14133 13880
rect 14091 13831 14133 13840
rect 15147 13880 15189 13889
rect 15147 13840 15148 13880
rect 15188 13840 15189 13880
rect 15147 13831 15189 13840
rect 17547 13880 17589 13889
rect 17547 13840 17548 13880
rect 17588 13840 17589 13880
rect 17547 13831 17589 13840
rect 21579 13880 21621 13889
rect 21579 13840 21580 13880
rect 21620 13840 21621 13880
rect 21579 13831 21621 13840
rect 24555 13880 24597 13889
rect 24555 13840 24556 13880
rect 24596 13840 24597 13880
rect 24555 13831 24597 13840
rect 24939 13880 24981 13889
rect 24939 13840 24940 13880
rect 24980 13840 24981 13880
rect 24939 13831 24981 13840
rect 27139 13880 27197 13881
rect 27139 13840 27148 13880
rect 27188 13840 27197 13880
rect 27139 13839 27197 13840
rect 32331 13880 32373 13889
rect 32331 13840 32332 13880
rect 32372 13840 32373 13880
rect 32331 13831 32373 13840
rect 32907 13880 32949 13889
rect 32907 13840 32908 13880
rect 32948 13840 32949 13880
rect 32907 13831 32949 13840
rect 33483 13880 33525 13889
rect 33483 13840 33484 13880
rect 33524 13840 33525 13880
rect 33483 13831 33525 13840
rect 35691 13880 35733 13889
rect 35691 13840 35692 13880
rect 35732 13840 35733 13880
rect 35691 13831 35733 13840
rect 39531 13880 39573 13889
rect 39531 13840 39532 13880
rect 39572 13840 39573 13880
rect 39531 13831 39573 13840
rect 3435 13796 3477 13805
rect 3435 13756 3436 13796
rect 3476 13756 3477 13796
rect 3435 13747 3477 13756
rect 14475 13796 14517 13805
rect 14475 13756 14476 13796
rect 14516 13756 14517 13796
rect 14475 13747 14517 13756
rect 16867 13796 16925 13797
rect 16867 13756 16876 13796
rect 16916 13756 16925 13796
rect 16867 13755 16925 13756
rect 18219 13796 18261 13805
rect 18219 13756 18220 13796
rect 18260 13756 18261 13796
rect 18219 13747 18261 13756
rect 20323 13796 20381 13797
rect 20323 13756 20332 13796
rect 20372 13756 20381 13796
rect 20323 13755 20381 13756
rect 25899 13796 25941 13805
rect 25899 13756 25900 13796
rect 25940 13756 25941 13796
rect 25899 13747 25941 13756
rect 31851 13796 31893 13805
rect 31851 13756 31852 13796
rect 31892 13756 31893 13796
rect 31851 13747 31893 13756
rect 36363 13796 36405 13805
rect 36363 13756 36364 13796
rect 36404 13756 36405 13796
rect 36363 13747 36405 13756
rect 37611 13796 37653 13805
rect 37611 13756 37612 13796
rect 37652 13756 37653 13796
rect 37611 13747 37653 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 23307 13460 23349 13469
rect 23307 13420 23308 13460
rect 23348 13420 23349 13460
rect 23307 13411 23349 13420
rect 25795 13460 25853 13461
rect 25795 13420 25804 13460
rect 25844 13420 25853 13460
rect 25795 13419 25853 13420
rect 30123 13460 30165 13469
rect 30123 13420 30124 13460
rect 30164 13420 30165 13460
rect 30123 13411 30165 13420
rect 30603 13460 30645 13469
rect 30603 13420 30604 13460
rect 30644 13420 30645 13460
rect 30603 13411 30645 13420
rect 31659 13460 31701 13469
rect 31659 13420 31660 13460
rect 31700 13420 31701 13460
rect 31659 13411 31701 13420
rect 32907 13460 32949 13469
rect 32907 13420 32908 13460
rect 32948 13420 32949 13460
rect 32907 13411 32949 13420
rect 3435 13376 3477 13385
rect 3435 13336 3436 13376
rect 3476 13336 3477 13376
rect 3435 13327 3477 13336
rect 5355 13376 5397 13385
rect 5355 13336 5356 13376
rect 5396 13336 5397 13376
rect 5355 13327 5397 13336
rect 12931 13376 12989 13377
rect 12931 13336 12940 13376
rect 12980 13336 12989 13376
rect 12931 13335 12989 13336
rect 17835 13376 17877 13385
rect 17835 13336 17836 13376
rect 17876 13336 17877 13376
rect 17835 13327 17877 13336
rect 19075 13376 19133 13377
rect 19075 13336 19084 13376
rect 19124 13336 19133 13376
rect 19075 13335 19133 13336
rect 19851 13376 19893 13385
rect 19851 13336 19852 13376
rect 19892 13336 19893 13376
rect 19851 13327 19893 13336
rect 20907 13376 20949 13385
rect 20907 13336 20908 13376
rect 20948 13336 20949 13376
rect 20907 13327 20949 13336
rect 28683 13376 28725 13385
rect 28683 13336 28684 13376
rect 28724 13336 28725 13376
rect 28683 13327 28725 13336
rect 29739 13376 29781 13385
rect 29739 13336 29740 13376
rect 29780 13336 29781 13376
rect 29739 13327 29781 13336
rect 32235 13376 32277 13385
rect 32235 13336 32236 13376
rect 32276 13336 32277 13376
rect 32235 13327 32277 13336
rect 42411 13376 42453 13385
rect 42411 13336 42412 13376
rect 42452 13336 42453 13376
rect 42411 13327 42453 13336
rect 17739 13292 17781 13301
rect 17739 13252 17740 13292
rect 17780 13252 17781 13292
rect 17739 13243 17781 13252
rect 17931 13292 17973 13301
rect 17931 13252 17932 13292
rect 17972 13252 17973 13292
rect 17931 13243 17973 13252
rect 19755 13292 19797 13301
rect 19755 13252 19756 13292
rect 19796 13252 19797 13292
rect 19755 13243 19797 13252
rect 19947 13292 19989 13301
rect 19947 13252 19948 13292
rect 19988 13252 19989 13292
rect 19947 13243 19989 13252
rect 22347 13292 22389 13301
rect 22347 13252 22348 13292
rect 22388 13252 22389 13292
rect 22347 13243 22389 13252
rect 32139 13292 32181 13301
rect 32139 13252 32140 13292
rect 32180 13252 32181 13292
rect 32139 13243 32181 13252
rect 32331 13292 32373 13301
rect 32331 13252 32332 13292
rect 32372 13252 32373 13292
rect 32331 13243 32373 13252
rect 42315 13292 42357 13301
rect 42315 13252 42316 13292
rect 42356 13252 42357 13292
rect 42315 13243 42357 13252
rect 42507 13292 42549 13301
rect 42507 13252 42508 13292
rect 42548 13252 42549 13292
rect 42507 13243 42549 13252
rect 30787 13222 30845 13223
rect 3819 13208 3861 13217
rect 3819 13168 3820 13208
rect 3860 13168 3861 13208
rect 3819 13159 3861 13168
rect 3915 13208 3957 13217
rect 3915 13168 3916 13208
rect 3956 13168 3957 13208
rect 3915 13159 3957 13168
rect 4011 13208 4053 13217
rect 4011 13168 4012 13208
rect 4052 13168 4053 13208
rect 4011 13159 4053 13168
rect 4963 13208 5021 13209
rect 4963 13168 4972 13208
rect 5012 13168 5021 13208
rect 4963 13167 5021 13168
rect 5547 13208 5589 13217
rect 5547 13168 5548 13208
rect 5588 13168 5589 13208
rect 5547 13159 5589 13168
rect 5643 13208 5685 13217
rect 5643 13168 5644 13208
rect 5684 13168 5685 13208
rect 5643 13159 5685 13168
rect 5739 13208 5781 13217
rect 5739 13168 5740 13208
rect 5780 13168 5781 13208
rect 5739 13159 5781 13168
rect 5835 13208 5877 13217
rect 5835 13168 5836 13208
rect 5876 13168 5877 13208
rect 5835 13159 5877 13168
rect 6691 13208 6749 13209
rect 6691 13168 6700 13208
rect 6740 13168 6749 13208
rect 6691 13167 6749 13168
rect 7843 13208 7901 13209
rect 7843 13168 7852 13208
rect 7892 13168 7901 13208
rect 7843 13167 7901 13168
rect 9283 13208 9341 13209
rect 9283 13168 9292 13208
rect 9332 13168 9341 13208
rect 9283 13167 9341 13168
rect 10147 13208 10205 13209
rect 10147 13168 10156 13208
rect 10196 13168 10205 13208
rect 10147 13167 10205 13168
rect 11395 13208 11453 13209
rect 11395 13168 11404 13208
rect 11444 13168 11453 13208
rect 11395 13167 11453 13168
rect 11875 13208 11933 13209
rect 11875 13168 11884 13208
rect 11924 13168 11933 13208
rect 11875 13167 11933 13168
rect 11979 13208 12021 13217
rect 11979 13168 11980 13208
rect 12020 13168 12021 13208
rect 11979 13159 12021 13168
rect 12171 13208 12213 13217
rect 12171 13168 12172 13208
rect 12212 13168 12213 13208
rect 12171 13159 12213 13168
rect 12355 13208 12413 13209
rect 12355 13168 12364 13208
rect 12404 13168 12413 13208
rect 12355 13167 12413 13168
rect 12459 13208 12501 13217
rect 12459 13168 12460 13208
rect 12500 13168 12501 13208
rect 12459 13159 12501 13168
rect 12651 13208 12693 13217
rect 12651 13168 12652 13208
rect 12692 13168 12693 13208
rect 12651 13159 12693 13168
rect 14083 13208 14141 13209
rect 14083 13168 14092 13208
rect 14132 13168 14141 13208
rect 14083 13167 14141 13168
rect 14947 13208 15005 13209
rect 14947 13168 14956 13208
rect 14996 13168 15005 13208
rect 14947 13167 15005 13168
rect 16195 13208 16253 13209
rect 16195 13168 16204 13208
rect 16244 13168 16253 13208
rect 16195 13167 16253 13168
rect 17635 13208 17693 13209
rect 17635 13168 17644 13208
rect 17684 13168 17693 13208
rect 17635 13167 17693 13168
rect 18027 13208 18069 13217
rect 18027 13168 18028 13208
rect 18068 13168 18069 13208
rect 18027 13159 18069 13168
rect 18403 13208 18461 13209
rect 18403 13168 18412 13208
rect 18452 13168 18461 13208
rect 18403 13167 18461 13168
rect 18699 13208 18741 13217
rect 18699 13168 18700 13208
rect 18740 13168 18741 13208
rect 18699 13159 18741 13168
rect 18795 13208 18837 13217
rect 18795 13168 18796 13208
rect 18836 13168 18837 13208
rect 18795 13159 18837 13168
rect 19275 13208 19317 13217
rect 19275 13168 19276 13208
rect 19316 13168 19317 13208
rect 19275 13159 19317 13168
rect 19467 13208 19509 13217
rect 19467 13168 19468 13208
rect 19508 13168 19509 13208
rect 19467 13159 19509 13168
rect 19651 13208 19709 13209
rect 19651 13168 19660 13208
rect 19700 13168 19709 13208
rect 19651 13167 19709 13168
rect 20043 13208 20085 13217
rect 20043 13168 20044 13208
rect 20084 13168 20085 13208
rect 20043 13159 20085 13168
rect 20419 13208 20477 13209
rect 20419 13168 20428 13208
rect 20468 13168 20477 13208
rect 20715 13208 20757 13217
rect 20419 13167 20477 13168
rect 20611 13193 20669 13194
rect 20611 13153 20620 13193
rect 20660 13153 20669 13193
rect 20715 13168 20716 13208
rect 20756 13168 20757 13208
rect 20715 13159 20757 13168
rect 20907 13208 20949 13217
rect 20907 13168 20908 13208
rect 20948 13168 20949 13208
rect 20907 13159 20949 13168
rect 21099 13208 21141 13217
rect 21099 13168 21100 13208
rect 21140 13168 21141 13208
rect 21099 13159 21141 13168
rect 21195 13208 21237 13217
rect 21195 13168 21196 13208
rect 21236 13168 21237 13208
rect 21195 13159 21237 13168
rect 21291 13208 21333 13217
rect 21291 13168 21292 13208
rect 21332 13168 21333 13208
rect 21291 13159 21333 13168
rect 21571 13208 21629 13209
rect 21571 13168 21580 13208
rect 21620 13168 21629 13208
rect 21571 13167 21629 13168
rect 21771 13208 21813 13217
rect 21771 13168 21772 13208
rect 21812 13168 21813 13208
rect 21771 13159 21813 13168
rect 22251 13208 22293 13217
rect 22251 13168 22252 13208
rect 22292 13168 22293 13208
rect 22251 13159 22293 13168
rect 22443 13208 22485 13217
rect 22443 13168 22444 13208
rect 22484 13168 22485 13208
rect 22443 13159 22485 13168
rect 22723 13208 22781 13209
rect 22723 13168 22732 13208
rect 22772 13168 22781 13208
rect 22723 13167 22781 13168
rect 23307 13208 23349 13217
rect 23307 13168 23308 13208
rect 23348 13168 23349 13208
rect 23307 13159 23349 13168
rect 23499 13208 23541 13217
rect 23499 13168 23500 13208
rect 23540 13168 23541 13208
rect 23499 13159 23541 13168
rect 24643 13208 24701 13209
rect 24643 13168 24652 13208
rect 24692 13168 24701 13208
rect 24643 13167 24701 13168
rect 25603 13208 25661 13209
rect 25603 13168 25612 13208
rect 25652 13168 25661 13208
rect 25603 13167 25661 13168
rect 26187 13208 26229 13217
rect 26187 13168 26188 13208
rect 26228 13168 26229 13208
rect 26187 13159 26229 13168
rect 26467 13208 26525 13209
rect 26467 13168 26476 13208
rect 26516 13168 26525 13208
rect 26467 13167 26525 13168
rect 26755 13208 26813 13209
rect 26755 13168 26764 13208
rect 26804 13168 26813 13208
rect 26755 13167 26813 13168
rect 26947 13208 27005 13209
rect 26947 13168 26956 13208
rect 26996 13168 27005 13208
rect 26947 13167 27005 13168
rect 27723 13208 27765 13217
rect 27723 13168 27724 13208
rect 27764 13168 27765 13208
rect 27723 13159 27765 13168
rect 27819 13208 27861 13217
rect 27819 13168 27820 13208
rect 27860 13168 27861 13208
rect 27819 13159 27861 13168
rect 27915 13208 27957 13217
rect 27915 13168 27916 13208
rect 27956 13168 27957 13208
rect 27915 13159 27957 13168
rect 28011 13208 28053 13217
rect 28011 13168 28012 13208
rect 28052 13168 28053 13208
rect 28011 13159 28053 13168
rect 28291 13208 28349 13209
rect 28291 13168 28300 13208
rect 28340 13168 28349 13208
rect 28291 13167 28349 13168
rect 28395 13208 28437 13217
rect 28395 13168 28396 13208
rect 28436 13168 28437 13208
rect 28395 13159 28437 13168
rect 29067 13208 29109 13217
rect 29067 13168 29068 13208
rect 29108 13168 29109 13208
rect 29067 13159 29109 13168
rect 29163 13208 29205 13217
rect 29163 13168 29164 13208
rect 29204 13168 29205 13208
rect 29163 13159 29205 13168
rect 29259 13208 29301 13217
rect 29259 13168 29260 13208
rect 29300 13168 29301 13208
rect 29259 13159 29301 13168
rect 29355 13208 29397 13217
rect 29355 13168 29356 13208
rect 29396 13168 29397 13208
rect 29355 13159 29397 13168
rect 29739 13208 29781 13217
rect 29739 13168 29740 13208
rect 29780 13168 29781 13208
rect 29739 13159 29781 13168
rect 30296 13208 30354 13209
rect 30296 13168 30305 13208
rect 30345 13168 30354 13208
rect 30296 13167 30354 13168
rect 30411 13208 30453 13217
rect 30411 13168 30412 13208
rect 30452 13168 30453 13208
rect 30411 13159 30453 13168
rect 30603 13208 30645 13217
rect 30603 13168 30604 13208
rect 30644 13168 30645 13208
rect 30787 13182 30796 13222
rect 30836 13182 30845 13222
rect 30787 13181 30845 13182
rect 30883 13208 30941 13209
rect 30603 13159 30645 13168
rect 30883 13168 30892 13208
rect 30932 13168 30941 13208
rect 30883 13167 30941 13168
rect 31555 13208 31613 13209
rect 31555 13168 31564 13208
rect 31604 13168 31613 13208
rect 31555 13167 31613 13168
rect 31755 13208 31797 13217
rect 31755 13168 31756 13208
rect 31796 13168 31797 13208
rect 31755 13159 31797 13168
rect 32043 13208 32085 13217
rect 32043 13168 32044 13208
rect 32084 13168 32085 13208
rect 32043 13159 32085 13168
rect 32419 13208 32477 13209
rect 32419 13168 32428 13208
rect 32468 13168 32477 13208
rect 32419 13167 32477 13168
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 32995 13208 33053 13209
rect 32995 13168 33004 13208
rect 33044 13168 33053 13208
rect 32995 13167 33053 13168
rect 33579 13208 33621 13217
rect 33579 13168 33580 13208
rect 33620 13168 33621 13208
rect 33579 13159 33621 13168
rect 33675 13208 33717 13217
rect 33675 13168 33676 13208
rect 33716 13168 33717 13208
rect 33675 13159 33717 13168
rect 34059 13208 34101 13217
rect 34059 13168 34060 13208
rect 34100 13168 34101 13208
rect 34059 13159 34101 13168
rect 34347 13208 34389 13217
rect 34347 13168 34348 13208
rect 34388 13168 34389 13208
rect 34347 13159 34389 13168
rect 34923 13208 34965 13217
rect 34923 13168 34924 13208
rect 34964 13168 34965 13208
rect 34923 13159 34965 13168
rect 35019 13208 35061 13217
rect 35019 13168 35020 13208
rect 35060 13168 35061 13208
rect 35019 13159 35061 13168
rect 35395 13208 35453 13209
rect 35395 13168 35404 13208
rect 35444 13168 35453 13208
rect 35395 13167 35453 13168
rect 35491 13208 35549 13209
rect 35491 13168 35500 13208
rect 35540 13168 35549 13208
rect 35491 13167 35549 13168
rect 35691 13208 35733 13217
rect 35691 13168 35692 13208
rect 35732 13168 35733 13208
rect 35691 13159 35733 13168
rect 35787 13208 35829 13217
rect 35787 13168 35788 13208
rect 35828 13168 35829 13208
rect 35787 13159 35829 13168
rect 35880 13208 35938 13209
rect 35880 13168 35889 13208
rect 35929 13168 35938 13208
rect 35880 13167 35938 13168
rect 36171 13208 36213 13217
rect 36171 13168 36172 13208
rect 36212 13168 36213 13208
rect 36171 13159 36213 13168
rect 36459 13208 36501 13217
rect 36459 13168 36460 13208
rect 36500 13168 36501 13208
rect 36459 13159 36501 13168
rect 37323 13208 37365 13217
rect 37323 13168 37324 13208
rect 37364 13168 37365 13208
rect 37323 13159 37365 13168
rect 37419 13208 37461 13217
rect 37419 13168 37420 13208
rect 37460 13168 37461 13208
rect 37419 13159 37461 13168
rect 37515 13208 37557 13217
rect 37515 13168 37516 13208
rect 37556 13168 37557 13208
rect 37515 13159 37557 13168
rect 37611 13208 37653 13217
rect 37611 13168 37612 13208
rect 37652 13168 37653 13208
rect 37611 13159 37653 13168
rect 37795 13208 37853 13209
rect 37795 13168 37804 13208
rect 37844 13168 37853 13208
rect 37795 13167 37853 13168
rect 38755 13208 38813 13209
rect 38755 13168 38764 13208
rect 38804 13168 38813 13208
rect 38755 13167 38813 13168
rect 39051 13208 39093 13217
rect 39051 13168 39052 13208
rect 39092 13168 39093 13208
rect 39051 13159 39093 13168
rect 39427 13208 39485 13209
rect 39427 13168 39436 13208
rect 39476 13168 39485 13208
rect 39427 13167 39485 13168
rect 40291 13208 40349 13209
rect 40291 13168 40300 13208
rect 40340 13168 40349 13208
rect 40291 13167 40349 13168
rect 41451 13208 41493 13217
rect 41451 13168 41452 13208
rect 41492 13168 41493 13208
rect 41451 13159 41493 13168
rect 41731 13208 41789 13209
rect 41731 13168 41740 13208
rect 41780 13168 41789 13208
rect 41731 13167 41789 13168
rect 41931 13208 41973 13217
rect 41931 13168 41932 13208
rect 41972 13168 41973 13208
rect 41931 13159 41973 13168
rect 42019 13208 42077 13209
rect 42019 13168 42028 13208
rect 42068 13168 42077 13208
rect 42019 13167 42077 13168
rect 42211 13208 42269 13209
rect 42211 13168 42220 13208
rect 42260 13168 42269 13208
rect 42211 13167 42269 13168
rect 42603 13208 42645 13217
rect 42603 13168 42604 13208
rect 42644 13168 42645 13208
rect 42603 13159 42645 13168
rect 42787 13208 42845 13209
rect 42787 13168 42796 13208
rect 42836 13168 42845 13208
rect 42787 13167 42845 13168
rect 43075 13208 43133 13209
rect 43075 13168 43084 13208
rect 43124 13168 43133 13208
rect 43075 13167 43133 13168
rect 43555 13208 43613 13209
rect 43555 13168 43564 13208
rect 43604 13168 43613 13208
rect 43555 13167 43613 13168
rect 44427 13208 44469 13217
rect 44427 13168 44428 13208
rect 44468 13168 44469 13208
rect 44427 13159 44469 13168
rect 44803 13208 44861 13209
rect 44803 13168 44812 13208
rect 44852 13168 44861 13208
rect 44803 13167 44861 13168
rect 45667 13208 45725 13209
rect 45667 13168 45676 13208
rect 45716 13168 45725 13208
rect 45667 13167 45725 13168
rect 46827 13208 46869 13217
rect 46827 13168 46828 13208
rect 46868 13168 46869 13208
rect 46827 13159 46869 13168
rect 47107 13208 47165 13209
rect 47107 13168 47116 13208
rect 47156 13168 47165 13208
rect 47107 13167 47165 13168
rect 47307 13208 47349 13217
rect 47307 13168 47308 13208
rect 47348 13168 47349 13208
rect 47307 13159 47349 13168
rect 47395 13208 47453 13209
rect 47395 13168 47404 13208
rect 47444 13168 47453 13208
rect 47395 13167 47453 13168
rect 20611 13152 20669 13153
rect 10539 13124 10581 13133
rect 10539 13084 10540 13124
rect 10580 13084 10581 13124
rect 10539 13075 10581 13084
rect 10731 13124 10773 13133
rect 10731 13084 10732 13124
rect 10772 13084 10773 13124
rect 10731 13075 10773 13084
rect 12555 13124 12597 13133
rect 12555 13084 12556 13124
rect 12596 13084 12597 13124
rect 12555 13075 12597 13084
rect 15339 13124 15381 13133
rect 15339 13084 15340 13124
rect 15380 13084 15381 13124
rect 15339 13075 15381 13084
rect 21675 13124 21717 13133
rect 21675 13084 21676 13124
rect 21716 13084 21717 13124
rect 21675 13075 21717 13084
rect 22915 13124 22973 13125
rect 22915 13084 22924 13124
rect 22964 13084 22973 13124
rect 22915 13083 22973 13084
rect 26091 13124 26133 13133
rect 26091 13084 26092 13124
rect 26132 13084 26133 13124
rect 26091 13075 26133 13084
rect 30211 13124 30269 13125
rect 30211 13084 30220 13124
rect 30260 13084 30269 13124
rect 30211 13083 30269 13084
rect 36363 13124 36405 13133
rect 36363 13084 36364 13124
rect 36404 13084 36405 13124
rect 36363 13075 36405 13084
rect 43267 13124 43325 13125
rect 43267 13084 43276 13124
rect 43316 13084 43325 13124
rect 43267 13083 43325 13084
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 4099 13040 4157 13041
rect 4099 13000 4108 13040
rect 4148 13000 4157 13040
rect 4099 12999 4157 13000
rect 4291 13040 4349 13041
rect 4291 13000 4300 13040
rect 4340 13000 4349 13040
rect 4291 12999 4349 13000
rect 6019 13040 6077 13041
rect 6019 13000 6028 13040
rect 6068 13000 6077 13040
rect 6019 12999 6077 13000
rect 7371 13040 7413 13049
rect 7371 13000 7372 13040
rect 7412 13000 7413 13040
rect 7371 12991 7413 13000
rect 8131 13040 8189 13041
rect 8131 13000 8140 13040
rect 8180 13000 8189 13040
rect 8131 12999 8189 13000
rect 12067 13040 12125 13041
rect 12067 13000 12076 13040
rect 12116 13000 12125 13040
rect 12067 12999 12125 13000
rect 15523 13040 15581 13041
rect 15523 13000 15532 13040
rect 15572 13000 15581 13040
rect 15523 12999 15581 13000
rect 19371 13040 19413 13049
rect 19371 13000 19372 13040
rect 19412 13000 19413 13040
rect 19371 12991 19413 13000
rect 20331 13040 20373 13049
rect 20331 13000 20332 13040
rect 20372 13000 20373 13040
rect 20331 12991 20373 13000
rect 21379 13040 21437 13041
rect 21379 13000 21388 13040
rect 21428 13000 21437 13040
rect 21379 12999 21437 13000
rect 22627 13040 22685 13041
rect 22627 13000 22636 13040
rect 22676 13000 22685 13040
rect 22627 12999 22685 13000
rect 29547 13040 29589 13049
rect 29547 13000 29548 13040
rect 29588 13000 29589 13040
rect 29547 12991 29589 13000
rect 30115 13040 30173 13041
rect 30115 13000 30124 13040
rect 30164 13000 30173 13040
rect 30115 12999 30173 13000
rect 33859 13040 33917 13041
rect 33859 13000 33868 13040
rect 33908 13000 33917 13040
rect 33859 12999 33917 13000
rect 34155 13040 34197 13049
rect 34155 13000 34156 13040
rect 34196 13000 34197 13040
rect 34155 12991 34197 13000
rect 35203 13040 35261 13041
rect 35203 13000 35212 13040
rect 35252 13000 35261 13040
rect 35203 12999 35261 13000
rect 35779 13040 35837 13041
rect 35779 13000 35788 13040
rect 35828 13000 35837 13040
rect 35779 12999 35837 13000
rect 41739 13040 41781 13049
rect 41739 13000 41740 13040
rect 41780 13000 41781 13040
rect 41739 12991 41781 13000
rect 44227 13040 44285 13041
rect 44227 13000 44236 13040
rect 44276 13000 44285 13040
rect 44227 12999 44285 13000
rect 47115 13040 47157 13049
rect 47115 13000 47116 13040
rect 47156 13000 47157 13040
rect 47115 12991 47157 13000
rect 28203 12982 28245 12991
rect 28203 12942 28204 12982
rect 28244 12942 28245 12982
rect 28203 12933 28245 12942
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 8803 12704 8861 12705
rect 8803 12664 8812 12704
rect 8852 12664 8861 12704
rect 8803 12663 8861 12664
rect 27531 12704 27573 12713
rect 27531 12664 27532 12704
rect 27572 12664 27573 12704
rect 27531 12655 27573 12664
rect 27811 12704 27869 12705
rect 27811 12664 27820 12704
rect 27860 12664 27869 12704
rect 27811 12663 27869 12664
rect 28483 12704 28541 12705
rect 28483 12664 28492 12704
rect 28532 12664 28541 12704
rect 28483 12663 28541 12664
rect 31843 12704 31901 12705
rect 31843 12664 31852 12704
rect 31892 12664 31901 12704
rect 31843 12663 31901 12664
rect 35403 12704 35445 12713
rect 35403 12664 35404 12704
rect 35444 12664 35445 12704
rect 35403 12655 35445 12664
rect 37987 12704 38045 12705
rect 37987 12664 37996 12704
rect 38036 12664 38045 12704
rect 37987 12663 38045 12664
rect 38467 12704 38525 12705
rect 38467 12664 38476 12704
rect 38516 12664 38525 12704
rect 38467 12663 38525 12664
rect 42115 12704 42173 12705
rect 42115 12664 42124 12704
rect 42164 12664 42173 12704
rect 42115 12663 42173 12664
rect 10539 12620 10581 12629
rect 10539 12580 10540 12620
rect 10580 12580 10581 12620
rect 10539 12571 10581 12580
rect 13611 12620 13653 12629
rect 13611 12580 13612 12620
rect 13652 12580 13653 12620
rect 13611 12571 13653 12580
rect 16683 12620 16725 12629
rect 16683 12580 16684 12620
rect 16724 12580 16725 12620
rect 16683 12571 16725 12580
rect 28971 12620 29013 12629
rect 28971 12580 28972 12620
rect 29012 12580 29013 12620
rect 17355 12563 17397 12572
rect 28971 12571 29013 12580
rect 32427 12620 32469 12629
rect 32427 12580 32428 12620
rect 32468 12580 32469 12620
rect 32427 12571 32469 12580
rect 40683 12620 40725 12629
rect 40683 12580 40684 12620
rect 40724 12580 40725 12620
rect 40683 12571 40725 12580
rect 42019 12620 42077 12621
rect 42019 12580 42028 12620
rect 42068 12580 42077 12620
rect 42019 12579 42077 12580
rect 43851 12620 43893 12629
rect 43851 12580 43852 12620
rect 43892 12580 43893 12620
rect 43851 12571 43893 12580
rect 2955 12536 2997 12545
rect 2955 12496 2956 12536
rect 2996 12496 2997 12536
rect 2955 12487 2997 12496
rect 3331 12536 3389 12537
rect 3331 12496 3340 12536
rect 3380 12496 3389 12536
rect 3331 12495 3389 12496
rect 4195 12536 4253 12537
rect 4195 12496 4204 12536
rect 4244 12496 4253 12536
rect 4195 12495 4253 12496
rect 5443 12536 5501 12537
rect 5443 12496 5452 12536
rect 5492 12496 5501 12536
rect 5443 12495 5501 12496
rect 5643 12536 5685 12545
rect 5643 12496 5644 12536
rect 5684 12496 5685 12536
rect 5643 12487 5685 12496
rect 6019 12536 6077 12537
rect 6019 12496 6028 12536
rect 6068 12496 6077 12536
rect 6019 12495 6077 12496
rect 6883 12536 6941 12537
rect 6883 12496 6892 12536
rect 6932 12496 6941 12536
rect 6883 12495 6941 12496
rect 8043 12536 8085 12545
rect 8043 12496 8044 12536
rect 8084 12496 8085 12536
rect 8043 12487 8085 12496
rect 8523 12536 8565 12545
rect 8523 12496 8524 12536
rect 8564 12496 8565 12536
rect 8523 12487 8565 12496
rect 8619 12536 8661 12545
rect 8619 12496 8620 12536
rect 8660 12496 8661 12536
rect 8619 12487 8661 12496
rect 8995 12536 9053 12537
rect 8995 12496 9004 12536
rect 9044 12496 9053 12536
rect 8995 12495 9053 12496
rect 9675 12536 9717 12545
rect 9675 12496 9676 12536
rect 9716 12496 9717 12536
rect 9675 12487 9717 12496
rect 9859 12536 9917 12537
rect 9859 12496 9868 12536
rect 9908 12496 9917 12536
rect 9859 12495 9917 12496
rect 10723 12536 10781 12537
rect 10723 12496 10732 12536
rect 10772 12496 10781 12536
rect 10723 12495 10781 12496
rect 11115 12536 11157 12545
rect 11115 12496 11116 12536
rect 11156 12496 11157 12536
rect 11115 12487 11157 12496
rect 11211 12536 11253 12545
rect 11211 12496 11212 12536
rect 11252 12496 11253 12536
rect 11211 12487 11253 12496
rect 11307 12536 11349 12545
rect 11307 12496 11308 12536
rect 11348 12496 11349 12536
rect 11307 12487 11349 12496
rect 11403 12536 11445 12545
rect 11403 12496 11404 12536
rect 11444 12496 11445 12536
rect 11403 12487 11445 12496
rect 11683 12536 11741 12537
rect 11683 12496 11692 12536
rect 11732 12496 11741 12536
rect 11683 12495 11741 12496
rect 12931 12536 12989 12537
rect 12931 12496 12940 12536
rect 12980 12496 12989 12536
rect 12931 12495 12989 12496
rect 14859 12536 14901 12545
rect 14859 12496 14860 12536
rect 14900 12496 14901 12536
rect 14859 12487 14901 12496
rect 16587 12536 16629 12545
rect 16587 12496 16588 12536
rect 16628 12496 16629 12536
rect 16587 12487 16629 12496
rect 16779 12536 16821 12545
rect 16779 12496 16780 12536
rect 16820 12496 16821 12536
rect 16779 12487 16821 12496
rect 17059 12536 17117 12537
rect 17059 12496 17068 12536
rect 17108 12496 17117 12536
rect 17355 12523 17356 12563
rect 17396 12523 17397 12563
rect 17355 12514 17397 12523
rect 17451 12536 17493 12545
rect 17059 12495 17117 12496
rect 17451 12496 17452 12536
rect 17492 12496 17493 12536
rect 17451 12487 17493 12496
rect 17923 12536 17981 12537
rect 17923 12496 17932 12536
rect 17972 12496 17981 12536
rect 17923 12495 17981 12496
rect 18315 12536 18357 12545
rect 18315 12496 18316 12536
rect 18356 12496 18357 12536
rect 18315 12487 18357 12496
rect 18507 12536 18549 12545
rect 18507 12496 18508 12536
rect 18548 12496 18549 12536
rect 18507 12487 18549 12496
rect 18603 12536 18645 12545
rect 18603 12496 18604 12536
rect 18644 12496 18645 12536
rect 18603 12487 18645 12496
rect 18699 12536 18741 12545
rect 18699 12496 18700 12536
rect 18740 12496 18741 12536
rect 18699 12487 18741 12496
rect 18795 12536 18837 12545
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 18795 12487 18837 12496
rect 19171 12536 19229 12537
rect 19171 12496 19180 12536
rect 19220 12496 19229 12536
rect 19171 12495 19229 12496
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19939 12536 19997 12537
rect 19939 12496 19948 12536
rect 19988 12496 19997 12536
rect 19939 12495 19997 12496
rect 20043 12536 20085 12545
rect 20043 12496 20044 12536
rect 20084 12496 20085 12536
rect 20043 12487 20085 12496
rect 20235 12536 20277 12545
rect 20235 12496 20236 12536
rect 20276 12496 20277 12536
rect 20235 12487 20277 12496
rect 20419 12536 20477 12537
rect 20419 12496 20428 12536
rect 20468 12496 20477 12536
rect 20419 12495 20477 12496
rect 20515 12536 20573 12537
rect 20515 12496 20524 12536
rect 20564 12496 20573 12536
rect 20515 12495 20573 12496
rect 20715 12536 20757 12545
rect 20715 12496 20716 12536
rect 20756 12496 20757 12536
rect 20715 12487 20757 12496
rect 20811 12536 20853 12545
rect 20811 12496 20812 12536
rect 20852 12496 20853 12536
rect 20811 12487 20853 12496
rect 20904 12536 20962 12537
rect 20904 12496 20913 12536
rect 20953 12496 20962 12536
rect 20904 12495 20962 12496
rect 21195 12536 21237 12545
rect 21195 12496 21196 12536
rect 21236 12496 21237 12536
rect 21195 12487 21237 12496
rect 21387 12536 21429 12545
rect 21387 12496 21388 12536
rect 21428 12496 21429 12536
rect 21387 12487 21429 12496
rect 21475 12536 21533 12537
rect 21475 12496 21484 12536
rect 21524 12496 21533 12536
rect 21475 12495 21533 12496
rect 21675 12536 21717 12545
rect 21675 12496 21676 12536
rect 21716 12496 21717 12536
rect 21675 12487 21717 12496
rect 21763 12536 21821 12537
rect 21763 12496 21772 12536
rect 21812 12496 21821 12536
rect 21763 12495 21821 12496
rect 22251 12536 22293 12545
rect 22251 12496 22252 12536
rect 22292 12496 22293 12536
rect 22251 12487 22293 12496
rect 22347 12536 22389 12545
rect 22347 12496 22348 12536
rect 22388 12496 22389 12536
rect 22347 12487 22389 12496
rect 22627 12536 22685 12537
rect 22627 12496 22636 12536
rect 22676 12496 22685 12536
rect 22627 12495 22685 12496
rect 26275 12536 26333 12537
rect 26275 12496 26284 12536
rect 26324 12496 26333 12536
rect 26275 12495 26333 12496
rect 27235 12536 27293 12537
rect 27235 12496 27244 12536
rect 27284 12496 27293 12536
rect 27235 12495 27293 12496
rect 27331 12536 27389 12537
rect 27331 12496 27340 12536
rect 27380 12496 27389 12536
rect 27331 12495 27389 12496
rect 27915 12536 27957 12545
rect 27915 12496 27916 12536
rect 27956 12496 27957 12536
rect 27915 12487 27957 12496
rect 28011 12536 28053 12545
rect 28011 12496 28012 12536
rect 28052 12496 28053 12536
rect 28011 12487 28053 12496
rect 28107 12536 28149 12545
rect 28107 12496 28108 12536
rect 28148 12496 28149 12536
rect 28107 12487 28149 12496
rect 28291 12536 28349 12537
rect 28291 12496 28300 12536
rect 28340 12496 28349 12536
rect 28291 12495 28349 12496
rect 28395 12536 28437 12545
rect 28395 12496 28396 12536
rect 28436 12496 28437 12536
rect 28395 12487 28437 12496
rect 28587 12536 28629 12545
rect 28587 12496 28588 12536
rect 28628 12496 28629 12536
rect 28587 12487 28629 12496
rect 28771 12536 28829 12537
rect 28771 12496 28780 12536
rect 28820 12496 28829 12536
rect 28771 12495 28829 12496
rect 28875 12536 28917 12545
rect 28875 12496 28876 12536
rect 28916 12496 28917 12536
rect 28875 12487 28917 12496
rect 29067 12536 29109 12545
rect 29067 12496 29068 12536
rect 29108 12496 29109 12536
rect 29067 12487 29109 12496
rect 29259 12536 29301 12545
rect 29259 12496 29260 12536
rect 29300 12496 29301 12536
rect 29259 12487 29301 12496
rect 29451 12536 29493 12545
rect 29451 12496 29452 12536
rect 29492 12496 29493 12536
rect 29451 12487 29493 12496
rect 30403 12536 30461 12537
rect 30403 12496 30412 12536
rect 30452 12496 30461 12536
rect 30403 12495 30461 12496
rect 30795 12536 30837 12545
rect 30795 12496 30796 12536
rect 30836 12496 30837 12536
rect 30795 12487 30837 12496
rect 30979 12536 31037 12537
rect 30979 12496 30988 12536
rect 31028 12496 31037 12536
rect 30979 12495 31037 12496
rect 31371 12536 31413 12545
rect 31371 12496 31372 12536
rect 31412 12496 31413 12536
rect 31371 12487 31413 12496
rect 31555 12536 31613 12537
rect 31555 12496 31564 12536
rect 31604 12496 31613 12536
rect 31555 12495 31613 12496
rect 31651 12536 31709 12537
rect 31651 12496 31660 12536
rect 31700 12496 31709 12536
rect 31651 12495 31709 12496
rect 31851 12536 31893 12545
rect 31851 12496 31852 12536
rect 31892 12496 31893 12536
rect 31851 12487 31893 12496
rect 31947 12536 31989 12545
rect 31947 12496 31948 12536
rect 31988 12496 31989 12536
rect 32331 12536 32373 12545
rect 31947 12487 31989 12496
rect 32104 12521 32146 12530
rect 32104 12481 32105 12521
rect 32145 12481 32146 12521
rect 32331 12496 32332 12536
rect 32372 12496 32373 12536
rect 32331 12487 32373 12496
rect 32515 12536 32573 12537
rect 32515 12496 32524 12536
rect 32564 12496 32573 12536
rect 32515 12495 32573 12496
rect 34051 12536 34109 12537
rect 34051 12496 34060 12536
rect 34100 12496 34109 12536
rect 34051 12495 34109 12496
rect 34147 12536 34205 12537
rect 34147 12496 34156 12536
rect 34196 12496 34205 12536
rect 34147 12495 34205 12496
rect 34347 12536 34389 12545
rect 34347 12496 34348 12536
rect 34388 12496 34389 12536
rect 34347 12487 34389 12496
rect 34443 12536 34485 12545
rect 34443 12496 34444 12536
rect 34484 12496 34485 12536
rect 34443 12487 34485 12496
rect 34590 12536 34648 12537
rect 34590 12496 34599 12536
rect 34639 12496 34648 12536
rect 34590 12495 34648 12496
rect 34827 12536 34869 12545
rect 34827 12496 34828 12536
rect 34868 12496 34869 12536
rect 34827 12487 34869 12496
rect 34915 12536 34973 12537
rect 34915 12496 34924 12536
rect 34964 12496 34973 12536
rect 34915 12495 34973 12496
rect 35307 12536 35349 12545
rect 35307 12496 35308 12536
rect 35348 12496 35349 12536
rect 35307 12487 35349 12496
rect 35595 12536 35637 12545
rect 35595 12496 35596 12536
rect 35636 12496 35637 12536
rect 35595 12487 35637 12496
rect 37035 12536 37077 12545
rect 37035 12496 37036 12536
rect 37076 12496 37077 12536
rect 37035 12487 37077 12496
rect 37227 12536 37269 12545
rect 37227 12496 37228 12536
rect 37268 12496 37269 12536
rect 37227 12487 37269 12496
rect 37315 12536 37373 12537
rect 37315 12496 37324 12536
rect 37364 12496 37373 12536
rect 37315 12495 37373 12496
rect 37515 12536 37557 12545
rect 37515 12496 37516 12536
rect 37556 12496 37557 12536
rect 37515 12487 37557 12496
rect 37803 12536 37845 12545
rect 37803 12496 37804 12536
rect 37844 12496 37845 12536
rect 37803 12487 37845 12496
rect 38187 12536 38229 12545
rect 38187 12496 38188 12536
rect 38228 12496 38229 12536
rect 38187 12487 38229 12496
rect 38283 12536 38325 12545
rect 38283 12496 38284 12536
rect 38324 12496 38325 12536
rect 38283 12487 38325 12496
rect 38667 12536 38709 12545
rect 38667 12496 38668 12536
rect 38708 12496 38709 12536
rect 38667 12487 38709 12496
rect 38763 12536 38805 12545
rect 38763 12496 38764 12536
rect 38804 12496 38805 12536
rect 38763 12487 38805 12496
rect 38955 12536 38997 12545
rect 38955 12496 38956 12536
rect 38996 12496 38997 12536
rect 38955 12487 38997 12496
rect 39243 12536 39285 12545
rect 39243 12496 39244 12536
rect 39284 12496 39285 12536
rect 39243 12487 39285 12496
rect 39627 12536 39669 12545
rect 39627 12496 39628 12536
rect 39668 12496 39669 12536
rect 39627 12487 39669 12496
rect 41347 12536 41405 12537
rect 41347 12496 41356 12536
rect 41396 12496 41405 12536
rect 41347 12495 41405 12496
rect 41835 12536 41877 12545
rect 41835 12496 41836 12536
rect 41876 12496 41877 12536
rect 41835 12487 41877 12496
rect 41931 12536 41973 12545
rect 41931 12496 41932 12536
rect 41972 12496 41973 12536
rect 41931 12487 41973 12496
rect 42603 12536 42645 12545
rect 42603 12496 42604 12536
rect 42644 12496 42645 12536
rect 42603 12487 42645 12496
rect 42691 12536 42749 12537
rect 42691 12496 42700 12536
rect 42740 12496 42749 12536
rect 42691 12495 42749 12496
rect 43171 12536 43229 12537
rect 43171 12496 43180 12536
rect 43220 12496 43229 12536
rect 43171 12495 43229 12496
rect 44043 12536 44085 12545
rect 44043 12496 44044 12536
rect 44084 12496 44085 12536
rect 44043 12487 44085 12496
rect 44419 12536 44477 12537
rect 44419 12496 44428 12536
rect 44468 12496 44477 12536
rect 44419 12495 44477 12496
rect 45283 12536 45341 12537
rect 45283 12496 45292 12536
rect 45332 12496 45341 12536
rect 45283 12495 45341 12496
rect 47587 12536 47645 12537
rect 47587 12496 47596 12536
rect 47636 12496 47645 12536
rect 47587 12495 47645 12496
rect 48643 12536 48701 12537
rect 48643 12496 48652 12536
rect 48692 12496 48701 12536
rect 48643 12495 48701 12496
rect 32104 12472 32146 12481
rect 18027 12452 18069 12461
rect 18027 12412 18028 12452
rect 18068 12412 18069 12452
rect 18027 12403 18069 12412
rect 18219 12452 18261 12461
rect 18219 12412 18220 12452
rect 18260 12412 18261 12452
rect 18219 12403 18261 12412
rect 19275 12452 19317 12461
rect 19275 12412 19276 12452
rect 19316 12412 19317 12452
rect 19275 12403 19317 12412
rect 19467 12452 19509 12461
rect 19467 12412 19468 12452
rect 19508 12412 19509 12452
rect 19467 12403 19509 12412
rect 29355 12452 29397 12461
rect 29355 12412 29356 12452
rect 29396 12412 29397 12452
rect 29355 12403 29397 12412
rect 30507 12452 30549 12461
rect 30507 12412 30508 12452
rect 30548 12412 30549 12452
rect 30507 12403 30549 12412
rect 30699 12452 30741 12461
rect 30699 12412 30700 12452
rect 30740 12412 30741 12452
rect 30699 12403 30741 12412
rect 31083 12452 31125 12461
rect 31083 12412 31084 12452
rect 31124 12412 31125 12452
rect 31083 12403 31125 12412
rect 31275 12452 31317 12461
rect 31275 12412 31276 12452
rect 31316 12412 31317 12452
rect 31275 12403 31317 12412
rect 37611 12452 37653 12461
rect 37611 12412 37612 12452
rect 37652 12412 37653 12452
rect 37611 12403 37653 12412
rect 18123 12368 18165 12377
rect 18123 12328 18124 12368
rect 18164 12328 18165 12368
rect 18123 12319 18165 12328
rect 19371 12368 19413 12377
rect 19371 12328 19372 12368
rect 19412 12328 19413 12368
rect 19371 12319 19413 12328
rect 20235 12368 20277 12377
rect 20235 12328 20236 12368
rect 20276 12328 20277 12368
rect 20235 12319 20277 12328
rect 21955 12368 22013 12369
rect 21955 12328 21964 12368
rect 22004 12328 22013 12368
rect 21955 12327 22013 12328
rect 30603 12368 30645 12377
rect 30603 12328 30604 12368
rect 30644 12328 30645 12368
rect 30603 12319 30645 12328
rect 31179 12368 31221 12377
rect 31179 12328 31180 12368
rect 31220 12328 31221 12368
rect 31179 12319 31221 12328
rect 42123 12368 42165 12377
rect 42123 12328 42124 12368
rect 42164 12328 42165 12368
rect 42123 12319 42165 12328
rect 42891 12368 42933 12377
rect 42891 12328 42892 12368
rect 42932 12328 42933 12368
rect 42891 12319 42933 12328
rect 10827 12284 10869 12293
rect 10827 12244 10828 12284
rect 10868 12244 10869 12284
rect 10827 12235 10869 12244
rect 12363 12284 12405 12293
rect 12363 12244 12364 12284
rect 12404 12244 12405 12284
rect 12363 12235 12405 12244
rect 14667 12284 14709 12293
rect 14667 12244 14668 12284
rect 14708 12244 14709 12284
rect 14667 12235 14709 12244
rect 17731 12284 17789 12285
rect 17731 12244 17740 12284
rect 17780 12244 17789 12284
rect 17731 12243 17789 12244
rect 20427 12284 20469 12293
rect 20427 12244 20428 12284
rect 20468 12244 20469 12284
rect 20427 12235 20469 12244
rect 21195 12284 21237 12293
rect 21195 12244 21196 12284
rect 21236 12244 21237 12284
rect 21195 12235 21237 12244
rect 25611 12284 25653 12293
rect 25611 12244 25612 12284
rect 25652 12244 25653 12284
rect 25611 12235 25653 12244
rect 34059 12284 34101 12293
rect 34059 12244 34060 12284
rect 34100 12244 34101 12284
rect 34059 12235 34101 12244
rect 37035 12284 37077 12293
rect 37035 12244 37036 12284
rect 37076 12244 37077 12284
rect 37035 12235 37077 12244
rect 38955 12284 38997 12293
rect 38955 12244 38956 12284
rect 38996 12244 38997 12284
rect 38955 12235 38997 12244
rect 40203 12284 40245 12293
rect 40203 12244 40204 12284
rect 40244 12244 40245 12284
rect 40203 12235 40245 12244
rect 41931 12284 41973 12293
rect 41931 12244 41932 12284
rect 41972 12244 41973 12284
rect 41931 12235 41973 12244
rect 46443 12284 46485 12293
rect 46443 12244 46444 12284
rect 46484 12244 46485 12284
rect 46443 12235 46485 12244
rect 46915 12284 46973 12285
rect 46915 12244 46924 12284
rect 46964 12244 46973 12284
rect 46915 12243 46973 12244
rect 47971 12284 48029 12285
rect 47971 12244 47980 12284
rect 48020 12244 48029 12284
rect 47971 12243 48029 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 6403 11948 6461 11949
rect 6403 11908 6412 11948
rect 6452 11908 6461 11948
rect 6403 11907 6461 11908
rect 10155 11948 10197 11957
rect 10155 11908 10156 11948
rect 10196 11908 10197 11948
rect 10155 11899 10197 11908
rect 12939 11948 12981 11957
rect 12939 11908 12940 11948
rect 12980 11908 12981 11948
rect 12939 11899 12981 11908
rect 17731 11948 17789 11949
rect 17731 11908 17740 11948
rect 17780 11908 17789 11948
rect 17731 11907 17789 11908
rect 27531 11948 27573 11957
rect 27531 11908 27532 11948
rect 27572 11908 27573 11948
rect 27531 11899 27573 11908
rect 44715 11948 44757 11957
rect 44715 11908 44716 11948
rect 44756 11908 44757 11948
rect 44715 11899 44757 11908
rect 45091 11948 45149 11949
rect 45091 11908 45100 11948
rect 45140 11908 45149 11948
rect 45091 11907 45149 11908
rect 49323 11948 49365 11957
rect 49323 11908 49324 11948
rect 49364 11908 49365 11948
rect 49323 11899 49365 11908
rect 4011 11864 4053 11873
rect 4011 11824 4012 11864
rect 4052 11824 4053 11864
rect 4011 11815 4053 11824
rect 11403 11864 11445 11873
rect 11403 11824 11404 11864
rect 11444 11824 11445 11864
rect 11403 11815 11445 11824
rect 14571 11864 14613 11873
rect 14571 11824 14572 11864
rect 14612 11824 14613 11864
rect 14571 11815 14613 11824
rect 14955 11864 14997 11873
rect 14955 11824 14956 11864
rect 14996 11824 14997 11864
rect 14955 11815 14997 11824
rect 16771 11864 16829 11865
rect 16771 11824 16780 11864
rect 16820 11824 16829 11864
rect 16771 11823 16829 11824
rect 18987 11864 19029 11873
rect 18987 11824 18988 11864
rect 19028 11824 19029 11864
rect 18987 11815 19029 11824
rect 31659 11864 31701 11873
rect 31659 11824 31660 11864
rect 31700 11824 31701 11864
rect 31659 11815 31701 11824
rect 32043 11864 32085 11873
rect 32043 11824 32044 11864
rect 32084 11824 32085 11864
rect 32043 11815 32085 11824
rect 6219 11780 6261 11789
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 18891 11780 18933 11789
rect 18891 11740 18892 11780
rect 18932 11740 18933 11780
rect 18891 11731 18933 11740
rect 19083 11780 19125 11789
rect 19083 11740 19084 11780
rect 19124 11740 19125 11780
rect 19083 11731 19125 11740
rect 24843 11780 24885 11789
rect 24843 11740 24844 11780
rect 24884 11740 24885 11780
rect 24843 11731 24885 11740
rect 26851 11780 26909 11781
rect 26851 11740 26860 11780
rect 26900 11740 26909 11780
rect 26851 11739 26909 11740
rect 46723 11780 46781 11781
rect 46723 11740 46732 11780
rect 46772 11740 46781 11780
rect 46723 11739 46781 11740
rect 20523 11711 20565 11720
rect 3715 11696 3773 11697
rect 3715 11656 3724 11696
rect 3764 11656 3773 11696
rect 3715 11655 3773 11656
rect 3819 11696 3861 11705
rect 3819 11656 3820 11696
rect 3860 11656 3861 11696
rect 3819 11647 3861 11656
rect 4011 11696 4053 11705
rect 4011 11656 4012 11696
rect 4052 11656 4053 11696
rect 4011 11647 4053 11656
rect 4203 11696 4245 11705
rect 4203 11656 4204 11696
rect 4244 11656 4245 11696
rect 4203 11647 4245 11656
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4395 11647 4437 11656
rect 4483 11696 4541 11697
rect 4483 11656 4492 11696
rect 4532 11656 4541 11696
rect 4483 11655 4541 11656
rect 4675 11696 4733 11697
rect 4675 11656 4684 11696
rect 4724 11656 4733 11696
rect 4675 11655 4733 11656
rect 5539 11696 5597 11697
rect 5539 11656 5548 11696
rect 5588 11656 5597 11696
rect 5539 11655 5597 11656
rect 6595 11696 6653 11697
rect 6595 11656 6604 11696
rect 6644 11656 6653 11696
rect 6595 11655 6653 11656
rect 7947 11696 7989 11705
rect 7947 11656 7948 11696
rect 7988 11656 7989 11696
rect 7947 11647 7989 11656
rect 8235 11696 8277 11705
rect 8235 11656 8236 11696
rect 8276 11656 8277 11696
rect 8235 11647 8277 11656
rect 8427 11696 8469 11705
rect 8427 11656 8428 11696
rect 8468 11656 8469 11696
rect 8427 11647 8469 11656
rect 8619 11696 8661 11705
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 8715 11696 8757 11705
rect 8715 11656 8716 11696
rect 8756 11656 8757 11696
rect 8715 11647 8757 11656
rect 8907 11696 8949 11705
rect 8907 11656 8908 11696
rect 8948 11656 8949 11696
rect 8907 11647 8949 11656
rect 9003 11696 9045 11705
rect 9003 11656 9004 11696
rect 9044 11656 9045 11696
rect 9003 11647 9045 11656
rect 9387 11696 9429 11705
rect 9387 11656 9388 11696
rect 9428 11656 9429 11696
rect 9387 11647 9429 11656
rect 9579 11696 9621 11705
rect 9579 11656 9580 11696
rect 9620 11656 9621 11696
rect 9579 11647 9621 11656
rect 9667 11696 9725 11697
rect 9667 11656 9676 11696
rect 9716 11656 9725 11696
rect 9667 11655 9725 11656
rect 9859 11696 9917 11697
rect 9859 11656 9868 11696
rect 9908 11656 9917 11696
rect 9859 11655 9917 11656
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10155 11696 10197 11705
rect 10155 11656 10156 11696
rect 10196 11656 10197 11696
rect 10155 11647 10197 11656
rect 11595 11696 11637 11705
rect 11595 11656 11596 11696
rect 11636 11656 11637 11696
rect 11595 11647 11637 11656
rect 11691 11696 11733 11705
rect 11691 11656 11692 11696
rect 11732 11656 11733 11696
rect 11691 11647 11733 11656
rect 11787 11696 11829 11705
rect 11787 11656 11788 11696
rect 11828 11656 11829 11696
rect 11787 11647 11829 11656
rect 11883 11696 11925 11705
rect 11883 11656 11884 11696
rect 11924 11656 11925 11696
rect 11883 11647 11925 11656
rect 12067 11696 12125 11697
rect 12067 11656 12076 11696
rect 12116 11656 12125 11696
rect 12067 11655 12125 11656
rect 13027 11696 13085 11697
rect 13027 11656 13036 11696
rect 13076 11656 13085 11696
rect 13027 11655 13085 11656
rect 13219 11696 13277 11697
rect 13219 11656 13228 11696
rect 13268 11656 13277 11696
rect 13219 11655 13277 11656
rect 14091 11696 14133 11705
rect 14091 11656 14092 11696
rect 14132 11656 14133 11696
rect 14091 11647 14133 11656
rect 14187 11696 14229 11705
rect 14187 11656 14188 11696
rect 14228 11656 14229 11696
rect 14187 11647 14229 11656
rect 14283 11696 14325 11705
rect 14283 11656 14284 11696
rect 14324 11656 14325 11696
rect 14283 11647 14325 11656
rect 14379 11696 14421 11705
rect 14379 11656 14380 11696
rect 14420 11656 14421 11696
rect 14379 11647 14421 11656
rect 16099 11696 16157 11697
rect 16099 11656 16108 11696
rect 16148 11656 16157 11696
rect 16099 11655 16157 11656
rect 16395 11696 16437 11705
rect 16395 11656 16396 11696
rect 16436 11656 16437 11696
rect 16395 11647 16437 11656
rect 17059 11696 17117 11697
rect 17059 11656 17068 11696
rect 17108 11656 17117 11696
rect 17059 11655 17117 11656
rect 17355 11696 17397 11705
rect 17355 11656 17356 11696
rect 17396 11656 17397 11696
rect 17355 11647 17397 11656
rect 17451 11696 17493 11705
rect 17451 11656 17452 11696
rect 17492 11656 17493 11696
rect 17451 11647 17493 11656
rect 18219 11696 18261 11705
rect 18219 11656 18220 11696
rect 18260 11656 18261 11696
rect 18219 11647 18261 11656
rect 18315 11696 18357 11705
rect 18315 11656 18316 11696
rect 18356 11656 18357 11696
rect 18315 11647 18357 11656
rect 18411 11696 18453 11705
rect 18411 11656 18412 11696
rect 18452 11656 18453 11696
rect 18411 11647 18453 11656
rect 18787 11696 18845 11697
rect 18787 11656 18796 11696
rect 18836 11656 18845 11696
rect 18787 11655 18845 11656
rect 19179 11696 19221 11705
rect 19179 11656 19180 11696
rect 19220 11656 19221 11696
rect 19179 11647 19221 11656
rect 19851 11696 19893 11705
rect 19851 11656 19852 11696
rect 19892 11656 19893 11696
rect 19851 11647 19893 11656
rect 19947 11696 19989 11705
rect 19947 11656 19948 11696
rect 19988 11656 19989 11696
rect 19947 11647 19989 11656
rect 20043 11696 20085 11705
rect 20043 11656 20044 11696
rect 20084 11656 20085 11696
rect 20043 11647 20085 11656
rect 20227 11696 20285 11697
rect 20227 11656 20236 11696
rect 20276 11656 20285 11696
rect 20227 11655 20285 11656
rect 20323 11696 20381 11697
rect 20323 11656 20332 11696
rect 20372 11656 20381 11696
rect 20523 11671 20524 11711
rect 20564 11671 20565 11711
rect 20776 11711 20818 11720
rect 20523 11662 20565 11671
rect 20619 11696 20661 11705
rect 20323 11655 20381 11656
rect 20619 11656 20620 11696
rect 20660 11656 20661 11696
rect 20776 11671 20777 11711
rect 20817 11671 20818 11711
rect 21640 11711 21682 11720
rect 20776 11662 20818 11671
rect 21091 11696 21149 11697
rect 20619 11647 20661 11656
rect 21091 11656 21100 11696
rect 21140 11656 21149 11696
rect 21091 11655 21149 11656
rect 21187 11696 21245 11697
rect 21187 11656 21196 11696
rect 21236 11656 21245 11696
rect 21187 11655 21245 11656
rect 21387 11696 21429 11705
rect 21387 11656 21388 11696
rect 21428 11656 21429 11696
rect 21387 11647 21429 11656
rect 21483 11696 21525 11705
rect 21483 11656 21484 11696
rect 21524 11656 21525 11696
rect 21640 11671 21641 11711
rect 21681 11671 21682 11711
rect 21640 11662 21682 11671
rect 23499 11696 23541 11705
rect 21483 11647 21525 11656
rect 23499 11656 23500 11696
rect 23540 11656 23541 11696
rect 23499 11647 23541 11656
rect 23595 11696 23637 11705
rect 23595 11656 23596 11696
rect 23636 11656 23637 11696
rect 23595 11647 23637 11656
rect 23683 11696 23741 11697
rect 23683 11656 23692 11696
rect 23732 11656 23741 11696
rect 23683 11655 23741 11656
rect 23971 11696 24029 11697
rect 23971 11656 23980 11696
rect 24020 11656 24029 11696
rect 23971 11655 24029 11656
rect 26563 11696 26621 11697
rect 26563 11656 26572 11696
rect 26612 11656 26621 11696
rect 26563 11655 26621 11656
rect 26659 11696 26717 11697
rect 26659 11656 26668 11696
rect 26708 11656 26717 11696
rect 26659 11655 26717 11656
rect 27043 11696 27101 11697
rect 27043 11656 27052 11696
rect 27092 11656 27101 11696
rect 27043 11655 27101 11656
rect 28003 11696 28061 11697
rect 28003 11656 28012 11696
rect 28052 11656 28061 11696
rect 28003 11655 28061 11656
rect 28299 11696 28341 11705
rect 28299 11656 28300 11696
rect 28340 11656 28341 11696
rect 28299 11647 28341 11656
rect 28491 11696 28533 11705
rect 28491 11656 28492 11696
rect 28532 11656 28533 11696
rect 28491 11647 28533 11656
rect 28875 11696 28917 11705
rect 28875 11656 28876 11696
rect 28916 11656 28917 11696
rect 28875 11647 28917 11656
rect 29067 11696 29109 11705
rect 29067 11656 29068 11696
rect 29108 11656 29109 11696
rect 29067 11647 29109 11656
rect 29155 11696 29213 11697
rect 29155 11656 29164 11696
rect 29204 11656 29213 11696
rect 29155 11655 29213 11656
rect 31459 11696 31517 11697
rect 31459 11656 31468 11696
rect 31508 11656 31517 11696
rect 31459 11655 31517 11656
rect 31651 11696 31709 11697
rect 31651 11656 31660 11696
rect 31700 11656 31709 11696
rect 31651 11655 31709 11656
rect 31947 11696 31989 11705
rect 31947 11656 31948 11696
rect 31988 11656 31989 11696
rect 31947 11647 31989 11656
rect 32139 11696 32181 11705
rect 32139 11656 32140 11696
rect 32180 11656 32181 11696
rect 32139 11647 32181 11656
rect 32235 11696 32277 11705
rect 32235 11656 32236 11696
rect 32276 11656 32277 11696
rect 32235 11647 32277 11656
rect 32427 11696 32469 11705
rect 32427 11656 32428 11696
rect 32468 11656 32469 11696
rect 32427 11647 32469 11656
rect 32523 11696 32565 11705
rect 32523 11656 32524 11696
rect 32564 11656 32565 11696
rect 32523 11647 32565 11656
rect 32619 11696 32661 11705
rect 32619 11656 32620 11696
rect 32660 11656 32661 11696
rect 32619 11647 32661 11656
rect 32907 11696 32949 11705
rect 32907 11656 32908 11696
rect 32948 11656 32949 11696
rect 32907 11647 32949 11656
rect 32995 11696 33053 11697
rect 32995 11656 33004 11696
rect 33044 11656 33053 11696
rect 32995 11655 33053 11656
rect 33771 11696 33813 11705
rect 33771 11656 33772 11696
rect 33812 11656 33813 11696
rect 33771 11647 33813 11656
rect 33867 11696 33909 11705
rect 33867 11656 33868 11696
rect 33908 11656 33909 11696
rect 33867 11647 33909 11656
rect 33963 11696 34005 11705
rect 33963 11656 33964 11696
rect 34004 11656 34005 11696
rect 33963 11647 34005 11656
rect 34155 11696 34197 11705
rect 34155 11656 34156 11696
rect 34196 11656 34197 11696
rect 34155 11647 34197 11656
rect 34251 11696 34293 11705
rect 34251 11656 34252 11696
rect 34292 11656 34293 11696
rect 34251 11647 34293 11656
rect 34731 11696 34773 11705
rect 34731 11656 34732 11696
rect 34772 11656 34773 11696
rect 34731 11647 34773 11656
rect 34827 11696 34869 11705
rect 34827 11656 34828 11696
rect 34868 11656 34869 11696
rect 34827 11647 34869 11656
rect 34923 11696 34965 11705
rect 34923 11656 34924 11696
rect 34964 11656 34965 11696
rect 34923 11647 34965 11656
rect 35203 11696 35261 11697
rect 35203 11656 35212 11696
rect 35252 11656 35261 11696
rect 35203 11655 35261 11656
rect 36259 11696 36317 11697
rect 36259 11656 36268 11696
rect 36308 11656 36317 11696
rect 36259 11655 36317 11656
rect 36555 11696 36597 11705
rect 36555 11656 36556 11696
rect 36596 11656 36597 11696
rect 36555 11647 36597 11656
rect 36651 11696 36693 11705
rect 36651 11656 36652 11696
rect 36692 11656 36693 11696
rect 36651 11647 36693 11656
rect 37419 11696 37461 11705
rect 37419 11656 37420 11696
rect 37460 11656 37461 11696
rect 37419 11647 37461 11656
rect 38563 11696 38621 11697
rect 38563 11656 38572 11696
rect 38612 11656 38621 11696
rect 38563 11655 38621 11656
rect 39243 11696 39285 11705
rect 39243 11656 39244 11696
rect 39284 11656 39285 11696
rect 39243 11647 39285 11656
rect 39435 11696 39477 11705
rect 39435 11656 39436 11696
rect 39476 11656 39477 11696
rect 39435 11647 39477 11656
rect 39531 11696 39573 11705
rect 39531 11656 39532 11696
rect 39572 11656 39573 11696
rect 39531 11647 39573 11656
rect 40387 11696 40445 11697
rect 40387 11656 40396 11696
rect 40436 11656 40445 11696
rect 40387 11655 40445 11656
rect 40483 11696 40541 11697
rect 40483 11656 40492 11696
rect 40532 11656 40541 11696
rect 40483 11655 40541 11656
rect 41251 11696 41309 11697
rect 41251 11656 41260 11696
rect 41300 11656 41309 11696
rect 41251 11655 41309 11656
rect 42115 11696 42173 11697
rect 42115 11656 42124 11696
rect 42164 11656 42173 11696
rect 42115 11655 42173 11656
rect 43459 11696 43517 11697
rect 43459 11656 43468 11696
rect 43508 11656 43517 11696
rect 43459 11655 43517 11656
rect 44331 11696 44373 11705
rect 44331 11656 44332 11696
rect 44372 11656 44373 11696
rect 44331 11647 44373 11656
rect 44803 11696 44861 11697
rect 44803 11656 44812 11696
rect 44852 11656 44861 11696
rect 44803 11655 44861 11656
rect 45763 11696 45821 11697
rect 45763 11656 45772 11696
rect 45812 11656 45821 11696
rect 45763 11655 45821 11656
rect 46435 11696 46493 11697
rect 46435 11656 46444 11696
rect 46484 11656 46493 11696
rect 46435 11655 46493 11656
rect 46531 11696 46589 11697
rect 46531 11656 46540 11696
rect 46580 11656 46589 11696
rect 46531 11655 46589 11656
rect 46923 11696 46965 11705
rect 46923 11656 46924 11696
rect 46964 11656 46965 11696
rect 46923 11647 46965 11656
rect 47299 11696 47357 11697
rect 47299 11656 47308 11696
rect 47348 11656 47357 11696
rect 47299 11655 47357 11656
rect 48163 11696 48221 11697
rect 48163 11656 48172 11696
rect 48212 11656 48221 11696
rect 48163 11655 48221 11656
rect 16491 11612 16533 11621
rect 16491 11572 16492 11612
rect 16532 11572 16533 11612
rect 16491 11563 16533 11572
rect 32715 11612 32757 11621
rect 32715 11572 32716 11612
rect 32756 11572 32757 11612
rect 32715 11563 32757 11572
rect 40875 11612 40917 11621
rect 40875 11572 40876 11612
rect 40916 11572 40917 11612
rect 40875 11563 40917 11572
rect 643 11528 701 11529
rect 643 11488 652 11528
rect 692 11488 701 11528
rect 643 11487 701 11488
rect 4291 11528 4349 11529
rect 4291 11488 4300 11528
rect 4340 11488 4349 11528
rect 4291 11487 4349 11488
rect 5347 11528 5405 11529
rect 5347 11488 5356 11528
rect 5396 11488 5405 11528
rect 5347 11487 5405 11488
rect 6691 11528 6749 11529
rect 6691 11488 6700 11528
rect 6740 11488 6749 11528
rect 6691 11487 6749 11488
rect 8139 11528 8181 11537
rect 8139 11488 8140 11528
rect 8180 11488 8181 11528
rect 8139 11479 8181 11488
rect 9187 11528 9245 11529
rect 9187 11488 9196 11528
rect 9236 11488 9245 11528
rect 9187 11487 9245 11488
rect 9475 11528 9533 11529
rect 9475 11488 9484 11528
rect 9524 11488 9533 11528
rect 9475 11487 9533 11488
rect 12739 11528 12797 11529
rect 12739 11488 12748 11528
rect 12788 11488 12797 11528
rect 12739 11487 12797 11488
rect 13891 11528 13949 11529
rect 13891 11488 13900 11528
rect 13940 11488 13949 11528
rect 13891 11487 13949 11488
rect 18115 11528 18173 11529
rect 18115 11488 18124 11528
rect 18164 11488 18173 11528
rect 18115 11487 18173 11488
rect 19747 11528 19805 11529
rect 19747 11488 19756 11528
rect 19796 11488 19805 11528
rect 19747 11487 19805 11488
rect 20419 11528 20477 11529
rect 20419 11488 20428 11528
rect 20468 11488 20477 11528
rect 20419 11487 20477 11488
rect 21379 11528 21437 11529
rect 21379 11488 21388 11528
rect 21428 11488 21437 11528
rect 21379 11487 21437 11488
rect 24459 11528 24501 11537
rect 24459 11488 24460 11528
rect 24500 11488 24501 11528
rect 24459 11479 24501 11488
rect 28395 11528 28437 11537
rect 28395 11488 28396 11528
rect 28436 11488 28437 11528
rect 28395 11479 28437 11488
rect 28963 11528 29021 11529
rect 28963 11488 28972 11528
rect 29012 11488 29021 11528
rect 28963 11487 29021 11488
rect 33667 11528 33725 11529
rect 33667 11488 33676 11528
rect 33716 11488 33725 11528
rect 33667 11487 33725 11488
rect 34435 11528 34493 11529
rect 34435 11488 34444 11528
rect 34484 11488 34493 11528
rect 34435 11487 34493 11488
rect 34627 11528 34685 11529
rect 34627 11488 34636 11528
rect 34676 11488 34685 11528
rect 34627 11487 34685 11488
rect 35307 11528 35349 11537
rect 35307 11488 35308 11528
rect 35348 11488 35349 11528
rect 35307 11479 35349 11488
rect 36171 11528 36213 11537
rect 36171 11488 36172 11528
rect 36212 11488 36213 11528
rect 36171 11479 36213 11488
rect 36835 11528 36893 11529
rect 36835 11488 36844 11528
rect 36884 11488 36893 11528
rect 36835 11487 36893 11488
rect 37131 11528 37173 11537
rect 37131 11488 37132 11528
rect 37172 11488 37173 11528
rect 37131 11479 37173 11488
rect 38091 11528 38133 11537
rect 38091 11488 38092 11528
rect 38132 11488 38133 11528
rect 38091 11479 38133 11488
rect 39523 11528 39581 11529
rect 39523 11488 39532 11528
rect 39572 11488 39581 11528
rect 39523 11487 39581 11488
rect 40683 11528 40725 11537
rect 40683 11488 40684 11528
rect 40724 11488 40725 11528
rect 40683 11479 40725 11488
rect 43267 11528 43325 11529
rect 43267 11488 43276 11528
rect 43316 11488 43325 11528
rect 43267 11487 43325 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 643 11192 701 11193
rect 643 11152 652 11192
rect 692 11152 701 11192
rect 643 11151 701 11152
rect 3715 11192 3773 11193
rect 3715 11152 3724 11192
rect 3764 11152 3773 11192
rect 3715 11151 3773 11152
rect 5539 11192 5597 11193
rect 5539 11152 5548 11192
rect 5588 11152 5597 11192
rect 5539 11151 5597 11152
rect 9099 11192 9141 11201
rect 9099 11152 9100 11192
rect 9140 11152 9141 11192
rect 9099 11143 9141 11152
rect 11299 11192 11357 11193
rect 11299 11152 11308 11192
rect 11348 11152 11357 11192
rect 11299 11151 11357 11152
rect 16291 11192 16349 11193
rect 16291 11152 16300 11192
rect 16340 11152 16349 11192
rect 16291 11151 16349 11152
rect 16771 11192 16829 11193
rect 16771 11152 16780 11192
rect 16820 11152 16829 11192
rect 16771 11151 16829 11152
rect 17059 11192 17117 11193
rect 17059 11152 17068 11192
rect 17108 11152 17117 11192
rect 17059 11151 17117 11152
rect 17251 11192 17309 11193
rect 17251 11152 17260 11192
rect 17300 11152 17309 11192
rect 17251 11151 17309 11152
rect 27051 11192 27093 11201
rect 27051 11152 27052 11192
rect 27092 11152 27093 11192
rect 27051 11143 27093 11152
rect 31747 11192 31805 11193
rect 31747 11152 31756 11192
rect 31796 11152 31805 11192
rect 31747 11151 31805 11152
rect 35203 11192 35261 11193
rect 35203 11152 35212 11192
rect 35252 11152 35261 11192
rect 35203 11151 35261 11152
rect 37507 11192 37565 11193
rect 37507 11152 37516 11192
rect 37556 11152 37565 11192
rect 37507 11151 37565 11152
rect 40003 11192 40061 11193
rect 40003 11152 40012 11192
rect 40052 11152 40061 11192
rect 40003 11151 40061 11152
rect 40867 11192 40925 11193
rect 40867 11152 40876 11192
rect 40916 11152 40925 11192
rect 40867 11151 40925 11152
rect 42403 11192 42461 11193
rect 42403 11152 42412 11192
rect 42452 11152 42461 11192
rect 42403 11151 42461 11152
rect 44227 11192 44285 11193
rect 44227 11152 44236 11192
rect 44276 11152 44285 11192
rect 44227 11151 44285 11152
rect 45091 11192 45149 11193
rect 45091 11152 45100 11192
rect 45140 11152 45149 11192
rect 45091 11151 45149 11152
rect 46635 11192 46677 11201
rect 46635 11152 46636 11192
rect 46676 11152 46677 11192
rect 46635 11143 46677 11152
rect 48547 11192 48605 11193
rect 48547 11152 48556 11192
rect 48596 11152 48605 11192
rect 48547 11151 48605 11152
rect 48835 11192 48893 11193
rect 48835 11152 48844 11192
rect 48884 11152 48893 11192
rect 48835 11151 48893 11152
rect 10155 11108 10197 11117
rect 10155 11068 10156 11108
rect 10196 11068 10197 11108
rect 10155 11059 10197 11068
rect 13707 11108 13749 11117
rect 13707 11068 13708 11108
rect 13748 11068 13749 11108
rect 13707 11059 13749 11068
rect 29163 11108 29205 11117
rect 29163 11068 29164 11108
rect 29204 11068 29205 11108
rect 29163 11059 29205 11068
rect 37803 11108 37845 11117
rect 37803 11068 37804 11108
rect 37844 11068 37845 11108
rect 37803 11059 37845 11068
rect 42307 11108 42365 11109
rect 42307 11068 42316 11108
rect 42356 11068 42365 11108
rect 42307 11067 42365 11068
rect 48451 11108 48509 11109
rect 48451 11068 48460 11108
rect 48500 11068 48509 11108
rect 48451 11067 48509 11068
rect 2571 11024 2613 11033
rect 2571 10984 2572 11024
rect 2612 10984 2613 11024
rect 2571 10975 2613 10984
rect 2667 11024 2709 11033
rect 2667 10984 2668 11024
rect 2708 10984 2709 11024
rect 2667 10975 2709 10984
rect 2859 11024 2901 11033
rect 2859 10984 2860 11024
rect 2900 10984 2901 11024
rect 2859 10975 2901 10984
rect 3619 11024 3677 11025
rect 3619 10984 3628 11024
rect 3668 10984 3677 11024
rect 3619 10983 3677 10984
rect 4291 11024 4349 11025
rect 4291 10984 4300 11024
rect 4340 10984 4349 11024
rect 4291 10983 4349 10984
rect 5251 11024 5309 11025
rect 5251 10984 5260 11024
rect 5300 10984 5309 11024
rect 5251 10983 5309 10984
rect 5739 11024 5781 11033
rect 5739 10984 5740 11024
rect 5780 10984 5781 11024
rect 5739 10975 5781 10984
rect 5835 11024 5877 11033
rect 5835 10984 5836 11024
rect 5876 10984 5877 11024
rect 5835 10975 5877 10984
rect 5931 11024 5973 11033
rect 5931 10984 5932 11024
rect 5972 10984 5973 11024
rect 5931 10975 5973 10984
rect 6027 11024 6069 11033
rect 6027 10984 6028 11024
rect 6068 10984 6069 11024
rect 6027 10975 6069 10984
rect 6979 11024 7037 11025
rect 6979 10984 6988 11024
rect 7028 10984 7037 11024
rect 6979 10983 7037 10984
rect 7659 11024 7701 11033
rect 7659 10984 7660 11024
rect 7700 10984 7701 11024
rect 7659 10975 7701 10984
rect 7755 11024 7797 11033
rect 7755 10984 7756 11024
rect 7796 10984 7797 11024
rect 7755 10975 7797 10984
rect 7851 11024 7893 11033
rect 7851 10984 7852 11024
rect 7892 10984 7893 11024
rect 7851 10975 7893 10984
rect 7947 11024 7989 11033
rect 7947 10984 7948 11024
rect 7988 10984 7989 11024
rect 7947 10975 7989 10984
rect 8139 11024 8181 11033
rect 8139 10984 8140 11024
rect 8180 10984 8181 11024
rect 8139 10975 8181 10984
rect 8427 11024 8469 11033
rect 8427 10984 8428 11024
rect 8468 10984 8469 11024
rect 8427 10975 8469 10984
rect 8619 11024 8661 11033
rect 8619 10984 8620 11024
rect 8660 10984 8661 11024
rect 8619 10975 8661 10984
rect 8907 11024 8949 11033
rect 8907 10984 8908 11024
rect 8948 10984 8949 11024
rect 8907 10975 8949 10984
rect 9283 11024 9341 11025
rect 9283 10984 9292 11024
rect 9332 10984 9341 11024
rect 9283 10983 9341 10984
rect 9379 11024 9437 11025
rect 9379 10984 9388 11024
rect 9428 10984 9437 11024
rect 9667 11024 9725 11025
rect 9379 10983 9437 10984
rect 9483 10982 9525 10991
rect 9667 10984 9676 11024
rect 9716 10984 9725 11024
rect 9667 10983 9725 10984
rect 9867 11024 9909 11033
rect 9867 10984 9868 11024
rect 9908 10984 9909 11024
rect 9483 10942 9484 10982
rect 9524 10942 9525 10982
rect 9867 10975 9909 10984
rect 9963 11024 10005 11033
rect 9963 10984 9964 11024
rect 10004 10984 10005 11024
rect 9963 10975 10005 10984
rect 10059 11024 10101 11033
rect 10059 10984 10060 11024
rect 10100 10984 10101 11024
rect 10059 10975 10101 10984
rect 12451 11024 12509 11025
rect 12451 10984 12460 11024
rect 12500 10984 12509 11024
rect 12451 10983 12509 10984
rect 13315 11024 13373 11025
rect 13315 10984 13324 11024
rect 13364 10984 13373 11024
rect 13315 10983 13373 10984
rect 13899 11024 13941 11033
rect 13899 10984 13900 11024
rect 13940 10984 13941 11024
rect 13899 10975 13941 10984
rect 14275 11024 14333 11025
rect 14275 10984 14284 11024
rect 14324 10984 14333 11024
rect 14275 10983 14333 10984
rect 15139 11024 15197 11025
rect 15139 10984 15148 11024
rect 15188 10984 15197 11024
rect 15139 10983 15197 10984
rect 16867 11024 16925 11025
rect 16867 10984 16876 11024
rect 16916 10984 16925 11024
rect 16867 10983 16925 10984
rect 17355 11024 17397 11033
rect 17355 10984 17356 11024
rect 17396 10984 17397 11024
rect 17355 10975 17397 10984
rect 17451 11024 17493 11033
rect 17451 10984 17452 11024
rect 17492 10984 17493 11024
rect 17451 10975 17493 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 18403 11024 18461 11025
rect 18403 10984 18412 11024
rect 18452 10984 18461 11024
rect 18403 10983 18461 10984
rect 18595 11024 18653 11025
rect 18595 10984 18604 11024
rect 18644 10984 18653 11024
rect 18595 10983 18653 10984
rect 19459 11024 19517 11025
rect 19459 10984 19468 11024
rect 19508 10984 19517 11024
rect 19459 10983 19517 10984
rect 19563 11024 19605 11033
rect 19563 10984 19564 11024
rect 19604 10984 19605 11024
rect 19563 10975 19605 10984
rect 19755 11024 19797 11033
rect 19755 10984 19756 11024
rect 19796 10984 19797 11024
rect 19755 10975 19797 10984
rect 20515 11024 20573 11025
rect 20515 10984 20524 11024
rect 20564 10984 20573 11024
rect 20515 10983 20573 10984
rect 20907 11024 20949 11033
rect 20907 10984 20908 11024
rect 20948 10984 20949 11024
rect 20907 10975 20949 10984
rect 23587 11024 23645 11025
rect 23587 10984 23596 11024
rect 23636 10984 23645 11024
rect 23587 10983 23645 10984
rect 23691 11024 23733 11033
rect 23691 10984 23692 11024
rect 23732 10984 23733 11024
rect 23691 10975 23733 10984
rect 23883 11024 23925 11033
rect 23883 10984 23884 11024
rect 23924 10984 23925 11024
rect 23883 10975 23925 10984
rect 24075 11024 24117 11033
rect 24075 10984 24076 11024
rect 24116 10984 24117 11024
rect 24075 10975 24117 10984
rect 24171 11024 24213 11033
rect 24171 10984 24172 11024
rect 24212 10984 24213 11024
rect 24171 10975 24213 10984
rect 24267 11024 24309 11033
rect 24267 10984 24268 11024
rect 24308 10984 24309 11024
rect 24267 10975 24309 10984
rect 24363 11024 24405 11033
rect 24363 10984 24364 11024
rect 24404 10984 24405 11024
rect 24363 10975 24405 10984
rect 24739 11024 24797 11025
rect 24739 10984 24748 11024
rect 24788 10984 24797 11024
rect 24739 10983 24797 10984
rect 24843 11024 24885 11033
rect 24843 10984 24844 11024
rect 24884 10984 24885 11024
rect 24843 10975 24885 10984
rect 27339 11024 27381 11033
rect 27339 10984 27340 11024
rect 27380 10984 27381 11024
rect 27339 10975 27381 10984
rect 27523 11024 27581 11025
rect 27523 10984 27532 11024
rect 27572 10984 27581 11024
rect 27523 10983 27581 10984
rect 27715 11024 27773 11025
rect 27715 10984 27724 11024
rect 27764 10984 27773 11024
rect 27715 10983 27773 10984
rect 28107 11024 28149 11033
rect 28107 10984 28108 11024
rect 28148 10984 28149 11024
rect 28107 10975 28149 10984
rect 29259 11024 29301 11033
rect 29259 10984 29260 11024
rect 29300 10984 29301 11024
rect 29259 10975 29301 10984
rect 29539 11024 29597 11025
rect 29539 10984 29548 11024
rect 29588 10984 29597 11024
rect 29539 10983 29597 10984
rect 30787 11024 30845 11025
rect 30787 10984 30796 11024
rect 30836 10984 30845 11024
rect 30787 10983 30845 10984
rect 31467 11024 31509 11033
rect 31467 10984 31468 11024
rect 31508 10984 31509 11024
rect 31467 10975 31509 10984
rect 31563 11024 31605 11033
rect 31563 10984 31564 11024
rect 31604 10984 31605 11024
rect 31563 10975 31605 10984
rect 31947 11024 31989 11033
rect 31947 10984 31948 11024
rect 31988 10984 31989 11024
rect 31947 10975 31989 10984
rect 32323 11024 32381 11025
rect 32323 10984 32332 11024
rect 32372 10984 32381 11024
rect 32323 10983 32381 10984
rect 32515 11024 32573 11025
rect 32515 10984 32524 11024
rect 32564 10984 32573 11024
rect 32515 10983 32573 10984
rect 32907 11024 32949 11033
rect 32907 10984 32908 11024
rect 32948 10984 32949 11024
rect 32213 10982 32271 10983
rect 9483 10933 9525 10942
rect 17739 10940 17781 10949
rect 17739 10900 17740 10940
rect 17780 10900 17781 10940
rect 17739 10891 17781 10900
rect 20619 10940 20661 10949
rect 20619 10900 20620 10940
rect 20660 10900 20661 10940
rect 20619 10891 20661 10900
rect 20811 10940 20853 10949
rect 20811 10900 20812 10940
rect 20852 10900 20853 10940
rect 20811 10891 20853 10900
rect 24939 10940 24981 10949
rect 24939 10900 24940 10940
rect 24980 10900 24981 10940
rect 24939 10891 24981 10900
rect 32043 10940 32085 10949
rect 32213 10942 32222 10982
rect 32262 10942 32271 10982
rect 32907 10975 32949 10984
rect 33099 11024 33141 11033
rect 33099 10984 33100 11024
rect 33140 10984 33141 11024
rect 33099 10975 33141 10984
rect 33195 11024 33237 11033
rect 33195 10984 33196 11024
rect 33236 10984 33237 11024
rect 33195 10975 33237 10984
rect 33291 11024 33333 11033
rect 33291 10984 33292 11024
rect 33332 10984 33333 11024
rect 33291 10975 33333 10984
rect 33387 11024 33429 11033
rect 33387 10984 33388 11024
rect 33428 10984 33429 11024
rect 33387 10975 33429 10984
rect 34923 11024 34965 11033
rect 34923 10984 34924 11024
rect 34964 10984 34965 11024
rect 34923 10975 34965 10984
rect 35019 11024 35061 11033
rect 35019 10984 35020 11024
rect 35060 10984 35061 11024
rect 35019 10975 35061 10984
rect 35499 11024 35541 11033
rect 35499 10984 35500 11024
rect 35540 10984 35541 11024
rect 35499 10975 35541 10984
rect 35595 11024 35637 11033
rect 35595 10984 35596 11024
rect 35636 10984 35637 11024
rect 35595 10975 35637 10984
rect 35691 11024 35733 11033
rect 35691 10984 35692 11024
rect 35732 10984 35733 11024
rect 35691 10975 35733 10984
rect 35787 11024 35829 11033
rect 35787 10984 35788 11024
rect 35828 10984 35829 11024
rect 35787 10975 35829 10984
rect 36171 11024 36213 11033
rect 36171 10984 36172 11024
rect 36212 10984 36213 11024
rect 36171 10975 36213 10984
rect 36267 11024 36309 11033
rect 36267 10984 36268 11024
rect 36308 10984 36309 11024
rect 36267 10975 36309 10984
rect 36363 11024 36405 11033
rect 36363 10984 36364 11024
rect 36404 10984 36405 11024
rect 36363 10975 36405 10984
rect 36459 11024 36501 11033
rect 36459 10984 36460 11024
rect 36500 10984 36501 11024
rect 36459 10975 36501 10984
rect 36643 11024 36701 11025
rect 36643 10984 36652 11024
rect 36692 10984 36701 11024
rect 36643 10983 36701 10984
rect 37035 11024 37077 11033
rect 37035 10984 37036 11024
rect 37076 10984 37077 11024
rect 37035 10975 37077 10984
rect 37227 11024 37269 11033
rect 37227 10984 37228 11024
rect 37268 10984 37269 11024
rect 37227 10975 37269 10984
rect 37323 11024 37365 11033
rect 37323 10984 37324 11024
rect 37364 10984 37365 11024
rect 37323 10975 37365 10984
rect 37707 11024 37749 11033
rect 37707 10984 37708 11024
rect 37748 10984 37749 11024
rect 37707 10975 37749 10984
rect 37899 11024 37941 11033
rect 37899 10984 37900 11024
rect 37940 10984 37941 11024
rect 37899 10975 37941 10984
rect 37987 11024 38045 11025
rect 37987 10984 37996 11024
rect 38036 10984 38045 11024
rect 37987 10983 38045 10984
rect 38187 11024 38229 11033
rect 38187 10984 38188 11024
rect 38228 10984 38229 11024
rect 38187 10975 38229 10984
rect 38379 11024 38421 11033
rect 38379 10984 38380 11024
rect 38420 10984 38421 11024
rect 38379 10975 38421 10984
rect 38467 11024 38525 11025
rect 38467 10984 38476 11024
rect 38516 10984 38525 11024
rect 38467 10983 38525 10984
rect 38659 11024 38717 11025
rect 38659 10984 38668 11024
rect 38708 10984 38717 11024
rect 38659 10983 38717 10984
rect 38763 11024 38805 11033
rect 38763 10984 38764 11024
rect 38804 10984 38805 11024
rect 38763 10975 38805 10984
rect 38947 11024 39005 11025
rect 38947 10984 38956 11024
rect 38996 10984 39005 11024
rect 38947 10983 39005 10984
rect 39811 11024 39869 11025
rect 39811 10984 39820 11024
rect 39860 10984 39869 11024
rect 39811 10983 39869 10984
rect 40675 11024 40733 11025
rect 40675 10984 40684 11024
rect 40724 10984 40733 11024
rect 40675 10983 40733 10984
rect 41539 11024 41597 11025
rect 41539 10984 41548 11024
rect 41588 10984 41597 11024
rect 41539 10983 41597 10984
rect 41739 11024 41781 11033
rect 41739 10984 41740 11024
rect 41780 10984 41781 11024
rect 41739 10975 41781 10984
rect 41931 11024 41973 11033
rect 41931 10984 41932 11024
rect 41972 10984 41973 11024
rect 41931 10975 41973 10984
rect 42123 11024 42165 11033
rect 42123 10984 42124 11024
rect 42164 10984 42165 11024
rect 42123 10975 42165 10984
rect 42219 11024 42261 11033
rect 42219 10984 42220 11024
rect 42260 10984 42261 11024
rect 42219 10975 42261 10984
rect 43651 11024 43709 11025
rect 43651 10984 43660 11024
rect 43700 10984 43709 11024
rect 43651 10983 43709 10984
rect 43939 11024 43997 11025
rect 43939 10984 43948 11024
rect 43988 10984 43997 11024
rect 43939 10983 43997 10984
rect 44899 11024 44957 11025
rect 44899 10984 44908 11024
rect 44948 10984 44957 11024
rect 44899 10983 44957 10984
rect 45763 11024 45821 11025
rect 45763 10984 45772 11024
rect 45812 10984 45821 11024
rect 45763 10983 45821 10984
rect 46147 11024 46205 11025
rect 46147 10984 46156 11024
rect 46196 10984 46205 11024
rect 46147 10983 46205 10984
rect 47395 11024 47453 11025
rect 47395 10984 47404 11024
rect 47444 10984 47453 11024
rect 47395 10983 47453 10984
rect 48267 11024 48309 11033
rect 48267 10984 48268 11024
rect 48308 10984 48309 11024
rect 48267 10975 48309 10984
rect 48363 11024 48405 11033
rect 48363 10984 48364 11024
rect 48404 10984 48405 11024
rect 48363 10975 48405 10984
rect 48931 11024 48989 11025
rect 48931 10984 48940 11024
rect 48980 10984 48989 11024
rect 48931 10983 48989 10984
rect 32213 10941 32271 10942
rect 32043 10900 32044 10940
rect 32084 10900 32085 10940
rect 32043 10891 32085 10900
rect 32619 10940 32661 10949
rect 32619 10900 32620 10940
rect 32660 10900 32661 10940
rect 32619 10891 32661 10900
rect 32811 10940 32853 10949
rect 32811 10900 32812 10940
rect 32852 10900 32853 10940
rect 32811 10891 32853 10900
rect 36747 10940 36789 10949
rect 36747 10900 36748 10940
rect 36788 10900 36789 10940
rect 36747 10891 36789 10900
rect 36939 10940 36981 10949
rect 36939 10900 36940 10940
rect 36980 10900 36981 10940
rect 36939 10891 36981 10900
rect 41835 10940 41877 10949
rect 41835 10900 41836 10940
rect 41876 10900 41877 10940
rect 41835 10891 41877 10900
rect 1995 10856 2037 10865
rect 1995 10816 1996 10856
rect 2036 10816 2037 10856
rect 1995 10807 2037 10816
rect 2563 10856 2621 10857
rect 2563 10816 2572 10856
rect 2612 10816 2621 10856
rect 2563 10815 2621 10816
rect 4107 10856 4149 10865
rect 4107 10816 4108 10856
rect 4148 10816 4149 10856
rect 4107 10807 4149 10816
rect 8427 10856 8469 10865
rect 8427 10816 8428 10856
rect 8468 10816 8469 10856
rect 8427 10807 8469 10816
rect 20715 10856 20757 10865
rect 20715 10816 20716 10856
rect 20756 10816 20757 10856
rect 20715 10807 20757 10816
rect 25035 10856 25077 10865
rect 25035 10816 25036 10856
rect 25076 10816 25077 10856
rect 25035 10807 25077 10816
rect 28011 10856 28053 10865
rect 28011 10816 28012 10856
rect 28052 10816 28053 10856
rect 28011 10807 28053 10816
rect 28867 10856 28925 10857
rect 28867 10816 28876 10856
rect 28916 10816 28925 10856
rect 28867 10815 28925 10816
rect 30123 10856 30165 10865
rect 30123 10816 30124 10856
rect 30164 10816 30165 10856
rect 32715 10856 32757 10865
rect 30123 10807 30165 10816
rect 32139 10814 32181 10823
rect 3427 10772 3485 10773
rect 3427 10732 3436 10772
rect 3476 10732 3485 10772
rect 3427 10731 3485 10732
rect 4971 10772 5013 10781
rect 4971 10732 4972 10772
rect 5012 10732 5013 10772
rect 4971 10723 5013 10732
rect 6307 10772 6365 10773
rect 6307 10732 6316 10772
rect 6356 10732 6365 10772
rect 6307 10731 6365 10732
rect 8907 10772 8949 10781
rect 8907 10732 8908 10772
rect 8948 10732 8949 10772
rect 8907 10723 8949 10732
rect 11299 10772 11357 10773
rect 11299 10732 11308 10772
rect 11348 10732 11357 10772
rect 11299 10731 11357 10732
rect 19267 10772 19325 10773
rect 19267 10732 19276 10772
rect 19316 10732 19325 10772
rect 19267 10731 19325 10732
rect 19755 10772 19797 10781
rect 19755 10732 19756 10772
rect 19796 10732 19797 10772
rect 19755 10723 19797 10732
rect 23883 10772 23925 10781
rect 23883 10732 23884 10772
rect 23924 10732 23925 10772
rect 23883 10723 23925 10732
rect 25131 10772 25173 10781
rect 25131 10732 25132 10772
rect 25172 10732 25173 10772
rect 32139 10774 32140 10814
rect 32180 10774 32181 10814
rect 32715 10816 32716 10856
rect 32756 10816 32757 10856
rect 32715 10807 32757 10816
rect 36843 10856 36885 10865
rect 36843 10816 36844 10856
rect 36884 10816 36885 10856
rect 36843 10807 36885 10816
rect 42987 10856 43029 10865
rect 42987 10816 42988 10856
rect 43028 10816 43029 10856
rect 42987 10807 43029 10816
rect 48355 10856 48413 10857
rect 48355 10816 48364 10856
rect 48404 10816 48413 10856
rect 48355 10815 48413 10816
rect 32139 10765 32181 10774
rect 38187 10772 38229 10781
rect 25131 10723 25173 10732
rect 38187 10732 38188 10772
rect 38228 10732 38229 10772
rect 38187 10723 38229 10732
rect 38763 10772 38805 10781
rect 38763 10732 38764 10772
rect 38804 10732 38805 10772
rect 38763 10723 38805 10732
rect 39139 10772 39197 10773
rect 39139 10732 39148 10772
rect 39188 10732 39197 10772
rect 39139 10731 39197 10732
rect 40003 10772 40061 10773
rect 40003 10732 40012 10772
rect 40052 10732 40061 10772
rect 40003 10731 40061 10732
rect 42411 10772 42453 10781
rect 42411 10732 42412 10772
rect 42452 10732 42453 10772
rect 42411 10723 42453 10732
rect 44043 10772 44085 10781
rect 44043 10732 44044 10772
rect 44084 10732 44085 10772
rect 44043 10723 44085 10732
rect 48067 10772 48125 10773
rect 48067 10732 48076 10772
rect 48116 10732 48125 10772
rect 48067 10731 48125 10732
rect 49123 10772 49181 10773
rect 49123 10732 49132 10772
rect 49172 10732 49181 10772
rect 49123 10731 49181 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 4195 10436 4253 10437
rect 4195 10396 4204 10436
rect 4244 10396 4253 10436
rect 4195 10395 4253 10396
rect 7467 10436 7509 10445
rect 7467 10396 7468 10436
rect 7508 10396 7509 10436
rect 7467 10387 7509 10396
rect 9579 10436 9621 10445
rect 9579 10396 9580 10436
rect 9620 10396 9621 10436
rect 9579 10387 9621 10396
rect 18211 10436 18269 10437
rect 18211 10396 18220 10436
rect 18260 10396 18269 10436
rect 18211 10395 18269 10396
rect 23979 10436 24021 10445
rect 23979 10396 23980 10436
rect 24020 10396 24021 10436
rect 23979 10387 24021 10396
rect 26275 10436 26333 10437
rect 26275 10396 26284 10436
rect 26324 10396 26333 10436
rect 26275 10395 26333 10396
rect 29355 10436 29397 10445
rect 29355 10396 29356 10436
rect 29396 10396 29397 10436
rect 29355 10387 29397 10396
rect 33483 10436 33525 10445
rect 33483 10396 33484 10436
rect 33524 10396 33525 10436
rect 33483 10387 33525 10396
rect 39147 10436 39189 10445
rect 39147 10396 39148 10436
rect 39188 10396 39189 10436
rect 39147 10387 39189 10396
rect 40203 10436 40245 10445
rect 40203 10396 40204 10436
rect 40244 10396 40245 10436
rect 40203 10387 40245 10396
rect 42891 10436 42933 10445
rect 42891 10396 42892 10436
rect 42932 10396 42933 10436
rect 42891 10387 42933 10396
rect 44227 10436 44285 10437
rect 44227 10396 44236 10436
rect 44276 10396 44285 10436
rect 44227 10395 44285 10396
rect 46347 10436 46389 10445
rect 46347 10396 46348 10436
rect 46388 10396 46389 10436
rect 46347 10387 46389 10396
rect 47019 10436 47061 10445
rect 47019 10396 47020 10436
rect 47060 10396 47061 10436
rect 47019 10387 47061 10396
rect 8235 10352 8277 10361
rect 8235 10312 8236 10352
rect 8276 10312 8277 10352
rect 8235 10303 8277 10312
rect 10251 10352 10293 10361
rect 10251 10312 10252 10352
rect 10292 10312 10293 10352
rect 10251 10303 10293 10312
rect 14091 10352 14133 10361
rect 14091 10312 14092 10352
rect 14132 10312 14133 10352
rect 14091 10303 14133 10312
rect 16011 10352 16053 10361
rect 16011 10312 16012 10352
rect 16052 10312 16053 10352
rect 16011 10303 16053 10312
rect 21187 10352 21245 10353
rect 21187 10312 21196 10352
rect 21236 10312 21245 10352
rect 21187 10311 21245 10312
rect 23011 10352 23069 10353
rect 23011 10312 23020 10352
rect 23060 10312 23069 10352
rect 23011 10311 23069 10312
rect 31563 10352 31605 10361
rect 31563 10312 31564 10352
rect 31604 10312 31605 10352
rect 31563 10303 31605 10312
rect 33099 10352 33141 10361
rect 33099 10312 33100 10352
rect 33140 10312 33141 10352
rect 33099 10303 33141 10312
rect 45291 10352 45333 10361
rect 45291 10312 45292 10352
rect 45332 10312 45333 10352
rect 45291 10303 45333 10312
rect 3915 10268 3957 10277
rect 3915 10228 3916 10268
rect 3956 10228 3957 10268
rect 3915 10219 3957 10228
rect 8331 10268 8373 10277
rect 8331 10228 8332 10268
rect 8372 10228 8373 10268
rect 8331 10219 8373 10228
rect 15435 10268 15477 10277
rect 15435 10228 15436 10268
rect 15476 10228 15477 10268
rect 15435 10219 15477 10228
rect 25035 10268 25077 10277
rect 25035 10228 25036 10268
rect 25076 10228 25077 10268
rect 25035 10219 25077 10228
rect 31467 10268 31509 10277
rect 31467 10228 31468 10268
rect 31508 10228 31509 10268
rect 31467 10219 31509 10228
rect 31659 10268 31701 10277
rect 31659 10228 31660 10268
rect 31700 10228 31701 10268
rect 31659 10219 31701 10228
rect 32811 10268 32853 10277
rect 32811 10228 32812 10268
rect 32852 10228 32853 10268
rect 32811 10219 32853 10228
rect 37707 10268 37749 10277
rect 37707 10228 37708 10268
rect 37748 10228 37749 10268
rect 37707 10219 37749 10228
rect 24520 10199 24562 10208
rect 1515 10184 1557 10193
rect 1515 10144 1516 10184
rect 1556 10144 1557 10184
rect 1515 10135 1557 10144
rect 1891 10184 1949 10185
rect 1891 10144 1900 10184
rect 1940 10144 1949 10184
rect 1891 10143 1949 10144
rect 2755 10184 2813 10185
rect 2755 10144 2764 10184
rect 2804 10144 2813 10184
rect 2755 10143 2813 10144
rect 4867 10184 4925 10185
rect 4867 10144 4876 10184
rect 4916 10144 4925 10184
rect 4867 10143 4925 10144
rect 5067 10184 5109 10193
rect 5067 10144 5068 10184
rect 5108 10144 5109 10184
rect 5067 10135 5109 10144
rect 5443 10184 5501 10185
rect 5443 10144 5452 10184
rect 5492 10144 5501 10184
rect 5443 10143 5501 10144
rect 6307 10184 6365 10185
rect 6307 10144 6316 10184
rect 6356 10144 6365 10184
rect 6307 10143 6365 10144
rect 8427 10184 8469 10193
rect 8427 10144 8428 10184
rect 8468 10144 8469 10184
rect 8427 10135 8469 10144
rect 8515 10184 8573 10185
rect 8515 10144 8524 10184
rect 8564 10144 8573 10184
rect 8515 10143 8573 10144
rect 9099 10184 9141 10193
rect 9099 10144 9100 10184
rect 9140 10144 9141 10184
rect 9099 10135 9141 10144
rect 9195 10184 9237 10193
rect 9195 10144 9196 10184
rect 9236 10144 9237 10184
rect 9195 10135 9237 10144
rect 9579 10184 9621 10193
rect 9579 10144 9580 10184
rect 9620 10144 9621 10184
rect 9579 10135 9621 10144
rect 9867 10184 9909 10193
rect 9867 10144 9868 10184
rect 9908 10144 9909 10184
rect 9867 10135 9909 10144
rect 10539 10184 10581 10193
rect 10539 10144 10540 10184
rect 10580 10144 10581 10184
rect 10539 10135 10581 10144
rect 10635 10184 10677 10193
rect 10635 10144 10636 10184
rect 10676 10144 10677 10184
rect 10635 10135 10677 10144
rect 10731 10184 10773 10193
rect 10731 10144 10732 10184
rect 10772 10144 10773 10184
rect 10731 10135 10773 10144
rect 11587 10184 11645 10185
rect 11587 10144 11596 10184
rect 11636 10144 11645 10184
rect 11587 10143 11645 10144
rect 11979 10184 12021 10193
rect 11979 10144 11980 10184
rect 12020 10144 12021 10184
rect 11979 10135 12021 10144
rect 12171 10184 12213 10193
rect 12171 10144 12172 10184
rect 12212 10144 12213 10184
rect 12171 10135 12213 10144
rect 12259 10184 12317 10185
rect 12259 10144 12268 10184
rect 12308 10144 12317 10184
rect 12259 10143 12317 10144
rect 13123 10184 13181 10185
rect 13123 10144 13132 10184
rect 13172 10144 13181 10184
rect 13123 10143 13181 10144
rect 13315 10184 13373 10185
rect 13315 10144 13324 10184
rect 13364 10144 13373 10184
rect 13315 10143 13373 10144
rect 13419 10184 13461 10193
rect 13419 10144 13420 10184
rect 13460 10144 13461 10184
rect 13419 10135 13461 10144
rect 16291 10184 16349 10185
rect 16291 10144 16300 10184
rect 16340 10144 16349 10184
rect 16291 10143 16349 10144
rect 16587 10184 16629 10193
rect 16587 10144 16588 10184
rect 16628 10144 16629 10184
rect 16587 10135 16629 10144
rect 17251 10184 17309 10185
rect 17251 10144 17260 10184
rect 17300 10144 17309 10184
rect 17251 10143 17309 10144
rect 17739 10184 17781 10193
rect 17739 10144 17740 10184
rect 17780 10144 17781 10184
rect 17739 10135 17781 10144
rect 17931 10184 17973 10193
rect 17931 10144 17932 10184
rect 17972 10144 17973 10184
rect 17931 10135 17973 10144
rect 18019 10184 18077 10185
rect 18019 10144 18028 10184
rect 18068 10144 18077 10184
rect 18019 10143 18077 10144
rect 18603 10184 18645 10193
rect 18603 10144 18604 10184
rect 18644 10144 18645 10184
rect 18603 10135 18645 10144
rect 18883 10184 18941 10185
rect 18883 10144 18892 10184
rect 18932 10144 18941 10184
rect 18883 10143 18941 10144
rect 19659 10184 19701 10193
rect 19659 10144 19660 10184
rect 19700 10144 19701 10184
rect 19659 10135 19701 10144
rect 20235 10184 20277 10193
rect 20235 10144 20236 10184
rect 20276 10144 20277 10184
rect 20235 10135 20277 10144
rect 20331 10184 20373 10193
rect 20331 10144 20332 10184
rect 20372 10144 20373 10184
rect 20331 10135 20373 10144
rect 20427 10184 20469 10193
rect 20427 10144 20428 10184
rect 20468 10144 20469 10184
rect 20427 10135 20469 10144
rect 20523 10184 20565 10193
rect 20523 10144 20524 10184
rect 20564 10144 20565 10184
rect 20523 10135 20565 10144
rect 20715 10184 20757 10193
rect 20715 10144 20716 10184
rect 20756 10144 20757 10184
rect 20715 10135 20757 10144
rect 20907 10184 20949 10193
rect 20907 10144 20908 10184
rect 20948 10144 20949 10184
rect 20907 10135 20949 10144
rect 20995 10184 21053 10185
rect 20995 10144 21004 10184
rect 21044 10144 21053 10184
rect 20995 10143 21053 10144
rect 21859 10184 21917 10185
rect 21859 10144 21868 10184
rect 21908 10144 21917 10184
rect 21859 10143 21917 10144
rect 22059 10184 22101 10193
rect 22059 10144 22060 10184
rect 22100 10144 22101 10184
rect 22059 10135 22101 10144
rect 22155 10184 22197 10193
rect 22155 10144 22156 10184
rect 22196 10144 22197 10184
rect 22155 10135 22197 10144
rect 22251 10184 22293 10193
rect 22251 10144 22252 10184
rect 22292 10144 22293 10184
rect 22251 10135 22293 10144
rect 22347 10184 22389 10193
rect 22347 10144 22348 10184
rect 22388 10144 22389 10184
rect 22347 10135 22389 10144
rect 22731 10184 22773 10193
rect 22731 10144 22732 10184
rect 22772 10144 22773 10184
rect 22731 10135 22773 10144
rect 22923 10184 22965 10193
rect 22923 10144 22924 10184
rect 22964 10144 22965 10184
rect 22923 10135 22965 10144
rect 23019 10184 23061 10193
rect 23019 10144 23020 10184
rect 23060 10144 23061 10184
rect 23019 10135 23061 10144
rect 23203 10184 23261 10185
rect 23203 10144 23212 10184
rect 23252 10144 23261 10184
rect 23203 10143 23261 10144
rect 23299 10184 23357 10185
rect 23299 10144 23308 10184
rect 23348 10144 23357 10184
rect 23299 10143 23357 10144
rect 23499 10184 23541 10193
rect 23499 10144 23500 10184
rect 23540 10144 23541 10184
rect 23499 10135 23541 10144
rect 23595 10184 23637 10193
rect 23595 10144 23596 10184
rect 23636 10144 23637 10184
rect 23595 10135 23637 10144
rect 23688 10184 23746 10185
rect 23688 10144 23697 10184
rect 23737 10144 23746 10184
rect 23688 10143 23746 10144
rect 23971 10184 24029 10185
rect 23971 10144 23980 10184
rect 24020 10144 24029 10184
rect 23971 10143 24029 10144
rect 24067 10184 24125 10185
rect 24067 10144 24076 10184
rect 24116 10144 24125 10184
rect 24067 10143 24125 10144
rect 24267 10184 24309 10193
rect 24267 10144 24268 10184
rect 24308 10144 24309 10184
rect 24267 10135 24309 10144
rect 24363 10184 24405 10193
rect 24363 10144 24364 10184
rect 24404 10144 24405 10184
rect 24520 10159 24521 10199
rect 24561 10159 24562 10199
rect 24520 10150 24562 10159
rect 24843 10184 24885 10193
rect 24363 10135 24405 10144
rect 24843 10144 24844 10184
rect 24884 10144 24885 10184
rect 24843 10135 24885 10144
rect 25131 10184 25173 10193
rect 25131 10144 25132 10184
rect 25172 10144 25173 10184
rect 25131 10135 25173 10144
rect 25419 10184 25461 10193
rect 25419 10144 25420 10184
rect 25460 10144 25461 10184
rect 25419 10135 25461 10144
rect 25515 10184 25557 10193
rect 25515 10144 25516 10184
rect 25556 10144 25557 10184
rect 25515 10135 25557 10144
rect 25611 10184 25653 10193
rect 25611 10144 25612 10184
rect 25652 10144 25653 10184
rect 25611 10135 25653 10144
rect 26667 10184 26709 10193
rect 26667 10144 26668 10184
rect 26708 10144 26709 10184
rect 26667 10135 26709 10144
rect 26947 10184 27005 10185
rect 26947 10144 26956 10184
rect 26996 10144 27005 10184
rect 26947 10143 27005 10144
rect 27715 10184 27773 10185
rect 27715 10144 27724 10184
rect 27764 10144 27773 10184
rect 27715 10143 27773 10144
rect 28003 10184 28061 10185
rect 28003 10144 28012 10184
rect 28052 10144 28061 10184
rect 28003 10143 28061 10144
rect 29443 10184 29501 10185
rect 29443 10144 29452 10184
rect 29492 10144 29501 10184
rect 29443 10143 29501 10144
rect 29643 10184 29685 10193
rect 29643 10144 29644 10184
rect 29684 10144 29685 10184
rect 29643 10135 29685 10144
rect 29835 10184 29877 10193
rect 29835 10144 29836 10184
rect 29876 10144 29877 10184
rect 29835 10135 29877 10144
rect 30211 10184 30269 10185
rect 30211 10144 30220 10184
rect 30260 10144 30269 10184
rect 30211 10143 30269 10144
rect 30403 10184 30461 10185
rect 30403 10144 30412 10184
rect 30452 10144 30461 10184
rect 30403 10143 30461 10144
rect 30691 10184 30749 10185
rect 30691 10144 30700 10184
rect 30740 10144 30749 10184
rect 30691 10143 30749 10144
rect 31363 10184 31421 10185
rect 31363 10144 31372 10184
rect 31412 10144 31421 10184
rect 31363 10143 31421 10144
rect 31755 10184 31797 10193
rect 31755 10144 31756 10184
rect 31796 10144 31797 10184
rect 31755 10135 31797 10144
rect 31981 10191 32023 10200
rect 35595 10199 35637 10208
rect 31981 10151 31982 10191
rect 32022 10151 32023 10191
rect 31981 10142 32023 10151
rect 32139 10184 32181 10193
rect 32139 10144 32140 10184
rect 32180 10144 32181 10184
rect 32139 10135 32181 10144
rect 32235 10184 32277 10193
rect 32235 10144 32236 10184
rect 32276 10144 32277 10184
rect 32235 10135 32277 10144
rect 32419 10184 32477 10185
rect 32419 10144 32428 10184
rect 32468 10144 32477 10184
rect 32419 10143 32477 10144
rect 32515 10184 32573 10185
rect 32515 10144 32524 10184
rect 32564 10144 32573 10184
rect 32515 10143 32573 10144
rect 32715 10184 32757 10193
rect 32715 10144 32716 10184
rect 32756 10144 32757 10184
rect 32715 10135 32757 10144
rect 32907 10184 32949 10193
rect 32907 10144 32908 10184
rect 32948 10144 32949 10184
rect 32907 10135 32949 10144
rect 33099 10184 33141 10193
rect 33099 10144 33100 10184
rect 33140 10144 33141 10184
rect 33099 10135 33141 10144
rect 33291 10184 33333 10193
rect 33291 10144 33292 10184
rect 33332 10144 33333 10184
rect 33291 10135 33333 10144
rect 33571 10184 33629 10185
rect 33571 10144 33580 10184
rect 33620 10144 33629 10184
rect 33571 10143 33629 10144
rect 33867 10184 33909 10193
rect 33867 10144 33868 10184
rect 33908 10144 33909 10184
rect 33867 10135 33909 10144
rect 34155 10184 34197 10193
rect 34155 10144 34156 10184
rect 34196 10144 34197 10184
rect 34155 10135 34197 10144
rect 34347 10184 34389 10193
rect 34347 10144 34348 10184
rect 34388 10144 34389 10184
rect 34347 10135 34389 10144
rect 34539 10184 34581 10193
rect 34539 10144 34540 10184
rect 34580 10144 34581 10184
rect 34539 10135 34581 10144
rect 34635 10184 34677 10193
rect 34635 10144 34636 10184
rect 34676 10144 34677 10184
rect 34635 10135 34677 10144
rect 34827 10184 34869 10193
rect 34827 10144 34828 10184
rect 34868 10144 34869 10184
rect 34827 10135 34869 10144
rect 34923 10184 34965 10193
rect 34923 10144 34924 10184
rect 34964 10144 34965 10184
rect 34923 10135 34965 10144
rect 35019 10184 35061 10193
rect 35019 10144 35020 10184
rect 35060 10144 35061 10184
rect 35019 10135 35061 10144
rect 35299 10184 35357 10185
rect 35299 10144 35308 10184
rect 35348 10144 35357 10184
rect 35299 10143 35357 10144
rect 35395 10184 35453 10185
rect 35395 10144 35404 10184
rect 35444 10144 35453 10184
rect 35595 10159 35596 10199
rect 35636 10159 35637 10199
rect 35595 10150 35637 10159
rect 35691 10184 35733 10193
rect 35395 10143 35453 10144
rect 35691 10144 35692 10184
rect 35732 10144 35733 10184
rect 35691 10135 35733 10144
rect 35784 10184 35842 10185
rect 35784 10144 35793 10184
rect 35833 10144 35842 10184
rect 35784 10143 35842 10144
rect 36267 10184 36309 10193
rect 36267 10144 36268 10184
rect 36308 10144 36309 10184
rect 36267 10135 36309 10144
rect 36363 10184 36405 10193
rect 36363 10144 36364 10184
rect 36404 10144 36405 10184
rect 36363 10135 36405 10144
rect 36555 10184 36597 10193
rect 36555 10144 36556 10184
rect 36596 10144 36597 10184
rect 36555 10135 36597 10144
rect 36747 10184 36789 10193
rect 36747 10144 36748 10184
rect 36788 10144 36789 10184
rect 36747 10135 36789 10144
rect 36843 10184 36885 10193
rect 36843 10144 36844 10184
rect 36884 10144 36885 10184
rect 36843 10135 36885 10144
rect 37131 10184 37173 10193
rect 37131 10144 37132 10184
rect 37172 10144 37173 10184
rect 37131 10135 37173 10144
rect 37227 10184 37269 10193
rect 37227 10144 37228 10184
rect 37268 10144 37269 10184
rect 37227 10135 37269 10144
rect 37323 10184 37365 10193
rect 37323 10144 37324 10184
rect 37364 10144 37365 10184
rect 37323 10135 37365 10144
rect 37515 10184 37557 10193
rect 37515 10144 37516 10184
rect 37556 10144 37557 10184
rect 37515 10135 37557 10144
rect 37803 10184 37845 10193
rect 37803 10144 37804 10184
rect 37844 10144 37845 10184
rect 37803 10135 37845 10144
rect 37987 10184 38045 10185
rect 37987 10144 37996 10184
rect 38036 10144 38045 10184
rect 37987 10143 38045 10144
rect 39811 10184 39869 10185
rect 39811 10144 39820 10184
rect 39860 10144 39869 10184
rect 39811 10143 39869 10144
rect 41347 10184 41405 10185
rect 41347 10144 41356 10184
rect 41396 10144 41405 10184
rect 41347 10143 41405 10144
rect 42211 10184 42269 10185
rect 42211 10144 42220 10184
rect 42260 10144 42269 10184
rect 42211 10143 42269 10144
rect 42603 10184 42645 10193
rect 42603 10144 42604 10184
rect 42644 10144 42645 10184
rect 42603 10135 42645 10144
rect 43179 10184 43221 10193
rect 43179 10144 43180 10184
rect 43220 10144 43221 10184
rect 43179 10135 43221 10144
rect 43267 10184 43325 10185
rect 43267 10144 43276 10184
rect 43316 10144 43325 10184
rect 43267 10143 43325 10144
rect 43555 10184 43613 10185
rect 43555 10144 43564 10184
rect 43604 10144 43613 10184
rect 43555 10143 43613 10144
rect 44419 10184 44477 10185
rect 44419 10144 44428 10184
rect 44468 10144 44477 10184
rect 44419 10143 44477 10144
rect 45291 10184 45333 10193
rect 45291 10144 45292 10184
rect 45332 10144 45333 10184
rect 45291 10135 45333 10144
rect 45483 10184 45525 10193
rect 45483 10144 45484 10184
rect 45524 10144 45525 10184
rect 45483 10135 45525 10144
rect 45667 10184 45725 10185
rect 45667 10144 45676 10184
rect 45716 10144 45725 10184
rect 45667 10143 45725 10144
rect 46627 10184 46685 10185
rect 46627 10144 46636 10184
rect 46676 10144 46685 10184
rect 46627 10143 46685 10144
rect 48163 10184 48221 10185
rect 48163 10144 48172 10184
rect 48212 10144 48221 10184
rect 48163 10143 48221 10144
rect 49027 10184 49085 10185
rect 49027 10144 49036 10184
rect 49076 10144 49085 10184
rect 49027 10143 49085 10144
rect 49419 10184 49461 10193
rect 49419 10144 49420 10184
rect 49460 10144 49461 10184
rect 49419 10135 49461 10144
rect 12075 10100 12117 10109
rect 12075 10060 12076 10100
rect 12116 10060 12117 10100
rect 12075 10051 12117 10060
rect 18507 10100 18549 10109
rect 18507 10060 18508 10100
rect 18548 10060 18549 10100
rect 18507 10051 18549 10060
rect 19371 10100 19413 10109
rect 19371 10060 19372 10100
rect 19412 10060 19413 10100
rect 19371 10051 19413 10060
rect 20811 10100 20853 10109
rect 20811 10060 20812 10100
rect 20852 10060 20853 10100
rect 20811 10051 20853 10060
rect 25323 10100 25365 10109
rect 25323 10060 25324 10100
rect 25364 10060 25365 10100
rect 25323 10051 25365 10060
rect 26571 10100 26613 10109
rect 26571 10060 26572 10100
rect 26612 10060 26613 10100
rect 26571 10051 26613 10060
rect 28195 10100 28253 10101
rect 28195 10060 28204 10100
rect 28244 10060 28253 10100
rect 28195 10059 28253 10060
rect 29739 10100 29781 10109
rect 29739 10060 29740 10100
rect 29780 10060 29781 10100
rect 29739 10051 29781 10060
rect 30507 10100 30549 10109
rect 30507 10060 30508 10100
rect 30548 10060 30549 10100
rect 30507 10051 30549 10060
rect 34059 10100 34101 10109
rect 34059 10060 34060 10100
rect 34100 10060 34101 10100
rect 34059 10051 34101 10060
rect 38667 10100 38709 10109
rect 38667 10060 38668 10100
rect 38708 10060 38709 10100
rect 38667 10051 38709 10060
rect 643 10016 701 10017
rect 643 9976 652 10016
rect 692 9976 701 10016
rect 643 9975 701 9976
rect 8427 10016 8469 10025
rect 8427 9976 8428 10016
rect 8468 9976 8469 10016
rect 8427 9967 8469 9976
rect 9379 10016 9437 10017
rect 9379 9976 9388 10016
rect 9428 9976 9437 10016
rect 9379 9975 9437 9976
rect 10435 10016 10493 10017
rect 10435 9976 10444 10016
rect 10484 9976 10493 10016
rect 10435 9975 10493 9976
rect 10915 10016 10973 10017
rect 10915 9976 10924 10016
rect 10964 9976 10973 10016
rect 10915 9975 10973 9976
rect 12451 10016 12509 10017
rect 12451 9976 12460 10016
rect 12500 9976 12509 10016
rect 12451 9975 12509 9976
rect 17827 10016 17885 10017
rect 17827 9976 17836 10016
rect 17876 9976 17885 10016
rect 17827 9975 17885 9976
rect 19171 10016 19229 10017
rect 19171 9976 19180 10016
rect 19220 9976 19229 10016
rect 19171 9975 19229 9976
rect 23395 10016 23453 10017
rect 23395 9976 23404 10016
rect 23444 9976 23453 10016
rect 23395 9975 23453 9976
rect 29355 10016 29397 10025
rect 29355 9976 29356 10016
rect 29396 9976 29397 10016
rect 29355 9967 29397 9976
rect 32035 10016 32093 10017
rect 32035 9976 32044 10016
rect 32084 9976 32093 10016
rect 32035 9975 32093 9976
rect 35107 10016 35165 10017
rect 35107 9976 35116 10016
rect 35156 9976 35165 10016
rect 35107 9975 35165 9976
rect 35587 10016 35645 10017
rect 35587 9976 35596 10016
rect 35636 9976 35645 10016
rect 35587 9975 35645 9976
rect 36067 10016 36125 10017
rect 36067 9976 36076 10016
rect 36116 9976 36125 10016
rect 36067 9975 36125 9976
rect 36651 10016 36693 10025
rect 36651 9976 36652 10016
rect 36692 9976 36693 10016
rect 36651 9967 36693 9976
rect 37027 10016 37085 10017
rect 37027 9976 37036 10016
rect 37076 9976 37085 10016
rect 37027 9975 37085 9976
rect 43371 10012 43413 10021
rect 43371 9972 43372 10012
rect 43412 9972 43413 10012
rect 45091 10016 45149 10017
rect 45091 9976 45100 10016
rect 45140 9976 45149 10016
rect 45091 9975 45149 9976
rect 43371 9963 43413 9972
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 643 9680 701 9681
rect 643 9640 652 9680
rect 692 9640 701 9680
rect 643 9639 701 9640
rect 5059 9680 5117 9681
rect 5059 9640 5068 9680
rect 5108 9640 5117 9680
rect 5059 9639 5117 9640
rect 7083 9680 7125 9689
rect 7083 9640 7084 9680
rect 7124 9640 7125 9680
rect 7083 9631 7125 9640
rect 9475 9680 9533 9681
rect 9475 9640 9484 9680
rect 9524 9640 9533 9680
rect 9475 9639 9533 9640
rect 9771 9680 9813 9689
rect 9771 9640 9772 9680
rect 9812 9640 9813 9680
rect 9771 9631 9813 9640
rect 12643 9680 12701 9681
rect 12643 9640 12652 9680
rect 12692 9640 12701 9680
rect 12643 9639 12701 9640
rect 16003 9680 16061 9681
rect 16003 9640 16012 9680
rect 16052 9640 16061 9680
rect 16003 9639 16061 9640
rect 16867 9680 16925 9681
rect 16867 9640 16876 9680
rect 16916 9640 16925 9680
rect 16867 9639 16925 9640
rect 21963 9680 22005 9689
rect 21963 9640 21964 9680
rect 22004 9640 22005 9680
rect 21963 9631 22005 9640
rect 24643 9680 24701 9681
rect 24643 9640 24652 9680
rect 24692 9640 24701 9680
rect 24643 9639 24701 9640
rect 25123 9680 25181 9681
rect 25123 9640 25132 9680
rect 25172 9640 25181 9680
rect 25123 9639 25181 9640
rect 27051 9680 27093 9689
rect 27051 9640 27052 9680
rect 27092 9640 27093 9680
rect 27051 9631 27093 9640
rect 30795 9680 30837 9689
rect 30795 9640 30796 9680
rect 30836 9640 30837 9680
rect 30795 9631 30837 9640
rect 37323 9680 37365 9689
rect 37323 9640 37324 9680
rect 37364 9640 37365 9680
rect 37323 9631 37365 9640
rect 44715 9680 44757 9689
rect 44715 9640 44716 9680
rect 44756 9640 44757 9680
rect 44715 9631 44757 9640
rect 48163 9680 48221 9681
rect 48163 9640 48172 9680
rect 48212 9640 48221 9680
rect 48163 9639 48221 9640
rect 9379 9596 9437 9597
rect 9379 9556 9388 9596
rect 9428 9556 9437 9596
rect 9379 9555 9437 9556
rect 10251 9596 10293 9605
rect 10251 9556 10252 9596
rect 10292 9556 10293 9596
rect 10251 9547 10293 9556
rect 16491 9596 16533 9605
rect 16491 9556 16492 9596
rect 16532 9556 16533 9596
rect 16491 9547 16533 9556
rect 23683 9596 23741 9597
rect 23683 9556 23692 9596
rect 23732 9556 23741 9596
rect 23683 9555 23741 9556
rect 27907 9596 27965 9597
rect 27907 9556 27916 9596
rect 27956 9556 27965 9596
rect 27907 9555 27965 9556
rect 29547 9596 29589 9605
rect 29547 9556 29548 9596
rect 29588 9556 29589 9596
rect 29547 9547 29589 9556
rect 30219 9596 30261 9605
rect 30219 9556 30220 9596
rect 30260 9556 30261 9596
rect 30219 9547 30261 9556
rect 1707 9512 1749 9521
rect 1707 9472 1708 9512
rect 1748 9472 1749 9512
rect 1707 9463 1749 9472
rect 1899 9512 1941 9521
rect 1899 9472 1900 9512
rect 1940 9472 1941 9512
rect 1899 9463 1941 9472
rect 2275 9512 2333 9513
rect 2275 9472 2284 9512
rect 2324 9472 2333 9512
rect 2275 9471 2333 9472
rect 2371 9512 2429 9513
rect 2371 9472 2380 9512
rect 2420 9472 2429 9512
rect 2371 9471 2429 9472
rect 3523 9512 3581 9513
rect 3523 9472 3532 9512
rect 3572 9472 3581 9512
rect 3523 9471 3581 9472
rect 4195 9512 4253 9513
rect 4195 9472 4204 9512
rect 4244 9472 4253 9512
rect 4195 9471 4253 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4779 9512 4821 9521
rect 4779 9472 4780 9512
rect 4820 9472 4821 9512
rect 4779 9463 4821 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 5731 9512 5789 9513
rect 5731 9472 5740 9512
rect 5780 9472 5789 9512
rect 5731 9471 5789 9472
rect 5931 9512 5973 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7179 9512 7221 9521
rect 7179 9472 7180 9512
rect 7220 9472 7221 9512
rect 7179 9463 7221 9472
rect 7275 9512 7317 9521
rect 7275 9472 7276 9512
rect 7316 9472 7317 9512
rect 7275 9463 7317 9472
rect 7459 9512 7517 9513
rect 7459 9472 7468 9512
rect 7508 9472 7517 9512
rect 7459 9471 7517 9472
rect 7563 9512 7605 9521
rect 7563 9472 7564 9512
rect 7604 9472 7605 9512
rect 7563 9463 7605 9472
rect 8331 9512 8373 9521
rect 8331 9472 8332 9512
rect 8372 9472 8373 9512
rect 8331 9463 8373 9472
rect 8995 9512 9053 9513
rect 8995 9472 9004 9512
rect 9044 9472 9053 9512
rect 8995 9471 9053 9472
rect 9195 9512 9237 9521
rect 9195 9472 9196 9512
rect 9236 9472 9237 9512
rect 9195 9463 9237 9472
rect 9291 9512 9333 9521
rect 9291 9472 9292 9512
rect 9332 9472 9333 9512
rect 9291 9463 9333 9472
rect 9763 9512 9821 9513
rect 9763 9472 9772 9512
rect 9812 9472 9821 9512
rect 9763 9471 9821 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10051 9512 10109 9513
rect 10051 9472 10060 9512
rect 10100 9472 10109 9512
rect 10051 9471 10109 9472
rect 10627 9512 10685 9513
rect 10627 9472 10636 9512
rect 10676 9472 10685 9512
rect 10627 9471 10685 9472
rect 11491 9512 11549 9513
rect 11491 9472 11500 9512
rect 11540 9472 11549 9512
rect 11491 9471 11549 9472
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13987 9512 14045 9513
rect 13987 9472 13996 9512
rect 14036 9472 14045 9512
rect 13987 9471 14045 9472
rect 14851 9512 14909 9513
rect 14851 9472 14860 9512
rect 14900 9472 14909 9512
rect 14851 9471 14909 9472
rect 16387 9512 16445 9513
rect 16387 9472 16396 9512
rect 16436 9472 16445 9512
rect 16387 9471 16445 9472
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 16779 9512 16821 9521
rect 16779 9472 16780 9512
rect 16820 9472 16821 9512
rect 16779 9463 16821 9472
rect 16971 9512 17013 9521
rect 16971 9472 16972 9512
rect 17012 9472 17013 9512
rect 16971 9463 17013 9472
rect 17059 9512 17117 9513
rect 17059 9472 17068 9512
rect 17108 9472 17117 9512
rect 17059 9471 17117 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17451 9512 17493 9521
rect 17451 9472 17452 9512
rect 17492 9472 17493 9512
rect 17451 9463 17493 9472
rect 17539 9512 17597 9513
rect 17539 9472 17548 9512
rect 17588 9472 17597 9512
rect 17539 9471 17597 9472
rect 17731 9512 17789 9513
rect 17731 9472 17740 9512
rect 17780 9472 17789 9512
rect 17731 9471 17789 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 19083 9512 19125 9521
rect 19083 9472 19084 9512
rect 19124 9472 19125 9512
rect 19083 9463 19125 9472
rect 20331 9512 20373 9521
rect 20331 9472 20332 9512
rect 20372 9472 20373 9512
rect 20331 9463 20373 9472
rect 20523 9512 20565 9521
rect 20523 9472 20524 9512
rect 20564 9472 20565 9512
rect 20523 9463 20565 9472
rect 20707 9512 20765 9513
rect 20707 9472 20716 9512
rect 20756 9472 20765 9512
rect 20707 9471 20765 9472
rect 20811 9512 20853 9521
rect 20811 9472 20812 9512
rect 20852 9472 20853 9512
rect 20811 9463 20853 9472
rect 21003 9512 21045 9521
rect 21003 9472 21004 9512
rect 21044 9472 21045 9512
rect 21003 9463 21045 9472
rect 21963 9512 22005 9521
rect 21963 9472 21964 9512
rect 22004 9472 22005 9512
rect 21963 9463 22005 9472
rect 22051 9512 22109 9513
rect 22051 9472 22060 9512
rect 22100 9472 22109 9512
rect 22051 9471 22109 9472
rect 22443 9512 22485 9521
rect 22443 9472 22444 9512
rect 22484 9472 22485 9512
rect 22443 9463 22485 9472
rect 22539 9512 22581 9521
rect 22539 9472 22540 9512
rect 22580 9472 22581 9512
rect 22539 9463 22581 9472
rect 22635 9512 22677 9521
rect 22635 9472 22636 9512
rect 22676 9472 22677 9512
rect 22635 9463 22677 9472
rect 22731 9512 22773 9521
rect 22731 9472 22732 9512
rect 22772 9472 22773 9512
rect 22731 9463 22773 9472
rect 23203 9512 23261 9513
rect 23203 9472 23212 9512
rect 23252 9472 23261 9512
rect 23203 9471 23261 9472
rect 23587 9512 23645 9513
rect 23587 9472 23596 9512
rect 23636 9472 23645 9512
rect 23587 9471 23645 9472
rect 23979 9512 24021 9521
rect 23979 9472 23980 9512
rect 24020 9472 24021 9512
rect 23979 9463 24021 9472
rect 24171 9512 24213 9521
rect 24171 9472 24172 9512
rect 24212 9472 24213 9512
rect 24171 9463 24213 9472
rect 24363 9512 24405 9521
rect 24363 9472 24364 9512
rect 24404 9472 24405 9512
rect 24363 9463 24405 9472
rect 24459 9512 24501 9521
rect 24459 9472 24460 9512
rect 24500 9472 24501 9512
rect 24459 9463 24501 9472
rect 24843 9512 24885 9521
rect 24843 9472 24844 9512
rect 24884 9472 24885 9512
rect 24843 9463 24885 9472
rect 24939 9512 24981 9521
rect 24939 9472 24940 9512
rect 24980 9472 24981 9512
rect 24939 9463 24981 9472
rect 25035 9512 25077 9521
rect 25035 9472 25036 9512
rect 25076 9472 25077 9512
rect 25035 9463 25077 9472
rect 25315 9512 25373 9513
rect 25315 9472 25324 9512
rect 25364 9472 25373 9512
rect 25315 9471 25373 9472
rect 25515 9512 25557 9521
rect 25515 9472 25516 9512
rect 25556 9472 25557 9512
rect 25515 9463 25557 9472
rect 26955 9512 26997 9521
rect 26955 9472 26956 9512
rect 26996 9472 26997 9512
rect 26955 9463 26997 9472
rect 27243 9512 27285 9521
rect 27243 9472 27244 9512
rect 27284 9472 27285 9512
rect 27243 9463 27285 9472
rect 27427 9512 27485 9513
rect 27427 9472 27436 9512
rect 27476 9472 27485 9512
rect 27427 9471 27485 9472
rect 27811 9512 27869 9513
rect 27811 9472 27820 9512
rect 27860 9472 27869 9512
rect 27811 9471 27869 9472
rect 28491 9512 28533 9521
rect 28491 9472 28492 9512
rect 28532 9472 28533 9512
rect 28491 9463 28533 9472
rect 28579 9512 28637 9513
rect 28579 9472 28588 9512
rect 28628 9472 28637 9512
rect 28579 9471 28637 9472
rect 29643 9512 29685 9521
rect 29643 9472 29644 9512
rect 29684 9472 29685 9512
rect 29643 9463 29685 9472
rect 29923 9512 29981 9513
rect 29923 9472 29932 9512
rect 29972 9472 29981 9512
rect 29923 9471 29981 9472
rect 30315 9512 30357 9521
rect 30315 9472 30316 9512
rect 30356 9472 30357 9512
rect 30315 9463 30357 9472
rect 30411 9512 30453 9521
rect 30411 9472 30412 9512
rect 30452 9472 30453 9512
rect 30411 9463 30453 9472
rect 30507 9512 30549 9521
rect 30507 9472 30508 9512
rect 30548 9472 30549 9512
rect 30507 9463 30549 9472
rect 30699 9512 30741 9521
rect 30699 9472 30700 9512
rect 30740 9472 30741 9512
rect 30699 9463 30741 9472
rect 30891 9512 30933 9521
rect 30891 9472 30892 9512
rect 30932 9472 30933 9512
rect 30891 9463 30933 9472
rect 31275 9512 31317 9521
rect 31275 9472 31276 9512
rect 31316 9472 31317 9512
rect 31275 9463 31317 9472
rect 31651 9512 31709 9513
rect 31651 9472 31660 9512
rect 31700 9472 31709 9512
rect 31651 9471 31709 9472
rect 31939 9512 31997 9513
rect 31939 9472 31948 9512
rect 31988 9472 31997 9512
rect 31939 9471 31997 9472
rect 34155 9512 34197 9521
rect 34155 9472 34156 9512
rect 34196 9472 34197 9512
rect 34155 9463 34197 9472
rect 34443 9512 34485 9521
rect 34443 9472 34444 9512
rect 34484 9472 34485 9512
rect 34443 9463 34485 9472
rect 34819 9512 34877 9513
rect 34819 9472 34828 9512
rect 34868 9472 34877 9512
rect 34819 9471 34877 9472
rect 34923 9512 34965 9521
rect 34923 9472 34924 9512
rect 34964 9472 34965 9512
rect 34923 9463 34965 9472
rect 35403 9512 35445 9521
rect 35403 9472 35404 9512
rect 35444 9472 35445 9512
rect 35403 9463 35445 9472
rect 35499 9512 35541 9521
rect 35499 9472 35500 9512
rect 35540 9472 35541 9512
rect 35499 9463 35541 9472
rect 35595 9512 35637 9521
rect 35595 9472 35596 9512
rect 35636 9472 35637 9512
rect 35595 9463 35637 9472
rect 35691 9512 35733 9521
rect 35691 9472 35692 9512
rect 35732 9472 35733 9512
rect 35691 9463 35733 9472
rect 35883 9512 35925 9521
rect 35883 9472 35884 9512
rect 35924 9472 35925 9512
rect 35883 9463 35925 9472
rect 36171 9512 36213 9521
rect 36171 9472 36172 9512
rect 36212 9472 36213 9512
rect 36171 9463 36213 9472
rect 37411 9512 37469 9513
rect 37411 9472 37420 9512
rect 37460 9472 37469 9512
rect 37411 9471 37469 9472
rect 38179 9512 38237 9513
rect 38179 9472 38188 9512
rect 38228 9472 38237 9512
rect 38179 9471 38237 9472
rect 38283 9512 38325 9521
rect 38283 9472 38284 9512
rect 38324 9472 38325 9512
rect 38283 9463 38325 9472
rect 38467 9512 38525 9513
rect 38467 9472 38476 9512
rect 38516 9472 38525 9512
rect 38467 9471 38525 9472
rect 38859 9512 38901 9521
rect 38859 9472 38860 9512
rect 38900 9472 38901 9512
rect 38859 9463 38901 9472
rect 39051 9512 39093 9521
rect 39051 9472 39052 9512
rect 39092 9472 39093 9512
rect 39051 9463 39093 9472
rect 39427 9512 39485 9513
rect 39427 9472 39436 9512
rect 39476 9472 39485 9512
rect 39427 9471 39485 9472
rect 40291 9512 40349 9513
rect 40291 9472 40300 9512
rect 40340 9472 40349 9512
rect 40291 9471 40349 9472
rect 41451 9512 41493 9521
rect 41451 9472 41452 9512
rect 41492 9472 41493 9512
rect 41451 9463 41493 9472
rect 42115 9512 42173 9513
rect 42115 9472 42124 9512
rect 42164 9472 42173 9512
rect 42115 9471 42173 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43083 9512 43125 9521
rect 43083 9472 43084 9512
rect 43124 9472 43125 9512
rect 43083 9463 43125 9472
rect 43275 9512 43317 9521
rect 43275 9472 43276 9512
rect 43316 9472 43317 9512
rect 43275 9463 43317 9472
rect 44131 9512 44189 9513
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44131 9471 44189 9472
rect 44419 9512 44477 9513
rect 44419 9472 44428 9512
rect 44468 9472 44477 9512
rect 44419 9471 44477 9472
rect 44611 9512 44669 9513
rect 44611 9472 44620 9512
rect 44660 9472 44669 9512
rect 44611 9471 44669 9472
rect 44899 9512 44957 9513
rect 44899 9472 44908 9512
rect 44948 9472 44957 9512
rect 44899 9471 44957 9472
rect 45187 9512 45245 9513
rect 45187 9472 45196 9512
rect 45236 9472 45245 9512
rect 45187 9471 45245 9472
rect 46051 9512 46109 9513
rect 46051 9472 46060 9512
rect 46100 9472 46109 9512
rect 46051 9471 46109 9472
rect 47787 9512 47829 9521
rect 47787 9472 47788 9512
rect 47828 9472 47829 9512
rect 47787 9463 47829 9472
rect 48835 9512 48893 9513
rect 48835 9472 48844 9512
rect 48884 9472 48893 9512
rect 48835 9471 48893 9472
rect 7659 9438 7701 9447
rect 2083 9428 2141 9429
rect 2083 9388 2092 9428
rect 2132 9388 2141 9428
rect 7659 9398 7660 9438
rect 7700 9398 7701 9438
rect 7659 9389 7701 9398
rect 21867 9428 21909 9437
rect 2083 9387 2141 9388
rect 21867 9388 21868 9428
rect 21908 9388 21909 9428
rect 21867 9379 21909 9388
rect 28395 9428 28437 9437
rect 28395 9388 28396 9428
rect 28436 9388 28437 9428
rect 28395 9379 28437 9388
rect 31371 9428 31413 9437
rect 31371 9388 31372 9428
rect 31412 9388 31413 9428
rect 31371 9379 31413 9388
rect 31563 9428 31605 9437
rect 31563 9388 31564 9428
rect 31604 9388 31605 9428
rect 31563 9379 31605 9388
rect 35019 9428 35061 9437
rect 35019 9388 35020 9428
rect 35060 9388 35061 9428
rect 35019 9379 35061 9388
rect 38571 9428 38613 9437
rect 38571 9388 38572 9428
rect 38612 9388 38613 9428
rect 38571 9379 38613 9388
rect 38763 9428 38805 9437
rect 38763 9388 38764 9428
rect 38804 9388 38805 9428
rect 38763 9379 38805 9388
rect 41731 9428 41789 9429
rect 41731 9388 41740 9428
rect 41780 9388 41789 9428
rect 41731 9387 41789 9388
rect 47019 9428 47061 9437
rect 47019 9388 47020 9428
rect 47060 9388 47061 9428
rect 47019 9379 47061 9388
rect 1515 9344 1557 9353
rect 1515 9304 1516 9344
rect 1556 9304 1557 9344
rect 1515 9295 1557 9304
rect 4011 9344 4053 9353
rect 4011 9304 4012 9344
rect 4052 9304 4053 9344
rect 4011 9295 4053 9304
rect 4867 9344 4925 9345
rect 4867 9304 4876 9344
rect 4916 9304 4925 9344
rect 4867 9303 4925 9304
rect 7755 9344 7797 9353
rect 7755 9304 7756 9344
rect 7796 9304 7797 9344
rect 7755 9295 7797 9304
rect 9283 9344 9341 9345
rect 9283 9304 9292 9344
rect 9332 9304 9341 9344
rect 9283 9303 9341 9304
rect 18027 9344 18069 9353
rect 18027 9304 18028 9344
rect 18068 9304 18069 9344
rect 18027 9295 18069 9304
rect 18891 9344 18933 9353
rect 18891 9304 18892 9344
rect 18932 9304 18933 9344
rect 18891 9295 18933 9304
rect 21771 9344 21813 9353
rect 21771 9304 21772 9344
rect 21812 9304 21813 9344
rect 21771 9295 21813 9304
rect 22243 9344 22301 9345
rect 22243 9304 22252 9344
rect 22292 9304 22301 9344
rect 22243 9303 22301 9304
rect 28203 9344 28245 9353
rect 28203 9304 28204 9344
rect 28244 9304 28245 9344
rect 28203 9295 28245 9304
rect 28299 9344 28341 9353
rect 28299 9304 28300 9344
rect 28340 9304 28341 9344
rect 28299 9295 28341 9304
rect 29251 9344 29309 9345
rect 29251 9304 29260 9344
rect 29300 9304 29309 9344
rect 29251 9303 29309 9304
rect 31467 9344 31509 9353
rect 31467 9304 31468 9344
rect 31508 9304 31509 9344
rect 31467 9295 31509 9304
rect 32235 9344 32277 9353
rect 32235 9304 32236 9344
rect 32276 9304 32277 9344
rect 32235 9295 32277 9304
rect 34443 9344 34485 9353
rect 34443 9304 34444 9344
rect 34484 9304 34485 9344
rect 34443 9295 34485 9304
rect 35115 9344 35157 9353
rect 35115 9304 35116 9344
rect 35156 9304 35157 9344
rect 35115 9295 35157 9304
rect 35883 9344 35925 9353
rect 35883 9304 35884 9344
rect 35924 9304 35925 9344
rect 35883 9295 35925 9304
rect 38667 9344 38709 9353
rect 38667 9304 38668 9344
rect 38708 9304 38709 9344
rect 38667 9295 38709 9304
rect 43179 9344 43221 9353
rect 43179 9304 43180 9344
rect 43220 9304 43221 9344
rect 43179 9295 43221 9304
rect 1899 9260 1941 9269
rect 1899 9220 1900 9260
rect 1940 9220 1941 9260
rect 1899 9211 1941 9220
rect 2851 9260 2909 9261
rect 2851 9220 2860 9260
rect 2900 9220 2909 9260
rect 2851 9219 2909 9220
rect 5931 9260 5973 9269
rect 5931 9220 5932 9260
rect 5972 9220 5973 9260
rect 5931 9211 5973 9220
rect 7851 9260 7893 9269
rect 7851 9220 7852 9260
rect 7892 9220 7893 9260
rect 7851 9211 7893 9220
rect 17259 9260 17301 9269
rect 17259 9220 17260 9260
rect 17300 9220 17301 9260
rect 17259 9211 17301 9220
rect 20331 9260 20373 9269
rect 20331 9220 20332 9260
rect 20372 9220 20373 9260
rect 20331 9211 20373 9220
rect 21003 9260 21045 9269
rect 21003 9220 21004 9260
rect 21044 9220 21045 9260
rect 21003 9211 21045 9220
rect 24171 9260 24213 9269
rect 24171 9220 24172 9260
rect 24212 9220 24213 9260
rect 24171 9211 24213 9220
rect 25419 9260 25461 9269
rect 25419 9220 25420 9260
rect 25460 9220 25461 9260
rect 25419 9211 25461 9220
rect 32427 9260 32469 9269
rect 32427 9220 32428 9260
rect 32468 9220 32469 9260
rect 32427 9211 32469 9220
rect 35211 9260 35253 9269
rect 35211 9220 35212 9260
rect 35252 9220 35253 9260
rect 35211 9211 35253 9220
rect 42787 9260 42845 9261
rect 42787 9220 42796 9260
rect 42836 9220 42845 9260
rect 42787 9219 42845 9220
rect 43459 9260 43517 9261
rect 43459 9220 43468 9260
rect 43508 9220 43517 9260
rect 43459 9219 43517 9220
rect 45859 9260 45917 9261
rect 45859 9220 45868 9260
rect 45908 9220 45917 9260
rect 45859 9219 45917 9220
rect 46723 9260 46781 9261
rect 46723 9220 46732 9260
rect 46772 9220 46781 9260
rect 46723 9219 46781 9220
rect 48163 9260 48221 9261
rect 48163 9220 48172 9260
rect 48212 9220 48221 9260
rect 48163 9219 48221 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 8907 8924 8949 8933
rect 8907 8884 8908 8924
rect 8948 8884 8949 8924
rect 8907 8875 8949 8884
rect 17163 8924 17205 8933
rect 17163 8884 17164 8924
rect 17204 8884 17205 8924
rect 17163 8875 17205 8884
rect 18315 8924 18357 8933
rect 18315 8884 18316 8924
rect 18356 8884 18357 8924
rect 18315 8875 18357 8884
rect 22827 8924 22869 8933
rect 22827 8884 22828 8924
rect 22868 8884 22869 8924
rect 22827 8875 22869 8884
rect 24939 8924 24981 8933
rect 24939 8884 24940 8924
rect 24980 8884 24981 8924
rect 24939 8875 24981 8884
rect 49035 8924 49077 8933
rect 49035 8884 49036 8924
rect 49076 8884 49077 8924
rect 49035 8875 49077 8884
rect 3723 8840 3765 8849
rect 3723 8800 3724 8840
rect 3764 8800 3765 8840
rect 3723 8791 3765 8800
rect 11403 8840 11445 8849
rect 11403 8800 11404 8840
rect 11444 8800 11445 8840
rect 11403 8791 11445 8800
rect 12171 8840 12213 8849
rect 12171 8800 12172 8840
rect 12212 8800 12213 8840
rect 12171 8791 12213 8800
rect 16491 8840 16533 8849
rect 16491 8800 16492 8840
rect 16532 8800 16533 8840
rect 16491 8791 16533 8800
rect 20427 8840 20469 8849
rect 20427 8800 20428 8840
rect 20468 8800 20469 8840
rect 20427 8791 20469 8800
rect 21963 8840 22005 8849
rect 21963 8800 21964 8840
rect 22004 8800 22005 8840
rect 21963 8791 22005 8800
rect 29259 8840 29301 8849
rect 29259 8800 29260 8840
rect 29300 8800 29301 8840
rect 29259 8791 29301 8800
rect 31563 8840 31605 8849
rect 31563 8800 31564 8840
rect 31604 8800 31605 8840
rect 31563 8791 31605 8800
rect 32235 8840 32277 8849
rect 32235 8800 32236 8840
rect 32276 8800 32277 8840
rect 32235 8791 32277 8800
rect 34059 8840 34101 8849
rect 34059 8800 34060 8840
rect 34100 8800 34101 8840
rect 34059 8791 34101 8800
rect 37899 8840 37941 8849
rect 37899 8800 37900 8840
rect 37940 8800 37941 8840
rect 37899 8791 37941 8800
rect 41067 8840 41109 8849
rect 41067 8800 41068 8840
rect 41108 8800 41109 8840
rect 41067 8791 41109 8800
rect 44323 8840 44381 8841
rect 44323 8800 44332 8840
rect 44372 8800 44381 8840
rect 44323 8799 44381 8800
rect 45771 8840 45813 8849
rect 45771 8800 45772 8840
rect 45812 8800 45813 8840
rect 45771 8791 45813 8800
rect 15627 8756 15669 8765
rect 15627 8716 15628 8756
rect 15668 8716 15669 8756
rect 15627 8707 15669 8716
rect 20331 8756 20373 8765
rect 20331 8716 20332 8756
rect 20372 8716 20373 8756
rect 20331 8707 20373 8716
rect 20523 8756 20565 8765
rect 20523 8716 20524 8756
rect 20564 8716 20565 8756
rect 20523 8707 20565 8716
rect 28491 8756 28533 8765
rect 28491 8716 28492 8756
rect 28532 8716 28533 8756
rect 28491 8707 28533 8716
rect 33771 8756 33813 8765
rect 33771 8716 33772 8756
rect 33812 8716 33813 8756
rect 33771 8707 33813 8716
rect 1035 8672 1077 8681
rect 1035 8632 1036 8672
rect 1076 8632 1077 8672
rect 1035 8623 1077 8632
rect 1411 8672 1469 8673
rect 1411 8632 1420 8672
rect 1460 8632 1469 8672
rect 1411 8631 1469 8632
rect 2275 8672 2333 8673
rect 2275 8632 2284 8672
rect 2324 8632 2333 8672
rect 2275 8631 2333 8632
rect 3435 8672 3477 8681
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 3915 8672 3957 8681
rect 3915 8632 3916 8672
rect 3956 8632 3957 8672
rect 3915 8623 3957 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4107 8623 4149 8632
rect 4483 8672 4541 8673
rect 4483 8632 4492 8672
rect 4532 8632 4541 8672
rect 4483 8631 4541 8632
rect 5347 8672 5405 8673
rect 5347 8632 5356 8672
rect 5396 8632 5405 8672
rect 5347 8631 5405 8632
rect 6595 8672 6653 8673
rect 6595 8632 6604 8672
rect 6644 8632 6653 8672
rect 6595 8631 6653 8632
rect 7459 8672 7517 8673
rect 7459 8632 7468 8672
rect 7508 8632 7517 8672
rect 7459 8631 7517 8632
rect 7651 8672 7709 8673
rect 7651 8632 7660 8672
rect 7700 8632 7709 8672
rect 7651 8631 7709 8632
rect 7755 8672 7797 8681
rect 7755 8632 7756 8672
rect 7796 8632 7797 8672
rect 7755 8623 7797 8632
rect 7939 8672 7997 8673
rect 7939 8632 7948 8672
rect 7988 8632 7997 8672
rect 7939 8631 7997 8632
rect 8227 8672 8285 8673
rect 8227 8632 8236 8672
rect 8276 8632 8285 8672
rect 8227 8631 8285 8632
rect 9667 8672 9725 8673
rect 9667 8632 9676 8672
rect 9716 8632 9725 8672
rect 9667 8631 9725 8632
rect 9867 8672 9909 8681
rect 9867 8632 9868 8672
rect 9908 8632 9909 8672
rect 9867 8623 9909 8632
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 10635 8672 10677 8681
rect 10635 8632 10636 8672
rect 10676 8632 10677 8672
rect 10635 8623 10677 8632
rect 11403 8672 11445 8681
rect 11403 8632 11404 8672
rect 11444 8632 11445 8672
rect 11403 8623 11445 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11683 8672 11741 8673
rect 11683 8632 11692 8672
rect 11732 8632 11741 8672
rect 11683 8631 11741 8632
rect 11971 8672 12029 8673
rect 11971 8632 11980 8672
rect 12020 8632 12029 8672
rect 11971 8631 12029 8632
rect 13411 8672 13469 8673
rect 13411 8632 13420 8672
rect 13460 8632 13469 8672
rect 13411 8631 13469 8632
rect 14371 8672 14429 8673
rect 14371 8632 14380 8672
rect 14420 8632 14429 8672
rect 14371 8631 14429 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15723 8672 15765 8681
rect 15723 8632 15724 8672
rect 15764 8632 15765 8672
rect 15723 8623 15765 8632
rect 16003 8672 16061 8673
rect 16003 8632 16012 8672
rect 16052 8632 16061 8672
rect 16003 8631 16061 8632
rect 17163 8672 17205 8681
rect 17163 8632 17164 8672
rect 17204 8632 17205 8672
rect 17163 8623 17205 8632
rect 17355 8672 17397 8681
rect 17355 8632 17356 8672
rect 17396 8632 17397 8672
rect 17355 8623 17397 8632
rect 17547 8672 17589 8681
rect 17547 8632 17548 8672
rect 17588 8632 17589 8672
rect 17547 8623 17589 8632
rect 17739 8672 17781 8681
rect 17739 8632 17740 8672
rect 17780 8632 17781 8672
rect 17739 8623 17781 8632
rect 17827 8672 17885 8673
rect 17827 8632 17836 8672
rect 17876 8632 17885 8672
rect 17827 8631 17885 8632
rect 18315 8672 18357 8681
rect 18315 8632 18316 8672
rect 18356 8632 18357 8672
rect 18315 8623 18357 8632
rect 18507 8672 18549 8681
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 18691 8672 18749 8673
rect 18691 8632 18700 8672
rect 18740 8632 18749 8672
rect 18691 8631 18749 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19851 8672 19893 8681
rect 19851 8632 19852 8672
rect 19892 8632 19893 8672
rect 19851 8623 19893 8632
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 20043 8672 20085 8681
rect 20043 8632 20044 8672
rect 20084 8632 20085 8672
rect 20043 8623 20085 8632
rect 20235 8672 20277 8681
rect 20235 8632 20236 8672
rect 20276 8632 20277 8672
rect 20235 8623 20277 8632
rect 20611 8672 20669 8673
rect 20611 8632 20620 8672
rect 20660 8632 20669 8672
rect 20611 8631 20669 8632
rect 20907 8672 20949 8681
rect 20907 8632 20908 8672
rect 20948 8632 20949 8672
rect 20907 8623 20949 8632
rect 21003 8672 21045 8681
rect 21003 8632 21004 8672
rect 21044 8632 21045 8672
rect 21003 8623 21045 8632
rect 21099 8672 21141 8681
rect 21099 8632 21100 8672
rect 21140 8632 21141 8672
rect 21099 8623 21141 8632
rect 21387 8672 21429 8681
rect 21387 8632 21388 8672
rect 21428 8632 21429 8672
rect 21387 8623 21429 8632
rect 21483 8672 21525 8681
rect 21483 8632 21484 8672
rect 21524 8632 21525 8672
rect 21483 8623 21525 8632
rect 21579 8672 21621 8681
rect 21579 8632 21580 8672
rect 21620 8632 21621 8672
rect 21579 8623 21621 8632
rect 21859 8672 21917 8673
rect 21859 8632 21868 8672
rect 21908 8632 21917 8672
rect 21859 8631 21917 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22731 8672 22773 8681
rect 22731 8632 22732 8672
rect 22772 8632 22773 8672
rect 23115 8672 23157 8681
rect 22731 8623 22773 8632
rect 22910 8651 22968 8652
rect 22910 8611 22919 8651
rect 22959 8611 22968 8651
rect 23115 8632 23116 8672
rect 23156 8632 23157 8672
rect 23115 8623 23157 8632
rect 23307 8672 23349 8681
rect 23307 8632 23308 8672
rect 23348 8632 23349 8672
rect 23307 8623 23349 8632
rect 23395 8672 23453 8673
rect 23395 8632 23404 8672
rect 23444 8632 23453 8672
rect 23395 8631 23453 8632
rect 23787 8672 23829 8681
rect 23787 8632 23788 8672
rect 23828 8632 23829 8672
rect 23787 8623 23829 8632
rect 23883 8672 23925 8681
rect 23883 8632 23884 8672
rect 23924 8632 23925 8672
rect 23883 8623 23925 8632
rect 24075 8672 24117 8681
rect 24075 8632 24076 8672
rect 24116 8632 24117 8672
rect 24075 8623 24117 8632
rect 24171 8672 24213 8681
rect 24171 8632 24172 8672
rect 24212 8632 24213 8672
rect 24171 8623 24213 8632
rect 24267 8672 24309 8681
rect 24267 8632 24268 8672
rect 24308 8632 24309 8672
rect 24267 8623 24309 8632
rect 24363 8672 24405 8681
rect 24363 8632 24364 8672
rect 24404 8632 24405 8672
rect 24363 8623 24405 8632
rect 24555 8672 24597 8681
rect 24555 8632 24556 8672
rect 24596 8632 24597 8672
rect 24555 8623 24597 8632
rect 24747 8672 24789 8681
rect 24747 8632 24748 8672
rect 24788 8632 24789 8672
rect 24747 8623 24789 8632
rect 25027 8672 25085 8673
rect 25027 8632 25036 8672
rect 25076 8632 25085 8672
rect 25027 8631 25085 8632
rect 25699 8672 25757 8673
rect 25699 8632 25708 8672
rect 25748 8632 25757 8672
rect 25699 8631 25757 8632
rect 26283 8672 26325 8681
rect 26283 8632 26284 8672
rect 26324 8632 26325 8672
rect 26283 8623 26325 8632
rect 26379 8672 26421 8681
rect 26379 8632 26380 8672
rect 26420 8632 26421 8672
rect 26379 8623 26421 8632
rect 26475 8672 26517 8681
rect 26475 8632 26476 8672
rect 26516 8632 26517 8672
rect 26475 8623 26517 8632
rect 27230 8672 27288 8673
rect 27230 8632 27239 8672
rect 27279 8632 27288 8672
rect 27230 8631 27288 8632
rect 27339 8672 27381 8681
rect 27339 8632 27340 8672
rect 27380 8632 27381 8672
rect 27339 8623 27381 8632
rect 27435 8672 27477 8681
rect 27435 8632 27436 8672
rect 27476 8632 27477 8672
rect 27435 8623 27477 8632
rect 27619 8672 27677 8673
rect 27619 8632 27628 8672
rect 27668 8632 27677 8672
rect 27619 8631 27677 8632
rect 27715 8672 27773 8673
rect 27715 8632 27724 8672
rect 27764 8632 27773 8672
rect 27715 8631 27773 8632
rect 27915 8668 27957 8677
rect 27915 8628 27916 8668
rect 27956 8628 27957 8668
rect 27915 8619 27957 8628
rect 28011 8672 28053 8681
rect 28210 8677 28252 8686
rect 28011 8632 28012 8672
rect 28052 8632 28053 8672
rect 28011 8623 28053 8632
rect 28114 8668 28156 8677
rect 28114 8628 28115 8668
rect 28155 8628 28156 8668
rect 28210 8637 28211 8677
rect 28251 8637 28252 8677
rect 28210 8628 28252 8637
rect 28395 8672 28437 8681
rect 28395 8632 28396 8672
rect 28436 8632 28437 8672
rect 28114 8619 28156 8628
rect 28395 8623 28437 8632
rect 28587 8672 28629 8681
rect 28587 8632 28588 8672
rect 28628 8632 28629 8672
rect 28587 8623 28629 8632
rect 28963 8672 29021 8673
rect 28963 8632 28972 8672
rect 29012 8632 29021 8672
rect 28963 8631 29021 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 29347 8672 29405 8673
rect 29347 8632 29356 8672
rect 29396 8632 29405 8672
rect 29347 8631 29405 8632
rect 29547 8672 29589 8681
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 29643 8672 29685 8681
rect 29643 8632 29644 8672
rect 29684 8632 29685 8672
rect 29643 8623 29685 8632
rect 29739 8672 29781 8681
rect 29739 8632 29740 8672
rect 29780 8632 29781 8672
rect 29739 8623 29781 8632
rect 29835 8672 29877 8681
rect 29835 8632 29836 8672
rect 29876 8632 29877 8672
rect 29835 8623 29877 8632
rect 30056 8672 30114 8673
rect 30056 8632 30065 8672
rect 30105 8632 30114 8672
rect 30056 8631 30114 8632
rect 30219 8672 30261 8681
rect 30219 8632 30220 8672
rect 30260 8632 30261 8672
rect 30219 8623 30261 8632
rect 30315 8672 30357 8681
rect 30315 8632 30316 8672
rect 30356 8632 30357 8672
rect 30315 8623 30357 8632
rect 30499 8672 30557 8673
rect 30499 8632 30508 8672
rect 30548 8632 30557 8672
rect 30499 8631 30557 8632
rect 30595 8672 30653 8673
rect 30595 8632 30604 8672
rect 30644 8632 30653 8672
rect 30595 8631 30653 8632
rect 31651 8672 31709 8673
rect 31651 8632 31660 8672
rect 31700 8632 31709 8672
rect 31651 8631 31709 8632
rect 31939 8672 31997 8673
rect 31939 8632 31948 8672
rect 31988 8632 31997 8672
rect 31939 8631 31997 8632
rect 33579 8672 33621 8681
rect 33579 8632 33580 8672
rect 33620 8632 33621 8672
rect 33579 8623 33621 8632
rect 33867 8672 33909 8681
rect 33867 8632 33868 8672
rect 33908 8632 33909 8672
rect 33867 8623 33909 8632
rect 34347 8672 34389 8681
rect 34347 8632 34348 8672
rect 34388 8632 34389 8672
rect 34347 8623 34389 8632
rect 34435 8672 34493 8673
rect 34435 8632 34444 8672
rect 34484 8632 34493 8672
rect 34435 8631 34493 8632
rect 34723 8672 34781 8673
rect 34723 8632 34732 8672
rect 34772 8632 34781 8672
rect 34723 8631 34781 8632
rect 35011 8672 35069 8673
rect 35011 8632 35020 8672
rect 35060 8632 35069 8672
rect 35011 8631 35069 8632
rect 35595 8672 35637 8681
rect 35595 8632 35596 8672
rect 35636 8632 35637 8672
rect 35595 8623 35637 8632
rect 35691 8672 35733 8681
rect 35691 8632 35692 8672
rect 35732 8632 35733 8672
rect 35691 8623 35733 8632
rect 35787 8672 35829 8681
rect 35787 8632 35788 8672
rect 35828 8632 35829 8672
rect 35787 8623 35829 8632
rect 35979 8672 36021 8681
rect 35979 8632 35980 8672
rect 36020 8632 36021 8672
rect 35979 8623 36021 8632
rect 36075 8672 36117 8681
rect 36075 8632 36076 8672
rect 36116 8632 36117 8672
rect 36075 8623 36117 8632
rect 37611 8672 37653 8681
rect 37611 8632 37612 8672
rect 37652 8632 37653 8672
rect 37611 8623 37653 8632
rect 37899 8672 37941 8681
rect 37899 8632 37900 8672
rect 37940 8632 37941 8672
rect 37899 8623 37941 8632
rect 38755 8672 38813 8673
rect 38755 8632 38764 8672
rect 38804 8632 38813 8672
rect 38755 8631 38813 8632
rect 38947 8672 39005 8673
rect 38947 8632 38956 8672
rect 38996 8632 39005 8672
rect 38947 8631 39005 8632
rect 39819 8672 39861 8681
rect 39819 8632 39820 8672
rect 39860 8632 39861 8672
rect 39819 8623 39861 8632
rect 40011 8672 40053 8681
rect 40011 8632 40012 8672
rect 40052 8632 40053 8672
rect 40011 8623 40053 8632
rect 40867 8672 40925 8673
rect 40867 8632 40876 8672
rect 40916 8632 40925 8672
rect 40867 8631 40925 8632
rect 41155 8672 41213 8673
rect 41155 8632 41164 8672
rect 41204 8632 41213 8672
rect 41155 8631 41213 8632
rect 41643 8672 41685 8681
rect 41643 8632 41644 8672
rect 41684 8632 41685 8672
rect 41643 8623 41685 8632
rect 41739 8672 41781 8681
rect 41739 8632 41740 8672
rect 41780 8632 41781 8672
rect 41739 8623 41781 8632
rect 42595 8672 42653 8673
rect 42595 8632 42604 8672
rect 42644 8632 42653 8672
rect 42595 8631 42653 8632
rect 42787 8672 42845 8673
rect 42787 8632 42796 8672
rect 42836 8632 42845 8672
rect 42787 8631 42845 8632
rect 43651 8672 43709 8673
rect 43651 8632 43660 8672
rect 43700 8632 43709 8672
rect 43651 8631 43709 8632
rect 45187 8672 45245 8673
rect 45187 8632 45196 8672
rect 45236 8632 45245 8672
rect 45187 8631 45245 8632
rect 45475 8672 45533 8673
rect 45475 8632 45484 8672
rect 45524 8632 45533 8672
rect 45475 8631 45533 8632
rect 46435 8672 46493 8673
rect 46435 8632 46444 8672
rect 46484 8632 46493 8672
rect 46435 8631 46493 8632
rect 46635 8672 46677 8681
rect 46635 8632 46636 8672
rect 46676 8632 46677 8672
rect 46635 8623 46677 8632
rect 47011 8672 47069 8673
rect 47011 8632 47020 8672
rect 47060 8632 47069 8672
rect 47011 8631 47069 8632
rect 47875 8672 47933 8673
rect 47875 8632 47884 8672
rect 47924 8632 47933 8672
rect 47875 8631 47933 8632
rect 22910 8610 22968 8611
rect 9091 8588 9149 8589
rect 9091 8548 9100 8588
rect 9140 8548 9149 8588
rect 9091 8547 9149 8548
rect 9771 8588 9813 8597
rect 9771 8548 9772 8588
rect 9812 8548 9813 8588
rect 9771 8539 9813 8548
rect 11883 8588 11925 8597
rect 11883 8548 11884 8588
rect 11924 8548 11925 8588
rect 11883 8539 11925 8548
rect 17643 8588 17685 8597
rect 17643 8548 17644 8588
rect 17684 8548 17685 8588
rect 17643 8539 17685 8548
rect 21675 8588 21717 8597
rect 21675 8548 21676 8588
rect 21716 8548 21717 8588
rect 21675 8539 21717 8548
rect 23211 8588 23253 8597
rect 23211 8548 23212 8588
rect 23252 8548 23253 8588
rect 23211 8539 23253 8548
rect 41539 8588 41597 8589
rect 41539 8548 41548 8588
rect 41588 8548 41597 8588
rect 41539 8547 41597 8548
rect 643 8504 701 8505
rect 643 8464 652 8504
rect 692 8464 701 8504
rect 643 8463 701 8464
rect 6787 8504 6845 8505
rect 6787 8464 6796 8504
rect 6836 8464 6845 8504
rect 6787 8463 6845 8464
rect 7947 8504 7989 8513
rect 7947 8464 7948 8504
rect 7988 8464 7989 8504
rect 7947 8455 7989 8464
rect 10723 8504 10781 8505
rect 10723 8464 10732 8504
rect 10772 8464 10781 8504
rect 10723 8463 10781 8464
rect 18795 8504 18837 8513
rect 18795 8464 18796 8504
rect 18836 8464 18837 8504
rect 18795 8455 18837 8464
rect 21187 8504 21245 8505
rect 21187 8464 21196 8504
rect 21236 8464 21245 8504
rect 21187 8463 21245 8464
rect 23587 8504 23645 8505
rect 23587 8464 23596 8504
rect 23636 8464 23645 8504
rect 23587 8463 23645 8464
rect 24651 8504 24693 8513
rect 24651 8464 24652 8504
rect 24692 8464 24693 8504
rect 24651 8455 24693 8464
rect 25803 8504 25845 8513
rect 25803 8464 25804 8504
rect 25844 8464 25845 8504
rect 25803 8455 25845 8464
rect 26179 8504 26237 8505
rect 26179 8464 26188 8504
rect 26228 8464 26237 8504
rect 26179 8463 26237 8464
rect 27523 8504 27581 8505
rect 27523 8464 27532 8504
rect 27572 8464 27581 8504
rect 27523 8463 27581 8464
rect 28875 8504 28917 8513
rect 28875 8464 28876 8504
rect 28916 8464 28917 8504
rect 28875 8455 28917 8464
rect 30403 8504 30461 8505
rect 30403 8464 30412 8504
rect 30452 8464 30461 8504
rect 30403 8463 30461 8464
rect 34539 8500 34581 8509
rect 34539 8460 34540 8500
rect 34580 8460 34581 8500
rect 34539 8451 34581 8460
rect 35211 8504 35253 8513
rect 35211 8464 35212 8504
rect 35252 8464 35253 8504
rect 35211 8455 35253 8464
rect 35491 8504 35549 8505
rect 35491 8464 35500 8504
rect 35540 8464 35549 8504
rect 35491 8463 35549 8464
rect 36259 8504 36317 8505
rect 36259 8464 36268 8504
rect 36308 8464 36317 8504
rect 36259 8463 36317 8464
rect 38083 8504 38141 8505
rect 38083 8464 38092 8504
rect 38132 8464 38141 8504
rect 38083 8463 38141 8464
rect 39619 8504 39677 8505
rect 39619 8464 39628 8504
rect 39668 8464 39677 8504
rect 39619 8463 39677 8464
rect 39915 8504 39957 8513
rect 39915 8464 39916 8504
rect 39956 8464 39957 8504
rect 39915 8455 39957 8464
rect 40195 8504 40253 8505
rect 40195 8464 40204 8504
rect 40244 8464 40253 8504
rect 40195 8463 40253 8464
rect 41355 8504 41397 8513
rect 41355 8464 41356 8504
rect 41396 8464 41397 8504
rect 41355 8455 41397 8464
rect 41443 8504 41501 8505
rect 41443 8464 41452 8504
rect 41492 8464 41501 8504
rect 41443 8463 41501 8464
rect 41923 8504 41981 8505
rect 41923 8464 41932 8504
rect 41972 8464 41981 8504
rect 41923 8463 41981 8464
rect 43459 8504 43517 8505
rect 43459 8464 43468 8504
rect 43508 8464 43517 8504
rect 43459 8463 43517 8464
rect 44515 8504 44573 8505
rect 44515 8464 44524 8504
rect 44564 8464 44573 8504
rect 44515 8463 44573 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 1507 8168 1565 8169
rect 1507 8128 1516 8168
rect 1556 8128 1565 8168
rect 1507 8127 1565 8128
rect 3715 8168 3773 8169
rect 3715 8128 3724 8168
rect 3764 8128 3773 8168
rect 3715 8127 3773 8128
rect 4875 8168 4917 8177
rect 4875 8128 4876 8168
rect 4916 8128 4917 8168
rect 4875 8119 4917 8128
rect 5547 8168 5589 8177
rect 5547 8128 5548 8168
rect 5588 8128 5589 8168
rect 5547 8119 5589 8128
rect 8131 8168 8189 8169
rect 8131 8128 8140 8168
rect 8180 8128 8189 8168
rect 8131 8127 8189 8128
rect 8235 8168 8277 8177
rect 8235 8128 8236 8168
rect 8276 8128 8277 8168
rect 8235 8119 8277 8128
rect 10819 8168 10877 8169
rect 10819 8128 10828 8168
rect 10868 8128 10877 8168
rect 10819 8127 10877 8128
rect 15915 8168 15957 8177
rect 15915 8128 15916 8168
rect 15956 8128 15957 8168
rect 15915 8119 15957 8128
rect 17347 8168 17405 8169
rect 17347 8128 17356 8168
rect 17396 8128 17405 8168
rect 17347 8127 17405 8128
rect 21187 8168 21245 8169
rect 21187 8128 21196 8168
rect 21236 8128 21245 8168
rect 21187 8127 21245 8128
rect 23491 8168 23549 8169
rect 23491 8128 23500 8168
rect 23540 8128 23549 8168
rect 23491 8127 23549 8128
rect 25219 8168 25277 8169
rect 25219 8128 25228 8168
rect 25268 8128 25277 8168
rect 25219 8127 25277 8128
rect 34915 8168 34973 8169
rect 34915 8128 34924 8168
rect 34964 8128 34973 8168
rect 34915 8127 34973 8128
rect 36355 8168 36413 8169
rect 36355 8128 36364 8168
rect 36404 8128 36413 8168
rect 36355 8127 36413 8128
rect 37795 8168 37853 8169
rect 37795 8128 37804 8168
rect 37844 8128 37853 8168
rect 37795 8127 37853 8128
rect 8035 8084 8093 8085
rect 8035 8044 8044 8084
rect 8084 8044 8093 8084
rect 8035 8043 8093 8044
rect 11107 8084 11165 8085
rect 11107 8044 11116 8084
rect 11156 8044 11165 8084
rect 11107 8043 11165 8044
rect 11691 8084 11733 8093
rect 11691 8044 11692 8084
rect 11732 8044 11733 8084
rect 11691 8035 11733 8044
rect 21579 8084 21621 8093
rect 21579 8044 21580 8084
rect 21620 8044 21621 8084
rect 21579 8035 21621 8044
rect 35307 8013 35349 8022
rect 843 8000 885 8009
rect 843 7960 844 8000
rect 884 7960 885 8000
rect 843 7951 885 7960
rect 1035 8000 1077 8009
rect 1035 7960 1036 8000
rect 1076 7960 1077 8000
rect 1035 7951 1077 7960
rect 1131 8000 1173 8009
rect 1131 7960 1132 8000
rect 1172 7960 1173 8000
rect 1131 7951 1173 7960
rect 1315 8000 1373 8001
rect 1315 7960 1324 8000
rect 1364 7960 1373 8000
rect 1315 7959 1373 7960
rect 1419 8000 1461 8009
rect 1419 7960 1420 8000
rect 1460 7960 1461 8000
rect 1419 7951 1461 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 2467 8000 2525 8001
rect 2467 7960 2476 8000
rect 2516 7960 2525 8000
rect 2467 7959 2525 7960
rect 3523 8000 3581 8001
rect 3523 7960 3532 8000
rect 3572 7960 3581 8000
rect 3523 7959 3581 7960
rect 4387 8000 4445 8001
rect 4387 7960 4396 8000
rect 4436 7960 4445 8000
rect 4387 7959 4445 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 5059 8000 5117 8001
rect 5059 7960 5068 8000
rect 5108 7960 5117 8000
rect 5059 7959 5117 7960
rect 5347 8000 5405 8001
rect 5347 7960 5356 8000
rect 5396 7960 5405 8000
rect 5347 7959 5405 7960
rect 5835 8000 5877 8009
rect 5835 7960 5836 8000
rect 5876 7960 5877 8000
rect 5835 7951 5877 7960
rect 6019 8000 6077 8001
rect 6019 7960 6028 8000
rect 6068 7960 6077 8000
rect 6019 7959 6077 7960
rect 7555 8000 7613 8001
rect 7555 7960 7564 8000
rect 7604 7960 7613 8000
rect 7555 7959 7613 7960
rect 7851 8000 7893 8009
rect 7851 7960 7852 8000
rect 7892 7960 7893 8000
rect 7851 7951 7893 7960
rect 7947 8000 7989 8009
rect 7947 7960 7948 8000
rect 7988 7960 7989 8000
rect 7947 7951 7989 7960
rect 9091 8000 9149 8001
rect 9091 7960 9100 8000
rect 9140 7960 9149 8000
rect 9091 7959 9149 7960
rect 9483 8000 9525 8009
rect 9483 7960 9484 8000
rect 9524 7960 9525 8000
rect 9483 7951 9525 7960
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 9675 8000 9717 8009
rect 9675 7960 9676 8000
rect 9716 7960 9717 8000
rect 9675 7951 9717 7960
rect 9771 8000 9813 8009
rect 9771 7960 9772 8000
rect 9812 7960 9813 8000
rect 9771 7951 9813 7960
rect 9955 8000 10013 8001
rect 9955 7960 9964 8000
rect 10004 7960 10013 8000
rect 9955 7959 10013 7960
rect 10155 8000 10197 8009
rect 10155 7960 10156 8000
rect 10196 7960 10197 8000
rect 10155 7951 10197 7960
rect 10243 8000 10301 8001
rect 10243 7960 10252 8000
rect 10292 7960 10301 8000
rect 10243 7959 10301 7960
rect 10827 8000 10869 8009
rect 10827 7960 10828 8000
rect 10868 7960 10869 8000
rect 10827 7951 10869 7960
rect 10923 8000 10965 8009
rect 10923 7960 10924 8000
rect 10964 7960 10965 8000
rect 10923 7951 10965 7960
rect 12067 8000 12125 8001
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 12067 7959 12125 7960
rect 12931 8000 12989 8001
rect 12931 7960 12940 8000
rect 12980 7960 12989 8000
rect 12931 7959 12989 7960
rect 15811 8000 15869 8001
rect 15811 7960 15820 8000
rect 15860 7960 15869 8000
rect 15811 7959 15869 7960
rect 16867 8000 16925 8001
rect 16867 7960 16876 8000
rect 16916 7960 16925 8000
rect 16867 7959 16925 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17163 8000 17205 8009
rect 17163 7960 17164 8000
rect 17204 7960 17205 8000
rect 17163 7951 17205 7960
rect 17259 8000 17301 8009
rect 17259 7960 17260 8000
rect 17300 7960 17301 8000
rect 17259 7951 17301 7960
rect 17827 8000 17885 8001
rect 17827 7960 17836 8000
rect 17876 7960 17885 8000
rect 17827 7959 17885 7960
rect 17931 8000 17973 8009
rect 17931 7960 17932 8000
rect 17972 7960 17973 8000
rect 17931 7951 17973 7960
rect 20323 8000 20381 8001
rect 20323 7960 20332 8000
rect 20372 7960 20381 8000
rect 20323 7959 20381 7960
rect 20707 8000 20765 8001
rect 20707 7960 20716 8000
rect 20756 7960 20765 8000
rect 20707 7959 20765 7960
rect 20803 8000 20861 8001
rect 20803 7960 20812 8000
rect 20852 7960 20861 8000
rect 20803 7959 20861 7960
rect 21003 8000 21045 8009
rect 21003 7960 21004 8000
rect 21044 7960 21045 8000
rect 21003 7951 21045 7960
rect 21099 8000 21141 8009
rect 21099 7960 21100 8000
rect 21140 7960 21141 8000
rect 21475 8000 21533 8001
rect 21099 7951 21141 7960
rect 21256 7985 21298 7994
rect 21256 7945 21257 7985
rect 21297 7945 21298 7985
rect 21475 7960 21484 8000
rect 21524 7960 21533 8000
rect 21475 7959 21533 7960
rect 21675 8000 21717 8009
rect 21675 7960 21676 8000
rect 21716 7960 21717 8000
rect 21675 7951 21717 7960
rect 22339 8000 22397 8001
rect 22339 7960 22348 8000
rect 22388 7960 22397 8000
rect 22339 7959 22397 7960
rect 22443 8000 22485 8009
rect 22443 7960 22444 8000
rect 22484 7960 22485 8000
rect 22443 7951 22485 7960
rect 22539 8000 22581 8009
rect 22539 7960 22540 8000
rect 22580 7960 22581 8000
rect 22539 7951 22581 7960
rect 22731 8000 22773 8009
rect 22731 7960 22732 8000
rect 22772 7960 22773 8000
rect 22731 7951 22773 7960
rect 22923 8000 22965 8009
rect 22923 7960 22924 8000
rect 22964 7960 22965 8000
rect 22923 7951 22965 7960
rect 23019 8000 23061 8009
rect 23019 7960 23020 8000
rect 23060 7960 23061 8000
rect 23019 7951 23061 7960
rect 23211 8000 23253 8009
rect 23211 7960 23212 8000
rect 23252 7960 23253 8000
rect 23211 7951 23253 7960
rect 23307 8000 23349 8009
rect 23307 7960 23308 8000
rect 23348 7960 23349 8000
rect 23307 7951 23349 7960
rect 23691 8000 23733 8009
rect 23691 7960 23692 8000
rect 23732 7960 23733 8000
rect 23691 7951 23733 7960
rect 23787 8000 23829 8009
rect 23787 7960 23788 8000
rect 23828 7960 23829 8000
rect 23787 7951 23829 7960
rect 23883 8000 23925 8009
rect 23883 7960 23884 8000
rect 23924 7960 23925 8000
rect 23883 7951 23925 7960
rect 23979 8000 24021 8009
rect 23979 7960 23980 8000
rect 24020 7960 24021 8000
rect 23979 7951 24021 7960
rect 24459 8000 24501 8009
rect 24459 7960 24460 8000
rect 24500 7960 24501 8000
rect 24459 7951 24501 7960
rect 24555 8000 24597 8009
rect 24555 7960 24556 8000
rect 24596 7960 24597 8000
rect 24555 7951 24597 7960
rect 24651 8000 24693 8009
rect 24651 7960 24652 8000
rect 24692 7960 24693 8000
rect 24651 7951 24693 7960
rect 24747 8000 24789 8009
rect 24747 7960 24748 8000
rect 24788 7960 24789 8000
rect 24747 7951 24789 7960
rect 24939 8000 24981 8009
rect 24939 7960 24940 8000
rect 24980 7960 24981 8000
rect 24939 7951 24981 7960
rect 25035 8000 25077 8009
rect 25035 7960 25036 8000
rect 25076 7960 25077 8000
rect 25035 7951 25077 7960
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 25611 8000 25653 8009
rect 25611 7960 25612 8000
rect 25652 7960 25653 8000
rect 25611 7951 25653 7960
rect 25707 8000 25749 8009
rect 25707 7960 25708 8000
rect 25748 7960 25749 8000
rect 25707 7951 25749 7960
rect 25982 8000 26040 8001
rect 25982 7960 25991 8000
rect 26031 7960 26040 8000
rect 25982 7959 26040 7960
rect 26091 8000 26133 8009
rect 26091 7960 26092 8000
rect 26132 7960 26133 8000
rect 26091 7951 26133 7960
rect 26187 8000 26229 8009
rect 26187 7960 26188 8000
rect 26228 7960 26229 8000
rect 26187 7951 26229 7960
rect 26371 8000 26429 8001
rect 26371 7960 26380 8000
rect 26420 7960 26429 8000
rect 26371 7959 26429 7960
rect 26467 8000 26525 8001
rect 26467 7960 26476 8000
rect 26516 7960 26525 8000
rect 26467 7959 26525 7960
rect 27051 8000 27093 8009
rect 27051 7960 27052 8000
rect 27092 7960 27093 8000
rect 27051 7951 27093 7960
rect 27147 8000 27189 8009
rect 27147 7960 27148 8000
rect 27188 7960 27189 8000
rect 27147 7951 27189 7960
rect 27243 8000 27285 8009
rect 27243 7960 27244 8000
rect 27284 7960 27285 8000
rect 27243 7951 27285 7960
rect 27339 8000 27381 8009
rect 27339 7960 27340 8000
rect 27380 7960 27381 8000
rect 27339 7951 27381 7960
rect 27531 8000 27573 8009
rect 27531 7960 27532 8000
rect 27572 7960 27573 8000
rect 27531 7951 27573 7960
rect 29835 8000 29877 8009
rect 29835 7960 29836 8000
rect 29876 7960 29877 8000
rect 29835 7951 29877 7960
rect 29931 8000 29973 8009
rect 29931 7960 29932 8000
rect 29972 7960 29973 8000
rect 29931 7951 29973 7960
rect 30027 8000 30069 8009
rect 30027 7960 30028 8000
rect 30068 7960 30069 8000
rect 30027 7951 30069 7960
rect 30123 8000 30165 8009
rect 30123 7960 30124 8000
rect 30164 7960 30165 8000
rect 30123 7951 30165 7960
rect 31267 8000 31325 8001
rect 31267 7960 31276 8000
rect 31316 7960 31325 8000
rect 31267 7959 31325 7960
rect 31459 8000 31517 8001
rect 31459 7960 31468 8000
rect 31508 7960 31517 8000
rect 31459 7959 31517 7960
rect 31843 8000 31901 8001
rect 31843 7960 31852 8000
rect 31892 7960 31901 8000
rect 31843 7959 31901 7960
rect 32235 8000 32277 8009
rect 32235 7960 32236 8000
rect 32276 7960 32277 8000
rect 32235 7951 32277 7960
rect 34059 8000 34101 8009
rect 34059 7960 34060 8000
rect 34100 7960 34101 8000
rect 34059 7951 34101 7960
rect 34251 8000 34293 8009
rect 34251 7960 34252 8000
rect 34292 7960 34293 8000
rect 34251 7951 34293 7960
rect 34347 8000 34389 8009
rect 34347 7960 34348 8000
rect 34388 7960 34389 8000
rect 34731 8000 34773 8009
rect 34347 7951 34389 7960
rect 34573 7985 34615 7994
rect 21256 7936 21298 7945
rect 34573 7945 34574 7985
rect 34614 7945 34615 7985
rect 34731 7960 34732 8000
rect 34772 7960 34773 8000
rect 34731 7951 34773 7960
rect 34827 8000 34869 8009
rect 34827 7960 34828 8000
rect 34868 7960 34869 8000
rect 34827 7951 34869 7960
rect 35011 8000 35069 8001
rect 35011 7960 35020 8000
rect 35060 7960 35069 8000
rect 35011 7959 35069 7960
rect 35107 8000 35165 8001
rect 35107 7960 35116 8000
rect 35156 7960 35165 8000
rect 35307 7973 35308 8013
rect 35348 7973 35349 8013
rect 35883 8021 35925 8030
rect 35307 7964 35349 7973
rect 35491 8000 35549 8001
rect 35107 7959 35165 7960
rect 35491 7960 35500 8000
rect 35540 7960 35549 8000
rect 35491 7959 35549 7960
rect 35691 8000 35733 8009
rect 35691 7960 35692 8000
rect 35732 7960 35733 8000
rect 35691 7951 35733 7960
rect 35787 8000 35829 8009
rect 35787 7960 35788 8000
rect 35828 7960 35829 8000
rect 35883 7981 35884 8021
rect 35924 7981 35925 8021
rect 35883 7972 35925 7981
rect 35979 8000 36021 8009
rect 35787 7951 35829 7960
rect 35979 7960 35980 8000
rect 36020 7960 36021 8000
rect 35979 7951 36021 7960
rect 36203 8000 36261 8001
rect 36203 7960 36212 8000
rect 36252 7960 36261 8000
rect 36203 7959 36261 7960
rect 36363 8000 36405 8009
rect 36363 7960 36364 8000
rect 36404 7960 36405 8000
rect 36363 7951 36405 7960
rect 36459 8000 36501 8009
rect 36459 7960 36460 8000
rect 36500 7960 36501 8000
rect 36459 7951 36501 7960
rect 36643 8000 36701 8001
rect 36643 7960 36652 8000
rect 36692 7960 36701 8000
rect 36643 7959 36701 7960
rect 36739 8000 36797 8001
rect 36739 7960 36748 8000
rect 36788 7960 36797 8000
rect 36739 7959 36797 7960
rect 36939 8000 36981 8009
rect 36939 7960 36940 8000
rect 36980 7960 36981 8000
rect 36939 7951 36981 7960
rect 37035 8000 37077 8009
rect 37035 7960 37036 8000
rect 37076 7960 37077 8000
rect 37035 7951 37077 7960
rect 37227 8000 37269 8009
rect 37227 7960 37228 8000
rect 37268 7960 37269 8000
rect 37227 7951 37269 7960
rect 37699 8000 37757 8001
rect 37699 7960 37708 8000
rect 37748 7960 37757 8000
rect 37699 7959 37757 7960
rect 37987 8000 38045 8001
rect 37987 7960 37996 8000
rect 38036 7960 38045 8000
rect 37987 7959 38045 7960
rect 38091 8000 38133 8009
rect 38091 7960 38092 8000
rect 38132 7960 38133 8000
rect 38091 7951 38133 7960
rect 38283 8000 38325 8009
rect 38283 7960 38284 8000
rect 38324 7960 38325 8000
rect 38283 7951 38325 7960
rect 38563 8000 38621 8001
rect 38563 7960 38572 8000
rect 38612 7960 38621 8000
rect 38563 7959 38621 7960
rect 38755 8000 38813 8001
rect 38755 7960 38764 8000
rect 38804 7960 38813 8000
rect 38755 7959 38813 7960
rect 38947 8000 39005 8001
rect 38947 7960 38956 8000
rect 38996 7960 39005 8000
rect 38947 7959 39005 7960
rect 40195 8000 40253 8001
rect 40195 7960 40204 8000
rect 40244 7960 40253 8000
rect 40195 7959 40253 7960
rect 41059 8000 41117 8001
rect 41059 7960 41068 8000
rect 41108 7960 41117 8000
rect 41059 7959 41117 7960
rect 41451 8000 41493 8009
rect 41451 7960 41452 8000
rect 41492 7960 41493 8000
rect 41451 7951 41493 7960
rect 41931 8000 41973 8009
rect 41931 7960 41932 8000
rect 41972 7960 41973 8000
rect 41931 7951 41973 7960
rect 43075 8000 43133 8001
rect 43075 7960 43084 8000
rect 43124 7960 43133 8000
rect 43075 7959 43133 7960
rect 43939 8000 43997 8001
rect 43939 7960 43948 8000
rect 43988 7960 43997 8000
rect 43939 7959 43997 7960
rect 44331 8000 44373 8009
rect 44331 7960 44332 8000
rect 44372 7960 44373 8000
rect 44331 7951 44373 7960
rect 44803 8000 44861 8001
rect 44803 7960 44812 8000
rect 44852 7960 44861 8000
rect 44803 7959 44861 7960
rect 46051 8000 46109 8001
rect 46051 7960 46060 8000
rect 46100 7960 46109 8000
rect 46051 7959 46109 7960
rect 46915 8000 46973 8001
rect 46915 7960 46924 8000
rect 46964 7960 46973 8000
rect 46915 7959 46973 7960
rect 47307 8000 47349 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 34573 7936 34615 7945
rect 17539 7916 17597 7917
rect 17539 7876 17548 7916
rect 17588 7876 17597 7916
rect 17539 7875 17597 7876
rect 18883 7916 18941 7917
rect 18883 7876 18892 7916
rect 18932 7876 18941 7916
rect 18883 7875 18941 7876
rect 31947 7916 31989 7925
rect 31947 7876 31948 7916
rect 31988 7876 31989 7916
rect 31947 7867 31989 7876
rect 32139 7916 32181 7925
rect 32139 7876 32140 7916
rect 32180 7876 32181 7916
rect 32139 7867 32181 7876
rect 1123 7832 1181 7833
rect 1123 7792 1132 7832
rect 1172 7792 1181 7832
rect 1123 7791 1181 7792
rect 4683 7832 4725 7841
rect 4683 7792 4684 7832
rect 4724 7792 4725 7832
rect 4683 7783 4725 7792
rect 6411 7832 6453 7841
rect 6411 7792 6412 7832
rect 6452 7792 6453 7832
rect 6411 7783 6453 7792
rect 10435 7832 10493 7833
rect 10435 7792 10444 7832
rect 10484 7792 10493 7832
rect 10435 7791 10493 7792
rect 14859 7832 14901 7841
rect 14859 7792 14860 7832
rect 14900 7792 14901 7832
rect 14859 7783 14901 7792
rect 20427 7832 20469 7841
rect 20427 7792 20428 7832
rect 20468 7792 20469 7832
rect 20427 7783 20469 7792
rect 23011 7832 23069 7833
rect 23011 7792 23020 7832
rect 23060 7792 23069 7832
rect 23011 7791 23069 7792
rect 25699 7832 25757 7833
rect 25699 7792 25708 7832
rect 25748 7792 25757 7832
rect 25699 7791 25757 7792
rect 31467 7832 31509 7841
rect 31467 7792 31468 7832
rect 31508 7792 31509 7832
rect 31467 7783 31509 7792
rect 32043 7832 32085 7841
rect 32043 7792 32044 7832
rect 32084 7792 32085 7832
rect 32043 7783 32085 7792
rect 34339 7832 34397 7833
rect 34339 7792 34348 7832
rect 34388 7792 34397 7832
rect 34339 7791 34397 7792
rect 36931 7832 36989 7833
rect 36931 7792 36940 7832
rect 36980 7792 36989 7832
rect 36931 7791 36989 7792
rect 38283 7832 38325 7841
rect 38283 7792 38284 7832
rect 38324 7792 38325 7832
rect 38283 7783 38325 7792
rect 1795 7748 1853 7749
rect 1795 7708 1804 7748
rect 1844 7708 1853 7748
rect 1795 7707 1853 7708
rect 2851 7748 2909 7749
rect 2851 7708 2860 7748
rect 2900 7708 2909 7748
rect 2851 7707 2909 7708
rect 3715 7748 3773 7749
rect 3715 7708 3724 7748
rect 3764 7708 3773 7748
rect 3715 7707 3773 7708
rect 5931 7748 5973 7757
rect 5931 7708 5932 7748
rect 5972 7708 5973 7748
rect 5931 7699 5973 7708
rect 7083 7748 7125 7757
rect 7083 7708 7084 7748
rect 7124 7708 7125 7748
rect 7083 7699 7125 7708
rect 8419 7748 8477 7749
rect 8419 7708 8428 7748
rect 8468 7708 8477 7748
rect 8419 7707 8477 7708
rect 14083 7748 14141 7749
rect 14083 7708 14092 7748
rect 14132 7708 14141 7748
rect 14083 7707 14141 7708
rect 16195 7748 16253 7749
rect 16195 7708 16204 7748
rect 16244 7708 16253 7748
rect 16195 7707 16253 7708
rect 19083 7748 19125 7757
rect 19083 7708 19084 7748
rect 19124 7708 19125 7748
rect 19083 7699 19125 7708
rect 26475 7748 26517 7757
rect 26475 7708 26476 7748
rect 26516 7708 26517 7748
rect 26475 7699 26517 7708
rect 27819 7748 27861 7757
rect 27819 7708 27820 7748
rect 27860 7708 27861 7748
rect 27819 7699 27861 7708
rect 35403 7748 35445 7757
rect 35403 7708 35404 7748
rect 35444 7708 35445 7748
rect 35403 7699 35445 7708
rect 37507 7748 37565 7749
rect 37507 7708 37516 7748
rect 37556 7708 37565 7748
rect 37507 7707 37565 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 8811 7412 8853 7421
rect 8811 7372 8812 7412
rect 8852 7372 8853 7412
rect 8811 7363 8853 7372
rect 23595 7412 23637 7421
rect 23595 7372 23596 7412
rect 23636 7372 23637 7412
rect 23595 7363 23637 7372
rect 25035 7412 25077 7421
rect 25035 7372 25036 7412
rect 25076 7372 25077 7412
rect 25035 7363 25077 7372
rect 25227 7412 25269 7421
rect 25227 7372 25228 7412
rect 25268 7372 25269 7412
rect 25227 7363 25269 7372
rect 26379 7412 26421 7421
rect 26379 7372 26380 7412
rect 26420 7372 26421 7412
rect 26379 7363 26421 7372
rect 27723 7412 27765 7421
rect 27723 7372 27724 7412
rect 27764 7372 27765 7412
rect 27723 7363 27765 7372
rect 34251 7412 34293 7421
rect 34251 7372 34252 7412
rect 34292 7372 34293 7412
rect 34251 7363 34293 7372
rect 34443 7412 34485 7421
rect 34443 7372 34444 7412
rect 34484 7372 34485 7412
rect 34443 7363 34485 7372
rect 37611 7412 37653 7421
rect 37611 7372 37612 7412
rect 37652 7372 37653 7412
rect 37611 7363 37653 7372
rect 40107 7412 40149 7421
rect 40107 7372 40108 7412
rect 40148 7372 40149 7412
rect 40107 7363 40149 7372
rect 43275 7412 43317 7421
rect 43275 7372 43276 7412
rect 43316 7372 43317 7412
rect 43275 7363 43317 7372
rect 4011 7328 4053 7337
rect 4011 7288 4012 7328
rect 4052 7288 4053 7328
rect 4011 7279 4053 7288
rect 9387 7328 9429 7337
rect 9387 7288 9388 7328
rect 9428 7288 9429 7328
rect 9387 7279 9429 7288
rect 10251 7328 10293 7337
rect 10251 7288 10252 7328
rect 10292 7288 10293 7328
rect 10251 7279 10293 7288
rect 21195 7328 21237 7337
rect 21195 7288 21196 7328
rect 21236 7288 21237 7328
rect 21195 7279 21237 7288
rect 23211 7328 23253 7337
rect 23211 7288 23212 7328
rect 23252 7288 23253 7328
rect 23211 7279 23253 7288
rect 29643 7328 29685 7337
rect 29643 7288 29644 7328
rect 29684 7288 29685 7328
rect 29643 7279 29685 7288
rect 30219 7328 30261 7337
rect 30219 7288 30220 7328
rect 30260 7288 30261 7328
rect 30219 7279 30261 7288
rect 31371 7328 31413 7337
rect 31371 7288 31372 7328
rect 31412 7288 31413 7328
rect 31371 7279 31413 7288
rect 32427 7328 32469 7337
rect 32427 7288 32428 7328
rect 32468 7288 32469 7328
rect 32427 7279 32469 7288
rect 33003 7328 33045 7337
rect 33003 7288 33004 7328
rect 33044 7288 33045 7328
rect 33003 7279 33045 7288
rect 35115 7328 35157 7337
rect 35115 7288 35116 7328
rect 35156 7288 35157 7328
rect 35115 7279 35157 7288
rect 42883 7328 42941 7329
rect 42883 7288 42892 7328
rect 42932 7288 42941 7328
rect 42883 7287 42941 7288
rect 23115 7244 23157 7253
rect 23115 7204 23116 7244
rect 23156 7204 23157 7244
rect 23115 7195 23157 7204
rect 23307 7244 23349 7253
rect 23307 7204 23308 7244
rect 23348 7204 23349 7244
rect 23307 7195 23349 7204
rect 27339 7244 27381 7253
rect 27339 7204 27340 7244
rect 27380 7204 27381 7244
rect 27339 7195 27381 7204
rect 29547 7244 29589 7253
rect 29547 7204 29548 7244
rect 29588 7204 29589 7244
rect 29547 7195 29589 7204
rect 29739 7244 29781 7253
rect 29739 7204 29740 7244
rect 29780 7204 29781 7244
rect 29739 7195 29781 7204
rect 30123 7244 30165 7253
rect 30123 7204 30124 7244
rect 30164 7204 30165 7244
rect 30123 7195 30165 7204
rect 30315 7244 30357 7253
rect 30315 7204 30316 7244
rect 30356 7204 30357 7244
rect 30315 7195 30357 7204
rect 32331 7244 32373 7253
rect 32331 7204 32332 7244
rect 32372 7204 32373 7244
rect 30691 7202 30749 7203
rect 843 7160 885 7169
rect 843 7120 844 7160
rect 884 7120 885 7160
rect 843 7111 885 7120
rect 1219 7160 1277 7161
rect 1219 7120 1228 7160
rect 1268 7120 1277 7160
rect 1219 7119 1277 7120
rect 2083 7160 2141 7161
rect 2083 7120 2092 7160
rect 2132 7120 2141 7160
rect 2083 7119 2141 7120
rect 3331 7160 3389 7161
rect 3331 7120 3340 7160
rect 3380 7120 3389 7160
rect 3331 7119 3389 7120
rect 3723 7160 3765 7169
rect 3723 7120 3724 7160
rect 3764 7120 3765 7160
rect 3723 7111 3765 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 4867 7160 4925 7161
rect 4867 7120 4876 7160
rect 4916 7120 4925 7160
rect 4867 7119 4925 7120
rect 5059 7160 5117 7161
rect 5059 7120 5068 7160
rect 5108 7120 5117 7160
rect 5059 7119 5117 7120
rect 6307 7160 6365 7161
rect 6307 7120 6316 7160
rect 6356 7120 6365 7160
rect 6307 7119 6365 7120
rect 7171 7160 7229 7161
rect 7171 7120 7180 7160
rect 7220 7120 7229 7160
rect 7171 7119 7229 7120
rect 8619 7160 8661 7169
rect 8619 7120 8620 7160
rect 8660 7120 8661 7160
rect 8619 7111 8661 7120
rect 8811 7160 8853 7169
rect 8811 7120 8812 7160
rect 8852 7120 8853 7160
rect 8811 7111 8853 7120
rect 8995 7160 9053 7161
rect 8995 7120 9004 7160
rect 9044 7120 9053 7160
rect 8995 7119 9053 7120
rect 9195 7160 9237 7169
rect 9195 7120 9196 7160
rect 9236 7120 9237 7160
rect 9195 7111 9237 7120
rect 9387 7160 9429 7169
rect 9387 7120 9388 7160
rect 9428 7120 9429 7160
rect 9387 7111 9429 7120
rect 9579 7160 9621 7169
rect 9579 7120 9580 7160
rect 9620 7120 9621 7160
rect 9579 7111 9621 7120
rect 9667 7160 9725 7161
rect 9667 7120 9676 7160
rect 9716 7120 9725 7160
rect 9667 7119 9725 7120
rect 11107 7160 11165 7161
rect 11107 7120 11116 7160
rect 11156 7120 11165 7160
rect 11107 7119 11165 7120
rect 12067 7160 12125 7161
rect 12067 7120 12076 7160
rect 12116 7120 12125 7160
rect 12067 7119 12125 7120
rect 13123 7160 13181 7161
rect 13123 7120 13132 7160
rect 13172 7120 13181 7160
rect 13123 7119 13181 7120
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13995 7111 14037 7120
rect 14379 7160 14421 7169
rect 14379 7120 14380 7160
rect 14420 7120 14421 7160
rect 14379 7111 14421 7120
rect 14755 7160 14813 7161
rect 14755 7120 14764 7160
rect 14804 7120 14813 7160
rect 14755 7119 14813 7120
rect 15619 7160 15677 7161
rect 15619 7120 15628 7160
rect 15668 7120 15677 7160
rect 15619 7119 15677 7120
rect 16867 7160 16925 7161
rect 16867 7120 16876 7160
rect 16916 7120 16925 7160
rect 16867 7119 16925 7120
rect 17347 7160 17405 7161
rect 17347 7120 17356 7160
rect 17396 7120 17405 7160
rect 17347 7119 17405 7120
rect 17635 7160 17693 7161
rect 17635 7120 17644 7160
rect 17684 7120 17693 7160
rect 17635 7119 17693 7120
rect 18499 7160 18557 7161
rect 18499 7120 18508 7160
rect 18548 7120 18557 7160
rect 18499 7119 18557 7120
rect 18691 7160 18749 7161
rect 18691 7120 18700 7160
rect 18740 7120 18749 7160
rect 18691 7119 18749 7120
rect 18795 7160 18837 7169
rect 18795 7120 18796 7160
rect 18836 7120 18837 7160
rect 18795 7111 18837 7120
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 20427 7160 20469 7169
rect 20427 7120 20428 7160
rect 20468 7120 20469 7160
rect 20427 7111 20469 7120
rect 20619 7160 20661 7169
rect 20619 7120 20620 7160
rect 20660 7120 20661 7160
rect 20619 7111 20661 7120
rect 20803 7160 20861 7161
rect 20803 7120 20812 7160
rect 20852 7120 20861 7160
rect 20803 7119 20861 7120
rect 20995 7160 21053 7161
rect 20995 7120 21004 7160
rect 21044 7120 21053 7160
rect 20995 7119 21053 7120
rect 21483 7160 21525 7169
rect 21483 7120 21484 7160
rect 21524 7120 21525 7160
rect 21483 7111 21525 7120
rect 21571 7160 21629 7161
rect 21571 7120 21580 7160
rect 21620 7120 21629 7160
rect 21571 7119 21629 7120
rect 22251 7160 22293 7169
rect 22251 7120 22252 7160
rect 22292 7120 22293 7160
rect 22251 7111 22293 7120
rect 22339 7160 22397 7161
rect 22339 7120 22348 7160
rect 22388 7120 22397 7160
rect 22339 7119 22397 7120
rect 22539 7160 22581 7169
rect 22539 7120 22540 7160
rect 22580 7120 22581 7160
rect 22539 7111 22581 7120
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 23011 7160 23069 7161
rect 23011 7120 23020 7160
rect 23060 7120 23069 7160
rect 23011 7119 23069 7120
rect 23403 7160 23445 7169
rect 23403 7120 23404 7160
rect 23444 7120 23445 7160
rect 23403 7111 23445 7120
rect 23587 7160 23645 7161
rect 23587 7120 23596 7160
rect 23636 7120 23645 7160
rect 23587 7119 23645 7120
rect 23683 7160 23741 7161
rect 23683 7120 23692 7160
rect 23732 7120 23741 7160
rect 23683 7119 23741 7120
rect 23883 7160 23925 7169
rect 23883 7120 23884 7160
rect 23924 7120 23925 7160
rect 23883 7111 23925 7120
rect 23979 7160 24021 7169
rect 23979 7120 23980 7160
rect 24020 7120 24021 7160
rect 23979 7111 24021 7120
rect 24072 7160 24130 7161
rect 24072 7120 24081 7160
rect 24121 7120 24130 7160
rect 24072 7119 24130 7120
rect 24363 7160 24405 7169
rect 24363 7120 24364 7160
rect 24404 7120 24405 7160
rect 24363 7111 24405 7120
rect 24459 7160 24501 7169
rect 24459 7120 24460 7160
rect 24500 7120 24501 7160
rect 24459 7111 24501 7120
rect 24555 7160 24597 7169
rect 24555 7120 24556 7160
rect 24596 7120 24597 7160
rect 24555 7111 24597 7120
rect 24651 7160 24693 7169
rect 24651 7120 24652 7160
rect 24692 7120 24693 7160
rect 24651 7111 24693 7120
rect 24843 7160 24885 7169
rect 24843 7120 24844 7160
rect 24884 7120 24885 7160
rect 24843 7111 24885 7120
rect 25035 7160 25077 7169
rect 25035 7120 25036 7160
rect 25076 7120 25077 7160
rect 25035 7111 25077 7120
rect 25315 7160 25373 7161
rect 25315 7120 25324 7160
rect 25364 7120 25373 7160
rect 25315 7119 25373 7120
rect 26379 7160 26421 7169
rect 26379 7120 26380 7160
rect 26420 7120 26421 7160
rect 26379 7111 26421 7120
rect 26571 7160 26613 7169
rect 26571 7120 26572 7160
rect 26612 7120 26613 7160
rect 26571 7111 26613 7120
rect 27147 7160 27189 7169
rect 27147 7120 27148 7160
rect 27188 7120 27189 7160
rect 27147 7111 27189 7120
rect 27435 7160 27477 7169
rect 27435 7120 27436 7160
rect 27476 7120 27477 7160
rect 27435 7111 27477 7120
rect 27619 7160 27677 7161
rect 27619 7120 27628 7160
rect 27668 7120 27677 7160
rect 27619 7119 27677 7120
rect 27819 7160 27861 7169
rect 27819 7120 27820 7160
rect 27860 7120 27861 7160
rect 27819 7111 27861 7120
rect 29059 7160 29117 7161
rect 29059 7120 29068 7160
rect 29108 7120 29117 7160
rect 29059 7119 29117 7120
rect 29251 7160 29309 7161
rect 29251 7120 29260 7160
rect 29300 7120 29309 7160
rect 29251 7119 29309 7120
rect 29443 7160 29501 7161
rect 29443 7120 29452 7160
rect 29492 7120 29501 7160
rect 29443 7119 29501 7120
rect 29835 7160 29877 7169
rect 29835 7120 29836 7160
rect 29876 7120 29877 7160
rect 29835 7111 29877 7120
rect 30019 7160 30077 7161
rect 30019 7120 30028 7160
rect 30068 7120 30077 7160
rect 30019 7119 30077 7120
rect 30411 7160 30453 7169
rect 30411 7120 30412 7160
rect 30452 7120 30453 7160
rect 30411 7111 30453 7120
rect 30603 7160 30645 7169
rect 30691 7162 30700 7202
rect 30740 7162 30749 7202
rect 32331 7195 32373 7204
rect 32523 7244 32565 7253
rect 32523 7204 32524 7244
rect 32564 7204 32565 7244
rect 32523 7195 32565 7204
rect 32907 7244 32949 7253
rect 32907 7204 32908 7244
rect 32948 7204 32949 7244
rect 32907 7195 32949 7204
rect 33099 7244 33141 7253
rect 33099 7204 33100 7244
rect 33140 7204 33141 7244
rect 33099 7195 33141 7204
rect 35019 7244 35061 7253
rect 35019 7204 35020 7244
rect 35060 7204 35061 7244
rect 35019 7195 35061 7204
rect 35211 7244 35253 7253
rect 35211 7204 35212 7244
rect 35252 7204 35253 7244
rect 35211 7195 35253 7204
rect 35683 7244 35741 7245
rect 35683 7204 35692 7244
rect 35732 7204 35741 7244
rect 35683 7203 35741 7204
rect 40587 7244 40629 7253
rect 40587 7204 40588 7244
rect 40628 7204 40629 7244
rect 40587 7195 40629 7204
rect 30691 7161 30749 7162
rect 30603 7120 30604 7160
rect 30644 7120 30645 7160
rect 30603 7111 30645 7120
rect 30795 7160 30837 7169
rect 30795 7120 30796 7160
rect 30836 7120 30837 7160
rect 30795 7111 30837 7120
rect 30891 7160 30933 7169
rect 30891 7120 30892 7160
rect 30932 7120 30933 7160
rect 30891 7111 30933 7120
rect 31659 7160 31701 7169
rect 31659 7120 31660 7160
rect 31700 7120 31701 7160
rect 31659 7111 31701 7120
rect 31747 7160 31805 7161
rect 31747 7120 31756 7160
rect 31796 7120 31805 7160
rect 31747 7119 31805 7120
rect 32235 7160 32277 7169
rect 32235 7120 32236 7160
rect 32276 7120 32277 7160
rect 32235 7111 32277 7120
rect 32611 7160 32669 7161
rect 32611 7120 32620 7160
rect 32660 7120 32669 7160
rect 32611 7119 32669 7120
rect 32803 7160 32861 7161
rect 32803 7120 32812 7160
rect 32852 7120 32861 7160
rect 32803 7119 32861 7120
rect 33195 7160 33237 7169
rect 33195 7120 33196 7160
rect 33236 7120 33237 7160
rect 33195 7111 33237 7120
rect 34147 7160 34205 7161
rect 34147 7120 34156 7160
rect 34196 7120 34205 7160
rect 34147 7119 34205 7120
rect 34443 7160 34485 7169
rect 34443 7120 34444 7160
rect 34484 7120 34485 7160
rect 34443 7111 34485 7120
rect 34635 7160 34677 7169
rect 34635 7120 34636 7160
rect 34676 7120 34677 7160
rect 34635 7111 34677 7120
rect 34915 7160 34973 7161
rect 34915 7120 34924 7160
rect 34964 7120 34973 7160
rect 34915 7119 34973 7120
rect 35307 7160 35349 7169
rect 35307 7120 35308 7160
rect 35348 7120 35349 7160
rect 35307 7111 35349 7120
rect 35875 7160 35933 7161
rect 35875 7120 35884 7160
rect 35924 7120 35933 7160
rect 35875 7119 35933 7120
rect 36835 7160 36893 7161
rect 36835 7120 36844 7160
rect 36884 7120 36893 7160
rect 36835 7119 36893 7120
rect 37315 7160 37373 7161
rect 37315 7120 37324 7160
rect 37364 7120 37373 7160
rect 37315 7119 37373 7120
rect 37419 7160 37461 7169
rect 37419 7120 37420 7160
rect 37460 7120 37461 7160
rect 37419 7111 37461 7120
rect 37603 7160 37661 7161
rect 37603 7120 37612 7160
rect 37652 7120 37661 7160
rect 37603 7119 37661 7120
rect 37803 7160 37845 7169
rect 37803 7120 37804 7160
rect 37844 7120 37845 7160
rect 37803 7111 37845 7120
rect 37995 7160 38037 7169
rect 37995 7120 37996 7160
rect 38036 7120 38037 7160
rect 37995 7111 38037 7120
rect 38091 7160 38133 7169
rect 38091 7120 38092 7160
rect 38132 7120 38133 7160
rect 38091 7111 38133 7120
rect 38467 7160 38525 7161
rect 38467 7120 38476 7160
rect 38516 7120 38525 7160
rect 38467 7119 38525 7120
rect 39427 7160 39485 7161
rect 39427 7120 39436 7160
rect 39476 7120 39485 7160
rect 39427 7119 39485 7120
rect 40387 7160 40445 7161
rect 40387 7120 40396 7160
rect 40436 7120 40445 7160
rect 40387 7119 40445 7120
rect 41251 7160 41309 7161
rect 41251 7120 41260 7160
rect 41300 7120 41309 7160
rect 41251 7119 41309 7120
rect 41443 7160 41501 7161
rect 41443 7120 41452 7160
rect 41492 7120 41501 7160
rect 41443 7119 41501 7120
rect 41827 7160 41885 7161
rect 41827 7120 41836 7160
rect 41876 7120 41885 7160
rect 41827 7119 41885 7120
rect 42211 7160 42269 7161
rect 42211 7120 42220 7160
rect 42260 7120 42269 7160
rect 42211 7119 42269 7120
rect 43179 7160 43221 7169
rect 43179 7120 43180 7160
rect 43220 7120 43221 7160
rect 43179 7111 43221 7120
rect 43275 7160 43317 7169
rect 43275 7120 43276 7160
rect 43316 7120 43317 7160
rect 43275 7111 43317 7120
rect 43747 7160 43805 7161
rect 43747 7120 43756 7160
rect 43796 7120 43805 7160
rect 43747 7119 43805 7120
rect 44611 7160 44669 7161
rect 44611 7120 44620 7160
rect 44660 7120 44669 7160
rect 44611 7119 44669 7120
rect 46243 7160 46301 7161
rect 46243 7120 46252 7160
rect 46292 7120 46301 7160
rect 46243 7119 46301 7120
rect 46627 7160 46685 7161
rect 46627 7120 46636 7160
rect 46676 7120 46685 7160
rect 46627 7119 46685 7120
rect 47011 7160 47069 7161
rect 47011 7120 47020 7160
rect 47060 7120 47069 7160
rect 47011 7119 47069 7120
rect 5931 7076 5973 7085
rect 5931 7036 5932 7076
rect 5972 7036 5973 7076
rect 5931 7027 5973 7036
rect 9099 7076 9141 7085
rect 9099 7036 9100 7076
rect 9140 7036 9141 7076
rect 9099 7027 9141 7036
rect 41923 7076 41981 7077
rect 41923 7036 41932 7076
rect 41972 7036 41981 7076
rect 41923 7035 41981 7036
rect 43363 7076 43421 7077
rect 43363 7036 43372 7076
rect 43412 7036 43421 7076
rect 43363 7035 43421 7036
rect 46531 7076 46589 7077
rect 46531 7036 46540 7076
rect 46580 7036 46589 7076
rect 46531 7035 46589 7036
rect 3715 6992 3773 6993
rect 3715 6952 3724 6992
rect 3764 6952 3773 6992
rect 3715 6951 3773 6952
rect 4195 6992 4253 6993
rect 4195 6952 4204 6992
rect 4244 6952 4253 6992
rect 4195 6951 4253 6952
rect 5731 6992 5789 6993
rect 5731 6952 5740 6992
rect 5780 6952 5789 6992
rect 5731 6951 5789 6952
rect 8323 6992 8381 6993
rect 8323 6952 8332 6992
rect 8372 6952 8381 6992
rect 8323 6951 8381 6952
rect 10435 6992 10493 6993
rect 10435 6952 10444 6992
rect 10484 6952 10493 6992
rect 10435 6951 10493 6952
rect 11395 6992 11453 6993
rect 11395 6952 11404 6992
rect 11444 6952 11453 6992
rect 11395 6951 11453 6952
rect 17163 6992 17205 7001
rect 17163 6952 17164 6992
rect 17204 6952 17205 6992
rect 17163 6943 17205 6952
rect 17827 6992 17885 6993
rect 17827 6952 17836 6992
rect 17876 6952 17885 6992
rect 17827 6951 17885 6952
rect 18883 6992 18941 6993
rect 18883 6952 18892 6992
rect 18932 6952 18941 6992
rect 18883 6951 18941 6952
rect 20523 6992 20565 7001
rect 20523 6952 20524 6992
rect 20564 6952 20565 6992
rect 20523 6943 20565 6952
rect 21675 6988 21717 6997
rect 21675 6948 21676 6988
rect 21716 6948 21717 6988
rect 22819 6992 22877 6993
rect 22819 6952 22828 6992
rect 22868 6952 22877 6992
rect 22819 6951 22877 6952
rect 31851 6988 31893 6997
rect 21675 6939 21717 6948
rect 31851 6948 31852 6988
rect 31892 6948 31893 6988
rect 31851 6939 31893 6948
rect 36363 6992 36405 7001
rect 36363 6952 36364 6992
rect 36404 6952 36405 6992
rect 36363 6943 36405 6952
rect 37611 6992 37653 7001
rect 37611 6952 37612 6992
rect 37652 6952 37653 6992
rect 37611 6943 37653 6952
rect 38083 6992 38141 6993
rect 38083 6952 38092 6992
rect 38132 6952 38141 6992
rect 38083 6951 38141 6952
rect 39139 6992 39197 6993
rect 39139 6952 39148 6992
rect 39188 6952 39197 6992
rect 39139 6951 39197 6952
rect 43459 6992 43517 6993
rect 43459 6952 43468 6992
rect 43508 6952 43517 6992
rect 43459 6951 43517 6952
rect 44419 6992 44477 6993
rect 44419 6952 44428 6992
rect 44468 6952 44477 6992
rect 44419 6951 44477 6952
rect 45283 6992 45341 6993
rect 45283 6952 45292 6992
rect 45332 6952 45341 6992
rect 45283 6951 45341 6952
rect 45571 6992 45629 6993
rect 45571 6952 45580 6992
rect 45620 6952 45629 6992
rect 45571 6951 45629 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 643 6656 701 6657
rect 643 6616 652 6656
rect 692 6616 701 6656
rect 643 6615 701 6616
rect 7747 6656 7805 6657
rect 7747 6616 7756 6656
rect 7796 6616 7805 6656
rect 7747 6615 7805 6616
rect 8331 6656 8373 6665
rect 8331 6616 8332 6656
rect 8372 6616 8373 6656
rect 8331 6607 8373 6616
rect 9483 6656 9525 6665
rect 9483 6616 9484 6656
rect 9524 6616 9525 6656
rect 9483 6607 9525 6616
rect 10147 6656 10205 6657
rect 10147 6616 10156 6656
rect 10196 6616 10205 6656
rect 10147 6615 10205 6616
rect 12835 6656 12893 6657
rect 12835 6616 12844 6656
rect 12884 6616 12893 6656
rect 12835 6615 12893 6616
rect 18211 6656 18269 6657
rect 18211 6616 18220 6656
rect 18260 6616 18269 6656
rect 18211 6615 18269 6616
rect 30115 6656 30173 6657
rect 30115 6616 30124 6656
rect 30164 6616 30173 6656
rect 30115 6615 30173 6616
rect 33195 6656 33237 6665
rect 33195 6616 33196 6656
rect 33236 6616 33237 6656
rect 33195 6607 33237 6616
rect 34059 6656 34101 6665
rect 34059 6616 34060 6656
rect 34100 6616 34101 6656
rect 34059 6607 34101 6616
rect 34635 6656 34677 6665
rect 34635 6616 34636 6656
rect 34676 6616 34677 6656
rect 34635 6607 34677 6616
rect 35299 6656 35357 6657
rect 35299 6616 35308 6656
rect 35348 6616 35357 6656
rect 35299 6615 35357 6616
rect 36075 6656 36117 6665
rect 36075 6616 36076 6656
rect 36116 6616 36117 6656
rect 36075 6607 36117 6616
rect 10443 6572 10485 6581
rect 10443 6532 10444 6572
rect 10484 6532 10485 6572
rect 10443 6523 10485 6532
rect 18115 6572 18173 6573
rect 18115 6532 18124 6572
rect 18164 6532 18173 6572
rect 31371 6572 31413 6581
rect 18115 6531 18173 6532
rect 18891 6530 18933 6539
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2755 6488 2813 6489
rect 2755 6448 2764 6488
rect 2804 6448 2813 6488
rect 2755 6447 2813 6448
rect 2851 6488 2909 6489
rect 2851 6448 2860 6488
rect 2900 6448 2909 6488
rect 2851 6447 2909 6448
rect 3619 6488 3677 6489
rect 3619 6448 3628 6488
rect 3668 6448 3677 6488
rect 3619 6447 3677 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 5155 6488 5213 6489
rect 5155 6448 5164 6488
rect 5204 6448 5213 6488
rect 5155 6447 5213 6448
rect 5443 6488 5501 6489
rect 5443 6448 5452 6488
rect 5492 6448 5501 6488
rect 5443 6447 5501 6448
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5739 6488 5781 6497
rect 5739 6448 5740 6488
rect 5780 6448 5781 6488
rect 5739 6439 5781 6448
rect 6595 6488 6653 6489
rect 6595 6448 6604 6488
rect 6644 6448 6653 6488
rect 6595 6447 6653 6448
rect 6787 6488 6845 6489
rect 6787 6448 6796 6488
rect 6836 6448 6845 6488
rect 6787 6447 6845 6448
rect 7083 6488 7125 6497
rect 7083 6448 7084 6488
rect 7124 6448 7125 6488
rect 7083 6439 7125 6448
rect 7267 6488 7325 6489
rect 7267 6448 7276 6488
rect 7316 6448 7325 6488
rect 7267 6447 7325 6448
rect 7467 6488 7509 6497
rect 7467 6448 7468 6488
rect 7508 6448 7509 6488
rect 7467 6439 7509 6448
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 8235 6488 8277 6497
rect 8235 6448 8236 6488
rect 8276 6448 8277 6488
rect 8235 6439 8277 6448
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8619 6488 8661 6497
rect 8619 6448 8620 6488
rect 8660 6448 8661 6488
rect 8619 6439 8661 6448
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 8995 6488 9053 6489
rect 8995 6448 9004 6488
rect 9044 6448 9053 6488
rect 8995 6447 9053 6448
rect 9195 6488 9237 6497
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 9379 6488 9437 6489
rect 9379 6448 9388 6488
rect 9428 6448 9437 6488
rect 9379 6447 9437 6448
rect 9763 6488 9821 6489
rect 9763 6448 9772 6488
rect 9812 6448 9821 6488
rect 9763 6447 9821 6448
rect 9955 6488 10013 6489
rect 9955 6448 9964 6488
rect 10004 6448 10013 6488
rect 9955 6447 10013 6448
rect 10059 6488 10101 6497
rect 10059 6448 10060 6488
rect 10100 6448 10101 6488
rect 10059 6439 10101 6448
rect 10251 6488 10293 6497
rect 10251 6448 10252 6488
rect 10292 6448 10293 6488
rect 10251 6439 10293 6448
rect 10819 6488 10877 6489
rect 10819 6448 10828 6488
rect 10868 6448 10877 6488
rect 10819 6447 10877 6448
rect 11683 6488 11741 6489
rect 11683 6448 11692 6488
rect 11732 6448 11741 6488
rect 11683 6447 11741 6448
rect 13611 6488 13653 6497
rect 13611 6448 13612 6488
rect 13652 6448 13653 6488
rect 13611 6439 13653 6448
rect 13899 6488 13941 6497
rect 13899 6448 13900 6488
rect 13940 6448 13941 6488
rect 13899 6439 13941 6448
rect 15523 6488 15581 6489
rect 15523 6448 15532 6488
rect 15572 6448 15581 6488
rect 15523 6447 15581 6448
rect 16395 6488 16437 6497
rect 16395 6448 16396 6488
rect 16436 6448 16437 6488
rect 16395 6439 16437 6448
rect 16779 6488 16821 6497
rect 16779 6448 16780 6488
rect 16820 6448 16821 6488
rect 16779 6439 16821 6448
rect 17443 6488 17501 6489
rect 17443 6448 17452 6488
rect 17492 6448 17501 6488
rect 17443 6447 17501 6448
rect 17931 6488 17973 6497
rect 17931 6448 17932 6488
rect 17972 6448 17973 6488
rect 17931 6439 17973 6448
rect 18027 6488 18069 6497
rect 18891 6490 18892 6530
rect 18932 6490 18933 6530
rect 22923 6530 22965 6539
rect 18027 6448 18028 6488
rect 18068 6448 18069 6488
rect 18027 6439 18069 6448
rect 18787 6488 18845 6489
rect 18787 6448 18796 6488
rect 18836 6448 18845 6488
rect 18891 6481 18933 6490
rect 19083 6488 19125 6497
rect 18787 6447 18845 6448
rect 19083 6448 19084 6488
rect 19124 6448 19125 6488
rect 19083 6439 19125 6448
rect 19275 6488 19317 6497
rect 19275 6448 19276 6488
rect 19316 6448 19317 6488
rect 19275 6439 19317 6448
rect 19371 6488 19413 6497
rect 19371 6448 19372 6488
rect 19412 6448 19413 6488
rect 19371 6439 19413 6448
rect 19467 6488 19509 6497
rect 19467 6448 19468 6488
rect 19508 6448 19509 6488
rect 19467 6439 19509 6448
rect 19563 6488 19605 6497
rect 19563 6448 19564 6488
rect 19604 6448 19605 6488
rect 19563 6439 19605 6448
rect 19755 6488 19797 6497
rect 19755 6448 19756 6488
rect 19796 6448 19797 6488
rect 19755 6439 19797 6448
rect 19851 6488 19893 6497
rect 19851 6448 19852 6488
rect 19892 6448 19893 6488
rect 19851 6439 19893 6448
rect 19947 6488 19989 6497
rect 19947 6448 19948 6488
rect 19988 6448 19989 6488
rect 19947 6439 19989 6448
rect 20043 6488 20085 6497
rect 22923 6490 22924 6530
rect 22964 6490 22965 6530
rect 31371 6532 31372 6572
rect 31412 6532 31413 6572
rect 31371 6523 31413 6532
rect 35587 6572 35645 6573
rect 35587 6532 35596 6572
rect 35636 6532 35645 6572
rect 35587 6531 35645 6532
rect 38755 6572 38813 6573
rect 38755 6532 38764 6572
rect 38804 6532 38813 6572
rect 38755 6531 38813 6532
rect 20043 6448 20044 6488
rect 20084 6448 20085 6488
rect 20043 6439 20085 6448
rect 22531 6488 22589 6489
rect 22531 6448 22540 6488
rect 22580 6448 22589 6488
rect 22923 6481 22965 6490
rect 23107 6488 23165 6489
rect 22531 6447 22589 6448
rect 23107 6448 23116 6488
rect 23156 6448 23165 6488
rect 23107 6447 23165 6448
rect 23499 6488 23541 6497
rect 23499 6448 23500 6488
rect 23540 6448 23541 6488
rect 23499 6439 23541 6448
rect 23683 6488 23741 6489
rect 23683 6448 23692 6488
rect 23732 6448 23741 6488
rect 23683 6447 23741 6448
rect 24075 6488 24117 6497
rect 24075 6448 24076 6488
rect 24116 6448 24117 6488
rect 24075 6439 24117 6448
rect 24267 6488 24309 6497
rect 24267 6448 24268 6488
rect 24308 6448 24309 6488
rect 24267 6439 24309 6448
rect 24459 6488 24501 6497
rect 24459 6448 24460 6488
rect 24500 6448 24501 6488
rect 24459 6439 24501 6448
rect 27243 6488 27285 6497
rect 27243 6448 27244 6488
rect 27284 6448 27285 6488
rect 27243 6439 27285 6448
rect 27619 6488 27677 6489
rect 27619 6448 27628 6488
rect 27668 6448 27677 6488
rect 27619 6447 27677 6448
rect 28203 6488 28245 6497
rect 28203 6448 28204 6488
rect 28244 6448 28245 6488
rect 28203 6439 28245 6448
rect 28395 6488 28437 6497
rect 28395 6448 28396 6488
rect 28436 6448 28437 6488
rect 28395 6439 28437 6448
rect 28587 6488 28629 6497
rect 28587 6448 28588 6488
rect 28628 6448 28629 6488
rect 28587 6439 28629 6448
rect 28779 6488 28821 6497
rect 28779 6448 28780 6488
rect 28820 6448 28821 6488
rect 28779 6439 28821 6448
rect 28971 6488 29013 6497
rect 28971 6448 28972 6488
rect 29012 6448 29013 6488
rect 28971 6439 29013 6448
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 29251 6488 29309 6489
rect 29251 6448 29260 6488
rect 29300 6448 29309 6488
rect 29251 6447 29309 6448
rect 29451 6488 29493 6497
rect 29451 6448 29452 6488
rect 29492 6448 29493 6488
rect 29451 6439 29493 6448
rect 29643 6488 29685 6497
rect 29643 6448 29644 6488
rect 29684 6448 29685 6488
rect 29643 6439 29685 6448
rect 29835 6488 29877 6497
rect 29835 6448 29836 6488
rect 29876 6448 29877 6488
rect 29835 6439 29877 6448
rect 29931 6488 29973 6497
rect 29931 6448 29932 6488
rect 29972 6448 29973 6488
rect 29931 6439 29973 6448
rect 31267 6488 31325 6489
rect 31267 6448 31276 6488
rect 31316 6448 31325 6488
rect 31267 6447 31325 6448
rect 31467 6488 31509 6497
rect 31467 6448 31468 6488
rect 31508 6448 31509 6488
rect 31467 6439 31509 6448
rect 31659 6488 31701 6497
rect 31659 6448 31660 6488
rect 31700 6448 31701 6488
rect 31659 6439 31701 6448
rect 31843 6488 31901 6489
rect 31843 6448 31852 6488
rect 31892 6448 31901 6488
rect 31843 6447 31901 6448
rect 32043 6488 32085 6497
rect 32043 6448 32044 6488
rect 32084 6448 32085 6488
rect 32043 6439 32085 6448
rect 32419 6488 32477 6489
rect 32419 6448 32428 6488
rect 32468 6448 32477 6488
rect 32419 6447 32477 6448
rect 32707 6488 32765 6489
rect 32707 6448 32716 6488
rect 32756 6448 32765 6488
rect 32707 6447 32765 6448
rect 33867 6488 33909 6497
rect 33867 6448 33868 6488
rect 33908 6448 33909 6488
rect 33867 6439 33909 6448
rect 34155 6488 34197 6497
rect 34155 6448 34156 6488
rect 34196 6448 34197 6488
rect 34155 6439 34197 6448
rect 34347 6488 34389 6497
rect 34347 6448 34348 6488
rect 34388 6448 34389 6488
rect 34347 6439 34389 6448
rect 35019 6488 35061 6497
rect 35019 6448 35020 6488
rect 35060 6448 35061 6488
rect 35019 6439 35061 6448
rect 35107 6488 35165 6489
rect 35107 6448 35116 6488
rect 35156 6448 35165 6488
rect 35107 6447 35165 6448
rect 35395 6488 35453 6489
rect 35395 6448 35404 6488
rect 35444 6448 35453 6488
rect 35395 6447 35453 6448
rect 35779 6488 35837 6489
rect 35779 6448 35788 6488
rect 35828 6448 35837 6488
rect 35779 6447 35837 6448
rect 35883 6488 35925 6497
rect 35883 6448 35884 6488
rect 35924 6448 35925 6488
rect 35883 6439 35925 6448
rect 36067 6488 36125 6489
rect 36067 6448 36076 6488
rect 36116 6448 36125 6488
rect 36067 6447 36125 6448
rect 36259 6488 36317 6489
rect 36259 6448 36268 6488
rect 36308 6448 36317 6488
rect 36259 6447 36317 6448
rect 37123 6488 37181 6489
rect 37123 6448 37132 6488
rect 37172 6448 37181 6488
rect 37123 6447 37181 6448
rect 37707 6488 37749 6497
rect 37707 6448 37708 6488
rect 37748 6448 37749 6488
rect 37707 6439 37749 6448
rect 37803 6488 37845 6497
rect 37803 6448 37804 6488
rect 37844 6448 37845 6488
rect 37803 6439 37845 6448
rect 37899 6488 37941 6497
rect 37899 6448 37900 6488
rect 37940 6448 37941 6488
rect 37899 6439 37941 6448
rect 37995 6488 38037 6497
rect 37995 6448 37996 6488
rect 38036 6448 38037 6488
rect 37995 6439 38037 6448
rect 38275 6488 38333 6489
rect 38275 6448 38284 6488
rect 38324 6448 38333 6488
rect 38275 6447 38333 6448
rect 38563 6488 38621 6489
rect 38563 6448 38572 6488
rect 38612 6448 38621 6488
rect 38563 6447 38621 6448
rect 39243 6488 39285 6497
rect 39243 6448 39244 6488
rect 39284 6448 39285 6488
rect 39243 6439 39285 6448
rect 39619 6488 39677 6489
rect 39619 6448 39628 6488
rect 39668 6448 39677 6488
rect 39619 6447 39677 6448
rect 40483 6488 40541 6489
rect 40483 6448 40492 6488
rect 40532 6448 40541 6488
rect 40483 6447 40541 6448
rect 41643 6488 41685 6497
rect 41643 6448 41644 6488
rect 41684 6448 41685 6488
rect 41643 6439 41685 6448
rect 43171 6488 43229 6489
rect 43171 6448 43180 6488
rect 43220 6448 43229 6488
rect 43171 6447 43229 6448
rect 44035 6488 44093 6489
rect 44035 6448 44044 6488
rect 44084 6448 44093 6488
rect 44035 6447 44093 6448
rect 44427 6488 44469 6497
rect 44427 6448 44428 6488
rect 44468 6448 44469 6488
rect 44427 6439 44469 6448
rect 44715 6488 44757 6497
rect 44715 6448 44716 6488
rect 44756 6448 44757 6488
rect 44715 6439 44757 6448
rect 45859 6488 45917 6489
rect 45859 6448 45868 6488
rect 45908 6448 45917 6488
rect 45859 6447 45917 6448
rect 46723 6488 46781 6489
rect 46723 6448 46732 6488
rect 46772 6448 46781 6488
rect 46723 6447 46781 6448
rect 47115 6488 47157 6497
rect 47115 6448 47116 6488
rect 47156 6448 47157 6488
rect 47115 6439 47157 6448
rect 2283 6404 2325 6413
rect 2283 6364 2284 6404
rect 2324 6364 2325 6404
rect 2283 6355 2325 6364
rect 2563 6404 2621 6405
rect 2563 6364 2572 6404
rect 2612 6364 2621 6404
rect 2563 6363 2621 6364
rect 22635 6404 22677 6413
rect 22635 6364 22636 6404
rect 22676 6364 22677 6404
rect 22635 6355 22677 6364
rect 22827 6404 22869 6413
rect 22827 6364 22828 6404
rect 22868 6364 22869 6404
rect 22827 6355 22869 6364
rect 23211 6404 23253 6413
rect 23211 6364 23212 6404
rect 23252 6364 23253 6404
rect 23211 6355 23253 6364
rect 23403 6404 23445 6413
rect 23403 6364 23404 6404
rect 23444 6364 23445 6404
rect 23403 6355 23445 6364
rect 23787 6404 23829 6413
rect 23787 6364 23788 6404
rect 23828 6364 23829 6404
rect 23787 6355 23829 6364
rect 23979 6404 24021 6413
rect 23979 6364 23980 6404
rect 24020 6364 24021 6404
rect 23979 6355 24021 6364
rect 27339 6404 27381 6413
rect 27339 6364 27340 6404
rect 27380 6364 27381 6404
rect 27339 6355 27381 6364
rect 27531 6404 27573 6413
rect 27531 6364 27532 6404
rect 27572 6364 27573 6404
rect 27531 6355 27573 6364
rect 29547 6404 29589 6413
rect 29547 6364 29548 6404
rect 29588 6364 29589 6404
rect 29547 6355 29589 6364
rect 32139 6404 32181 6413
rect 32139 6364 32140 6404
rect 32180 6364 32181 6404
rect 32139 6355 32181 6364
rect 32331 6404 32373 6413
rect 32331 6364 32332 6404
rect 32372 6364 32373 6404
rect 32331 6355 32373 6364
rect 42027 6404 42069 6413
rect 42027 6364 42028 6404
rect 42068 6364 42069 6404
rect 42027 6355 42069 6364
rect 1323 6320 1365 6329
rect 1323 6280 1324 6320
rect 1364 6280 1365 6320
rect 1323 6271 1365 6280
rect 5739 6320 5781 6329
rect 5739 6280 5740 6320
rect 5780 6280 5781 6320
rect 5739 6271 5781 6280
rect 8811 6320 8853 6329
rect 8811 6280 8812 6320
rect 8852 6280 8853 6320
rect 8811 6271 8853 6280
rect 9099 6320 9141 6329
rect 9099 6280 9100 6320
rect 9140 6280 9141 6320
rect 9099 6271 9141 6280
rect 9675 6320 9717 6329
rect 9675 6280 9676 6320
rect 9716 6280 9717 6320
rect 9675 6271 9717 6280
rect 14091 6320 14133 6329
rect 14091 6280 14092 6320
rect 14132 6280 14133 6320
rect 14091 6271 14133 6280
rect 16203 6320 16245 6329
rect 16203 6280 16204 6320
rect 16244 6280 16245 6320
rect 16203 6271 16245 6280
rect 19083 6320 19125 6329
rect 19083 6280 19084 6320
rect 19124 6280 19125 6320
rect 19083 6271 19125 6280
rect 22731 6320 22773 6329
rect 22731 6280 22732 6320
rect 22772 6280 22773 6320
rect 22731 6271 22773 6280
rect 23307 6320 23349 6329
rect 23307 6280 23308 6320
rect 23348 6280 23349 6320
rect 23307 6271 23349 6280
rect 23883 6320 23925 6329
rect 23883 6280 23884 6320
rect 23924 6280 23925 6320
rect 23883 6271 23925 6280
rect 27435 6320 27477 6329
rect 27435 6280 27436 6320
rect 27476 6280 27477 6320
rect 27435 6271 27477 6280
rect 32235 6278 32277 6287
rect 4291 6236 4349 6237
rect 4291 6196 4300 6236
rect 4340 6196 4349 6236
rect 4291 6195 4349 6196
rect 5923 6236 5981 6237
rect 5923 6196 5932 6236
rect 5972 6196 5981 6236
rect 5923 6195 5981 6196
rect 7179 6236 7221 6245
rect 7179 6196 7180 6236
rect 7220 6196 7221 6236
rect 7179 6187 7221 6196
rect 13611 6236 13653 6245
rect 13611 6196 13612 6236
rect 13652 6196 13653 6236
rect 13611 6187 13653 6196
rect 18219 6236 18261 6245
rect 18219 6196 18220 6236
rect 18260 6196 18261 6236
rect 18219 6187 18261 6196
rect 24267 6236 24309 6245
rect 24267 6196 24268 6236
rect 24308 6196 24309 6236
rect 24267 6187 24309 6196
rect 28203 6236 28245 6245
rect 28203 6196 28204 6236
rect 28244 6196 28245 6236
rect 28203 6187 28245 6196
rect 28587 6236 28629 6245
rect 28587 6196 28588 6236
rect 28628 6196 28629 6236
rect 28587 6187 28629 6196
rect 28971 6236 29013 6245
rect 28971 6196 28972 6236
rect 29012 6196 29013 6236
rect 28971 6187 29013 6196
rect 31755 6236 31797 6245
rect 31755 6196 31756 6236
rect 31796 6196 31797 6236
rect 32235 6238 32236 6278
rect 32276 6238 32277 6278
rect 32235 6229 32277 6238
rect 36931 6236 36989 6237
rect 31755 6187 31797 6196
rect 36931 6196 36940 6236
rect 36980 6196 36989 6236
rect 36931 6195 36989 6196
rect 37227 6236 37269 6245
rect 37227 6196 37228 6236
rect 37268 6196 37269 6236
rect 37227 6187 37269 6196
rect 37507 6236 37565 6237
rect 37507 6196 37516 6236
rect 37556 6196 37565 6236
rect 37507 6195 37565 6196
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 6795 5900 6837 5909
rect 6795 5860 6796 5900
rect 6836 5860 6837 5900
rect 6795 5851 6837 5860
rect 8907 5900 8949 5909
rect 8907 5860 8908 5900
rect 8948 5860 8949 5900
rect 8907 5851 8949 5860
rect 15819 5900 15861 5909
rect 15819 5860 15820 5900
rect 15860 5860 15861 5900
rect 15819 5851 15861 5860
rect 17067 5900 17109 5909
rect 17067 5860 17068 5900
rect 17108 5860 17109 5900
rect 17067 5851 17109 5860
rect 22059 5900 22101 5909
rect 22059 5860 22060 5900
rect 22100 5860 22101 5900
rect 22059 5851 22101 5860
rect 27147 5900 27189 5909
rect 27147 5860 27148 5900
rect 27188 5860 27189 5900
rect 27147 5851 27189 5860
rect 34539 5900 34581 5909
rect 34539 5860 34540 5900
rect 34580 5860 34581 5900
rect 34539 5851 34581 5860
rect 2283 5816 2325 5825
rect 2283 5776 2284 5816
rect 2324 5776 2325 5816
rect 2283 5767 2325 5776
rect 21387 5816 21429 5825
rect 21387 5776 21388 5816
rect 21428 5776 21429 5816
rect 21387 5767 21429 5776
rect 31563 5816 31605 5825
rect 31563 5776 31564 5816
rect 31604 5776 31605 5816
rect 31563 5767 31605 5776
rect 32235 5816 32277 5825
rect 32235 5776 32236 5816
rect 32276 5776 32277 5816
rect 32235 5767 32277 5776
rect 36363 5816 36405 5825
rect 36363 5776 36364 5816
rect 36404 5776 36405 5816
rect 36363 5767 36405 5776
rect 37131 5816 37173 5825
rect 37131 5776 37132 5816
rect 37172 5776 37173 5816
rect 37131 5767 37173 5776
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 24843 5732 24885 5741
rect 24843 5692 24844 5732
rect 24884 5692 24885 5732
rect 24843 5683 24885 5692
rect 35787 5732 35829 5741
rect 35787 5692 35788 5732
rect 35828 5692 35829 5732
rect 35787 5683 35829 5692
rect 37035 5732 37077 5741
rect 37035 5692 37036 5732
rect 37076 5692 37077 5732
rect 37035 5683 37077 5692
rect 37227 5732 37269 5741
rect 37227 5692 37228 5732
rect 37268 5692 37269 5732
rect 37227 5683 37269 5692
rect 3531 5648 3573 5657
rect 3531 5608 3532 5648
rect 3572 5608 3573 5648
rect 3531 5599 3573 5608
rect 3723 5648 3765 5657
rect 3723 5608 3724 5648
rect 3764 5608 3765 5648
rect 3723 5599 3765 5608
rect 3907 5648 3965 5649
rect 3907 5608 3916 5648
rect 3956 5608 3965 5648
rect 3907 5607 3965 5608
rect 4011 5648 4053 5657
rect 4011 5608 4012 5648
rect 4052 5608 4053 5648
rect 4011 5599 4053 5608
rect 4195 5648 4253 5649
rect 4195 5608 4204 5648
rect 4244 5608 4253 5648
rect 4195 5607 4253 5608
rect 4395 5648 4437 5657
rect 4395 5608 4396 5648
rect 4436 5608 4437 5648
rect 4395 5599 4437 5608
rect 4771 5648 4829 5649
rect 4771 5608 4780 5648
rect 4820 5608 4829 5648
rect 4771 5607 4829 5608
rect 5635 5648 5693 5649
rect 5635 5608 5644 5648
rect 5684 5608 5693 5648
rect 5635 5607 5693 5608
rect 7371 5648 7413 5657
rect 7371 5608 7372 5648
rect 7412 5608 7413 5648
rect 7371 5599 7413 5608
rect 7467 5648 7509 5657
rect 7467 5608 7468 5648
rect 7508 5608 7509 5648
rect 7467 5599 7509 5608
rect 7659 5648 7701 5657
rect 7659 5608 7660 5648
rect 7700 5608 7701 5648
rect 7659 5599 7701 5608
rect 7755 5648 7797 5657
rect 7755 5608 7756 5648
rect 7796 5608 7797 5648
rect 7755 5599 7797 5608
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8235 5648 8277 5657
rect 8235 5608 8236 5648
rect 8276 5608 8277 5648
rect 8235 5599 8277 5608
rect 8899 5648 8957 5649
rect 8899 5608 8908 5648
rect 8948 5608 8957 5648
rect 8899 5607 8957 5608
rect 8995 5648 9053 5649
rect 8995 5608 9004 5648
rect 9044 5608 9053 5648
rect 8995 5607 9053 5608
rect 9195 5648 9237 5657
rect 9195 5608 9196 5648
rect 9236 5608 9237 5648
rect 9195 5599 9237 5608
rect 9291 5648 9333 5657
rect 9291 5608 9292 5648
rect 9332 5608 9333 5648
rect 9291 5599 9333 5608
rect 9384 5648 9442 5649
rect 9384 5608 9393 5648
rect 9433 5608 9442 5648
rect 9384 5607 9442 5608
rect 9675 5648 9717 5657
rect 9675 5608 9676 5648
rect 9716 5608 9717 5648
rect 9675 5599 9717 5608
rect 9867 5648 9909 5657
rect 9867 5608 9868 5648
rect 9908 5608 9909 5648
rect 9867 5599 9909 5608
rect 11883 5648 11925 5657
rect 11883 5608 11884 5648
rect 11924 5608 11925 5648
rect 11883 5599 11925 5608
rect 11979 5648 12021 5657
rect 11979 5608 11980 5648
rect 12020 5608 12021 5648
rect 11979 5599 12021 5608
rect 12075 5648 12117 5657
rect 12075 5608 12076 5648
rect 12116 5608 12117 5648
rect 12075 5599 12117 5608
rect 12171 5648 12213 5657
rect 12171 5608 12172 5648
rect 12212 5608 12213 5648
rect 12171 5599 12213 5608
rect 12939 5648 12981 5657
rect 12939 5608 12940 5648
rect 12980 5608 12981 5648
rect 12939 5599 12981 5608
rect 13035 5648 13077 5657
rect 13035 5608 13036 5648
rect 13076 5608 13077 5648
rect 13035 5599 13077 5608
rect 13131 5648 13173 5657
rect 13131 5608 13132 5648
rect 13172 5608 13173 5648
rect 13131 5599 13173 5608
rect 13227 5648 13269 5657
rect 13227 5608 13228 5648
rect 13268 5608 13269 5648
rect 13227 5599 13269 5608
rect 13419 5648 13461 5657
rect 13419 5608 13420 5648
rect 13460 5608 13461 5648
rect 13419 5599 13461 5608
rect 13795 5648 13853 5649
rect 13795 5608 13804 5648
rect 13844 5608 13853 5648
rect 13795 5607 13853 5608
rect 14659 5648 14717 5649
rect 14659 5608 14668 5648
rect 14708 5608 14717 5648
rect 14659 5607 14717 5608
rect 16099 5648 16157 5649
rect 16099 5608 16108 5648
rect 16148 5608 16157 5648
rect 16099 5607 16157 5608
rect 16203 5648 16245 5657
rect 16203 5608 16204 5648
rect 16244 5608 16245 5648
rect 16203 5599 16245 5608
rect 16395 5648 16437 5657
rect 16395 5608 16396 5648
rect 16436 5608 16437 5648
rect 16395 5599 16437 5608
rect 16587 5648 16629 5657
rect 16587 5608 16588 5648
rect 16628 5608 16629 5648
rect 16587 5599 16629 5608
rect 16683 5648 16725 5657
rect 16683 5608 16684 5648
rect 16724 5608 16725 5648
rect 16683 5599 16725 5608
rect 16779 5648 16821 5657
rect 16779 5608 16780 5648
rect 16820 5608 16821 5648
rect 16779 5599 16821 5608
rect 16875 5648 16917 5657
rect 16875 5608 16876 5648
rect 16916 5608 16917 5648
rect 16875 5599 16917 5608
rect 17067 5648 17109 5657
rect 17067 5608 17068 5648
rect 17108 5608 17109 5648
rect 17067 5599 17109 5608
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 17347 5648 17405 5649
rect 17347 5608 17356 5648
rect 17396 5608 17405 5648
rect 17347 5607 17405 5608
rect 17827 5648 17885 5649
rect 17827 5608 17836 5648
rect 17876 5608 17885 5648
rect 17827 5607 17885 5608
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 17931 5599 17973 5608
rect 18795 5648 18837 5657
rect 18795 5608 18796 5648
rect 18836 5608 18837 5648
rect 18795 5599 18837 5608
rect 18891 5648 18933 5657
rect 18891 5608 18892 5648
rect 18932 5608 18933 5648
rect 18891 5599 18933 5608
rect 19363 5648 19421 5649
rect 19363 5608 19372 5648
rect 19412 5608 19421 5648
rect 19363 5607 19421 5608
rect 19651 5648 19709 5649
rect 19651 5608 19660 5648
rect 19700 5608 19709 5648
rect 19651 5607 19709 5608
rect 19939 5648 19997 5649
rect 19939 5608 19948 5648
rect 19988 5608 19997 5648
rect 19939 5607 19997 5608
rect 20131 5648 20189 5649
rect 20131 5608 20140 5648
rect 20180 5608 20189 5648
rect 20131 5607 20189 5608
rect 20715 5648 20757 5657
rect 20715 5608 20716 5648
rect 20756 5608 20757 5648
rect 20715 5599 20757 5608
rect 20811 5648 20853 5657
rect 20811 5608 20812 5648
rect 20852 5608 20853 5648
rect 20811 5599 20853 5608
rect 21283 5648 21341 5649
rect 21283 5608 21292 5648
rect 21332 5608 21341 5648
rect 21283 5607 21341 5608
rect 21483 5648 21525 5657
rect 21483 5608 21484 5648
rect 21524 5608 21525 5648
rect 21483 5599 21525 5608
rect 22347 5648 22389 5657
rect 22347 5608 22348 5648
rect 22388 5608 22389 5648
rect 22347 5599 22389 5608
rect 22435 5648 22493 5649
rect 22435 5608 22444 5648
rect 22484 5608 22493 5648
rect 22435 5607 22493 5608
rect 23019 5648 23061 5657
rect 23019 5608 23020 5648
rect 23060 5608 23061 5648
rect 23019 5599 23061 5608
rect 23211 5648 23253 5657
rect 23211 5608 23212 5648
rect 23252 5608 23253 5648
rect 23211 5599 23253 5608
rect 23299 5648 23357 5649
rect 23299 5608 23308 5648
rect 23348 5608 23357 5648
rect 23299 5607 23357 5608
rect 23491 5648 23549 5649
rect 23491 5608 23500 5648
rect 23540 5608 23549 5648
rect 23491 5607 23549 5608
rect 23595 5648 23637 5657
rect 23595 5608 23596 5648
rect 23636 5608 23637 5648
rect 23595 5599 23637 5608
rect 23787 5648 23829 5657
rect 23787 5608 23788 5648
rect 23828 5608 23829 5648
rect 23787 5599 23829 5608
rect 23971 5648 24029 5649
rect 23971 5608 23980 5648
rect 24020 5608 24029 5648
rect 23971 5607 24029 5608
rect 24075 5648 24117 5657
rect 24075 5608 24076 5648
rect 24116 5608 24117 5648
rect 24075 5599 24117 5608
rect 24171 5648 24213 5657
rect 24171 5608 24172 5648
rect 24212 5608 24213 5648
rect 24171 5599 24213 5608
rect 24363 5648 24405 5657
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 24555 5648 24597 5657
rect 24555 5608 24556 5648
rect 24596 5608 24597 5648
rect 24555 5599 24597 5608
rect 24739 5648 24797 5649
rect 24739 5608 24748 5648
rect 24788 5608 24797 5648
rect 24739 5607 24797 5608
rect 24939 5648 24981 5657
rect 24939 5608 24940 5648
rect 24980 5608 24981 5648
rect 26571 5648 26613 5657
rect 26379 5634 26421 5643
rect 24939 5599 24981 5608
rect 26276 5633 26334 5634
rect 26276 5593 26285 5633
rect 26325 5593 26334 5633
rect 26276 5592 26334 5593
rect 26379 5594 26380 5634
rect 26420 5594 26421 5634
rect 26571 5608 26572 5648
rect 26612 5608 26613 5648
rect 26571 5599 26613 5608
rect 26851 5648 26909 5649
rect 26851 5608 26860 5648
rect 26900 5608 26909 5648
rect 26851 5607 26909 5608
rect 27811 5648 27869 5649
rect 27811 5608 27820 5648
rect 27860 5608 27869 5648
rect 27811 5607 27869 5608
rect 28203 5648 28245 5657
rect 28203 5608 28204 5648
rect 28244 5608 28245 5648
rect 28203 5599 28245 5608
rect 28395 5648 28437 5657
rect 28395 5608 28396 5648
rect 28436 5608 28437 5648
rect 28395 5599 28437 5608
rect 28483 5648 28541 5649
rect 28483 5608 28492 5648
rect 28532 5608 28541 5648
rect 28483 5607 28541 5608
rect 28875 5648 28917 5657
rect 28875 5608 28876 5648
rect 28916 5608 28917 5648
rect 28875 5599 28917 5608
rect 28963 5648 29021 5649
rect 28963 5608 28972 5648
rect 29012 5608 29021 5648
rect 28963 5607 29021 5608
rect 29643 5648 29685 5657
rect 29643 5608 29644 5648
rect 29684 5608 29685 5648
rect 29643 5599 29685 5608
rect 29739 5648 29781 5657
rect 29739 5608 29740 5648
rect 29780 5608 29781 5648
rect 29739 5599 29781 5608
rect 29835 5648 29877 5657
rect 29835 5608 29836 5648
rect 29876 5608 29877 5648
rect 29835 5599 29877 5608
rect 31083 5648 31125 5657
rect 31083 5608 31084 5648
rect 31124 5608 31125 5648
rect 31083 5599 31125 5608
rect 31371 5648 31413 5657
rect 31371 5608 31372 5648
rect 31412 5608 31413 5648
rect 31371 5599 31413 5608
rect 31851 5648 31893 5657
rect 31851 5608 31852 5648
rect 31892 5608 31893 5648
rect 31851 5599 31893 5608
rect 31939 5648 31997 5649
rect 31939 5608 31948 5648
rect 31988 5608 31997 5648
rect 31939 5607 31997 5608
rect 32523 5648 32565 5657
rect 32523 5608 32524 5648
rect 32564 5608 32565 5648
rect 32523 5599 32565 5608
rect 32611 5648 32669 5649
rect 32611 5608 32620 5648
rect 32660 5608 32669 5648
rect 32611 5607 32669 5608
rect 32899 5648 32957 5649
rect 32899 5608 32908 5648
rect 32948 5608 32957 5648
rect 32899 5607 32957 5608
rect 33003 5648 33045 5657
rect 33003 5608 33004 5648
rect 33044 5608 33045 5648
rect 33003 5599 33045 5608
rect 33099 5648 33141 5657
rect 33099 5608 33100 5648
rect 33140 5608 33141 5648
rect 33099 5599 33141 5608
rect 33291 5648 33333 5657
rect 33291 5608 33292 5648
rect 33332 5608 33333 5648
rect 33291 5599 33333 5608
rect 33483 5648 33525 5657
rect 33483 5608 33484 5648
rect 33524 5608 33525 5648
rect 33483 5599 33525 5608
rect 34435 5648 34493 5649
rect 34435 5608 34444 5648
rect 34484 5608 34493 5648
rect 34435 5607 34493 5608
rect 34731 5648 34773 5657
rect 34731 5608 34732 5648
rect 34772 5608 34773 5648
rect 34731 5599 34773 5608
rect 34827 5648 34869 5657
rect 34827 5608 34828 5648
rect 34868 5608 34869 5648
rect 34827 5599 34869 5608
rect 34923 5648 34965 5657
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 35403 5648 35445 5657
rect 35403 5608 35404 5648
rect 35444 5608 35445 5648
rect 35403 5599 35445 5608
rect 35499 5648 35541 5657
rect 35499 5608 35500 5648
rect 35540 5608 35541 5648
rect 35499 5599 35541 5608
rect 36643 5648 36701 5649
rect 36643 5608 36652 5648
rect 36692 5608 36701 5648
rect 36643 5607 36701 5608
rect 36931 5648 36989 5649
rect 36931 5608 36940 5648
rect 36980 5608 36989 5648
rect 36931 5607 36989 5608
rect 37323 5648 37365 5657
rect 37323 5608 37324 5648
rect 37364 5608 37365 5648
rect 37323 5599 37365 5608
rect 37603 5648 37661 5649
rect 37603 5608 37612 5648
rect 37652 5608 37661 5648
rect 37603 5607 37661 5608
rect 38563 5648 38621 5649
rect 38563 5608 38572 5648
rect 38612 5608 38621 5648
rect 38563 5607 38621 5608
rect 38667 5648 38709 5657
rect 38667 5608 38668 5648
rect 38708 5608 38709 5648
rect 38667 5599 38709 5608
rect 39523 5648 39581 5649
rect 39523 5608 39532 5648
rect 39572 5608 39581 5648
rect 39523 5607 39581 5608
rect 40483 5648 40541 5649
rect 40483 5608 40492 5648
rect 40532 5608 40541 5648
rect 40483 5607 40541 5608
rect 40683 5648 40725 5657
rect 40683 5608 40684 5648
rect 40724 5608 40725 5648
rect 40683 5599 40725 5608
rect 40875 5648 40917 5657
rect 40875 5608 40876 5648
rect 40916 5608 40917 5648
rect 40875 5599 40917 5608
rect 40963 5648 41021 5649
rect 40963 5608 40972 5648
rect 41012 5608 41021 5648
rect 40963 5607 41021 5608
rect 42219 5648 42261 5657
rect 42219 5608 42220 5648
rect 42260 5608 42261 5648
rect 42219 5599 42261 5608
rect 42411 5648 42453 5657
rect 42411 5608 42412 5648
rect 42452 5608 42453 5648
rect 42411 5599 42453 5608
rect 42595 5648 42653 5649
rect 42595 5608 42604 5648
rect 42644 5608 42653 5648
rect 42595 5607 42653 5608
rect 42699 5648 42741 5657
rect 42699 5608 42700 5648
rect 42740 5608 42741 5648
rect 42699 5599 42741 5608
rect 42891 5648 42933 5657
rect 42891 5608 42892 5648
rect 42932 5608 42933 5648
rect 42891 5599 42933 5608
rect 43939 5648 43997 5649
rect 43939 5608 43948 5648
rect 43988 5608 43997 5648
rect 43939 5607 43997 5608
rect 44227 5648 44285 5649
rect 44227 5608 44236 5648
rect 44276 5608 44285 5648
rect 44227 5607 44285 5608
rect 44715 5648 44757 5657
rect 44715 5608 44716 5648
rect 44756 5608 44757 5648
rect 44715 5599 44757 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 44995 5648 45053 5649
rect 44995 5608 45004 5648
rect 45044 5608 45053 5648
rect 44995 5607 45053 5608
rect 26379 5585 26421 5594
rect 8323 5564 8381 5565
rect 8323 5524 8332 5564
rect 8372 5524 8381 5564
rect 8323 5523 8381 5524
rect 16299 5564 16341 5573
rect 16299 5524 16300 5564
rect 16340 5524 16341 5564
rect 16299 5515 16341 5524
rect 18691 5564 18749 5565
rect 18691 5524 18700 5564
rect 18740 5524 18749 5564
rect 18691 5523 18749 5524
rect 19171 5564 19229 5565
rect 19171 5524 19180 5564
rect 19220 5524 19229 5564
rect 19171 5523 19229 5524
rect 20515 5564 20573 5565
rect 20515 5524 20524 5564
rect 20564 5524 20573 5564
rect 20515 5523 20573 5524
rect 38859 5564 38901 5573
rect 38859 5524 38860 5564
rect 38900 5524 38901 5564
rect 38859 5515 38901 5524
rect 40779 5564 40821 5573
rect 40779 5524 40780 5564
rect 40820 5524 40821 5564
rect 40779 5515 40821 5524
rect 42795 5564 42837 5573
rect 42795 5524 42796 5564
rect 42836 5524 42837 5564
rect 42795 5515 42837 5524
rect 44419 5564 44477 5565
rect 44419 5524 44428 5564
rect 44468 5524 44477 5564
rect 44419 5523 44477 5524
rect 44811 5564 44853 5573
rect 44811 5524 44812 5564
rect 44852 5524 44853 5564
rect 44811 5515 44853 5524
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 1027 5480 1085 5481
rect 1027 5440 1036 5480
rect 1076 5440 1085 5480
rect 1027 5439 1085 5440
rect 4203 5480 4245 5489
rect 4203 5440 4204 5480
rect 4244 5440 4245 5480
rect 4203 5431 4245 5440
rect 7171 5480 7229 5481
rect 7171 5440 7180 5480
rect 7220 5440 7229 5480
rect 7171 5439 7229 5440
rect 7939 5480 7997 5481
rect 7939 5440 7948 5480
rect 7988 5440 7997 5480
rect 7939 5439 7997 5440
rect 8419 5480 8477 5481
rect 8419 5440 8428 5480
rect 8468 5440 8477 5480
rect 8419 5439 8477 5440
rect 8523 5480 8565 5489
rect 8523 5440 8524 5480
rect 8564 5440 8565 5480
rect 8523 5431 8565 5440
rect 9771 5480 9813 5489
rect 9771 5440 9772 5480
rect 9812 5440 9813 5480
rect 9771 5431 9813 5440
rect 17547 5480 17589 5489
rect 17547 5440 17548 5480
rect 17588 5440 17589 5480
rect 17547 5431 17589 5440
rect 18507 5480 18549 5489
rect 18507 5440 18508 5480
rect 18548 5440 18549 5480
rect 18507 5431 18549 5440
rect 18595 5480 18653 5481
rect 18595 5440 18604 5480
rect 18644 5440 18653 5480
rect 18595 5439 18653 5440
rect 20803 5480 20861 5481
rect 20803 5440 20812 5480
rect 20852 5440 20861 5480
rect 20803 5439 20861 5440
rect 22539 5476 22581 5485
rect 22539 5436 22540 5476
rect 22580 5436 22581 5476
rect 23107 5480 23165 5481
rect 23107 5440 23116 5480
rect 23156 5440 23165 5480
rect 23107 5439 23165 5440
rect 23683 5480 23741 5481
rect 23683 5440 23692 5480
rect 23732 5440 23741 5480
rect 23683 5439 23741 5440
rect 24459 5480 24501 5489
rect 24459 5440 24460 5480
rect 24500 5440 24501 5480
rect 22539 5427 22581 5436
rect 24459 5431 24501 5440
rect 26467 5480 26525 5481
rect 26467 5440 26476 5480
rect 26516 5440 26525 5480
rect 26467 5439 26525 5440
rect 28291 5480 28349 5481
rect 28291 5440 28300 5480
rect 28340 5440 28349 5480
rect 28291 5439 28349 5440
rect 29259 5480 29301 5489
rect 29259 5440 29260 5480
rect 29300 5440 29301 5480
rect 29259 5431 29301 5440
rect 29923 5480 29981 5481
rect 29923 5440 29932 5480
rect 29972 5440 29981 5480
rect 29923 5439 29981 5440
rect 31275 5480 31317 5489
rect 31275 5440 31276 5480
rect 31316 5440 31317 5480
rect 31275 5431 31317 5440
rect 32043 5476 32085 5485
rect 32043 5436 32044 5476
rect 32084 5436 32085 5476
rect 32043 5427 32085 5436
rect 32715 5476 32757 5485
rect 32715 5436 32716 5476
rect 32756 5436 32757 5476
rect 32715 5427 32757 5436
rect 33387 5480 33429 5489
rect 33387 5440 33388 5480
rect 33428 5440 33429 5480
rect 33387 5431 33429 5440
rect 35011 5480 35069 5481
rect 35011 5440 35020 5480
rect 35060 5440 35069 5480
rect 35011 5439 35069 5440
rect 35203 5480 35261 5481
rect 35203 5440 35212 5480
rect 35252 5440 35261 5480
rect 35203 5439 35261 5440
rect 38275 5480 38333 5481
rect 38275 5440 38284 5480
rect 38324 5440 38333 5480
rect 38275 5439 38333 5440
rect 39811 5480 39869 5481
rect 39811 5440 39820 5480
rect 39860 5440 39869 5480
rect 39811 5439 39869 5440
rect 42315 5480 42357 5489
rect 42315 5440 42316 5480
rect 42356 5440 42357 5480
rect 42315 5431 42357 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 643 5144 701 5145
rect 643 5104 652 5144
rect 692 5104 701 5144
rect 643 5103 701 5104
rect 7939 5144 7997 5145
rect 7939 5104 7948 5144
rect 7988 5104 7997 5144
rect 7939 5103 7997 5104
rect 8715 5144 8757 5153
rect 8715 5104 8716 5144
rect 8756 5104 8757 5144
rect 8715 5095 8757 5104
rect 9675 5148 9717 5157
rect 9675 5108 9676 5148
rect 9716 5108 9717 5148
rect 9675 5099 9717 5108
rect 12075 5144 12117 5153
rect 12075 5104 12076 5144
rect 12116 5104 12117 5144
rect 12075 5095 12117 5104
rect 21475 5144 21533 5145
rect 21475 5104 21484 5144
rect 21524 5104 21533 5144
rect 21475 5103 21533 5104
rect 24259 5144 24317 5145
rect 24259 5104 24268 5144
rect 24308 5104 24317 5144
rect 24259 5103 24317 5104
rect 27043 5144 27101 5145
rect 27043 5104 27052 5144
rect 27092 5104 27101 5144
rect 27043 5103 27101 5104
rect 29251 5144 29309 5145
rect 29251 5104 29260 5144
rect 29300 5104 29309 5144
rect 29251 5103 29309 5104
rect 30219 5144 30261 5153
rect 30219 5104 30220 5144
rect 30260 5104 30261 5144
rect 30219 5095 30261 5104
rect 30307 5144 30365 5145
rect 30307 5104 30316 5144
rect 30356 5104 30365 5144
rect 30307 5103 30365 5104
rect 30883 5144 30941 5145
rect 30883 5104 30892 5144
rect 30932 5104 30941 5144
rect 30883 5103 30941 5104
rect 4779 5060 4821 5069
rect 4779 5020 4780 5060
rect 4820 5020 4821 5060
rect 4779 5011 4821 5020
rect 5163 5060 5205 5069
rect 5163 5020 5164 5060
rect 5204 5020 5205 5060
rect 5163 5011 5205 5020
rect 16011 5060 16053 5069
rect 16011 5020 16012 5060
rect 16052 5020 16053 5060
rect 16011 5011 16053 5020
rect 16387 5060 16445 5061
rect 16387 5020 16396 5060
rect 16436 5020 16445 5060
rect 16387 5019 16445 5020
rect 21571 5060 21629 5061
rect 21571 5020 21580 5060
rect 21620 5020 21629 5060
rect 21571 5019 21629 5020
rect 23883 5060 23925 5069
rect 23883 5020 23884 5060
rect 23924 5020 23925 5060
rect 23883 5011 23925 5020
rect 24355 5060 24413 5061
rect 24355 5020 24364 5060
rect 24404 5020 24413 5060
rect 24355 5019 24413 5020
rect 28779 5060 28821 5069
rect 28779 5020 28780 5060
rect 28820 5020 28821 5060
rect 28779 5011 28821 5020
rect 30403 5060 30461 5061
rect 30403 5020 30412 5060
rect 30452 5020 30461 5060
rect 30403 5019 30461 5020
rect 30979 5060 31037 5061
rect 30979 5020 30988 5060
rect 31028 5020 31037 5060
rect 30979 5019 31037 5020
rect 1707 4976 1749 4985
rect 1707 4936 1708 4976
rect 1748 4936 1749 4976
rect 1707 4927 1749 4936
rect 2083 4976 2141 4977
rect 2083 4936 2092 4976
rect 2132 4936 2141 4976
rect 2083 4935 2141 4936
rect 2947 4976 3005 4977
rect 2947 4936 2956 4976
rect 2996 4936 3005 4976
rect 2947 4935 3005 4936
rect 4195 4976 4253 4977
rect 4195 4936 4204 4976
rect 4244 4936 4253 4976
rect 4195 4935 4253 4936
rect 4579 4976 4637 4977
rect 4579 4936 4588 4976
rect 4628 4936 4637 4976
rect 4579 4935 4637 4936
rect 4683 4976 4725 4985
rect 4683 4936 4684 4976
rect 4724 4936 4725 4976
rect 4683 4927 4725 4936
rect 4875 4976 4917 4985
rect 4875 4936 4876 4976
rect 4916 4936 4917 4976
rect 4875 4927 4917 4936
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 5251 4976 5309 4977
rect 5251 4936 5260 4976
rect 5300 4936 5309 4976
rect 5251 4935 5309 4936
rect 6595 4976 6653 4977
rect 6595 4936 6604 4976
rect 6644 4936 6653 4976
rect 6595 4935 6653 4936
rect 7459 4976 7517 4977
rect 7459 4936 7468 4976
rect 7508 4936 7517 4976
rect 7459 4935 7517 4936
rect 7659 4976 7701 4985
rect 7659 4936 7660 4976
rect 7700 4936 7701 4976
rect 7659 4927 7701 4936
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 8611 4976 8669 4977
rect 8611 4936 8620 4976
rect 8660 4936 8669 4976
rect 8611 4935 8669 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 9483 4976 9525 4985
rect 9483 4936 9484 4976
rect 9524 4936 9525 4976
rect 9483 4927 9525 4936
rect 9571 4976 9629 4977
rect 9571 4936 9580 4976
rect 9620 4936 9629 4976
rect 9571 4935 9629 4936
rect 9867 4976 9909 4985
rect 9867 4936 9868 4976
rect 9908 4936 9909 4976
rect 9867 4927 9909 4936
rect 10059 4976 10101 4985
rect 10059 4936 10060 4976
rect 10100 4936 10101 4976
rect 10059 4927 10101 4936
rect 10147 4976 10205 4977
rect 10147 4936 10156 4976
rect 10196 4936 10205 4976
rect 10147 4935 10205 4936
rect 10347 4976 10389 4985
rect 10347 4936 10348 4976
rect 10388 4936 10389 4976
rect 10347 4927 10389 4936
rect 10539 4976 10581 4985
rect 10539 4936 10540 4976
rect 10580 4936 10581 4976
rect 10539 4927 10581 4936
rect 11587 4976 11645 4977
rect 11587 4936 11596 4976
rect 11636 4936 11645 4976
rect 11587 4935 11645 4936
rect 14659 4976 14717 4977
rect 14659 4936 14668 4976
rect 14708 4936 14717 4976
rect 14659 4935 14717 4936
rect 15915 4976 15957 4985
rect 15915 4936 15916 4976
rect 15956 4936 15957 4976
rect 15915 4927 15957 4936
rect 16099 4976 16157 4977
rect 16099 4936 16108 4976
rect 16148 4936 16157 4976
rect 16099 4935 16157 4936
rect 17251 4976 17309 4977
rect 17251 4936 17260 4976
rect 17300 4936 17309 4976
rect 17251 4935 17309 4936
rect 17547 4976 17589 4985
rect 17547 4936 17548 4976
rect 17588 4936 17589 4976
rect 17547 4927 17589 4936
rect 17739 4976 17781 4985
rect 17739 4936 17740 4976
rect 17780 4936 17781 4976
rect 17739 4927 17781 4936
rect 17827 4976 17885 4977
rect 17827 4936 17836 4976
rect 17876 4936 17885 4976
rect 17827 4935 17885 4936
rect 18019 4976 18077 4977
rect 18019 4936 18028 4976
rect 18068 4936 18077 4976
rect 18019 4935 18077 4936
rect 19083 4976 19125 4985
rect 19083 4936 19084 4976
rect 19124 4936 19125 4976
rect 19083 4927 19125 4936
rect 19179 4976 19221 4985
rect 19179 4936 19180 4976
rect 19220 4936 19221 4976
rect 19179 4927 19221 4936
rect 19275 4976 19317 4985
rect 19275 4936 19276 4976
rect 19316 4936 19317 4976
rect 19275 4927 19317 4936
rect 19371 4976 19413 4985
rect 19371 4936 19372 4976
rect 19412 4936 19413 4976
rect 19371 4927 19413 4936
rect 20043 4976 20085 4985
rect 20043 4936 20044 4976
rect 20084 4936 20085 4976
rect 20043 4927 20085 4936
rect 20227 4976 20285 4977
rect 20227 4936 20236 4976
rect 20276 4936 20285 4976
rect 20227 4935 20285 4936
rect 20427 4976 20469 4985
rect 20427 4936 20428 4976
rect 20468 4936 20469 4976
rect 20427 4927 20469 4936
rect 20523 4976 20565 4985
rect 20523 4936 20524 4976
rect 20564 4936 20565 4976
rect 20523 4927 20565 4936
rect 20619 4976 20661 4985
rect 20619 4936 20620 4976
rect 20660 4936 20661 4976
rect 20619 4927 20661 4936
rect 20715 4976 20757 4985
rect 20715 4936 20716 4976
rect 20756 4936 20757 4976
rect 20715 4927 20757 4936
rect 21675 4976 21717 4985
rect 21675 4936 21676 4976
rect 21716 4936 21717 4976
rect 21675 4927 21717 4936
rect 21771 4976 21813 4985
rect 21771 4936 21772 4976
rect 21812 4936 21813 4976
rect 21771 4927 21813 4936
rect 22731 4976 22773 4985
rect 22731 4936 22732 4976
rect 22772 4936 22773 4976
rect 22731 4927 22773 4936
rect 22923 4976 22965 4985
rect 22923 4936 22924 4976
rect 22964 4936 22965 4976
rect 22923 4927 22965 4936
rect 23107 4976 23165 4977
rect 23107 4936 23116 4976
rect 23156 4936 23165 4976
rect 23107 4935 23165 4936
rect 23307 4976 23349 4985
rect 23307 4936 23308 4976
rect 23348 4936 23349 4976
rect 23307 4927 23349 4936
rect 23395 4976 23453 4977
rect 23395 4936 23404 4976
rect 23444 4936 23453 4976
rect 23395 4935 23453 4936
rect 23683 4976 23741 4977
rect 23683 4936 23692 4976
rect 23732 4936 23741 4976
rect 23683 4935 23741 4936
rect 23787 4976 23829 4985
rect 23787 4936 23788 4976
rect 23828 4936 23829 4976
rect 23787 4927 23829 4936
rect 23979 4976 24021 4985
rect 23979 4936 23980 4976
rect 24020 4936 24021 4976
rect 23979 4927 24021 4936
rect 24459 4976 24501 4985
rect 24459 4936 24460 4976
rect 24500 4936 24501 4976
rect 24459 4927 24501 4936
rect 24555 4976 24597 4985
rect 24555 4936 24556 4976
rect 24596 4936 24597 4976
rect 24555 4927 24597 4936
rect 24747 4976 24789 4985
rect 24747 4936 24748 4976
rect 24788 4936 24789 4976
rect 24747 4927 24789 4936
rect 25035 4976 25077 4985
rect 25035 4936 25036 4976
rect 25076 4936 25077 4976
rect 25035 4927 25077 4936
rect 26091 4976 26133 4985
rect 26091 4936 26092 4976
rect 26132 4936 26133 4976
rect 26091 4927 26133 4936
rect 26187 4976 26229 4985
rect 26187 4936 26188 4976
rect 26228 4936 26229 4976
rect 26187 4927 26229 4936
rect 26283 4976 26325 4985
rect 26283 4936 26284 4976
rect 26324 4936 26325 4976
rect 26283 4927 26325 4936
rect 26379 4976 26421 4985
rect 26379 4936 26380 4976
rect 26420 4936 26421 4976
rect 26379 4927 26421 4936
rect 26571 4976 26613 4985
rect 26571 4936 26572 4976
rect 26612 4936 26613 4976
rect 26571 4927 26613 4936
rect 26667 4976 26709 4985
rect 26667 4936 26668 4976
rect 26708 4936 26709 4976
rect 26667 4927 26709 4936
rect 26763 4976 26805 4985
rect 26763 4936 26764 4976
rect 26804 4936 26805 4976
rect 26763 4927 26805 4936
rect 26859 4976 26901 4985
rect 26859 4936 26860 4976
rect 26900 4936 26901 4976
rect 26859 4927 26901 4936
rect 27243 4976 27285 4985
rect 27243 4936 27244 4976
rect 27284 4936 27285 4976
rect 27243 4927 27285 4936
rect 27339 4976 27381 4985
rect 27339 4936 27340 4976
rect 27380 4936 27381 4976
rect 27339 4927 27381 4936
rect 27531 4976 27573 4985
rect 27531 4936 27532 4976
rect 27572 4936 27573 4976
rect 27531 4927 27573 4936
rect 27907 4976 27965 4977
rect 27907 4936 27916 4976
rect 27956 4936 27965 4976
rect 27907 4935 27965 4936
rect 28683 4976 28725 4985
rect 28683 4936 28684 4976
rect 28724 4936 28725 4976
rect 28683 4927 28725 4936
rect 28875 4976 28917 4985
rect 28875 4936 28876 4976
rect 28916 4936 28917 4976
rect 28875 4927 28917 4936
rect 28963 4976 29021 4977
rect 28963 4936 28972 4976
rect 29012 4936 29021 4976
rect 28963 4935 29021 4936
rect 29163 4976 29205 4985
rect 29163 4936 29164 4976
rect 29204 4936 29205 4976
rect 29163 4927 29205 4936
rect 29355 4976 29397 4985
rect 29355 4936 29356 4976
rect 29396 4936 29397 4976
rect 29355 4927 29397 4936
rect 29443 4976 29501 4977
rect 29443 4936 29452 4976
rect 29492 4936 29501 4976
rect 29443 4935 29501 4936
rect 29643 4976 29685 4985
rect 29643 4936 29644 4976
rect 29684 4936 29685 4976
rect 29643 4927 29685 4936
rect 29739 4976 29781 4985
rect 29739 4936 29740 4976
rect 29780 4936 29781 4976
rect 29739 4927 29781 4936
rect 29835 4976 29877 4985
rect 29835 4936 29836 4976
rect 29876 4936 29877 4976
rect 29835 4927 29877 4936
rect 29931 4976 29973 4985
rect 29931 4936 29932 4976
rect 29972 4936 29973 4976
rect 29931 4927 29973 4936
rect 30507 4976 30549 4985
rect 30507 4936 30508 4976
rect 30548 4936 30549 4976
rect 30507 4927 30549 4936
rect 30603 4976 30645 4985
rect 30603 4936 30604 4976
rect 30644 4936 30645 4976
rect 30603 4927 30645 4936
rect 31083 4976 31125 4985
rect 31083 4936 31084 4976
rect 31124 4936 31125 4976
rect 31083 4927 31125 4936
rect 31179 4976 31221 4985
rect 31179 4936 31180 4976
rect 31220 4936 31221 4976
rect 31179 4927 31221 4936
rect 31563 4976 31605 4985
rect 31563 4936 31564 4976
rect 31604 4936 31605 4976
rect 31563 4927 31605 4936
rect 32611 4976 32669 4977
rect 32611 4936 32620 4976
rect 32660 4936 32669 4976
rect 32611 4935 32669 4936
rect 32715 4976 32757 4985
rect 32715 4936 32716 4976
rect 32756 4936 32757 4976
rect 32715 4927 32757 4936
rect 32907 4976 32949 4985
rect 32907 4936 32908 4976
rect 32948 4936 32949 4976
rect 32907 4927 32949 4936
rect 34251 4976 34293 4985
rect 34251 4936 34252 4976
rect 34292 4936 34293 4976
rect 34251 4927 34293 4936
rect 35107 4976 35165 4977
rect 35107 4936 35116 4976
rect 35156 4936 35165 4976
rect 35107 4935 35165 4936
rect 35299 4976 35357 4977
rect 35299 4936 35308 4976
rect 35348 4936 35357 4976
rect 35299 4935 35357 4936
rect 36547 4976 36605 4977
rect 36547 4936 36556 4976
rect 36596 4936 36605 4976
rect 36547 4935 36605 4936
rect 37411 4976 37469 4977
rect 37411 4936 37420 4976
rect 37460 4936 37469 4976
rect 37411 4935 37469 4936
rect 37803 4976 37845 4985
rect 37803 4936 37804 4976
rect 37844 4936 37845 4976
rect 37803 4927 37845 4936
rect 38179 4976 38237 4977
rect 38179 4936 38188 4976
rect 38228 4936 38237 4976
rect 38179 4935 38237 4936
rect 38371 4976 38429 4977
rect 38371 4936 38380 4976
rect 38420 4936 38429 4976
rect 38371 4935 38429 4936
rect 39243 4976 39285 4985
rect 39243 4936 39244 4976
rect 39284 4936 39285 4976
rect 39243 4927 39285 4936
rect 39619 4976 39677 4977
rect 39619 4936 39628 4976
rect 39668 4936 39677 4976
rect 39619 4935 39677 4936
rect 40483 4976 40541 4977
rect 40483 4936 40492 4976
rect 40532 4936 40541 4976
rect 40483 4935 40541 4936
rect 41643 4976 41685 4985
rect 41643 4936 41644 4976
rect 41684 4936 41685 4976
rect 41643 4927 41685 4936
rect 8811 4892 8853 4901
rect 8811 4852 8812 4892
rect 8852 4852 8853 4892
rect 8811 4843 8853 4852
rect 10443 4892 10485 4901
rect 10443 4852 10444 4892
rect 10484 4852 10485 4892
rect 8899 4850 8957 4851
rect 5451 4808 5493 4817
rect 8899 4810 8908 4850
rect 8948 4810 8957 4850
rect 10443 4843 10485 4852
rect 20139 4892 20181 4901
rect 20139 4852 20140 4892
rect 20180 4852 20181 4892
rect 20139 4843 20181 4852
rect 28099 4892 28157 4893
rect 28099 4852 28108 4892
rect 28148 4852 28157 4892
rect 28099 4851 28157 4852
rect 33859 4892 33917 4893
rect 33859 4852 33868 4892
rect 33908 4852 33917 4892
rect 33859 4851 33917 4852
rect 8899 4809 8957 4810
rect 5451 4768 5452 4808
rect 5492 4768 5493 4808
rect 5451 4759 5493 4768
rect 9195 4808 9237 4817
rect 9195 4768 9196 4808
rect 9236 4768 9237 4808
rect 9195 4759 9237 4768
rect 12747 4808 12789 4817
rect 12747 4768 12748 4808
rect 12788 4768 12789 4808
rect 12747 4759 12789 4768
rect 15051 4808 15093 4817
rect 15051 4768 15052 4808
rect 15092 4768 15093 4808
rect 15051 4759 15093 4768
rect 24451 4808 24509 4809
rect 24451 4768 24460 4808
rect 24500 4768 24509 4808
rect 24451 4767 24509 4768
rect 27627 4808 27669 4817
rect 27627 4768 27628 4808
rect 27668 4768 27669 4808
rect 27627 4759 27669 4768
rect 33675 4808 33717 4817
rect 33675 4768 33676 4808
rect 33716 4768 33717 4808
rect 33675 4759 33717 4768
rect 5923 4724 5981 4725
rect 5923 4684 5932 4724
rect 5972 4684 5981 4724
rect 5923 4683 5981 4684
rect 6787 4724 6845 4725
rect 6787 4684 6796 4724
rect 6836 4684 6845 4724
rect 6787 4683 6845 4684
rect 9867 4724 9909 4733
rect 9867 4684 9868 4724
rect 9908 4684 9909 4724
rect 9867 4675 9909 4684
rect 11883 4724 11925 4733
rect 11883 4684 11884 4724
rect 11924 4684 11925 4724
rect 11883 4675 11925 4684
rect 13987 4724 14045 4725
rect 13987 4684 13996 4724
rect 14036 4684 14045 4724
rect 13987 4683 14045 4684
rect 17547 4724 17589 4733
rect 17547 4684 17548 4724
rect 17588 4684 17589 4724
rect 17547 4675 17589 4684
rect 18691 4724 18749 4725
rect 18691 4684 18700 4724
rect 18740 4684 18749 4724
rect 18691 4683 18749 4684
rect 21675 4724 21717 4733
rect 21675 4684 21676 4724
rect 21716 4684 21717 4724
rect 21675 4675 21717 4684
rect 22731 4724 22773 4733
rect 22731 4684 22732 4724
rect 22772 4684 22773 4724
rect 22731 4675 22773 4684
rect 23115 4724 23157 4733
rect 23115 4684 23116 4724
rect 23156 4684 23157 4724
rect 23115 4675 23157 4684
rect 25035 4724 25077 4733
rect 25035 4684 25036 4724
rect 25076 4684 25077 4724
rect 25035 4675 25077 4684
rect 31083 4724 31125 4733
rect 31083 4684 31084 4724
rect 31124 4684 31125 4724
rect 31083 4675 31125 4684
rect 31947 4724 31989 4733
rect 31947 4684 31948 4724
rect 31988 4684 31989 4724
rect 31947 4675 31989 4684
rect 32907 4724 32949 4733
rect 32907 4684 32908 4724
rect 32948 4684 32949 4724
rect 32907 4675 32949 4684
rect 34443 4724 34485 4733
rect 34443 4684 34444 4724
rect 34484 4684 34485 4724
rect 34443 4675 34485 4684
rect 38091 4724 38133 4733
rect 38091 4684 38092 4724
rect 38132 4684 38133 4724
rect 38091 4675 38133 4684
rect 39043 4724 39101 4725
rect 39043 4684 39052 4724
rect 39092 4684 39101 4724
rect 39043 4683 39101 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 14187 4388 14229 4397
rect 14187 4348 14188 4388
rect 14228 4348 14229 4388
rect 14187 4339 14229 4348
rect 23499 4388 23541 4397
rect 23499 4348 23500 4388
rect 23540 4348 23541 4388
rect 23499 4339 23541 4348
rect 24555 4388 24597 4397
rect 24555 4348 24556 4388
rect 24596 4348 24597 4388
rect 24555 4339 24597 4348
rect 26379 4388 26421 4397
rect 26379 4348 26380 4388
rect 26420 4348 26421 4388
rect 26379 4339 26421 4348
rect 34243 4388 34301 4389
rect 34243 4348 34252 4388
rect 34292 4348 34301 4388
rect 34243 4347 34301 4348
rect 40779 4388 40821 4397
rect 40779 4348 40780 4388
rect 40820 4348 40821 4388
rect 40779 4339 40821 4348
rect 9195 4304 9237 4313
rect 9195 4264 9196 4304
rect 9236 4264 9237 4304
rect 9195 4255 9237 4264
rect 13131 4304 13173 4313
rect 13131 4264 13132 4304
rect 13172 4264 13173 4304
rect 13131 4255 13173 4264
rect 22251 4304 22293 4313
rect 22251 4264 22252 4304
rect 22292 4264 22293 4304
rect 22251 4255 22293 4264
rect 26667 4304 26709 4313
rect 26667 4264 26668 4304
rect 26708 4264 26709 4304
rect 26667 4255 26709 4264
rect 27619 4304 27677 4305
rect 27619 4264 27628 4304
rect 27668 4264 27677 4304
rect 27619 4263 27677 4264
rect 28299 4304 28341 4313
rect 28299 4264 28300 4304
rect 28340 4264 28341 4304
rect 28299 4255 28341 4264
rect 9579 4220 9621 4229
rect 9579 4180 9580 4220
rect 9620 4180 9621 4220
rect 9579 4171 9621 4180
rect 18315 4220 18357 4229
rect 18315 4180 18316 4220
rect 18356 4180 18357 4220
rect 18315 4171 18357 4180
rect 22923 4220 22965 4229
rect 22923 4180 22924 4220
rect 22964 4180 22965 4220
rect 22923 4171 22965 4180
rect 34539 4220 34581 4229
rect 34539 4180 34540 4220
rect 34580 4180 34581 4220
rect 34539 4171 34581 4180
rect 4299 4136 4341 4145
rect 4299 4096 4300 4136
rect 4340 4096 4341 4136
rect 4299 4087 4341 4096
rect 4675 4136 4733 4137
rect 4675 4096 4684 4136
rect 4724 4096 4733 4136
rect 4675 4095 4733 4096
rect 5539 4136 5597 4137
rect 5539 4096 5548 4136
rect 5588 4096 5597 4136
rect 5539 4095 5597 4096
rect 7651 4136 7709 4137
rect 7651 4096 7660 4136
rect 7700 4096 7709 4136
rect 7651 4095 7709 4096
rect 7939 4136 7997 4137
rect 7939 4096 7948 4136
rect 7988 4096 7997 4136
rect 7939 4095 7997 4096
rect 8139 4136 8181 4145
rect 8139 4096 8140 4136
rect 8180 4096 8181 4136
rect 8139 4087 8181 4096
rect 8803 4136 8861 4137
rect 8803 4096 8812 4136
rect 8852 4096 8861 4136
rect 8803 4095 8861 4096
rect 9387 4136 9429 4145
rect 9387 4096 9388 4136
rect 9428 4096 9429 4136
rect 9387 4087 9429 4096
rect 9675 4136 9717 4145
rect 9675 4096 9676 4136
rect 9716 4096 9717 4136
rect 9675 4087 9717 4096
rect 9859 4136 9917 4137
rect 9859 4096 9868 4136
rect 9908 4096 9917 4136
rect 9859 4095 9917 4096
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 10155 4087 10197 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 10443 4136 10485 4145
rect 10443 4096 10444 4136
rect 10484 4096 10485 4136
rect 10443 4087 10485 4096
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11019 4136 11061 4145
rect 11019 4096 11020 4136
rect 11060 4096 11061 4136
rect 11019 4087 11061 4096
rect 11115 4136 11157 4145
rect 11115 4096 11116 4136
rect 11156 4096 11157 4136
rect 11115 4087 11157 4096
rect 11403 4136 11445 4145
rect 11403 4096 11404 4136
rect 11444 4096 11445 4136
rect 11403 4087 11445 4096
rect 11499 4136 11541 4145
rect 11499 4096 11500 4136
rect 11540 4096 11541 4136
rect 11499 4087 11541 4096
rect 11595 4136 11637 4145
rect 11595 4096 11596 4136
rect 11636 4096 11637 4136
rect 11595 4087 11637 4096
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12931 4136 12989 4137
rect 12931 4096 12940 4136
rect 12980 4096 12989 4136
rect 12931 4095 12989 4096
rect 13131 4136 13173 4145
rect 13131 4096 13132 4136
rect 13172 4096 13173 4136
rect 13131 4087 13173 4096
rect 13323 4136 13365 4145
rect 13323 4096 13324 4136
rect 13364 4096 13365 4136
rect 13323 4087 13365 4096
rect 13411 4136 13469 4137
rect 13411 4096 13420 4136
rect 13460 4096 13469 4136
rect 13411 4095 13469 4096
rect 13603 4136 13661 4137
rect 13603 4096 13612 4136
rect 13652 4096 13661 4136
rect 13603 4095 13661 4096
rect 13795 4136 13853 4137
rect 13795 4096 13804 4136
rect 13844 4096 13853 4136
rect 13795 4095 13853 4096
rect 15331 4136 15389 4137
rect 15331 4096 15340 4136
rect 15380 4096 15389 4136
rect 15331 4095 15389 4096
rect 16195 4136 16253 4137
rect 16195 4096 16204 4136
rect 16244 4096 16253 4136
rect 16195 4095 16253 4096
rect 16587 4136 16629 4145
rect 16587 4096 16588 4136
rect 16628 4096 16629 4136
rect 16587 4087 16629 4096
rect 16971 4136 17013 4145
rect 16971 4096 16972 4136
rect 17012 4096 17013 4136
rect 16971 4087 17013 4096
rect 17067 4136 17109 4145
rect 17067 4096 17068 4136
rect 17108 4096 17109 4136
rect 17067 4087 17109 4096
rect 17163 4136 17205 4145
rect 17163 4096 17164 4136
rect 17204 4096 17205 4136
rect 17163 4087 17205 4096
rect 17259 4136 17301 4145
rect 17259 4096 17260 4136
rect 17300 4096 17301 4136
rect 17259 4087 17301 4096
rect 17635 4136 17693 4137
rect 17635 4096 17644 4136
rect 17684 4096 17693 4136
rect 17635 4095 17693 4096
rect 17739 4136 17781 4145
rect 17739 4096 17740 4136
rect 17780 4096 17781 4136
rect 17739 4087 17781 4096
rect 17931 4136 17973 4145
rect 17931 4096 17932 4136
rect 17972 4096 17973 4136
rect 17931 4087 17973 4096
rect 18123 4136 18165 4145
rect 18123 4096 18124 4136
rect 18164 4096 18165 4136
rect 18123 4087 18165 4096
rect 18411 4136 18453 4145
rect 18411 4096 18412 4136
rect 18452 4096 18453 4136
rect 18411 4087 18453 4096
rect 18603 4136 18645 4145
rect 18603 4096 18604 4136
rect 18644 4096 18645 4136
rect 18603 4087 18645 4096
rect 18699 4136 18741 4145
rect 18699 4096 18700 4136
rect 18740 4096 18741 4136
rect 18699 4087 18741 4096
rect 18795 4136 18837 4145
rect 18795 4096 18796 4136
rect 18836 4096 18837 4136
rect 18795 4087 18837 4096
rect 18891 4136 18933 4145
rect 18891 4096 18892 4136
rect 18932 4096 18933 4136
rect 18891 4087 18933 4096
rect 19363 4136 19421 4137
rect 19363 4096 19372 4136
rect 19412 4096 19421 4136
rect 19363 4095 19421 4096
rect 20323 4136 20381 4137
rect 20323 4096 20332 4136
rect 20372 4096 20381 4136
rect 20323 4095 20381 4096
rect 20803 4136 20861 4137
rect 20803 4096 20812 4136
rect 20852 4096 20861 4136
rect 20803 4095 20861 4096
rect 20899 4136 20957 4137
rect 20899 4096 20908 4136
rect 20948 4096 20957 4136
rect 20899 4095 20957 4096
rect 23779 4136 23837 4137
rect 23779 4096 23788 4136
rect 23828 4096 23837 4136
rect 23779 4095 23837 4096
rect 24163 4136 24221 4137
rect 24163 4096 24172 4136
rect 24212 4096 24221 4136
rect 24163 4095 24221 4096
rect 24267 4136 24309 4145
rect 24267 4096 24268 4136
rect 24308 4096 24309 4136
rect 24267 4087 24309 4096
rect 25131 4136 25173 4145
rect 25131 4096 25132 4136
rect 25172 4096 25173 4136
rect 25131 4087 25173 4096
rect 25227 4136 25269 4145
rect 25227 4096 25228 4136
rect 25268 4096 25269 4136
rect 25227 4087 25269 4096
rect 25323 4136 25365 4145
rect 25323 4096 25324 4136
rect 25364 4096 25365 4136
rect 25323 4087 25365 4096
rect 25419 4136 25461 4145
rect 25419 4096 25420 4136
rect 25460 4096 25461 4136
rect 25419 4087 25461 4096
rect 25611 4136 25653 4145
rect 25611 4096 25612 4136
rect 25652 4096 25653 4136
rect 25611 4087 25653 4096
rect 25803 4136 25845 4145
rect 25803 4096 25804 4136
rect 25844 4096 25845 4136
rect 25803 4087 25845 4096
rect 25891 4136 25949 4137
rect 25891 4096 25900 4136
rect 25940 4096 25949 4136
rect 25891 4095 25949 4096
rect 26083 4136 26141 4137
rect 26083 4096 26092 4136
rect 26132 4096 26141 4136
rect 26083 4095 26141 4096
rect 26187 4136 26229 4145
rect 26187 4096 26188 4136
rect 26228 4096 26229 4136
rect 26187 4087 26229 4096
rect 26379 4136 26421 4145
rect 26379 4096 26380 4136
rect 26420 4096 26421 4136
rect 26379 4087 26421 4096
rect 26755 4136 26813 4137
rect 26755 4096 26764 4136
rect 26804 4096 26813 4136
rect 26755 4095 26813 4096
rect 26851 4136 26909 4137
rect 26851 4096 26860 4136
rect 26900 4096 26909 4136
rect 26851 4095 26909 4096
rect 27339 4136 27381 4145
rect 27339 4096 27340 4136
rect 27380 4096 27381 4136
rect 27339 4087 27381 4096
rect 27531 4136 27573 4145
rect 27531 4096 27532 4136
rect 27572 4096 27573 4136
rect 27531 4087 27573 4096
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 27811 4136 27869 4137
rect 27811 4096 27820 4136
rect 27860 4096 27869 4136
rect 27811 4095 27869 4096
rect 27915 4136 27957 4145
rect 27915 4096 27916 4136
rect 27956 4096 27957 4136
rect 27915 4087 27957 4096
rect 28107 4136 28149 4145
rect 28107 4096 28108 4136
rect 28148 4096 28149 4136
rect 28107 4087 28149 4096
rect 28587 4136 28629 4145
rect 28587 4096 28588 4136
rect 28628 4096 28629 4136
rect 28587 4087 28629 4096
rect 28675 4136 28733 4137
rect 28675 4096 28684 4136
rect 28724 4096 28733 4136
rect 28675 4095 28733 4096
rect 29251 4136 29309 4137
rect 29251 4096 29260 4136
rect 29300 4096 29309 4136
rect 29251 4095 29309 4096
rect 29539 4136 29597 4137
rect 29539 4096 29548 4136
rect 29588 4096 29597 4136
rect 29539 4095 29597 4096
rect 31371 4136 31413 4145
rect 31371 4096 31372 4136
rect 31412 4096 31413 4136
rect 31371 4087 31413 4096
rect 31467 4136 31509 4145
rect 31467 4096 31468 4136
rect 31508 4096 31509 4136
rect 31467 4087 31509 4096
rect 31563 4136 31605 4145
rect 31563 4096 31564 4136
rect 31604 4096 31605 4136
rect 31563 4087 31605 4096
rect 31659 4136 31701 4145
rect 31659 4096 31660 4136
rect 31700 4096 31701 4136
rect 31659 4087 31701 4096
rect 31851 4136 31893 4145
rect 31851 4096 31852 4136
rect 31892 4096 31893 4136
rect 31851 4087 31893 4096
rect 32227 4136 32285 4137
rect 32227 4096 32236 4136
rect 32276 4096 32285 4136
rect 32227 4095 32285 4096
rect 33091 4136 33149 4137
rect 33091 4096 33100 4136
rect 33140 4096 33149 4136
rect 33091 4095 33149 4096
rect 35307 4136 35349 4145
rect 35307 4096 35308 4136
rect 35348 4096 35349 4136
rect 35307 4087 35349 4096
rect 35875 4136 35933 4137
rect 35875 4096 35884 4136
rect 35924 4096 35933 4136
rect 35875 4095 35933 4096
rect 36259 4136 36317 4137
rect 36259 4096 36268 4136
rect 36308 4096 36317 4136
rect 36259 4095 36317 4096
rect 36651 4136 36693 4145
rect 36651 4096 36652 4136
rect 36692 4096 36693 4136
rect 36651 4087 36693 4096
rect 37315 4136 37373 4137
rect 37315 4096 37324 4136
rect 37364 4096 37373 4136
rect 37315 4095 37373 4096
rect 37507 4136 37565 4137
rect 37507 4096 37516 4136
rect 37556 4096 37565 4136
rect 37507 4095 37565 4096
rect 38187 4136 38229 4145
rect 38187 4096 38188 4136
rect 38228 4096 38229 4136
rect 38187 4087 38229 4096
rect 38379 4136 38421 4145
rect 38379 4096 38380 4136
rect 38420 4096 38421 4136
rect 38379 4087 38421 4096
rect 38755 4136 38813 4137
rect 38755 4096 38764 4136
rect 38804 4096 38813 4136
rect 38755 4095 38813 4096
rect 39619 4136 39677 4137
rect 39619 4096 39628 4136
rect 39668 4096 39677 4136
rect 39619 4095 39677 4096
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 36355 4052 36413 4053
rect 36355 4012 36364 4052
rect 36404 4012 36413 4052
rect 36355 4011 36413 4012
rect 643 3968 701 3969
rect 643 3928 652 3968
rect 692 3928 701 3968
rect 643 3927 701 3928
rect 6691 3968 6749 3969
rect 6691 3928 6700 3968
rect 6740 3928 6749 3968
rect 6691 3927 6749 3928
rect 6979 3968 7037 3969
rect 6979 3928 6988 3968
rect 7028 3928 7037 3968
rect 6979 3927 7037 3928
rect 7851 3968 7893 3977
rect 7851 3928 7852 3968
rect 7892 3928 7893 3968
rect 7851 3919 7893 3928
rect 10051 3968 10109 3969
rect 10051 3928 10060 3968
rect 10100 3928 10109 3968
rect 10051 3927 10109 3928
rect 10819 3968 10877 3969
rect 10819 3928 10828 3968
rect 10868 3928 10877 3968
rect 10819 3927 10877 3928
rect 11299 3968 11357 3969
rect 11299 3928 11308 3968
rect 11348 3928 11357 3968
rect 11299 3927 11357 3928
rect 12259 3968 12317 3969
rect 12259 3928 12268 3968
rect 12308 3928 12317 3968
rect 12259 3927 12317 3928
rect 17827 3968 17885 3969
rect 17827 3928 17836 3968
rect 17876 3928 17885 3968
rect 17827 3927 17885 3928
rect 20619 3968 20661 3977
rect 20619 3928 20620 3968
rect 20660 3928 20661 3968
rect 20619 3919 20661 3928
rect 24075 3964 24117 3973
rect 24075 3924 24076 3964
rect 24116 3924 24117 3964
rect 25699 3968 25757 3969
rect 25699 3928 25708 3968
rect 25748 3928 25757 3968
rect 25699 3927 25757 3928
rect 29067 3968 29109 3977
rect 29067 3928 29068 3968
rect 29108 3928 29109 3968
rect 24075 3915 24117 3924
rect 29067 3919 29109 3928
rect 34243 3968 34301 3969
rect 34243 3928 34252 3968
rect 34292 3928 34301 3968
rect 34243 3927 34301 3928
rect 28779 3910 28821 3919
rect 28779 3870 28780 3910
rect 28820 3870 28821 3910
rect 28779 3861 28821 3870
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 643 3632 701 3633
rect 643 3592 652 3632
rect 692 3592 701 3632
rect 643 3591 701 3592
rect 7747 3632 7805 3633
rect 7747 3592 7756 3632
rect 7796 3592 7805 3632
rect 7747 3591 7805 3592
rect 8131 3632 8189 3633
rect 8131 3592 8140 3632
rect 8180 3592 8189 3632
rect 8131 3591 8189 3592
rect 8811 3632 8853 3641
rect 8811 3592 8812 3632
rect 8852 3592 8853 3632
rect 8811 3583 8853 3592
rect 10155 3632 10197 3641
rect 10155 3592 10156 3632
rect 10196 3592 10197 3632
rect 10155 3583 10197 3592
rect 14083 3632 14141 3633
rect 14083 3592 14092 3632
rect 14132 3592 14141 3632
rect 14083 3591 14141 3592
rect 15811 3632 15869 3633
rect 15811 3592 15820 3632
rect 15860 3592 15869 3632
rect 15811 3591 15869 3592
rect 16771 3632 16829 3633
rect 16771 3592 16780 3632
rect 16820 3592 16829 3632
rect 16771 3591 16829 3592
rect 17539 3632 17597 3633
rect 17539 3592 17548 3632
rect 17588 3592 17597 3632
rect 17539 3591 17597 3592
rect 17731 3632 17789 3633
rect 17731 3592 17740 3632
rect 17780 3592 17789 3632
rect 17731 3591 17789 3592
rect 20611 3632 20669 3633
rect 20611 3592 20620 3632
rect 20660 3592 20669 3632
rect 20611 3591 20669 3592
rect 23779 3632 23837 3633
rect 23779 3592 23788 3632
rect 23828 3592 23837 3632
rect 23779 3591 23837 3592
rect 23971 3632 24029 3633
rect 23971 3592 23980 3632
rect 24020 3592 24029 3632
rect 23971 3591 24029 3592
rect 25515 3632 25557 3641
rect 25515 3592 25516 3632
rect 25556 3592 25557 3632
rect 25515 3583 25557 3592
rect 28579 3632 28637 3633
rect 28579 3592 28588 3632
rect 28628 3592 28637 3632
rect 28579 3591 28637 3592
rect 28867 3632 28925 3633
rect 28867 3592 28876 3632
rect 28916 3592 28925 3632
rect 28867 3591 28925 3592
rect 29155 3632 29213 3633
rect 29155 3592 29164 3632
rect 29204 3592 29213 3632
rect 29155 3591 29213 3592
rect 32899 3632 32957 3633
rect 32899 3592 32908 3632
rect 32948 3592 32957 3632
rect 32899 3591 32957 3592
rect 35011 3632 35069 3633
rect 35011 3592 35020 3632
rect 35060 3592 35069 3632
rect 35011 3591 35069 3592
rect 5355 3548 5397 3557
rect 5355 3508 5356 3548
rect 5396 3508 5397 3548
rect 5355 3499 5397 3508
rect 11691 3548 11733 3557
rect 11691 3508 11692 3548
rect 11732 3508 11733 3548
rect 11691 3499 11733 3508
rect 17059 3548 17117 3549
rect 17059 3508 17068 3548
rect 17108 3508 17117 3548
rect 17059 3507 17117 3508
rect 19747 3548 19805 3549
rect 19747 3508 19756 3548
rect 19796 3508 19805 3548
rect 19747 3507 19805 3508
rect 29251 3548 29309 3549
rect 29251 3508 29260 3548
rect 29300 3508 29309 3548
rect 29251 3507 29309 3508
rect 29739 3548 29781 3557
rect 29739 3508 29740 3548
rect 29780 3508 29781 3548
rect 29739 3499 29781 3508
rect 35299 3548 35357 3549
rect 35299 3508 35308 3548
rect 35348 3508 35357 3548
rect 35299 3507 35357 3508
rect 5731 3464 5789 3465
rect 5731 3424 5740 3464
rect 5780 3424 5789 3464
rect 5731 3423 5789 3424
rect 6595 3464 6653 3465
rect 6595 3424 6604 3464
rect 6644 3424 6653 3464
rect 6595 3423 6653 3424
rect 7939 3464 7997 3465
rect 7939 3424 7948 3464
rect 7988 3424 7997 3464
rect 7939 3423 7997 3424
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 8043 3415 8085 3424
rect 8235 3464 8277 3473
rect 8235 3424 8236 3464
rect 8276 3424 8277 3464
rect 8235 3415 8277 3424
rect 8715 3464 8757 3473
rect 8715 3424 8716 3464
rect 8756 3424 8757 3464
rect 8715 3415 8757 3424
rect 8907 3464 8949 3473
rect 8907 3424 8908 3464
rect 8948 3424 8949 3464
rect 8907 3415 8949 3424
rect 9003 3464 9045 3473
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9187 3464 9245 3465
rect 9187 3424 9196 3464
rect 9236 3424 9245 3464
rect 9187 3423 9245 3424
rect 9867 3464 9909 3473
rect 9867 3424 9868 3464
rect 9908 3424 9909 3464
rect 9867 3415 9909 3424
rect 10051 3464 10109 3465
rect 10051 3424 10060 3464
rect 10100 3424 10109 3464
rect 10051 3423 10109 3424
rect 11299 3464 11357 3465
rect 11299 3424 11308 3464
rect 11348 3424 11357 3464
rect 11299 3423 11357 3424
rect 12067 3464 12125 3465
rect 12067 3424 12076 3464
rect 12116 3424 12125 3464
rect 12067 3423 12125 3424
rect 12931 3464 12989 3465
rect 12931 3424 12940 3464
rect 12980 3424 12989 3464
rect 12931 3423 12989 3424
rect 15907 3464 15965 3465
rect 15907 3424 15916 3464
rect 15956 3424 15965 3464
rect 15907 3423 15965 3424
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 16299 3415 16341 3424
rect 16395 3464 16437 3473
rect 16395 3424 16396 3464
rect 16436 3424 16437 3464
rect 16395 3415 16437 3424
rect 16491 3464 16533 3473
rect 16491 3424 16492 3464
rect 16532 3424 16533 3464
rect 16491 3415 16533 3424
rect 16587 3464 16629 3473
rect 16587 3424 16588 3464
rect 16628 3424 16629 3464
rect 16587 3415 16629 3424
rect 16867 3464 16925 3465
rect 16867 3424 16876 3464
rect 16916 3424 16925 3464
rect 16867 3423 16925 3424
rect 17259 3464 17301 3473
rect 17259 3424 17260 3464
rect 17300 3424 17301 3464
rect 17259 3415 17301 3424
rect 17355 3464 17397 3473
rect 17355 3424 17356 3464
rect 17396 3424 17397 3464
rect 17355 3415 17397 3424
rect 17451 3464 17493 3473
rect 17451 3424 17452 3464
rect 17492 3424 17493 3464
rect 17451 3415 17493 3424
rect 17835 3464 17877 3473
rect 17835 3424 17836 3464
rect 17876 3424 17877 3464
rect 17835 3415 17877 3424
rect 17931 3464 17973 3473
rect 17931 3424 17932 3464
rect 17972 3424 17973 3464
rect 17931 3415 17973 3424
rect 18027 3464 18069 3473
rect 18027 3424 18028 3464
rect 18068 3424 18069 3464
rect 18027 3415 18069 3424
rect 19267 3464 19325 3465
rect 19267 3424 19276 3464
rect 19316 3424 19325 3464
rect 19267 3423 19325 3424
rect 19555 3464 19613 3465
rect 19555 3424 19564 3464
rect 19604 3424 19613 3464
rect 19555 3423 19613 3424
rect 20331 3464 20373 3473
rect 20331 3424 20332 3464
rect 20372 3424 20373 3464
rect 20331 3415 20373 3424
rect 20427 3464 20469 3473
rect 20427 3424 20428 3464
rect 20468 3424 20469 3464
rect 20427 3415 20469 3424
rect 20523 3464 20565 3473
rect 20523 3424 20524 3464
rect 20564 3424 20565 3464
rect 20523 3415 20565 3424
rect 20811 3464 20853 3473
rect 20811 3424 20812 3464
rect 20852 3424 20853 3464
rect 20811 3415 20853 3424
rect 20907 3464 20949 3473
rect 20907 3424 20908 3464
rect 20948 3424 20949 3464
rect 20907 3415 20949 3424
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 21099 3464 21141 3473
rect 21099 3424 21100 3464
rect 21140 3424 21141 3464
rect 21099 3415 21141 3424
rect 21291 3464 21333 3473
rect 21291 3424 21292 3464
rect 21332 3424 21333 3464
rect 21291 3415 21333 3424
rect 21387 3464 21429 3473
rect 21387 3424 21388 3464
rect 21428 3424 21429 3464
rect 21387 3415 21429 3424
rect 21483 3464 21525 3473
rect 21483 3424 21484 3464
rect 21524 3424 21525 3464
rect 21483 3415 21525 3424
rect 21579 3464 21621 3473
rect 21579 3424 21580 3464
rect 21620 3424 21621 3464
rect 21579 3415 21621 3424
rect 22435 3464 22493 3465
rect 22435 3424 22444 3464
rect 22484 3424 22493 3464
rect 22435 3423 22493 3424
rect 22627 3464 22685 3465
rect 22627 3424 22636 3464
rect 22676 3424 22685 3464
rect 22627 3423 22685 3424
rect 22731 3464 22773 3473
rect 22731 3424 22732 3464
rect 22772 3424 22773 3464
rect 22731 3415 22773 3424
rect 22923 3464 22965 3473
rect 22923 3424 22924 3464
rect 22964 3424 22965 3464
rect 22923 3415 22965 3424
rect 23499 3464 23541 3473
rect 23499 3424 23500 3464
rect 23540 3424 23541 3464
rect 23499 3415 23541 3424
rect 23595 3464 23637 3473
rect 23595 3424 23596 3464
rect 23636 3424 23637 3464
rect 23595 3415 23637 3424
rect 23691 3464 23733 3473
rect 23691 3424 23692 3464
rect 23732 3424 23733 3464
rect 23691 3415 23733 3424
rect 24075 3464 24117 3473
rect 24075 3424 24076 3464
rect 24116 3424 24117 3464
rect 24075 3415 24117 3424
rect 24171 3464 24213 3473
rect 24171 3424 24172 3464
rect 24212 3424 24213 3464
rect 24171 3415 24213 3424
rect 24267 3464 24309 3473
rect 24267 3424 24268 3464
rect 24308 3424 24309 3464
rect 24267 3415 24309 3424
rect 24451 3464 24509 3465
rect 24451 3424 24460 3464
rect 24500 3424 24509 3464
rect 24451 3423 24509 3424
rect 26371 3464 26429 3465
rect 26371 3424 26380 3464
rect 26420 3424 26429 3464
rect 26371 3423 26429 3424
rect 26763 3464 26805 3473
rect 26763 3424 26764 3464
rect 26804 3424 26805 3464
rect 26763 3415 26805 3424
rect 27427 3464 27485 3465
rect 27427 3424 27436 3464
rect 27476 3424 27485 3464
rect 27427 3423 27485 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 27907 3464 27965 3465
rect 27907 3424 27916 3464
rect 27956 3424 27965 3464
rect 27907 3423 27965 3424
rect 28107 3464 28149 3473
rect 28107 3424 28108 3464
rect 28148 3424 28149 3464
rect 28107 3415 28149 3424
rect 28203 3464 28245 3473
rect 28203 3424 28204 3464
rect 28244 3424 28245 3464
rect 28203 3415 28245 3424
rect 28299 3464 28341 3473
rect 28299 3424 28300 3464
rect 28340 3424 28341 3464
rect 28299 3415 28341 3424
rect 28395 3464 28437 3473
rect 28395 3424 28396 3464
rect 28436 3424 28437 3464
rect 28395 3415 28437 3424
rect 28675 3464 28733 3465
rect 28675 3424 28684 3464
rect 28724 3424 28733 3464
rect 28675 3423 28733 3424
rect 29355 3464 29397 3473
rect 29355 3424 29356 3464
rect 29396 3424 29397 3464
rect 29355 3415 29397 3424
rect 29451 3464 29493 3473
rect 29451 3424 29452 3464
rect 29492 3424 29493 3464
rect 29451 3415 29493 3424
rect 29635 3464 29693 3465
rect 29635 3424 29644 3464
rect 29684 3424 29693 3464
rect 29635 3423 29693 3424
rect 29835 3464 29877 3473
rect 29835 3424 29836 3464
rect 29876 3424 29877 3464
rect 29835 3415 29877 3424
rect 31275 3464 31317 3473
rect 31275 3424 31276 3464
rect 31316 3424 31317 3464
rect 31275 3415 31317 3424
rect 31371 3464 31413 3473
rect 31371 3424 31372 3464
rect 31412 3424 31413 3464
rect 31371 3415 31413 3424
rect 31467 3464 31509 3473
rect 31467 3424 31468 3464
rect 31508 3424 31509 3464
rect 31467 3415 31509 3424
rect 31563 3464 31605 3473
rect 31563 3424 31564 3464
rect 31604 3424 31605 3464
rect 31563 3415 31605 3424
rect 31755 3464 31797 3473
rect 31755 3424 31756 3464
rect 31796 3424 31797 3464
rect 31755 3415 31797 3424
rect 32043 3464 32085 3473
rect 32043 3424 32044 3464
rect 32084 3424 32085 3464
rect 32043 3415 32085 3424
rect 33571 3464 33629 3465
rect 33571 3424 33580 3464
rect 33620 3424 33629 3464
rect 33571 3423 33629 3424
rect 34339 3464 34397 3465
rect 34339 3424 34348 3464
rect 34388 3424 34397 3464
rect 34339 3423 34397 3424
rect 36163 3464 36221 3465
rect 36163 3424 36172 3464
rect 36212 3424 36221 3464
rect 36163 3423 36221 3424
rect 37227 3464 37269 3473
rect 37227 3424 37228 3464
rect 37268 3424 37269 3464
rect 37227 3415 37269 3424
rect 38371 3464 38429 3465
rect 38371 3424 38380 3464
rect 38420 3424 38429 3464
rect 38371 3423 38429 3424
rect 39235 3464 39293 3465
rect 39235 3424 39244 3464
rect 39284 3424 39293 3464
rect 39235 3423 39293 3424
rect 39627 3464 39669 3473
rect 39627 3424 39628 3464
rect 39668 3424 39669 3464
rect 39627 3415 39669 3424
rect 25315 3380 25373 3381
rect 25315 3340 25324 3380
rect 25364 3340 25373 3380
rect 25315 3339 25373 3340
rect 4779 3296 4821 3305
rect 4779 3256 4780 3296
rect 4820 3256 4821 3296
rect 4779 3247 4821 3256
rect 32331 3296 32373 3305
rect 32331 3256 32332 3296
rect 32372 3256 32373 3296
rect 32331 3247 32373 3256
rect 33771 3296 33813 3305
rect 33771 3256 33772 3296
rect 33812 3256 33813 3296
rect 33771 3247 33813 3256
rect 10627 3212 10685 3213
rect 10627 3172 10636 3212
rect 10676 3172 10685 3212
rect 10627 3171 10685 3172
rect 16099 3212 16157 3213
rect 16099 3172 16108 3212
rect 16148 3172 16157 3212
rect 16099 3171 16157 3172
rect 21763 3212 21821 3213
rect 21763 3172 21772 3212
rect 21812 3172 21821 3212
rect 21763 3171 21821 3172
rect 22923 3212 22965 3221
rect 22923 3172 22924 3212
rect 22964 3172 22965 3212
rect 22923 3163 22965 3172
rect 25123 3212 25181 3213
rect 25123 3172 25132 3212
rect 25172 3172 25181 3212
rect 25123 3171 25181 3172
rect 25699 3212 25757 3213
rect 25699 3172 25708 3212
rect 25748 3172 25757 3212
rect 25699 3171 25757 3172
rect 27627 3212 27669 3221
rect 27627 3172 27628 3212
rect 27668 3172 27669 3212
rect 27627 3163 27669 3172
rect 29163 3212 29205 3221
rect 29163 3172 29164 3212
rect 29204 3172 29205 3212
rect 29163 3163 29205 3172
rect 32043 3212 32085 3221
rect 32043 3172 32044 3212
rect 32084 3172 32085 3212
rect 32043 3163 32085 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 7371 2876 7413 2885
rect 7371 2836 7372 2876
rect 7412 2836 7413 2876
rect 7371 2827 7413 2836
rect 8227 2876 8285 2877
rect 8227 2836 8236 2876
rect 8276 2836 8285 2876
rect 8227 2835 8285 2836
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 16779 2876 16821 2885
rect 16779 2836 16780 2876
rect 16820 2836 16821 2876
rect 16779 2827 16821 2836
rect 20427 2876 20469 2885
rect 20427 2836 20428 2876
rect 20468 2836 20469 2876
rect 20427 2827 20469 2836
rect 24163 2876 24221 2877
rect 24163 2836 24172 2876
rect 24212 2836 24221 2876
rect 24163 2835 24221 2836
rect 25131 2876 25173 2885
rect 25131 2836 25132 2876
rect 25172 2836 25173 2876
rect 25131 2827 25173 2836
rect 26571 2876 26613 2885
rect 26571 2836 26572 2876
rect 26612 2836 26613 2876
rect 26571 2827 26613 2836
rect 27051 2876 27093 2885
rect 27051 2836 27052 2876
rect 27092 2836 27093 2876
rect 27051 2827 27093 2836
rect 35683 2876 35741 2877
rect 35683 2836 35692 2876
rect 35732 2836 35741 2876
rect 35683 2835 35741 2836
rect 36643 2876 36701 2877
rect 36643 2836 36652 2876
rect 36692 2836 36701 2876
rect 36643 2835 36701 2836
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 5835 2792 5877 2801
rect 5835 2752 5836 2792
rect 5876 2752 5877 2792
rect 5835 2743 5877 2752
rect 32427 2792 32469 2801
rect 32427 2752 32428 2792
rect 32468 2752 32469 2792
rect 32427 2743 32469 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 20619 2708 20661 2717
rect 20619 2668 20620 2708
rect 20660 2668 20661 2708
rect 20619 2659 20661 2668
rect 7075 2624 7133 2625
rect 7075 2584 7084 2624
rect 7124 2584 7133 2624
rect 7075 2583 7133 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7371 2624 7413 2633
rect 7371 2584 7372 2624
rect 7412 2584 7413 2624
rect 7371 2575 7413 2584
rect 7563 2624 7605 2633
rect 7563 2584 7564 2624
rect 7604 2584 7605 2624
rect 7563 2575 7605 2584
rect 7651 2624 7709 2625
rect 7651 2584 7660 2624
rect 7700 2584 7709 2624
rect 7651 2583 7709 2584
rect 9379 2624 9437 2625
rect 9379 2584 9388 2624
rect 9428 2584 9437 2624
rect 9379 2583 9437 2584
rect 10243 2624 10301 2625
rect 10243 2584 10252 2624
rect 10292 2584 10301 2624
rect 10243 2583 10301 2584
rect 10635 2624 10677 2633
rect 10635 2584 10636 2624
rect 10676 2584 10677 2624
rect 10635 2575 10677 2584
rect 15819 2624 15861 2633
rect 15819 2584 15820 2624
rect 15860 2584 15861 2624
rect 15819 2575 15861 2584
rect 15915 2624 15957 2633
rect 15915 2584 15916 2624
rect 15956 2584 15957 2624
rect 15915 2575 15957 2584
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 16107 2624 16149 2633
rect 16107 2584 16108 2624
rect 16148 2584 16149 2624
rect 16107 2575 16149 2584
rect 16299 2624 16341 2633
rect 16299 2584 16300 2624
rect 16340 2584 16341 2624
rect 16299 2575 16341 2584
rect 16491 2624 16533 2633
rect 17163 2626 17205 2635
rect 16491 2584 16492 2624
rect 16532 2584 16533 2624
rect 16491 2575 16533 2584
rect 16579 2624 16637 2625
rect 16579 2584 16588 2624
rect 16628 2584 16637 2624
rect 16579 2583 16637 2584
rect 16963 2624 17021 2625
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 16963 2583 17021 2584
rect 17059 2624 17117 2625
rect 17059 2584 17068 2624
rect 17108 2584 17117 2624
rect 17059 2583 17117 2584
rect 17163 2586 17164 2626
rect 17204 2586 17205 2626
rect 17163 2577 17205 2586
rect 17347 2624 17405 2625
rect 17347 2584 17356 2624
rect 17396 2584 17405 2624
rect 17347 2583 17405 2584
rect 17539 2624 17597 2625
rect 17539 2584 17548 2624
rect 17588 2584 17597 2624
rect 17539 2583 17597 2584
rect 17827 2624 17885 2625
rect 17827 2584 17836 2624
rect 17876 2584 17885 2624
rect 17827 2583 17885 2584
rect 18315 2624 18357 2633
rect 18315 2584 18316 2624
rect 18356 2584 18357 2624
rect 18315 2575 18357 2584
rect 18411 2624 18453 2633
rect 18411 2584 18412 2624
rect 18452 2584 18453 2624
rect 18411 2575 18453 2584
rect 18507 2624 18549 2633
rect 18507 2584 18508 2624
rect 18548 2584 18549 2624
rect 18507 2575 18549 2584
rect 19275 2624 19317 2633
rect 19275 2584 19276 2624
rect 19316 2584 19317 2624
rect 19275 2575 19317 2584
rect 19371 2624 19413 2633
rect 19371 2584 19372 2624
rect 19412 2584 19413 2624
rect 19371 2575 19413 2584
rect 19467 2624 19509 2633
rect 19467 2584 19468 2624
rect 19508 2584 19509 2624
rect 19467 2575 19509 2584
rect 19851 2624 19893 2633
rect 19851 2584 19852 2624
rect 19892 2584 19893 2624
rect 19851 2575 19893 2584
rect 19947 2624 19989 2633
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 20131 2624 20189 2625
rect 20131 2584 20140 2624
rect 20180 2584 20189 2624
rect 20131 2583 20189 2584
rect 20235 2624 20277 2633
rect 20235 2584 20236 2624
rect 20276 2584 20277 2624
rect 20235 2575 20277 2584
rect 20427 2624 20469 2633
rect 20427 2584 20428 2624
rect 20468 2584 20469 2624
rect 20427 2575 20469 2584
rect 21283 2624 21341 2625
rect 21283 2584 21292 2624
rect 21332 2584 21341 2624
rect 21283 2583 21341 2584
rect 21771 2624 21813 2633
rect 21771 2584 21772 2624
rect 21812 2584 21813 2624
rect 21771 2575 21813 2584
rect 22147 2624 22205 2625
rect 22147 2584 22156 2624
rect 22196 2584 22205 2624
rect 22147 2583 22205 2584
rect 23011 2624 23069 2625
rect 23011 2584 23020 2624
rect 23060 2584 23069 2624
rect 23011 2583 23069 2584
rect 25323 2624 25365 2633
rect 25323 2584 25324 2624
rect 25364 2584 25365 2624
rect 25323 2575 25365 2584
rect 25891 2624 25949 2625
rect 25891 2584 25900 2624
rect 25940 2584 25949 2624
rect 25891 2583 25949 2584
rect 27139 2624 27197 2625
rect 27139 2584 27148 2624
rect 27188 2584 27197 2624
rect 27139 2583 27197 2584
rect 27523 2624 27581 2625
rect 27523 2584 27532 2624
rect 27572 2584 27581 2624
rect 27523 2583 27581 2584
rect 27907 2624 27965 2625
rect 27907 2584 27916 2624
rect 27956 2584 27965 2624
rect 27907 2583 27965 2584
rect 28099 2624 28157 2625
rect 28099 2584 28108 2624
rect 28148 2584 28157 2624
rect 28099 2583 28157 2584
rect 28483 2624 28541 2625
rect 28483 2584 28492 2624
rect 28532 2584 28541 2624
rect 28483 2583 28541 2584
rect 29163 2624 29205 2633
rect 29163 2584 29164 2624
rect 29204 2584 29205 2624
rect 29163 2575 29205 2584
rect 29355 2624 29397 2633
rect 29355 2584 29356 2624
rect 29396 2584 29397 2624
rect 29355 2575 29397 2584
rect 29451 2624 29493 2633
rect 29451 2584 29452 2624
rect 29492 2584 29493 2624
rect 29451 2575 29493 2584
rect 29643 2624 29685 2633
rect 29643 2584 29644 2624
rect 29684 2584 29685 2624
rect 29643 2575 29685 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 29835 2624 29877 2633
rect 29835 2584 29836 2624
rect 29876 2584 29877 2624
rect 29835 2575 29877 2584
rect 29931 2624 29973 2633
rect 29931 2584 29932 2624
rect 29972 2584 29973 2624
rect 29931 2575 29973 2584
rect 30307 2624 30365 2625
rect 30307 2584 30316 2624
rect 30356 2584 30365 2624
rect 30307 2583 30365 2584
rect 31267 2624 31325 2625
rect 31267 2584 31276 2624
rect 31316 2584 31325 2624
rect 31267 2583 31325 2584
rect 31563 2624 31605 2633
rect 31563 2584 31564 2624
rect 31604 2584 31605 2624
rect 33291 2624 33333 2633
rect 31563 2575 31605 2584
rect 32227 2591 32285 2592
rect 32227 2551 32236 2591
rect 32276 2551 32285 2591
rect 33291 2584 33292 2624
rect 33332 2584 33333 2624
rect 33291 2575 33333 2584
rect 33667 2624 33725 2625
rect 33667 2584 33676 2624
rect 33716 2584 33725 2624
rect 33667 2583 33725 2584
rect 34531 2624 34589 2625
rect 34531 2584 34540 2624
rect 34580 2584 34589 2624
rect 34531 2583 34589 2584
rect 35971 2624 36029 2625
rect 35971 2584 35980 2624
rect 36020 2584 36029 2624
rect 35971 2583 36029 2584
rect 37507 2624 37565 2625
rect 37507 2584 37516 2624
rect 37556 2584 37565 2624
rect 37507 2583 37565 2584
rect 37611 2624 37653 2633
rect 37611 2584 37612 2624
rect 37652 2584 37653 2624
rect 37611 2575 37653 2584
rect 37803 2624 37845 2633
rect 37803 2584 37804 2624
rect 37844 2584 37845 2624
rect 37803 2575 37845 2584
rect 37987 2624 38045 2625
rect 37987 2584 37996 2624
rect 38036 2584 38045 2624
rect 37987 2583 38045 2584
rect 38187 2624 38229 2633
rect 38187 2584 38188 2624
rect 38228 2584 38229 2624
rect 38187 2575 38229 2584
rect 38275 2624 38333 2625
rect 38275 2584 38284 2624
rect 38324 2584 38333 2624
rect 38275 2583 38333 2584
rect 32227 2550 32285 2551
rect 18019 2540 18077 2541
rect 18019 2500 18028 2540
rect 18068 2500 18077 2540
rect 18019 2499 18077 2500
rect 18603 2540 18645 2549
rect 18603 2500 18604 2540
rect 18644 2500 18645 2540
rect 18603 2491 18645 2500
rect 27427 2540 27485 2541
rect 27427 2500 27436 2540
rect 27476 2500 27485 2540
rect 27427 2499 27485 2500
rect 28579 2540 28637 2541
rect 28579 2500 28588 2540
rect 28628 2500 28637 2540
rect 28579 2499 28637 2500
rect 37707 2540 37749 2549
rect 37707 2500 37708 2540
rect 37748 2500 37749 2540
rect 37707 2491 37749 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 19171 2456 19229 2457
rect 19171 2416 19180 2456
rect 19220 2416 19229 2456
rect 19171 2415 19229 2416
rect 19651 2456 19709 2457
rect 19651 2416 19660 2456
rect 19700 2416 19709 2456
rect 19651 2415 19709 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 17443 2120 17501 2121
rect 17443 2080 17452 2120
rect 17492 2080 17501 2120
rect 17443 2079 17501 2080
rect 21771 2120 21813 2129
rect 21771 2080 21772 2120
rect 21812 2080 21813 2120
rect 21771 2071 21813 2080
rect 22539 2036 22581 2045
rect 22539 1996 22540 2036
rect 22580 1996 22581 2036
rect 22539 1987 22581 1996
rect 22923 2036 22965 2045
rect 22923 1996 22924 2036
rect 22964 1996 22965 2036
rect 22923 1987 22965 1996
rect 16963 1962 17021 1963
rect 16299 1952 16341 1961
rect 16299 1912 16300 1952
rect 16340 1912 16341 1952
rect 16299 1903 16341 1912
rect 16491 1952 16533 1961
rect 16491 1912 16492 1952
rect 16532 1912 16533 1952
rect 16491 1903 16533 1912
rect 16875 1952 16917 1961
rect 16875 1912 16876 1952
rect 16916 1912 16917 1952
rect 16963 1922 16972 1962
rect 17012 1922 17021 1962
rect 16963 1921 17021 1922
rect 17547 1952 17589 1961
rect 16875 1903 16917 1912
rect 17547 1912 17548 1952
rect 17588 1912 17589 1952
rect 17547 1903 17589 1912
rect 17643 1952 17685 1961
rect 17643 1912 17644 1952
rect 17684 1912 17685 1952
rect 17643 1903 17685 1912
rect 17739 1952 17781 1961
rect 17739 1912 17740 1952
rect 17780 1912 17781 1952
rect 17739 1903 17781 1912
rect 17923 1952 17981 1953
rect 17923 1912 17932 1952
rect 17972 1912 17981 1952
rect 17923 1911 17981 1912
rect 18027 1952 18069 1961
rect 18027 1912 18028 1952
rect 18068 1912 18069 1952
rect 18027 1903 18069 1912
rect 18219 1952 18261 1961
rect 18219 1912 18220 1952
rect 18260 1912 18261 1952
rect 18219 1903 18261 1912
rect 18987 1952 19029 1961
rect 18987 1912 18988 1952
rect 19028 1912 19029 1952
rect 18987 1903 19029 1912
rect 19363 1952 19421 1953
rect 19363 1912 19372 1952
rect 19412 1912 19421 1952
rect 19363 1911 19421 1912
rect 20227 1952 20285 1953
rect 20227 1912 20236 1952
rect 20276 1912 20285 1952
rect 20227 1911 20285 1912
rect 21475 1952 21533 1953
rect 21475 1912 21484 1952
rect 21524 1912 21533 1952
rect 21475 1911 21533 1912
rect 21675 1952 21717 1961
rect 21675 1912 21676 1952
rect 21716 1912 21717 1952
rect 21675 1903 21717 1912
rect 21963 1952 22005 1961
rect 21963 1912 21964 1952
rect 22004 1912 22005 1952
rect 21963 1903 22005 1912
rect 22443 1952 22485 1961
rect 22443 1912 22444 1952
rect 22484 1912 22485 1952
rect 22443 1903 22485 1912
rect 22635 1952 22677 1961
rect 22635 1912 22636 1952
rect 22676 1912 22677 1952
rect 22635 1903 22677 1912
rect 23299 1952 23357 1953
rect 23299 1912 23308 1952
rect 23348 1912 23357 1952
rect 23299 1911 23357 1912
rect 24163 1952 24221 1953
rect 24163 1912 24172 1952
rect 24212 1912 24221 1952
rect 24163 1911 24221 1912
rect 25611 1952 25653 1961
rect 25611 1912 25612 1952
rect 25652 1912 25653 1952
rect 25611 1903 25653 1912
rect 25987 1952 26045 1953
rect 25987 1912 25996 1952
rect 26036 1912 26045 1952
rect 25987 1911 26045 1912
rect 26851 1952 26909 1953
rect 26851 1912 26860 1952
rect 26900 1912 26909 1952
rect 26851 1911 26909 1912
rect 28011 1952 28053 1961
rect 28011 1912 28012 1952
rect 28052 1912 28053 1952
rect 28011 1903 28053 1912
rect 28875 1952 28917 1961
rect 28875 1912 28876 1952
rect 28916 1912 28917 1952
rect 28875 1903 28917 1912
rect 29251 1952 29309 1953
rect 29251 1912 29260 1952
rect 29300 1912 29309 1952
rect 29251 1911 29309 1912
rect 30115 1952 30173 1953
rect 30115 1912 30124 1952
rect 30164 1912 30173 1952
rect 30115 1911 30173 1912
rect 31275 1952 31317 1961
rect 31275 1912 31276 1952
rect 31316 1912 31317 1952
rect 31275 1903 31317 1912
rect 31563 1952 31605 1961
rect 31563 1912 31564 1952
rect 31604 1912 31605 1952
rect 31563 1903 31605 1912
rect 31939 1952 31997 1953
rect 31939 1912 31948 1952
rect 31988 1912 31997 1952
rect 31939 1911 31997 1912
rect 32803 1952 32861 1953
rect 32803 1912 32812 1952
rect 32852 1912 32861 1952
rect 32803 1911 32861 1912
rect 34051 1952 34109 1953
rect 34051 1912 34060 1952
rect 34100 1912 34109 1952
rect 34051 1911 34109 1912
rect 17163 1784 17205 1793
rect 17163 1744 17164 1784
rect 17204 1744 17205 1784
rect 17163 1735 17205 1744
rect 18219 1784 18261 1793
rect 18219 1744 18220 1784
rect 18260 1744 18261 1784
rect 18219 1735 18261 1744
rect 18795 1784 18837 1793
rect 18795 1744 18796 1784
rect 18836 1744 18837 1784
rect 18795 1735 18837 1744
rect 16491 1700 16533 1709
rect 16491 1660 16492 1700
rect 16532 1660 16533 1700
rect 16491 1651 16533 1660
rect 25315 1700 25373 1701
rect 25315 1660 25324 1700
rect 25364 1660 25373 1700
rect 25315 1659 25373 1660
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 23403 1280 23445 1289
rect 23403 1240 23404 1280
rect 23444 1240 23445 1280
rect 23403 1231 23445 1240
rect 26091 1280 26133 1289
rect 26091 1240 26092 1280
rect 26132 1240 26133 1280
rect 26091 1231 26133 1240
rect 29643 1280 29685 1289
rect 29643 1240 29644 1280
rect 29684 1240 29685 1280
rect 29643 1231 29685 1240
rect 17355 1196 17397 1205
rect 17355 1156 17356 1196
rect 17396 1156 17397 1196
rect 17355 1147 17397 1156
rect 17259 1112 17301 1121
rect 17259 1072 17260 1112
rect 17300 1072 17301 1112
rect 17259 1063 17301 1072
rect 17451 1112 17493 1121
rect 17451 1072 17452 1112
rect 17492 1072 17493 1112
rect 17451 1063 17493 1072
rect 19275 1112 19317 1121
rect 19275 1072 19276 1112
rect 19316 1072 19317 1112
rect 19275 1063 19317 1072
rect 19467 1112 19509 1121
rect 19467 1072 19468 1112
rect 19508 1072 19509 1112
rect 19467 1063 19509 1072
rect 19555 1112 19613 1113
rect 19555 1072 19564 1112
rect 19604 1072 19613 1112
rect 19555 1071 19613 1072
rect 26659 1112 26717 1113
rect 26659 1072 26668 1112
rect 26708 1072 26717 1112
rect 26659 1071 26717 1072
rect 26851 1112 26909 1113
rect 26851 1072 26860 1112
rect 26900 1072 26909 1112
rect 26851 1071 26909 1072
rect 19363 944 19421 945
rect 19363 904 19372 944
rect 19412 904 19421 944
rect 19363 903 19421 904
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 9676 38368 9716 38408
rect 9580 38200 9620 38240
rect 9868 38200 9908 38240
rect 10540 38200 10580 38240
rect 10732 38200 10772 38240
rect 11596 38200 11636 38240
rect 11788 38200 11828 38240
rect 11884 38200 11924 38240
rect 8044 38032 8084 38072
rect 11596 38032 11636 38072
rect 12268 38032 12308 38072
rect 11404 37948 11444 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 9868 37612 9908 37652
rect 7084 37360 7124 37400
rect 7852 37360 7892 37400
rect 8716 37360 8756 37400
rect 10060 37360 10100 37400
rect 11596 37360 11636 37400
rect 12460 37360 12500 37400
rect 12844 37360 12884 37400
rect 13996 37360 14036 37400
rect 16396 37360 16436 37400
rect 7468 37276 7508 37316
rect 6988 37192 7028 37232
rect 9868 37192 9908 37232
rect 10156 37192 10196 37232
rect 10444 37192 10484 37232
rect 14668 37192 14708 37232
rect 15724 37192 15764 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 9964 36856 10004 36896
rect 15532 36856 15572 36896
rect 16492 36772 16532 36812
rect 6508 36688 6548 36728
rect 7180 36688 7220 36728
rect 7564 36688 7604 36728
rect 8428 36688 8468 36728
rect 10636 36688 10676 36728
rect 11116 36688 11156 36728
rect 11212 36688 11252 36728
rect 11404 36688 11444 36728
rect 11788 36688 11828 36728
rect 14860 36688 14900 36728
rect 14956 36688 14996 36728
rect 15340 36688 15380 36728
rect 15436 36688 15476 36728
rect 15628 36688 15668 36728
rect 15820 36688 15860 36728
rect 16684 36688 16724 36728
rect 16780 36688 16820 36728
rect 16876 36688 16916 36728
rect 16972 36688 17012 36728
rect 17548 36688 17588 36728
rect 6604 36604 6644 36644
rect 9580 36604 9620 36644
rect 4300 36520 4340 36560
rect 4684 36520 4724 36560
rect 6988 36520 7028 36560
rect 11404 36520 11444 36560
rect 12652 36520 12692 36560
rect 17164 36520 17204 36560
rect 9964 36436 10004 36476
rect 12460 36436 12500 36476
rect 17644 36436 17684 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 6892 36100 6932 36140
rect 8332 36100 8372 36140
rect 8524 36016 8564 36056
rect 11116 36016 11156 36056
rect 14572 36016 14612 36056
rect 19180 36016 19220 36056
rect 4300 35848 4340 35888
rect 5164 35848 5204 35888
rect 6604 35848 6644 35888
rect 6700 35848 6740 35888
rect 6892 35848 6932 35888
rect 7756 35848 7796 35888
rect 8044 35848 8084 35888
rect 8140 35848 8180 35888
rect 8332 35848 8372 35888
rect 9004 35848 9044 35888
rect 9100 35848 9140 35888
rect 9196 35848 9236 35888
rect 9388 35848 9428 35888
rect 9484 35848 9524 35888
rect 9580 35848 9620 35888
rect 9676 35848 9716 35888
rect 9868 35848 9908 35888
rect 9964 35848 10004 35888
rect 10060 35848 10100 35888
rect 10156 35848 10196 35888
rect 10444 35848 10484 35888
rect 10732 35848 10772 35888
rect 10828 35848 10868 35888
rect 11596 35848 11636 35888
rect 11788 35848 11828 35888
rect 11980 35848 12020 35888
rect 12364 35848 12404 35888
rect 13228 35848 13268 35888
rect 14860 35848 14900 35888
rect 14956 35848 14996 35888
rect 15244 35848 15284 35888
rect 15628 35848 15668 35888
rect 16012 35848 16052 35888
rect 16876 35848 16916 35888
rect 18316 35848 18356 35888
rect 21100 35848 21140 35888
rect 3916 35764 3956 35804
rect 8908 35764 8948 35804
rect 6316 35680 6356 35720
rect 7084 35680 7124 35720
rect 14380 35680 14420 35720
rect 18028 35680 18068 35720
rect 18988 35680 19028 35720
rect 21196 35680 21236 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 8524 35344 8564 35384
rect 9196 35344 9236 35384
rect 21100 35344 21140 35384
rect 3436 35260 3476 35300
rect 10924 35260 10964 35300
rect 16876 35260 16916 35300
rect 17164 35260 17204 35300
rect 18220 35260 18260 35300
rect 18412 35260 18452 35300
rect 3244 35176 3284 35216
rect 3340 35176 3380 35216
rect 3532 35176 3572 35216
rect 3724 35176 3764 35216
rect 3820 35176 3860 35216
rect 3916 35176 3956 35216
rect 4012 35176 4052 35216
rect 4204 35176 4244 35216
rect 4588 35176 4628 35216
rect 5452 35176 5492 35216
rect 6796 35176 6836 35216
rect 7660 35176 7700 35216
rect 8044 35176 8084 35216
rect 9580 35176 9620 35216
rect 9676 35176 9716 35216
rect 9772 35176 9812 35216
rect 9868 35176 9908 35216
rect 10732 35176 10772 35216
rect 11020 35176 11060 35216
rect 11116 35176 11156 35216
rect 11212 35176 11252 35216
rect 11404 35176 11444 35216
rect 12364 35176 12404 35216
rect 13420 35176 13460 35216
rect 13612 35176 13652 35216
rect 14092 35176 14132 35216
rect 15340 35176 15380 35216
rect 16204 35176 16244 35216
rect 16588 35176 16628 35216
rect 16684 35176 16724 35216
rect 16780 35176 16820 35216
rect 17068 35176 17108 35216
rect 17260 35176 17300 35216
rect 17356 35176 17396 35216
rect 17548 35176 17588 35216
rect 18796 35176 18836 35216
rect 19660 35176 19700 35216
rect 21772 35176 21812 35216
rect 24076 35176 24116 35216
rect 26476 35176 26516 35216
rect 30220 35176 30260 35216
rect 32140 35176 32180 35216
rect 6604 35092 6644 35132
rect 9388 35092 9428 35132
rect 1996 35008 2036 35048
rect 13228 35008 13268 35048
rect 21964 35008 22004 35048
rect 26668 35008 26708 35048
rect 29356 35008 29396 35048
rect 32716 35008 32756 35048
rect 7468 34924 7508 34964
rect 7756 34924 7796 34964
rect 8716 34924 8756 34964
rect 10060 34924 10100 34964
rect 14764 34924 14804 34964
rect 20812 34924 20852 34964
rect 23404 34924 23444 34964
rect 25804 34924 25844 34964
rect 29548 34924 29588 34964
rect 31468 34924 31508 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 5452 34588 5492 34628
rect 6796 34588 6836 34628
rect 10156 34588 10196 34628
rect 13324 34588 13364 34628
rect 31660 34588 31700 34628
rect 1324 34504 1364 34544
rect 10732 34504 10772 34544
rect 18316 34504 18356 34544
rect 18796 34504 18836 34544
rect 24844 34504 24884 34544
rect 35500 34504 35540 34544
rect 37996 34504 38036 34544
rect 1900 34336 1940 34376
rect 2764 34336 2804 34376
rect 4492 34336 4532 34376
rect 4588 34336 4628 34376
rect 4684 34336 4724 34376
rect 4780 34336 4820 34376
rect 5068 34336 5108 34376
rect 5164 34336 5204 34376
rect 5260 34381 5300 34421
rect 6124 34336 6164 34376
rect 6316 34336 6356 34376
rect 6412 34336 6452 34376
rect 6508 34336 6548 34376
rect 6604 34336 6644 34376
rect 6796 34336 6836 34376
rect 6988 34336 7028 34376
rect 7084 34336 7124 34376
rect 7276 34336 7316 34376
rect 7372 34336 7412 34376
rect 7564 34336 7604 34376
rect 8140 34336 8180 34376
rect 9004 34336 9044 34376
rect 10444 34336 10484 34376
rect 10540 34336 10580 34376
rect 10732 34336 10772 34376
rect 10924 34336 10964 34376
rect 11980 34336 12020 34376
rect 13036 34336 13076 34376
rect 13996 34336 14036 34376
rect 14380 34336 14420 34376
rect 14956 34336 14996 34376
rect 15820 34336 15860 34376
rect 17836 34336 17876 34376
rect 18508 34336 18548 34376
rect 18604 34336 18644 34376
rect 18796 34336 18836 34376
rect 19660 34336 19700 34376
rect 19852 34336 19892 34376
rect 19948 34336 19988 34376
rect 20044 34336 20084 34376
rect 20140 34315 20180 34355
rect 21196 34336 21236 34376
rect 21772 34336 21812 34376
rect 22636 34336 22676 34376
rect 24652 34336 24692 34376
rect 25612 34336 25652 34376
rect 26188 34336 26228 34376
rect 27052 34336 27092 34376
rect 29068 34336 29108 34376
rect 29260 34336 29300 34376
rect 29644 34336 29684 34376
rect 30508 34336 30548 34376
rect 32620 34336 32660 34376
rect 33484 34336 33524 34376
rect 36364 34336 36404 34376
rect 36556 34336 36596 34376
rect 36652 34336 36692 34376
rect 36748 34336 36788 34376
rect 37036 34336 37076 34376
rect 37228 34336 37268 34376
rect 1516 34252 1556 34292
rect 7756 34252 7796 34292
rect 14572 34252 14612 34292
rect 21388 34252 21428 34292
rect 25804 34252 25844 34292
rect 32236 34252 32276 34292
rect 37132 34252 37172 34292
rect 3916 34168 3956 34208
rect 4972 34168 5012 34208
rect 7468 34168 7508 34208
rect 10156 34168 10196 34208
rect 11596 34168 11636 34208
rect 12364 34168 12404 34208
rect 14284 34168 14324 34208
rect 16972 34168 17012 34208
rect 17164 34168 17204 34208
rect 18988 34168 19028 34208
rect 20524 34168 20564 34208
rect 23788 34168 23828 34208
rect 23980 34168 24020 34208
rect 25516 34168 25556 34208
rect 28204 34168 28244 34208
rect 28396 34168 28436 34208
rect 34636 34168 34676 34208
rect 35692 34168 35732 34208
rect 36844 34168 36884 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 6124 33832 6164 33872
rect 9388 33832 9428 33872
rect 13708 33832 13748 33872
rect 14956 33832 14996 33872
rect 18316 33832 18356 33872
rect 21388 33832 21428 33872
rect 22156 33832 22196 33872
rect 23116 33832 23156 33872
rect 26092 33832 26132 33872
rect 28972 33832 29012 33872
rect 30796 33832 30836 33872
rect 32236 33832 32276 33872
rect 37804 33832 37844 33872
rect 8140 33748 8180 33788
rect 11020 33748 11060 33788
rect 11308 33748 11348 33788
rect 16108 33748 16148 33788
rect 18988 33748 19028 33788
rect 23404 33748 23444 33788
rect 27148 33748 27188 33788
rect 35404 33748 35444 33788
rect 1228 33664 1268 33704
rect 1612 33664 1652 33704
rect 2476 33664 2516 33704
rect 3820 33664 3860 33704
rect 4012 33664 4052 33704
rect 4108 33664 4148 33704
rect 4300 33664 4340 33704
rect 4492 33664 4532 33704
rect 4588 33664 4628 33704
rect 4780 33664 4820 33704
rect 4876 33664 4916 33704
rect 4972 33664 5012 33704
rect 5068 33664 5108 33704
rect 5452 33664 5492 33704
rect 6412 33664 6452 33704
rect 6508 33684 6548 33724
rect 6892 33664 6932 33704
rect 6988 33664 7028 33704
rect 7468 33664 7508 33704
rect 7948 33650 7988 33690
rect 9484 33664 9524 33704
rect 10156 33664 10196 33704
rect 11692 33664 11732 33704
rect 12556 33664 12596 33704
rect 14764 33664 14804 33704
rect 15628 33664 15668 33704
rect 16780 33664 16820 33704
rect 17356 33664 17396 33704
rect 3628 33580 3668 33620
rect 16252 33622 16292 33662
rect 17740 33664 17780 33704
rect 17836 33664 17876 33704
rect 18220 33664 18260 33704
rect 18508 33664 18548 33704
rect 18700 33664 18740 33704
rect 18796 33664 18836 33704
rect 19372 33664 19412 33704
rect 20236 33664 20276 33704
rect 21580 33664 21620 33704
rect 21676 33664 21716 33704
rect 21772 33664 21812 33704
rect 21868 33664 21908 33704
rect 22060 33664 22100 33704
rect 22252 33664 22292 33704
rect 22348 33664 22388 33704
rect 22924 33664 22964 33704
rect 23020 33664 23060 33704
rect 23212 33664 23252 33704
rect 23788 33664 23828 33704
rect 24652 33664 24692 33704
rect 25996 33664 26036 33704
rect 26188 33664 26228 33704
rect 26284 33664 26324 33704
rect 26764 33664 26804 33704
rect 27052 33664 27092 33704
rect 28108 33664 28148 33704
rect 28204 33664 28244 33704
rect 28780 33664 28820 33704
rect 28876 33664 28916 33704
rect 29068 33664 29108 33704
rect 29932 33664 29972 33704
rect 30892 33664 30932 33704
rect 31084 33664 31124 33704
rect 31180 33664 31220 33704
rect 31276 33664 31316 33704
rect 31372 33664 31412 33704
rect 31564 33664 31604 33704
rect 31660 33664 31700 33704
rect 31756 33664 31796 33704
rect 31852 33664 31892 33704
rect 32044 33664 32084 33704
rect 32140 33664 32180 33704
rect 32332 33664 32372 33704
rect 32524 33664 32564 33704
rect 32908 33664 32948 33704
rect 33772 33664 33812 33704
rect 35212 33664 35252 33704
rect 35788 33664 35828 33704
rect 36652 33664 36692 33704
rect 37996 33664 38036 33704
rect 17260 33580 17300 33620
rect 25804 33580 25844 33620
rect 9868 33496 9908 33536
rect 28588 33496 28628 33536
rect 3820 33412 3860 33452
rect 4300 33412 4340 33452
rect 6124 33412 6164 33452
rect 14092 33412 14132 33452
rect 18508 33412 18548 33452
rect 21388 33412 21428 33452
rect 27436 33412 27476 33452
rect 29260 33412 29300 33452
rect 34924 33412 34964 33452
rect 35116 33412 35156 33452
rect 38668 33412 38708 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 2380 33076 2420 33116
rect 3244 33076 3284 33116
rect 5644 33076 5684 33116
rect 6220 33076 6260 33116
rect 19852 33076 19892 33116
rect 23500 33076 23540 33116
rect 24844 33076 24884 33116
rect 31948 33076 31988 33116
rect 34156 33076 34196 33116
rect 34348 33076 34388 33116
rect 35212 33076 35252 33116
rect 1612 32992 1652 33032
rect 6700 32992 6740 33032
rect 10636 32992 10676 33032
rect 19660 32992 19700 33032
rect 21292 32992 21332 33032
rect 33004 32992 33044 33032
rect 33676 32992 33716 33032
rect 36460 32992 36500 33032
rect 9292 32908 9332 32948
rect 12748 32908 12788 32948
rect 16396 32908 16436 32948
rect 19276 32908 19316 32948
rect 28588 32908 28628 32948
rect 33484 32908 33524 32948
rect 2476 32824 2516 32864
rect 2668 32824 2708 32864
rect 2764 32824 2804 32864
rect 2956 32824 2996 32864
rect 3052 32824 3092 32864
rect 3244 32824 3284 32864
rect 3532 32824 3572 32864
rect 3724 32824 3764 32864
rect 3916 32824 3956 32864
rect 4780 32824 4820 32864
rect 5644 32824 5684 32864
rect 5836 32824 5876 32864
rect 5932 32824 5972 32864
rect 6124 32824 6164 32864
rect 7276 32824 7316 32864
rect 8140 32824 8180 32864
rect 9964 32824 10004 32864
rect 10252 32824 10292 32864
rect 10348 32824 10388 32864
rect 10828 32824 10868 32864
rect 10924 32824 10964 32864
rect 11116 32824 11156 32864
rect 11404 32824 11444 32864
rect 11500 32824 11540 32864
rect 11596 32824 11636 32864
rect 11692 32824 11732 32864
rect 11884 32824 11924 32864
rect 11980 32824 12020 32864
rect 12076 32824 12116 32864
rect 12172 32824 12212 32864
rect 12556 32824 12596 32864
rect 13804 32824 13844 32864
rect 13996 32824 14036 32864
rect 14380 32824 14420 32864
rect 15244 32824 15284 32864
rect 16684 32824 16724 32864
rect 16780 32824 16820 32864
rect 16876 32824 16916 32864
rect 17548 32824 17588 32864
rect 18412 32824 18452 32864
rect 18604 32824 18644 32864
rect 19948 32824 19988 32864
rect 21580 32824 21620 32864
rect 21676 32824 21716 32864
rect 21964 32824 22004 32864
rect 23596 32824 23636 32864
rect 23788 32824 23828 32864
rect 23884 32824 23924 32864
rect 23980 32824 24020 32864
rect 24076 32824 24116 32864
rect 24364 32824 24404 32864
rect 25324 32824 25364 32864
rect 25708 32824 25748 32864
rect 25804 32824 25844 32864
rect 25900 32824 25940 32864
rect 25996 32824 26036 32864
rect 26572 32824 26612 32864
rect 27436 32824 27476 32864
rect 28780 32824 28820 32864
rect 29164 32824 29204 32864
rect 30028 32824 30068 32864
rect 31660 32824 31700 32864
rect 31756 32824 31796 32864
rect 31948 32824 31988 32864
rect 32140 32824 32180 32864
rect 33868 32824 33908 32864
rect 33964 32824 34004 32864
rect 34156 32824 34196 32864
rect 35020 32824 35060 32864
rect 35884 32824 35924 32864
rect 36172 32824 36212 32864
rect 36268 32824 36308 32864
rect 36460 32824 36500 32864
rect 36652 32824 36692 32864
rect 37900 32824 37940 32864
rect 38764 32824 38804 32864
rect 4588 32740 4628 32780
rect 5452 32740 5492 32780
rect 6892 32740 6932 32780
rect 11020 32740 11060 32780
rect 26188 32740 26228 32780
rect 37324 32740 37364 32780
rect 37516 32740 37556 32780
rect 12460 32656 12500 32696
rect 13132 32656 13172 32696
rect 16588 32656 16628 32696
rect 31180 32656 31220 32696
rect 32812 32656 32852 32696
rect 39916 32656 39956 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3724 32320 3764 32360
rect 5260 32320 5300 32360
rect 6412 32320 6452 32360
rect 6796 32320 6836 32360
rect 7276 32320 7316 32360
rect 13612 32320 13652 32360
rect 18124 32320 18164 32360
rect 22156 32320 22196 32360
rect 26380 32320 26420 32360
rect 31948 32320 31988 32360
rect 32428 32320 32468 32360
rect 33196 32320 33236 32360
rect 35788 32320 35828 32360
rect 36268 32320 36308 32360
rect 1132 32236 1172 32276
rect 31468 32236 31508 32276
rect 1516 32152 1556 32192
rect 2380 32152 2420 32192
rect 4396 32152 4436 32192
rect 5740 32152 5780 32192
rect 6124 32152 6164 32192
rect 6316 32152 6356 32192
rect 6700 32152 6740 32192
rect 7180 32152 7220 32192
rect 7372 32152 7412 32192
rect 7468 32152 7508 32192
rect 7948 32152 7988 32192
rect 8044 32152 8084 32192
rect 8140 32152 8180 32192
rect 8236 32152 8276 32192
rect 9580 32152 9620 32192
rect 10252 32152 10292 32192
rect 11116 32152 11156 32192
rect 11980 32152 12020 32192
rect 12172 32152 12212 32192
rect 12364 32152 12404 32192
rect 12748 32152 12788 32192
rect 13036 32152 13076 32192
rect 13132 32152 13172 32192
rect 14284 32152 14324 32192
rect 14476 32152 14516 32192
rect 14572 32152 14612 32192
rect 14668 32152 14708 32192
rect 14764 32152 14804 32192
rect 16012 32152 16052 32192
rect 16396 32152 16436 32192
rect 16588 32152 16628 32192
rect 17452 32152 17492 32192
rect 17836 32152 17876 32192
rect 17932 32152 17972 32192
rect 18028 32152 18068 32192
rect 18412 32152 18452 32192
rect 19660 32152 19700 32192
rect 20524 32152 20564 32192
rect 20908 32152 20948 32192
rect 22540 32152 22580 32192
rect 23212 32152 23252 32192
rect 25612 32152 25652 32192
rect 25900 32152 25940 32192
rect 25996 32152 26036 32192
rect 26188 32152 26228 32192
rect 27052 32152 27092 32192
rect 27244 32152 27284 32192
rect 27340 32152 27380 32192
rect 27436 32152 27476 32192
rect 27532 32152 27572 32192
rect 28780 32152 28820 32192
rect 28972 32152 29012 32192
rect 29644 32152 29684 32192
rect 30028 32152 30068 32192
rect 30124 32152 30164 32192
rect 30220 32152 30260 32192
rect 30316 32152 30356 32192
rect 30508 32152 30548 32192
rect 30700 32152 30740 32192
rect 30796 32152 30836 32192
rect 31084 32152 31124 32192
rect 31372 32152 31412 32192
rect 32044 32152 32084 32192
rect 32140 32152 32180 32192
rect 32236 32152 32276 32192
rect 32812 32152 32852 32192
rect 32908 32152 32948 32192
rect 33100 32152 33140 32192
rect 33772 32152 33812 32192
rect 34540 32152 34580 32192
rect 35692 32152 35732 32192
rect 35980 32152 36020 32192
rect 36076 32152 36116 32192
rect 36172 32152 36212 32192
rect 36460 32152 36500 32192
rect 36556 32152 36596 32192
rect 36652 32152 36692 32192
rect 36748 32152 36788 32192
rect 36940 32152 36980 32192
rect 37612 32152 37652 32192
rect 38092 32152 38132 32192
rect 39628 32152 39668 32192
rect 40588 32152 40628 32192
rect 32620 32068 32660 32108
rect 39724 32068 39764 32108
rect 6028 31984 6068 32024
rect 9388 31984 9428 32024
rect 14956 31984 14996 32024
rect 24268 31984 24308 32024
rect 26188 31984 26228 32024
rect 27724 31984 27764 32024
rect 34252 31984 34292 32024
rect 34828 31984 34868 32024
rect 38764 31984 38804 32024
rect 39244 31984 39284 32024
rect 3532 31900 3572 31940
rect 10444 31900 10484 31940
rect 11308 31900 11348 31940
rect 12268 31900 12308 31940
rect 13420 31900 13460 31940
rect 15340 31900 15380 31940
rect 16300 31900 16340 31940
rect 23788 31900 23828 31940
rect 24940 31900 24980 31940
rect 28684 31900 28724 31940
rect 30508 31900 30548 31940
rect 31756 31900 31796 31940
rect 33868 31900 33908 31940
rect 38572 31900 38612 31940
rect 39916 31900 39956 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 13996 31564 14036 31604
rect 15148 31564 15188 31604
rect 26188 31564 26228 31604
rect 29644 31564 29684 31604
rect 32428 31564 32468 31604
rect 37132 31564 37172 31604
rect 1324 31480 1364 31520
rect 3916 31480 3956 31520
rect 6316 31480 6356 31520
rect 6892 31480 6932 31520
rect 9772 31480 9812 31520
rect 12364 31480 12404 31520
rect 18220 31480 18260 31520
rect 18412 31480 18452 31520
rect 21676 31480 21716 31520
rect 26476 31480 26516 31520
rect 28300 31480 28340 31520
rect 41932 31480 41972 31520
rect 4876 31396 4916 31436
rect 1900 31312 1940 31352
rect 2764 31312 2804 31352
rect 4396 31312 4436 31352
rect 4492 31312 4532 31352
rect 4972 31312 5012 31352
rect 5452 31312 5492 31352
rect 5932 31317 5972 31357
rect 6412 31312 6452 31352
rect 7084 31312 7124 31352
rect 7756 31312 7796 31352
rect 8812 31312 8852 31352
rect 9676 31312 9716 31352
rect 9964 31312 10004 31352
rect 10348 31312 10388 31352
rect 11212 31312 11252 31352
rect 12556 31312 12596 31352
rect 12652 31312 12692 31352
rect 12748 31312 12788 31352
rect 13228 31312 13268 31352
rect 13324 31312 13364 31352
rect 13516 31312 13556 31352
rect 13612 31312 13652 31352
rect 13804 31312 13844 31352
rect 13996 31312 14036 31352
rect 14188 31312 14228 31352
rect 14284 31312 14324 31352
rect 14668 31312 14708 31352
rect 14860 31312 14900 31352
rect 14956 31312 14996 31352
rect 15148 31312 15188 31352
rect 15340 31312 15380 31352
rect 15436 31312 15476 31352
rect 15532 31312 15572 31352
rect 15628 31312 15668 31352
rect 15820 31312 15860 31352
rect 16012 31312 16052 31352
rect 16108 31312 16148 31352
rect 16300 31312 16340 31352
rect 17164 31312 17204 31352
rect 17836 31312 17876 31352
rect 20716 31312 20756 31352
rect 20908 31312 20948 31352
rect 22540 31312 22580 31352
rect 22732 31312 22772 31352
rect 22828 31312 22868 31352
rect 22924 31312 22964 31352
rect 24172 31312 24212 31352
rect 25036 31312 25076 31352
rect 26380 31312 26420 31352
rect 28108 31312 28148 31352
rect 29356 31312 29396 31352
rect 29452 31312 29492 31352
rect 29644 31312 29684 31352
rect 30508 31312 30548 31352
rect 30700 31312 30740 31352
rect 31660 31312 31700 31352
rect 31948 31312 31988 31352
rect 32908 31312 32948 31352
rect 33388 31312 33428 31352
rect 35116 31312 35156 31352
rect 35980 31312 36020 31352
rect 38188 31312 38228 31352
rect 38764 31312 38804 31352
rect 39628 31312 39668 31352
rect 43276 31312 43316 31352
rect 1516 31228 1556 31268
rect 8044 31228 8084 31268
rect 13708 31228 13748 31268
rect 15916 31228 15956 31268
rect 23788 31228 23828 31268
rect 34732 31228 34772 31268
rect 38380 31228 38420 31268
rect 6124 31144 6164 31184
rect 12844 31144 12884 31184
rect 14572 31144 14612 31184
rect 16972 31144 17012 31184
rect 21868 31144 21908 31184
rect 23020 31144 23060 31184
rect 27436 31144 27476 31184
rect 29836 31144 29876 31184
rect 33772 31144 33812 31184
rect 37516 31144 37556 31184
rect 40780 31144 40820 31184
rect 43180 31144 43220 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3916 30808 3956 30848
rect 4780 30808 4820 30848
rect 7564 30808 7604 30848
rect 10924 30808 10964 30848
rect 12844 30808 12884 30848
rect 16492 30808 16532 30848
rect 32236 30808 32276 30848
rect 33292 30808 33332 30848
rect 35596 30808 35636 30848
rect 38956 30808 38996 30848
rect 9964 30724 10004 30764
rect 13516 30724 13556 30764
rect 18892 30724 18932 30764
rect 21388 30724 21428 30764
rect 25996 30724 26036 30764
rect 26764 30724 26804 30764
rect 27436 30724 27476 30764
rect 36652 30724 36692 30764
rect 3724 30640 3764 30680
rect 4588 30640 4628 30680
rect 4876 30640 4916 30680
rect 4972 30640 5012 30680
rect 5068 30640 5108 30680
rect 5836 30640 5876 30680
rect 6028 30640 6068 30680
rect 6220 30640 6260 30680
rect 6316 30640 6356 30680
rect 6412 30640 6452 30680
rect 6508 30640 6548 30680
rect 8716 30640 8756 30680
rect 9580 30640 9620 30680
rect 10732 30640 10772 30680
rect 10828 30640 10868 30680
rect 11020 30640 11060 30680
rect 12076 30640 12116 30680
rect 12556 30640 12596 30680
rect 12652 30640 12692 30680
rect 12748 30640 12788 30680
rect 13132 30640 13172 30680
rect 13420 30640 13460 30680
rect 13996 30640 14036 30680
rect 15532 30640 15572 30680
rect 15820 30640 15860 30680
rect 15916 30640 15956 30680
rect 17644 30640 17684 30680
rect 18508 30640 18548 30680
rect 19084 30640 19124 30680
rect 19180 30640 19220 30680
rect 19276 30640 19316 30680
rect 19372 30640 19412 30680
rect 19660 30640 19700 30680
rect 19756 30640 19796 30680
rect 19852 30640 19892 30680
rect 20140 30640 20180 30680
rect 21100 30640 21140 30680
rect 21772 30640 21812 30680
rect 22636 30640 22676 30680
rect 25036 30640 25076 30680
rect 19948 30595 19988 30635
rect 25132 30640 25172 30680
rect 25228 30640 25268 30680
rect 25324 30640 25364 30680
rect 25612 30640 25652 30680
rect 25900 30640 25940 30680
rect 26476 30640 26516 30680
rect 26572 30640 26612 30680
rect 26668 30640 26708 30680
rect 26956 30640 26996 30680
rect 27052 30640 27092 30680
rect 27244 30640 27284 30680
rect 27820 30640 27860 30680
rect 28684 30640 28724 30680
rect 30028 30640 30068 30680
rect 31564 30640 31604 30680
rect 31756 30640 31796 30680
rect 31948 30640 31988 30680
rect 32044 30640 32084 30680
rect 32332 30640 32372 30680
rect 32428 30640 32468 30680
rect 32524 30640 32564 30680
rect 33676 30640 33716 30680
rect 34060 30640 34100 30680
rect 34252 30640 34292 30680
rect 34540 30640 34580 30680
rect 34636 30640 34676 30680
rect 34732 30640 34772 30680
rect 34828 30640 34868 30680
rect 35020 30640 35060 30680
rect 35116 30640 35156 30680
rect 35212 30640 35252 30680
rect 35308 30640 35348 30680
rect 35500 30640 35540 30680
rect 35692 30640 35732 30680
rect 35788 30640 35828 30680
rect 36460 30640 36500 30680
rect 36556 30640 36596 30680
rect 36748 30640 36788 30680
rect 36940 30640 36980 30680
rect 37036 30640 37076 30680
rect 37132 30640 37172 30680
rect 37228 30640 37268 30680
rect 37420 30640 37460 30680
rect 38284 30640 38324 30680
rect 39148 30640 39188 30680
rect 39244 30640 39284 30680
rect 39340 30640 39380 30680
rect 39436 30640 39476 30680
rect 40108 30640 40148 30680
rect 41452 30640 41492 30680
rect 41836 30640 41876 30680
rect 42700 30640 42740 30680
rect 44812 30640 44852 30680
rect 45484 30640 45524 30680
rect 45676 30640 45716 30680
rect 39628 30556 39668 30596
rect 1804 30472 1844 30512
rect 5356 30472 5396 30512
rect 11500 30472 11540 30512
rect 15052 30472 15092 30512
rect 27244 30472 27284 30512
rect 36172 30472 36212 30512
rect 44428 30472 44468 30512
rect 3052 30388 3092 30428
rect 13804 30388 13844 30428
rect 14668 30388 14708 30428
rect 16204 30388 16244 30428
rect 20620 30388 20660 30428
rect 23788 30388 23828 30428
rect 26284 30388 26324 30428
rect 29836 30388 29876 30428
rect 30700 30388 30740 30428
rect 30892 30388 30932 30428
rect 31756 30388 31796 30428
rect 38092 30388 38132 30428
rect 40012 30388 40052 30428
rect 43852 30388 43892 30428
rect 45772 30388 45812 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 3724 30052 3764 30092
rect 4876 30052 4916 30092
rect 6508 30052 6548 30092
rect 12460 30052 12500 30092
rect 13420 30052 13460 30092
rect 16492 30052 16532 30092
rect 22252 30052 22292 30092
rect 26764 30052 26804 30092
rect 36076 30052 36116 30092
rect 41644 30052 41684 30092
rect 7852 29968 7892 30008
rect 9868 29968 9908 30008
rect 20716 29968 20756 30008
rect 27724 29968 27764 30008
rect 29260 29968 29300 30008
rect 33388 29968 33428 30008
rect 40492 29968 40532 30008
rect 46636 29968 46676 30008
rect 37420 29884 37460 29924
rect 1324 29800 1364 29840
rect 1708 29800 1748 29840
rect 2572 29800 2612 29840
rect 4204 29800 4244 29840
rect 4300 29800 4340 29840
rect 4396 29800 4436 29840
rect 4588 29800 4628 29840
rect 4684 29800 4724 29840
rect 4876 29800 4916 29840
rect 5068 29800 5108 29840
rect 5164 29800 5204 29840
rect 5260 29800 5300 29840
rect 5356 29800 5396 29840
rect 6316 29800 6356 29840
rect 7180 29800 7220 29840
rect 7468 29800 7508 29840
rect 8044 29800 8084 29840
rect 8140 29800 8180 29840
rect 8236 29800 8276 29840
rect 8332 29800 8372 29840
rect 8524 29800 8564 29840
rect 8716 29800 8756 29840
rect 8812 29800 8852 29840
rect 9676 29800 9716 29840
rect 10924 29800 10964 29840
rect 11884 29800 11924 29840
rect 12172 29800 12212 29840
rect 13036 29800 13076 29840
rect 14572 29800 14612 29840
rect 15436 29800 15476 29840
rect 15820 29800 15860 29840
rect 16876 29800 16916 29840
rect 17260 29800 17300 29840
rect 18508 29800 18548 29840
rect 19372 29800 19412 29840
rect 21772 29800 21812 29840
rect 21964 29800 22004 29840
rect 22060 29800 22100 29840
rect 22252 29800 22292 29840
rect 22924 29800 22964 29840
rect 23788 29800 23828 29840
rect 25228 29800 25268 29840
rect 25420 29800 25460 29840
rect 25516 29800 25556 29840
rect 25708 29800 25748 29840
rect 26668 29800 26708 29840
rect 27052 29800 27092 29840
rect 27340 29800 27380 29840
rect 27436 29800 27476 29840
rect 29836 29800 29876 29840
rect 30700 29800 30740 29840
rect 32716 29800 32756 29840
rect 32908 29800 32948 29840
rect 33004 29800 33044 29840
rect 33100 29800 33140 29840
rect 33196 29800 33236 29840
rect 33964 29800 34004 29840
rect 34636 29800 34676 29840
rect 35020 29800 35060 29840
rect 35212 29800 35252 29840
rect 35308 29800 35348 29840
rect 35692 29800 35732 29840
rect 35884 29800 35924 29840
rect 36748 29800 36788 29840
rect 36940 29800 36980 29840
rect 37132 29800 37172 29840
rect 37228 29785 37268 29825
rect 38572 29800 38612 29840
rect 39436 29800 39476 29840
rect 39820 29800 39860 29840
rect 40684 29800 40724 29840
rect 40780 29800 40820 29840
rect 40972 29800 41012 29840
rect 41164 29800 41204 29840
rect 41260 29800 41300 29840
rect 41356 29800 41396 29840
rect 41452 29800 41492 29840
rect 42316 29800 42356 29840
rect 42604 29800 42644 29840
rect 42700 29800 42740 29840
rect 42796 29800 42836 29840
rect 43180 29800 43220 29840
rect 44428 29800 44468 29840
rect 45292 29800 45332 29840
rect 47884 29800 47924 29840
rect 8620 29716 8660 29756
rect 17932 29716 17972 29756
rect 18124 29716 18164 29756
rect 22540 29716 22580 29756
rect 25324 29716 25364 29756
rect 29452 29716 29492 29756
rect 35788 29716 35828 29756
rect 37036 29716 37076 29756
rect 43852 29716 43892 29756
rect 44044 29716 44084 29756
rect 4108 29632 4148 29672
rect 5644 29632 5684 29672
rect 6508 29632 6548 29672
rect 7372 29632 7412 29672
rect 9004 29632 9044 29672
rect 20524 29632 20564 29672
rect 21676 29632 21716 29672
rect 24940 29632 24980 29672
rect 26380 29632 26420 29672
rect 31852 29632 31892 29672
rect 32044 29632 32084 29672
rect 35116 29632 35156 29672
rect 40876 29632 40916 29672
rect 42508 29632 42548 29672
rect 46444 29632 46484 29672
rect 47788 29632 47828 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3724 29296 3764 29336
rect 7948 29296 7988 29336
rect 11788 29296 11828 29336
rect 16684 29296 16724 29336
rect 18700 29296 18740 29336
rect 23116 29296 23156 29336
rect 26572 29296 26612 29336
rect 34252 29296 34292 29336
rect 43756 29296 43796 29336
rect 48460 29296 48500 29336
rect 1324 29212 1364 29252
rect 3916 29212 3956 29252
rect 4876 29212 4916 29252
rect 8716 29212 8756 29252
rect 16972 29212 17012 29252
rect 23500 29212 23540 29252
rect 25900 29212 25940 29252
rect 26860 29212 26900 29252
rect 30988 29212 31028 29252
rect 31852 29212 31892 29252
rect 40396 29212 40436 29252
rect 1708 29128 1748 29168
rect 2572 29128 2612 29168
rect 4588 29128 4628 29168
rect 5260 29128 5300 29168
rect 6124 29128 6164 29168
rect 8428 29128 8468 29168
rect 9100 29128 9140 29168
rect 9964 29128 10004 29168
rect 12460 29128 12500 29168
rect 13516 29128 13556 29168
rect 13708 29128 13748 29168
rect 14572 29128 14612 29168
rect 14860 29128 14900 29168
rect 16108 29128 16148 29168
rect 16492 29128 16532 29168
rect 16588 29128 16628 29168
rect 16780 29128 16820 29168
rect 17644 29128 17684 29168
rect 17836 29128 17876 29168
rect 19372 29128 19412 29168
rect 19564 29128 19604 29168
rect 19756 29128 19796 29168
rect 19852 29128 19892 29168
rect 20620 29128 20660 29168
rect 21484 29128 21524 29168
rect 22540 29128 22580 29168
rect 22636 29128 22676 29168
rect 22732 29128 22772 29168
rect 22828 29128 22868 29168
rect 23020 29128 23060 29168
rect 23212 29128 23252 29168
rect 23308 29128 23348 29168
rect 24172 29128 24212 29168
rect 24940 29128 24980 29168
rect 25036 29128 25076 29168
rect 25132 29128 25172 29168
rect 25228 29128 25268 29168
rect 25516 29128 25556 29168
rect 25804 29128 25844 29168
rect 26668 29128 26708 29168
rect 27532 29128 27572 29168
rect 27724 29128 27764 29168
rect 28108 29128 28148 29168
rect 28204 29128 28244 29168
rect 28300 29128 28340 29168
rect 28396 29128 28436 29168
rect 29260 29128 29300 29168
rect 29452 29128 29492 29168
rect 30412 29128 30452 29168
rect 31084 29128 31124 29168
rect 31372 29128 31412 29168
rect 32236 29128 32276 29168
rect 33100 29128 33140 29168
rect 34444 29128 34484 29168
rect 35692 29128 35732 29168
rect 36556 29128 36596 29168
rect 36940 29128 36980 29168
rect 37228 29128 37268 29168
rect 37324 29128 37364 29168
rect 37420 29128 37460 29168
rect 37516 29128 37556 29168
rect 39532 29128 39572 29168
rect 40780 29128 40820 29168
rect 41644 29128 41684 29168
rect 43084 29128 43124 29168
rect 44044 29128 44084 29168
rect 44140 29128 44180 29168
rect 44236 29128 44276 29168
rect 44332 29128 44372 29168
rect 45484 29128 45524 29168
rect 45868 29128 45908 29168
rect 46252 29128 46292 29168
rect 47116 29128 47156 29168
rect 49132 29128 49172 29168
rect 7276 29044 7316 29084
rect 27820 29044 27860 29084
rect 29164 29044 29204 29084
rect 48268 29044 48308 29084
rect 1132 28960 1172 29000
rect 15916 28960 15956 29000
rect 24748 28960 24788 29000
rect 30700 28960 30740 29000
rect 38092 28960 38132 29000
rect 40204 28960 40244 29000
rect 42796 28960 42836 29000
rect 45196 28960 45236 29000
rect 11116 28876 11156 28916
rect 13612 28876 13652 28916
rect 14476 28876 14516 28916
rect 14764 28876 14804 28916
rect 18508 28876 18548 28916
rect 19564 28876 19604 28916
rect 20812 28876 20852 28916
rect 26188 28876 26228 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 2572 28540 2612 28580
rect 3532 28540 3572 28580
rect 6124 28540 6164 28580
rect 15244 28540 15284 28580
rect 18412 28540 18452 28580
rect 18604 28540 18644 28580
rect 22252 28540 22292 28580
rect 26860 28540 26900 28580
rect 30604 28540 30644 28580
rect 32524 28540 32564 28580
rect 35116 28540 35156 28580
rect 37036 28540 37076 28580
rect 40780 28540 40820 28580
rect 43180 28540 43220 28580
rect 1708 28456 1748 28496
rect 13612 28456 13652 28496
rect 23500 28456 23540 28496
rect 32908 28456 32948 28496
rect 33388 28456 33428 28496
rect 37708 28456 37748 28496
rect 41836 28456 41876 28496
rect 45580 28456 45620 28496
rect 48748 28456 48788 28496
rect 49228 28456 49268 28496
rect 7852 28372 7892 28412
rect 30220 28372 30260 28412
rect 2668 28288 2708 28328
rect 2860 28288 2900 28328
rect 3820 28288 3860 28328
rect 4780 28288 4820 28328
rect 4972 28288 5012 28328
rect 5068 28288 5108 28328
rect 5164 28288 5204 28328
rect 5452 28288 5492 28328
rect 5836 28288 5876 28328
rect 6124 28288 6164 28328
rect 6316 28288 6356 28328
rect 6412 28288 6452 28328
rect 7564 28288 7604 28328
rect 8524 28288 8564 28328
rect 8716 28288 8756 28328
rect 10348 28288 10388 28328
rect 11692 28288 11732 28328
rect 12556 28288 12596 28328
rect 14188 28288 14228 28328
rect 15724 28288 15764 28328
rect 16396 28288 16436 28328
rect 17260 28288 17300 28328
rect 18700 28288 18740 28328
rect 18988 28288 19028 28328
rect 20236 28288 20276 28328
rect 21100 28288 21140 28328
rect 24844 28288 24884 28328
rect 25708 28288 25748 28328
rect 27340 28288 27380 28328
rect 27436 28288 27476 28328
rect 27628 28288 27668 28328
rect 28204 28288 28244 28328
rect 29068 28288 29108 28328
rect 31276 28288 31316 28328
rect 31468 28288 31508 28328
rect 31564 28288 31604 28328
rect 31756 28288 31796 28328
rect 31948 28288 31988 28328
rect 32044 28288 32084 28328
rect 32140 28288 32180 28328
rect 32236 28288 32276 28328
rect 32428 28288 32468 28328
rect 33100 28273 33140 28313
rect 33196 28288 33236 28328
rect 33388 28288 33428 28328
rect 33580 28288 33620 28328
rect 34444 28288 34484 28328
rect 35404 28288 35444 28328
rect 35692 28288 35732 28328
rect 35884 28288 35924 28328
rect 36844 28288 36884 28328
rect 37132 28288 37172 28328
rect 38380 28288 38420 28328
rect 40300 28288 40340 28328
rect 40492 28288 40532 28328
rect 40588 28288 40628 28328
rect 40780 28288 40820 28328
rect 40972 28288 41012 28328
rect 42124 28288 42164 28328
rect 42220 28288 42260 28328
rect 42508 28288 42548 28328
rect 42892 28288 42932 28328
rect 42988 28288 43028 28328
rect 43180 28288 43220 28328
rect 43372 28288 43412 28328
rect 43468 28288 43508 28328
rect 43660 28288 43700 28328
rect 43852 28288 43892 28328
rect 43948 28288 43988 28328
rect 44044 28288 44084 28328
rect 44140 28333 44180 28373
rect 44332 28288 44372 28328
rect 45196 28288 45236 28328
rect 46156 28288 46196 28328
rect 46444 28288 46484 28328
rect 47116 28288 47156 28328
rect 47404 28288 47444 28328
rect 47500 28288 47540 28328
rect 47596 28288 47636 28328
rect 47692 28288 47732 28328
rect 48556 28288 48596 28328
rect 48748 28288 48788 28328
rect 48940 28288 48980 28328
rect 49036 28288 49076 28328
rect 50572 28288 50612 28328
rect 6700 28204 6740 28244
rect 12940 28204 12980 28244
rect 16012 28204 16052 28244
rect 19660 28204 19700 28244
rect 19852 28204 19892 28244
rect 24460 28204 24500 28244
rect 27820 28204 27860 28244
rect 39244 28204 39284 28244
rect 43564 28204 43604 28244
rect 4108 28120 4148 28160
rect 5260 28120 5300 28160
rect 5548 28120 5588 28160
rect 5740 28120 5780 28160
rect 9388 28120 9428 28160
rect 9676 28120 9716 28160
rect 10540 28120 10580 28160
rect 27532 28120 27572 28160
rect 31660 28120 31700 28160
rect 34252 28120 34292 28160
rect 36172 28120 36212 28160
rect 39628 28120 39668 28160
rect 41644 28120 41684 28160
rect 46060 28120 46100 28160
rect 47884 28120 47924 28160
rect 49900 28120 49940 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 23596 27784 23636 27824
rect 33676 27784 33716 27824
rect 5260 27700 5300 27740
rect 9676 27700 9716 27740
rect 11596 27700 11636 27740
rect 15340 27700 15380 27740
rect 17452 27700 17492 27740
rect 20716 27700 20756 27740
rect 25996 27700 26036 27740
rect 29836 27700 29876 27740
rect 31276 27700 31316 27740
rect 34156 27700 34196 27740
rect 39532 27700 39572 27740
rect 42220 27700 42260 27740
rect 47884 27700 47924 27740
rect 1228 27616 1268 27656
rect 1612 27616 1652 27656
rect 2476 27616 2516 27656
rect 3820 27616 3860 27656
rect 3916 27616 3956 27656
rect 4108 27616 4148 27656
rect 4492 27616 4532 27656
rect 5644 27616 5684 27656
rect 5932 27616 5972 27656
rect 6028 27616 6068 27656
rect 6604 27616 6644 27656
rect 6796 27616 6836 27656
rect 6892 27616 6932 27656
rect 6988 27616 7028 27656
rect 7084 27616 7124 27656
rect 8428 27616 8468 27656
rect 9292 27616 9332 27656
rect 10924 27616 10964 27656
rect 11212 27616 11252 27656
rect 11500 27616 11540 27656
rect 12076 27616 12116 27656
rect 13036 27616 13076 27656
rect 13324 27616 13364 27656
rect 14188 27616 14228 27656
rect 14572 27616 14612 27656
rect 14764 27616 14804 27656
rect 14860 27616 14900 27656
rect 15436 27616 15476 27656
rect 15724 27616 15764 27656
rect 17356 27616 17396 27656
rect 17548 27616 17588 27656
rect 17644 27616 17684 27656
rect 18124 27616 18164 27656
rect 18220 27616 18260 27656
rect 18508 27616 18548 27656
rect 18796 27616 18836 27656
rect 18892 27616 18932 27656
rect 18988 27616 19028 27656
rect 19084 27616 19124 27656
rect 19564 27616 19604 27656
rect 20524 27616 20564 27656
rect 20812 27616 20852 27656
rect 21004 27616 21044 27656
rect 21676 27616 21716 27656
rect 21868 27616 21908 27656
rect 22828 27616 22868 27656
rect 23980 27616 24020 27656
rect 24748 27616 24788 27656
rect 24844 27616 24884 27656
rect 25036 27616 25076 27656
rect 25228 27616 25268 27656
rect 25324 27616 25364 27656
rect 25612 27616 25652 27656
rect 25900 27616 25940 27656
rect 27820 27616 27860 27656
rect 27916 27616 27956 27656
rect 28108 27616 28148 27656
rect 29740 27616 29780 27656
rect 30028 27616 30068 27656
rect 30124 27616 30164 27656
rect 30220 27616 30260 27656
rect 30316 27616 30356 27656
rect 30508 27616 30548 27656
rect 30700 27616 30740 27656
rect 30796 27616 30836 27656
rect 31372 27616 31412 27656
rect 31660 27616 31700 27656
rect 32620 27616 32660 27656
rect 33388 27616 33428 27656
rect 33772 27616 33812 27656
rect 33868 27616 33908 27656
rect 33964 27616 34004 27656
rect 34540 27616 34580 27656
rect 35404 27616 35444 27656
rect 36940 27616 36980 27656
rect 37324 27616 37364 27656
rect 38188 27616 38228 27656
rect 39916 27616 39956 27656
rect 40780 27616 40820 27656
rect 42124 27616 42164 27656
rect 43756 27616 43796 27656
rect 44140 27616 44180 27656
rect 44524 27616 44564 27656
rect 45388 27616 45428 27656
rect 46828 27616 46868 27656
rect 47692 27616 47732 27656
rect 48268 27616 48308 27656
rect 49132 27616 49172 27656
rect 51148 27616 51188 27656
rect 3628 27532 3668 27572
rect 28684 27532 28724 27572
rect 39340 27532 39380 27572
rect 50284 27532 50324 27572
rect 4108 27448 4148 27488
rect 10060 27448 10100 27488
rect 16492 27448 16532 27488
rect 23788 27448 23828 27488
rect 25036 27448 25076 27488
rect 28876 27448 28916 27488
rect 32812 27448 32852 27488
rect 36556 27448 36596 27488
rect 41932 27448 41972 27488
rect 4684 27364 4724 27404
rect 6316 27364 6356 27404
rect 6508 27364 6548 27404
rect 7276 27364 7316 27404
rect 10252 27364 10292 27404
rect 11884 27364 11924 27404
rect 12364 27364 12404 27404
rect 14572 27364 14612 27404
rect 15052 27364 15092 27404
rect 17836 27364 17876 27404
rect 19852 27364 19892 27404
rect 26284 27364 26324 27404
rect 28108 27364 28148 27404
rect 28492 27364 28532 27404
rect 30508 27364 30548 27404
rect 30988 27364 31028 27404
rect 31948 27364 31988 27404
rect 33292 27364 33332 27404
rect 43564 27364 43604 27404
rect 46540 27364 46580 27404
rect 46732 27364 46772 27404
rect 47020 27364 47060 27404
rect 50476 27364 50516 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 2764 27028 2804 27068
rect 4876 27028 4916 27068
rect 8428 27028 8468 27068
rect 9292 27028 9332 27068
rect 12460 27028 12500 27068
rect 17740 27028 17780 27068
rect 20524 27028 20564 27068
rect 24076 27028 24116 27068
rect 30988 27028 31028 27068
rect 34252 27028 34292 27068
rect 37708 27028 37748 27068
rect 39436 27028 39476 27068
rect 40492 27028 40532 27068
rect 42988 27028 43028 27068
rect 45100 27028 45140 27068
rect 45580 27028 45620 27068
rect 46540 27028 46580 27068
rect 51724 27028 51764 27068
rect 2188 26944 2228 26984
rect 9100 26944 9140 26984
rect 11500 26944 11540 26984
rect 13228 26944 13268 26984
rect 23404 26944 23444 26984
rect 38476 26944 38516 26984
rect 40012 26944 40052 26984
rect 27436 26860 27476 26900
rect 30124 26860 30164 26900
rect 2860 26776 2900 26816
rect 3148 26776 3188 26816
rect 3340 26776 3380 26816
rect 3436 26776 3476 26816
rect 3628 26776 3668 26816
rect 3916 26776 3956 26816
rect 4012 26776 4052 26816
rect 4108 26776 4148 26816
rect 4396 26776 4436 26816
rect 4492 26776 4532 26816
rect 4588 26776 4628 26816
rect 4684 26776 4724 26816
rect 5548 26776 5588 26816
rect 5740 26776 5780 26816
rect 5932 26776 5972 26816
rect 6028 26776 6068 26816
rect 6220 26776 6260 26816
rect 6412 26776 6452 26816
rect 7564 26776 7604 26816
rect 7852 26776 7892 26816
rect 7948 26776 7988 26816
rect 8140 26776 8180 26816
rect 8332 26776 8372 26816
rect 8524 26776 8564 26816
rect 9292 26776 9332 26816
rect 9484 26776 9524 26816
rect 9580 26776 9620 26816
rect 9772 26776 9812 26816
rect 9868 26776 9908 26816
rect 9964 26776 10004 26816
rect 10252 26776 10292 26816
rect 10348 26776 10388 26816
rect 10444 26776 10484 26816
rect 10540 26776 10580 26816
rect 10828 26776 10868 26816
rect 11116 26776 11156 26816
rect 11692 26776 11732 26816
rect 12460 26776 12500 26816
rect 12652 26776 12692 26816
rect 12748 26776 12788 26816
rect 12940 26776 12980 26816
rect 13036 26776 13076 26816
rect 13228 26776 13268 26816
rect 13420 26776 13460 26816
rect 13516 26776 13556 26816
rect 13708 26776 13748 26816
rect 13804 26776 13844 26816
rect 13961 26791 14001 26831
rect 14188 26776 14228 26816
rect 14284 26776 14324 26816
rect 14476 26776 14516 26816
rect 14572 26776 14612 26816
rect 14727 26776 14767 26816
rect 14956 26776 14996 26816
rect 15148 26776 15188 26816
rect 15340 26776 15380 26816
rect 15436 26776 15476 26816
rect 15628 26776 15668 26816
rect 16012 26776 16052 26816
rect 16108 26776 16148 26816
rect 16300 26776 16340 26816
rect 16588 26776 16628 26816
rect 16780 26776 16820 26816
rect 16972 26776 17012 26816
rect 17164 26776 17204 26816
rect 17836 26776 17876 26816
rect 18124 26776 18164 26816
rect 18220 26776 18260 26816
rect 18316 26776 18356 26816
rect 18604 26776 18644 26816
rect 18700 26776 18740 26816
rect 18796 26776 18836 26816
rect 19084 26776 19124 26816
rect 19276 26776 19316 26816
rect 19372 26776 19412 26816
rect 19564 26776 19604 26816
rect 20236 26776 20276 26816
rect 21676 26776 21716 26816
rect 22540 26776 22580 26816
rect 24460 26776 24500 26816
rect 24940 26776 24980 26816
rect 25036 26776 25076 26816
rect 25132 26776 25172 26816
rect 25420 26776 25460 26816
rect 25612 26776 25652 26816
rect 25708 26776 25748 26816
rect 26572 26776 26612 26816
rect 26956 26776 26996 26816
rect 27052 26776 27092 26816
rect 27532 26776 27572 26816
rect 28012 26776 28052 26816
rect 28492 26781 28532 26821
rect 28876 26776 28916 26816
rect 29068 26776 29108 26816
rect 29164 26776 29204 26816
rect 29548 26776 29588 26816
rect 29644 26776 29684 26816
rect 30508 26776 30548 26816
rect 30604 26776 30644 26816
rect 30700 26776 30740 26816
rect 30988 26776 31028 26816
rect 31180 26776 31220 26816
rect 31276 26776 31316 26816
rect 31852 26776 31892 26816
rect 32236 26776 32276 26816
rect 33100 26776 33140 26816
rect 34636 26776 34676 26816
rect 34732 26776 34772 26816
rect 34924 26776 34964 26816
rect 35404 26776 35444 26816
rect 35596 26776 35636 26816
rect 35788 26776 35828 26816
rect 38188 26776 38228 26816
rect 38764 26776 38804 26816
rect 38860 26776 38900 26816
rect 39148 26776 39188 26816
rect 39436 26776 39476 26816
rect 39628 26776 39668 26816
rect 39724 26776 39764 26816
rect 40396 26776 40436 26816
rect 41068 26776 41108 26816
rect 42028 26776 42068 26816
rect 42700 26776 42740 26816
rect 42796 26776 42836 26816
rect 42988 26776 43028 26816
rect 43180 26776 43220 26816
rect 43276 26776 43316 26816
rect 43372 26776 43412 26816
rect 43468 26776 43508 26816
rect 43660 26776 43700 26816
rect 43756 26776 43796 26816
rect 43948 26776 43988 26816
rect 44812 26776 44852 26816
rect 45004 26776 45044 26816
rect 45292 26776 45332 26816
rect 45388 26776 45428 26816
rect 45580 26776 45620 26816
rect 45868 26776 45908 26816
rect 47884 26776 47924 26816
rect 48172 26776 48212 26816
rect 49708 26776 49748 26816
rect 50572 26776 50612 26816
rect 3820 26692 3860 26732
rect 5836 26692 5876 26732
rect 6316 26692 6356 26732
rect 6700 26692 6740 26732
rect 8044 26692 8084 26732
rect 11212 26692 11252 26732
rect 11788 26692 11828 26732
rect 15052 26692 15092 26732
rect 15532 26692 15572 26732
rect 17068 26692 17108 26732
rect 22924 26692 22964 26732
rect 28972 26692 29012 26732
rect 35692 26692 35732 26732
rect 49036 26692 49076 26732
rect 49324 26692 49364 26732
rect 3052 26608 3092 26648
rect 3532 26608 3572 26648
rect 7084 26608 7124 26648
rect 10060 26608 10100 26648
rect 13804 26608 13844 26648
rect 14380 26608 14420 26648
rect 16204 26608 16244 26648
rect 18028 26608 18068 26648
rect 18892 26608 18932 26648
rect 19180 26608 19220 26648
rect 24844 26608 24884 26648
rect 25516 26608 25556 26648
rect 25900 26608 25940 26648
rect 28684 26608 28724 26648
rect 29356 26608 29396 26648
rect 29932 26608 29972 26648
rect 30796 26608 30836 26648
rect 34828 26608 34868 26648
rect 35308 26608 35348 26648
rect 43852 26608 43892 26648
rect 44140 26608 44180 26648
rect 47212 26608 47252 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 30796 26330 30836 26370
rect 11212 26272 11252 26312
rect 11404 26272 11444 26312
rect 14764 26272 14804 26312
rect 21100 26272 21140 26312
rect 25996 26272 26036 26312
rect 29164 26272 29204 26312
rect 35500 26272 35540 26312
rect 36556 26272 36596 26312
rect 38380 26272 38420 26312
rect 39052 26272 39092 26312
rect 42796 26272 42836 26312
rect 47404 26272 47444 26312
rect 48940 26272 48980 26312
rect 51244 26272 51284 26312
rect 1708 26188 1748 26228
rect 8812 26188 8852 26228
rect 17644 26188 17684 26228
rect 20140 26188 20180 26228
rect 37324 26188 37364 26228
rect 37804 26188 37844 26228
rect 41932 26188 41972 26228
rect 44236 26188 44276 26228
rect 45004 26188 45044 26228
rect 2092 26104 2132 26144
rect 2956 26104 2996 26144
rect 4396 26104 4436 26144
rect 4684 26104 4724 26144
rect 5356 26104 5396 26144
rect 5836 26104 5876 26144
rect 6124 26104 6164 26144
rect 6220 26104 6260 26144
rect 6892 26104 6932 26144
rect 7756 26104 7796 26144
rect 7948 26104 7988 26144
rect 8044 26104 8084 26144
rect 9196 26104 9236 26144
rect 10060 26104 10100 26144
rect 12076 26104 12116 26144
rect 13612 26104 13652 26144
rect 13804 26104 13844 26144
rect 13900 26104 13940 26144
rect 14092 26104 14132 26144
rect 14188 26104 14228 26144
rect 14380 26104 14420 26144
rect 14572 26104 14612 26144
rect 14668 26104 14708 26144
rect 14860 26104 14900 26144
rect 15244 26104 15284 26144
rect 15340 26104 15380 26144
rect 15436 26104 15476 26144
rect 15724 26104 15764 26144
rect 15820 26104 15860 26144
rect 16012 26104 16052 26144
rect 16108 26104 16148 26144
rect 16209 26104 16249 26144
rect 16588 26104 16628 26144
rect 16684 26104 16724 26144
rect 16780 26104 16820 26144
rect 16876 26104 16916 26144
rect 17068 26104 17108 26144
rect 17164 26104 17204 26144
rect 17260 26104 17300 26144
rect 17356 26104 17396 26144
rect 17548 26104 17588 26144
rect 17740 26104 17780 26144
rect 17836 26104 17876 26144
rect 18700 26104 18740 26144
rect 19084 26104 19124 26144
rect 19372 26104 19412 26144
rect 19468 26104 19508 26144
rect 19948 26104 19988 26144
rect 20044 26104 20084 26144
rect 20236 26104 20276 26144
rect 20428 26104 20468 26144
rect 21964 26104 22004 26144
rect 22156 26104 22196 26144
rect 23596 26104 23636 26144
rect 23980 26104 24020 26144
rect 24844 26104 24884 26144
rect 26380 26104 26420 26144
rect 26476 26104 26516 26144
rect 26572 26104 26612 26144
rect 26668 26104 26708 26144
rect 26956 26104 26996 26144
rect 27916 26104 27956 26144
rect 28492 26104 28532 26144
rect 28588 26099 28628 26139
rect 28684 26104 28724 26144
rect 29068 26104 29108 26144
rect 29260 26104 29300 26144
rect 29356 26104 29396 26144
rect 29644 26104 29684 26144
rect 29836 26104 29876 26144
rect 29932 26104 29972 26144
rect 30604 26104 30644 26144
rect 30700 26104 30740 26144
rect 31372 26093 31412 26133
rect 31564 26104 31604 26144
rect 31660 26104 31700 26144
rect 31852 26104 31892 26144
rect 32812 26104 32852 26144
rect 33100 26104 33140 26144
rect 33964 26104 34004 26144
rect 35020 26104 35060 26144
rect 35212 26104 35252 26144
rect 35308 26104 35348 26144
rect 35404 26104 35444 26144
rect 36172 26104 36212 26144
rect 37036 26104 37076 26144
rect 37228 26104 37268 26144
rect 37420 26104 37460 26144
rect 37900 26104 37940 26144
rect 37996 26104 38036 26144
rect 38092 26104 38132 26144
rect 38284 26104 38324 26144
rect 38476 26104 38516 26144
rect 38572 26104 38612 26144
rect 38764 26104 38804 26144
rect 38860 26104 38900 26144
rect 38956 26104 38996 26144
rect 40492 26104 40532 26144
rect 40588 26104 40628 26144
rect 40780 26104 40820 26144
rect 41164 26104 41204 26144
rect 41260 26104 41300 26144
rect 41356 26104 41396 26144
rect 41452 26104 41492 26144
rect 42028 26104 42068 26144
rect 42316 26104 42356 26144
rect 42892 26104 42932 26144
rect 43084 26104 43124 26144
rect 43756 26104 43796 26144
rect 44332 26104 44372 26144
rect 44620 26104 44660 26144
rect 45388 26104 45428 26144
rect 46252 26104 46292 26144
rect 47788 26104 47828 26144
rect 47884 26090 47924 26130
rect 48076 26104 48116 26144
rect 48268 26104 48308 26144
rect 49132 26104 49172 26144
rect 50764 26104 50804 26144
rect 50956 26104 50996 26144
rect 51052 26104 51092 26144
rect 51148 26104 51188 26144
rect 4108 26020 4148 26060
rect 1516 25936 1556 25976
rect 6508 25936 6548 25976
rect 7756 25936 7796 25976
rect 8428 25936 8468 25976
rect 12460 25936 12500 25976
rect 19756 25936 19796 25976
rect 21484 25936 21524 25976
rect 31372 25936 31412 25976
rect 40300 25936 40340 25976
rect 41644 25936 41684 25976
rect 43948 25936 43988 25976
rect 48076 25936 48116 25976
rect 51436 25936 51476 25976
rect 4492 25852 4532 25892
rect 7564 25852 7604 25892
rect 13612 25852 13652 25892
rect 14380 25852 14420 25892
rect 15724 25852 15764 25892
rect 18028 25852 18068 25892
rect 22060 25852 22100 25892
rect 27244 25852 27284 25892
rect 28204 25852 28244 25892
rect 29644 25852 29684 25892
rect 30316 25852 30356 25892
rect 34348 25852 34388 25892
rect 40780 25852 40820 25892
rect 49804 25852 49844 25892
rect 50092 25852 50132 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 3436 25516 3476 25556
rect 6316 25516 6356 25556
rect 13708 25516 13748 25556
rect 15244 25516 15284 25556
rect 17836 25516 17876 25556
rect 20428 25516 20468 25556
rect 20620 25516 20660 25556
rect 27916 25516 27956 25556
rect 32044 25516 32084 25556
rect 36172 25516 36212 25556
rect 39340 25516 39380 25556
rect 42700 25516 42740 25556
rect 43756 25516 43796 25556
rect 11884 25432 11924 25472
rect 16396 25432 16436 25472
rect 22636 25432 22676 25472
rect 30508 25432 30548 25472
rect 45100 25432 45140 25472
rect 9292 25348 9332 25388
rect 12652 25348 12692 25388
rect 26860 25348 26900 25388
rect 1420 25264 1460 25304
rect 2284 25264 2324 25304
rect 4300 25264 4340 25304
rect 4588 25264 4628 25304
rect 5452 25264 5492 25304
rect 5932 25264 5972 25304
rect 6028 25264 6068 25304
rect 7852 25264 7892 25304
rect 8716 25264 8756 25304
rect 9100 25264 9140 25304
rect 9388 25264 9428 25304
rect 9676 25264 9716 25304
rect 9964 25264 10004 25304
rect 10060 25264 10100 25304
rect 10156 25264 10196 25304
rect 10540 25264 10580 25304
rect 10636 25264 10676 25304
rect 10732 25264 10772 25304
rect 10828 25264 10868 25304
rect 11020 25264 11060 25304
rect 11884 25264 11924 25304
rect 12076 25264 12116 25304
rect 12172 25264 12212 25304
rect 12556 25264 12596 25304
rect 12748 25287 12788 25327
rect 13223 25264 13263 25304
rect 13324 25264 13364 25304
rect 13420 25264 13460 25304
rect 13612 25264 13652 25304
rect 13708 25264 13748 25304
rect 13900 25264 13940 25304
rect 14956 25264 14996 25304
rect 15052 25264 15092 25304
rect 15244 25264 15284 25304
rect 16108 25264 16148 25304
rect 16204 25264 16244 25304
rect 16396 25264 16436 25304
rect 17548 25264 17588 25304
rect 17644 25264 17684 25304
rect 17836 25264 17876 25304
rect 18028 25264 18068 25304
rect 18412 25264 18452 25304
rect 19276 25264 19316 25304
rect 20716 25264 20756 25304
rect 20908 25264 20948 25304
rect 21580 25264 21620 25304
rect 22156 25264 22196 25304
rect 22252 25299 22292 25339
rect 37612 25348 37652 25388
rect 37708 25348 37748 25388
rect 46924 25348 46964 25388
rect 47020 25348 47060 25388
rect 49420 25348 49460 25388
rect 22348 25264 22388 25304
rect 22732 25264 22772 25304
rect 23500 25264 23540 25304
rect 23596 25269 23636 25309
rect 23692 25264 23732 25304
rect 24652 25264 24692 25304
rect 24844 25264 24884 25304
rect 24940 25264 24980 25304
rect 26476 25264 26516 25304
rect 26572 25299 26612 25339
rect 26668 25264 26708 25304
rect 27244 25264 27284 25304
rect 28204 25264 28244 25304
rect 28876 25264 28916 25304
rect 29836 25264 29876 25304
rect 30316 25264 30356 25304
rect 32620 25264 32660 25304
rect 33004 25264 33044 25304
rect 33388 25264 33428 25304
rect 34252 25264 34292 25304
rect 35596 25264 35636 25304
rect 35692 25264 35732 25304
rect 35788 25264 35828 25304
rect 35884 25264 35924 25304
rect 36268 25264 36308 25304
rect 36652 25278 36692 25318
rect 37132 25264 37172 25304
rect 38092 25264 38132 25304
rect 38188 25264 38228 25304
rect 39148 25264 39188 25304
rect 40300 25264 40340 25304
rect 40684 25264 40724 25304
rect 41548 25264 41588 25304
rect 42892 25264 42932 25304
rect 43852 25264 43892 25304
rect 44524 25264 44564 25304
rect 44620 25264 44660 25304
rect 44716 25264 44756 25304
rect 44812 25264 44852 25304
rect 45580 25264 45620 25304
rect 45964 25278 46004 25318
rect 46444 25264 46484 25304
rect 47404 25264 47444 25304
rect 47500 25264 47540 25304
rect 47788 25264 47828 25304
rect 47884 25264 47924 25304
rect 48076 25264 48116 25304
rect 48172 25264 48212 25304
rect 48268 25264 48308 25304
rect 48556 25264 48596 25304
rect 50572 25264 50612 25304
rect 51436 25264 51476 25304
rect 51820 25264 51860 25304
rect 1036 25180 1076 25220
rect 3628 25180 3668 25220
rect 24748 25180 24788 25220
rect 26188 25180 26228 25220
rect 36460 25180 36500 25220
rect 43564 25180 43604 25220
rect 45772 25180 45812 25220
rect 6700 25096 6740 25136
rect 9580 25096 9620 25136
rect 9868 25096 9908 25136
rect 11692 25096 11732 25136
rect 14572 25096 14612 25136
rect 21868 25096 21908 25136
rect 23212 25096 23252 25136
rect 35404 25096 35444 25136
rect 45484 25096 45524 25136
rect 48364 25096 48404 25136
rect 49228 25096 49268 25136
rect 5836 25038 5876 25078
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 844 24760 884 24800
rect 1996 24760 2036 24800
rect 4204 24760 4244 24800
rect 6700 24760 6740 24800
rect 9676 24760 9716 24800
rect 10828 24760 10868 24800
rect 17068 24760 17108 24800
rect 24076 24760 24116 24800
rect 25324 24760 25364 24800
rect 26380 24760 26420 24800
rect 27052 24760 27092 24800
rect 31276 24760 31316 24800
rect 35404 24760 35444 24800
rect 41644 24760 41684 24800
rect 41932 24760 41972 24800
rect 46252 24760 46292 24800
rect 47020 24760 47060 24800
rect 48652 24760 48692 24800
rect 49036 24760 49076 24800
rect 4396 24676 4436 24716
rect 6124 24676 6164 24716
rect 10348 24676 10388 24716
rect 13228 24676 13268 24716
rect 27436 24676 27476 24716
rect 33004 24676 33044 24716
rect 38860 24676 38900 24716
rect 44332 24676 44372 24716
rect 49324 24676 49364 24716
rect 940 24592 980 24632
rect 1900 24592 1940 24632
rect 2092 24592 2132 24632
rect 2188 24592 2228 24632
rect 2380 24592 2420 24632
rect 2476 24592 2516 24632
rect 2572 24592 2612 24632
rect 2668 24592 2708 24632
rect 3532 24592 3572 24632
rect 3916 24592 3956 24632
rect 4012 24592 4052 24632
rect 4108 24592 4148 24632
rect 5068 24592 5108 24632
rect 5452 24592 5492 24632
rect 5548 24592 5588 24632
rect 5644 24592 5684 24632
rect 5740 24592 5780 24632
rect 5932 24592 5972 24632
rect 6028 24592 6068 24632
rect 6220 24592 6260 24632
rect 6412 24592 6452 24632
rect 6508 24592 6548 24632
rect 6604 24592 6644 24632
rect 7564 24592 7604 24632
rect 7756 24592 7796 24632
rect 7948 24592 7988 24632
rect 8620 24592 8660 24632
rect 8812 24592 8852 24632
rect 9004 24592 9044 24632
rect 9964 24592 10004 24632
rect 10252 24592 10292 24632
rect 11980 24592 12020 24632
rect 12844 24592 12884 24632
rect 13516 24592 13556 24632
rect 13804 24592 13844 24632
rect 13900 24592 13940 24632
rect 14476 24592 14516 24632
rect 15436 24592 15476 24632
rect 15532 24592 15572 24632
rect 15724 24592 15764 24632
rect 15916 24592 15956 24632
rect 16012 24592 16052 24632
rect 16108 24592 16148 24632
rect 16204 24592 16244 24632
rect 16972 24592 17012 24632
rect 17260 24592 17300 24632
rect 17932 24592 17972 24632
rect 18124 24592 18164 24632
rect 18220 24592 18260 24632
rect 18316 24592 18356 24632
rect 18412 24592 18452 24632
rect 18700 24592 18740 24632
rect 20908 24592 20948 24632
rect 21004 24592 21044 24632
rect 21100 24592 21140 24632
rect 21196 24592 21236 24632
rect 21772 24592 21812 24632
rect 21868 24587 21908 24627
rect 21964 24592 22004 24632
rect 22252 24592 22292 24632
rect 24556 24592 24596 24632
rect 25708 24592 25748 24632
rect 26092 24592 26132 24632
rect 26188 24592 26228 24632
rect 26476 24592 26516 24632
rect 26956 24592 26996 24632
rect 27148 24592 27188 24632
rect 27244 24592 27284 24632
rect 28108 24592 28148 24632
rect 29260 24592 29300 24632
rect 29644 24592 29684 24632
rect 29836 24592 29876 24632
rect 30028 24592 30068 24632
rect 30124 24605 30164 24645
rect 30316 24592 30356 24632
rect 30796 24592 30836 24632
rect 31660 24592 31700 24632
rect 32140 24592 32180 24632
rect 32908 24592 32948 24632
rect 33100 24592 33140 24632
rect 33292 24592 33332 24632
rect 33964 24592 34004 24632
rect 34252 24592 34292 24632
rect 35212 24592 35252 24632
rect 36076 24592 36116 24632
rect 37708 24592 37748 24632
rect 38572 24592 38612 24632
rect 39052 24587 39092 24627
rect 39532 24592 39572 24632
rect 40108 24592 40148 24632
rect 40492 24592 40532 24632
rect 40588 24592 40628 24632
rect 40972 24592 41012 24632
rect 41068 24592 41108 24632
rect 41164 24592 41204 24632
rect 41260 24592 41300 24632
rect 41452 24592 41492 24632
rect 41548 24592 41588 24632
rect 41740 24592 41780 24632
rect 43084 24592 43124 24632
rect 43948 24592 43988 24632
rect 44716 24592 44756 24632
rect 45676 24592 45716 24632
rect 46348 24592 46388 24632
rect 46444 24592 46484 24632
rect 46540 24592 46580 24632
rect 46732 24592 46772 24632
rect 46828 24592 46868 24632
rect 46924 24592 46964 24632
rect 47212 24592 47252 24632
rect 47308 24592 47348 24632
rect 47500 24592 47540 24632
rect 47692 24592 47732 24632
rect 48556 24592 48596 24632
rect 48748 24592 48788 24632
rect 48844 24592 48884 24632
rect 49132 24592 49172 24632
rect 49708 24592 49748 24632
rect 50572 24592 50612 24632
rect 7852 24508 7892 24548
rect 23116 24508 23156 24548
rect 40012 24508 40052 24548
rect 1324 24424 1364 24464
rect 1708 24424 1748 24464
rect 8140 24424 8180 24464
rect 8716 24424 8756 24464
rect 10636 24424 10676 24464
rect 14188 24424 14228 24464
rect 14764 24424 14804 24464
rect 15724 24424 15764 24464
rect 18892 24424 18932 24464
rect 19276 24424 19316 24464
rect 30316 24424 30356 24464
rect 32716 24424 32756 24464
rect 47500 24424 47540 24464
rect 2860 24340 2900 24380
rect 6892 24340 6932 24380
rect 14380 24340 14420 24380
rect 18604 24340 18644 24380
rect 21484 24340 21524 24380
rect 28588 24340 28628 24380
rect 29740 24340 29780 24380
rect 32044 24340 32084 24380
rect 35404 24340 35444 24380
rect 48364 24340 48404 24380
rect 51724 24340 51764 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 17740 24004 17780 24044
rect 40012 24004 40052 24044
rect 40780 24004 40820 24044
rect 46252 24004 46292 24044
rect 46732 24004 46772 24044
rect 4012 23920 4052 23960
rect 6124 23920 6164 23960
rect 9292 23920 9332 23960
rect 9676 23920 9716 23960
rect 14092 23920 14132 23960
rect 16684 23920 16724 23960
rect 21388 23920 21428 23960
rect 25132 23920 25172 23960
rect 26764 23920 26804 23960
rect 30796 23920 30836 23960
rect 31276 23920 31316 23960
rect 40492 23920 40532 23960
rect 43660 23920 43700 23960
rect 44908 23920 44948 23960
rect 49612 23920 49652 23960
rect 50860 23920 50900 23960
rect 3532 23836 3572 23876
rect 10444 23836 10484 23876
rect 23788 23836 23828 23876
rect 33004 23836 33044 23876
rect 1516 23752 1556 23792
rect 2380 23752 2420 23792
rect 3724 23752 3764 23792
rect 3820 23752 3860 23792
rect 4012 23752 4052 23792
rect 4204 23752 4244 23792
rect 4300 23752 4340 23792
rect 4588 23752 4628 23792
rect 4780 23752 4820 23792
rect 4876 23752 4916 23792
rect 5164 23752 5204 23792
rect 5260 23752 5300 23792
rect 5356 23752 5396 23792
rect 5452 23752 5492 23792
rect 6604 23752 6644 23792
rect 6892 23752 6932 23792
rect 7276 23752 7316 23792
rect 8140 23752 8180 23792
rect 9964 23752 10004 23792
rect 10060 23752 10100 23792
rect 10156 23752 10196 23792
rect 11212 23752 11252 23792
rect 12748 23752 12788 23792
rect 13804 23752 13844 23792
rect 13900 23752 13940 23792
rect 14092 23752 14132 23792
rect 14284 23752 14324 23792
rect 14668 23752 14708 23792
rect 15532 23752 15572 23792
rect 16972 23752 17012 23792
rect 17068 23752 17108 23792
rect 17452 23752 17492 23792
rect 17548 23752 17588 23792
rect 17740 23763 17780 23803
rect 17932 23752 17972 23792
rect 19468 23752 19508 23792
rect 20716 23752 20756 23792
rect 21580 23752 21620 23792
rect 23020 23752 23060 23792
rect 24364 23752 24404 23792
rect 24460 23752 24500 23792
rect 24652 23752 24692 23792
rect 25612 23752 25652 23792
rect 25900 23752 25940 23792
rect 26572 23752 26612 23792
rect 28204 23752 28244 23792
rect 29452 23752 29492 23792
rect 29740 23752 29780 23792
rect 30412 23752 30452 23792
rect 30988 23752 31028 23792
rect 31084 23752 31124 23792
rect 31276 23752 31316 23792
rect 32140 23752 32180 23792
rect 32332 23752 32372 23792
rect 32428 23752 32468 23792
rect 32524 23752 32564 23792
rect 32620 23752 32660 23792
rect 33388 23752 33428 23792
rect 33484 23752 33524 23792
rect 33580 23752 33620 23792
rect 33676 23752 33716 23792
rect 33868 23752 33908 23792
rect 33964 23752 34004 23792
rect 34060 23752 34100 23792
rect 34156 23752 34196 23792
rect 34348 23752 34388 23792
rect 34444 23752 34484 23792
rect 36700 23794 36740 23834
rect 37804 23836 37844 23876
rect 46540 23836 46580 23876
rect 47884 23836 47924 23876
rect 34636 23752 34676 23792
rect 35500 23752 35540 23792
rect 36364 23752 36404 23792
rect 37228 23752 37268 23792
rect 37708 23752 37748 23792
rect 38188 23752 38228 23792
rect 38284 23752 38324 23792
rect 39244 23752 39284 23792
rect 40108 23752 40148 23792
rect 40876 23752 40916 23792
rect 41740 23752 41780 23792
rect 41932 23752 41972 23792
rect 42028 23752 42068 23792
rect 42124 23752 42164 23792
rect 43276 23752 43316 23792
rect 45772 23752 45812 23792
rect 45868 23752 45908 23792
rect 45964 23752 46004 23792
rect 46156 23752 46196 23792
rect 46348 23752 46388 23792
rect 47596 23752 47636 23792
rect 48748 23752 48788 23792
rect 49132 23752 49172 23792
rect 49804 23752 49844 23792
rect 50476 23752 50516 23792
rect 1132 23668 1172 23708
rect 4684 23668 4724 23708
rect 11980 23668 12020 23708
rect 27340 23668 27380 23708
rect 34540 23668 34580 23708
rect 36556 23668 36596 23708
rect 42604 23668 42644 23708
rect 9868 23584 9908 23624
rect 17260 23584 17300 23624
rect 18604 23584 18644 23624
rect 18796 23584 18836 23624
rect 23404 23584 23444 23624
rect 24172 23584 24212 23624
rect 28972 23584 29012 23624
rect 31468 23584 31508 23624
rect 33196 23584 33236 23624
rect 34828 23584 34868 23624
rect 35692 23584 35732 23624
rect 38572 23584 38612 23624
rect 41068 23584 41108 23624
rect 42220 23584 42260 23624
rect 45676 23584 45716 23624
rect 46924 23584 46964 23624
rect 49036 23584 49076 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3820 23248 3860 23288
rect 5644 23248 5684 23288
rect 5932 23248 5972 23288
rect 18028 23248 18068 23288
rect 20812 23248 20852 23288
rect 22156 23248 22196 23288
rect 33484 23248 33524 23288
rect 33676 23248 33716 23288
rect 37324 23248 37364 23288
rect 38668 23248 38708 23288
rect 39532 23248 39572 23288
rect 43372 23248 43412 23288
rect 46828 23248 46868 23288
rect 50188 23248 50228 23288
rect 1420 23164 1460 23204
rect 12844 23164 12884 23204
rect 16492 23164 16532 23204
rect 18412 23164 18452 23204
rect 28876 23164 28916 23204
rect 31084 23164 31124 23204
rect 34924 23164 34964 23204
rect 40684 23164 40724 23204
rect 47788 23164 47828 23204
rect 1804 23080 1844 23120
rect 2668 23080 2708 23120
rect 4108 23080 4148 23120
rect 4972 23080 5012 23120
rect 5836 23080 5876 23120
rect 6124 23080 6164 23120
rect 7180 23080 7220 23120
rect 8044 23080 8084 23120
rect 8716 23080 8756 23120
rect 8812 23080 8852 23120
rect 9004 23080 9044 23120
rect 9868 23080 9908 23120
rect 10732 23080 10772 23120
rect 11596 23080 11636 23120
rect 11884 23080 11924 23120
rect 13708 23080 13748 23120
rect 14476 23080 14516 23120
rect 15148 23080 15188 23120
rect 15436 23080 15476 23120
rect 15532 23080 15572 23120
rect 15628 23080 15668 23120
rect 15724 23080 15764 23120
rect 16396 23080 16436 23120
rect 16588 23080 16628 23120
rect 16780 23080 16820 23120
rect 16876 23080 16916 23120
rect 17068 23080 17108 23120
rect 17452 23080 17492 23120
rect 17548 23101 17588 23141
rect 17644 23080 17684 23120
rect 17740 23080 17780 23120
rect 17932 23080 17972 23120
rect 18124 23080 18164 23120
rect 18220 23080 18260 23120
rect 18796 23080 18836 23120
rect 19660 23080 19700 23120
rect 22540 23080 22580 23120
rect 22924 23080 22964 23120
rect 23308 23080 23348 23120
rect 24172 23080 24212 23120
rect 25420 23080 25460 23120
rect 25804 23080 25844 23120
rect 26188 23080 26228 23120
rect 27052 23080 27092 23120
rect 28204 23080 28244 23120
rect 29644 23080 29684 23120
rect 30316 23080 30356 23120
rect 30412 23080 30452 23120
rect 30700 23080 30740 23120
rect 31468 23080 31508 23120
rect 32332 23080 32372 23120
rect 34348 23080 34388 23120
rect 35308 23080 35348 23120
rect 36172 23080 36212 23120
rect 38572 23080 38612 23120
rect 38956 23080 38996 23120
rect 39052 23080 39092 23120
rect 39148 23080 39188 23120
rect 39244 23080 39284 23120
rect 39436 23080 39476 23120
rect 39724 23080 39764 23120
rect 40396 23080 40436 23120
rect 41068 23080 41108 23120
rect 41932 23080 41972 23120
rect 43468 23080 43508 23120
rect 43564 23080 43604 23120
rect 43660 23080 43700 23120
rect 43948 23080 43988 23120
rect 44236 23080 44276 23120
rect 44428 23080 44468 23120
rect 44812 23080 44852 23120
rect 45676 23080 45716 23120
rect 47212 23080 47252 23120
rect 47308 23080 47348 23120
rect 47404 23080 47444 23120
rect 47500 23080 47540 23120
rect 48172 23080 48212 23120
rect 49036 23080 49076 23120
rect 652 22996 692 23036
rect 16108 22996 16148 23036
rect 9004 22912 9044 22952
rect 14284 22912 14324 22952
rect 15916 22912 15956 22952
rect 30028 22912 30068 22952
rect 34732 22912 34772 22952
rect 37804 22912 37844 22952
rect 43084 22912 43124 22952
rect 844 22828 884 22868
rect 4780 22828 4820 22868
rect 5644 22828 5684 22868
rect 6508 22828 6548 22868
rect 7372 22828 7412 22868
rect 9196 22828 9236 22868
rect 10060 22828 10100 22868
rect 10924 22828 10964 22868
rect 12556 22828 12596 22868
rect 17068 22828 17108 22868
rect 43852 22828 43892 22868
rect 44140 22828 44180 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4108 22492 4148 22532
rect 6412 22492 6452 22532
rect 8524 22492 8564 22532
rect 11980 22492 12020 22532
rect 14188 22492 14228 22532
rect 14860 22492 14900 22532
rect 16300 22492 16340 22532
rect 22348 22492 22388 22532
rect 29164 22492 29204 22532
rect 34252 22492 34292 22532
rect 39724 22492 39764 22532
rect 41452 22492 41492 22532
rect 43084 22492 43124 22532
rect 48364 22492 48404 22532
rect 1516 22408 1556 22448
rect 5932 22408 5972 22448
rect 12940 22408 12980 22448
rect 19756 22408 19796 22448
rect 23404 22408 23444 22448
rect 27244 22408 27284 22448
rect 47596 22408 47636 22448
rect 51628 22408 51668 22448
rect 34444 22324 34484 22364
rect 40396 22324 40436 22364
rect 2092 22240 2132 22280
rect 2956 22240 2996 22280
rect 4300 22240 4340 22280
rect 4396 22240 4436 22280
rect 4492 22240 4532 22280
rect 4588 22240 4628 22280
rect 4780 22240 4820 22280
rect 4972 22240 5012 22280
rect 5068 22240 5108 22280
rect 5548 22240 5588 22280
rect 6124 22240 6164 22280
rect 6220 22240 6260 22280
rect 6412 22240 6452 22280
rect 7276 22240 7316 22280
rect 7468 22240 7508 22280
rect 7564 22240 7604 22280
rect 7852 22240 7892 22280
rect 8140 22240 8180 22280
rect 9292 22240 9332 22280
rect 9580 22240 9620 22280
rect 9964 22240 10004 22280
rect 10828 22240 10868 22280
rect 12268 22240 12308 22280
rect 12556 22240 12596 22280
rect 12652 22240 12692 22280
rect 13516 22240 13556 22280
rect 13804 22240 13844 22280
rect 14572 22240 14612 22280
rect 14668 22240 14708 22280
rect 14860 22240 14900 22280
rect 15148 22240 15188 22280
rect 16108 22240 16148 22280
rect 16396 22240 16436 22280
rect 16588 22240 16628 22280
rect 17260 22240 17300 22280
rect 17452 22240 17492 22280
rect 17548 22240 17588 22280
rect 17644 22240 17684 22280
rect 17740 22240 17780 22280
rect 18220 22240 18260 22280
rect 20332 22240 20372 22280
rect 21196 22240 21236 22280
rect 23212 22240 23252 22280
rect 24364 22240 24404 22280
rect 30316 22240 30356 22280
rect 31180 22240 31220 22280
rect 32428 22240 32468 22280
rect 32620 22240 32660 22280
rect 32812 22240 32852 22280
rect 32908 22240 32948 22280
rect 33772 22240 33812 22280
rect 34156 22240 34196 22280
rect 34540 22240 34580 22280
rect 34828 22240 34868 22280
rect 35692 22240 35732 22280
rect 37708 22240 37748 22280
rect 38572 22240 38612 22280
rect 40204 22240 40244 22280
rect 40780 22240 40820 22280
rect 40876 22240 40916 22280
rect 40972 22240 41012 22280
rect 41164 22240 41204 22280
rect 41260 22240 41300 22280
rect 41452 22240 41492 22280
rect 41644 22240 41684 22280
rect 41740 22240 41780 22280
rect 41836 22240 41876 22280
rect 41932 22240 41972 22280
rect 42796 22240 42836 22280
rect 42988 22240 43028 22280
rect 43180 22240 43220 22280
rect 43372 22240 43412 22280
rect 43468 22240 43508 22280
rect 43660 22240 43700 22280
rect 43852 22240 43892 22280
rect 43948 22240 43988 22280
rect 44044 22240 44084 22280
rect 44140 22240 44180 22280
rect 44332 22240 44372 22280
rect 44428 22240 44468 22280
rect 44524 22240 44564 22280
rect 44812 22240 44852 22280
rect 45004 22240 45044 22280
rect 45388 22240 45428 22280
rect 45580 22240 45620 22280
rect 45772 22240 45812 22280
rect 45868 22240 45908 22280
rect 46060 22240 46100 22280
rect 46156 22240 46196 22280
rect 46252 22240 46292 22280
rect 46348 22240 46388 22280
rect 47212 22240 47252 22280
rect 47788 22240 47828 22280
rect 47884 22240 47924 22280
rect 48076 22240 48116 22280
rect 49036 22240 49076 22280
rect 49612 22240 49652 22280
rect 50476 22240 50516 22280
rect 1708 22156 1748 22196
rect 4876 22156 4916 22196
rect 8236 22156 8276 22196
rect 13900 22156 13940 22196
rect 19948 22156 19988 22196
rect 31564 22156 31604 22196
rect 31756 22156 31796 22196
rect 32716 22156 32756 22196
rect 37324 22156 37364 22196
rect 40108 22156 40148 22196
rect 45676 22156 45716 22196
rect 46540 22156 46580 22196
rect 47980 22156 48020 22196
rect 49228 22156 49268 22196
rect 652 22072 692 22112
rect 5452 22072 5492 22112
rect 6604 22072 6644 22112
rect 9388 22072 9428 22112
rect 18700 22072 18740 22112
rect 22540 22072 22580 22112
rect 24172 22072 24212 22112
rect 24460 22072 24500 22112
rect 33100 22072 33140 22112
rect 42124 22072 42164 22112
rect 43564 22072 43604 22112
rect 44620 22072 44660 22112
rect 45292 22072 45332 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4492 21736 4532 21776
rect 5548 21736 5588 21776
rect 16396 21736 16436 21776
rect 18988 21736 19028 21776
rect 19468 21736 19508 21776
rect 22636 21736 22676 21776
rect 25900 21736 25940 21776
rect 26476 21736 26516 21776
rect 29164 21736 29204 21776
rect 32620 21736 32660 21776
rect 35212 21736 35252 21776
rect 39340 21736 39380 21776
rect 41260 21736 41300 21776
rect 42604 21736 42644 21776
rect 45196 21736 45236 21776
rect 46156 21736 46196 21776
rect 6124 21652 6164 21692
rect 13996 21652 14036 21692
rect 16588 21652 16628 21692
rect 26764 21652 26804 21692
rect 32812 21652 32852 21692
rect 38380 21652 38420 21692
rect 47596 21652 47636 21692
rect 2092 21568 2132 21608
rect 2476 21568 2516 21608
rect 3340 21568 3380 21608
rect 4876 21568 4916 21608
rect 5068 21568 5108 21608
rect 5260 21568 5300 21608
rect 5356 21568 5396 21608
rect 5644 21568 5684 21608
rect 5740 21568 5780 21608
rect 5836 21568 5876 21608
rect 6508 21568 6548 21608
rect 7372 21568 7412 21608
rect 9580 21568 9620 21608
rect 9676 21568 9716 21608
rect 9772 21568 9812 21608
rect 9868 21568 9908 21608
rect 10156 21568 10196 21608
rect 11308 21568 11348 21608
rect 11404 21568 11444 21608
rect 11500 21568 11540 21608
rect 11596 21568 11636 21608
rect 11788 21568 11828 21608
rect 13036 21568 13076 21608
rect 14380 21568 14420 21608
rect 15244 21568 15284 21608
rect 16972 21568 17012 21608
rect 17836 21568 17876 21608
rect 21004 21568 21044 21608
rect 21196 21568 21236 21608
rect 21292 21568 21332 21608
rect 21388 21568 21428 21608
rect 21484 21568 21524 21608
rect 22540 21568 22580 21608
rect 22732 21568 22772 21608
rect 22924 21568 22964 21608
rect 23596 21568 23636 21608
rect 23788 21568 23828 21608
rect 23980 21568 24020 21608
rect 24844 21568 24884 21608
rect 24940 21568 24980 21608
rect 25036 21568 25076 21608
rect 25132 21568 25172 21608
rect 25324 21568 25364 21608
rect 25420 21568 25460 21608
rect 25516 21568 25556 21608
rect 25612 21568 25652 21608
rect 25804 21568 25844 21608
rect 25996 21568 26036 21608
rect 26092 21568 26132 21608
rect 26380 21568 26420 21608
rect 26572 21568 26612 21608
rect 27148 21568 27188 21608
rect 28012 21568 28052 21608
rect 30988 21568 31028 21608
rect 31084 21568 31124 21608
rect 31276 21568 31316 21608
rect 31468 21568 31508 21608
rect 31564 21568 31604 21608
rect 31660 21568 31700 21608
rect 31756 21568 31796 21608
rect 32332 21568 32372 21608
rect 32428 21568 32468 21608
rect 32524 21568 32564 21608
rect 33196 21568 33236 21608
rect 34060 21568 34100 21608
rect 35596 21568 35636 21608
rect 37420 21568 37460 21608
rect 37900 21568 37940 21608
rect 37996 21568 38036 21608
rect 38092 21568 38132 21608
rect 38188 21568 38228 21608
rect 39052 21568 39092 21608
rect 39244 21568 39284 21608
rect 39436 21568 39476 21608
rect 39532 21568 39572 21608
rect 40300 21568 40340 21608
rect 40396 21568 40436 21608
rect 40492 21568 40532 21608
rect 40588 21568 40628 21608
rect 40780 21568 40820 21608
rect 40972 21568 41012 21608
rect 41068 21568 41108 21608
rect 41932 21568 41972 21608
rect 42124 21568 42164 21608
rect 43084 21568 43124 21608
rect 43372 21568 43412 21608
rect 44044 21568 44084 21608
rect 44236 21568 44276 21608
rect 44332 21568 44372 21608
rect 44524 21568 44564 21608
rect 45580 21568 45620 21608
rect 47020 21568 47060 21608
rect 47116 21568 47156 21608
rect 47212 21568 47252 21608
rect 47308 21568 47348 21608
rect 47500 21568 47540 21608
rect 47692 21568 47732 21608
rect 47788 21568 47828 21608
rect 47980 21568 48020 21608
rect 8524 21484 8564 21524
rect 20140 21509 20180 21549
rect 21868 21484 21908 21524
rect 23884 21484 23924 21524
rect 36460 21484 36500 21524
rect 46348 21484 46388 21524
rect 48652 21484 48692 21524
rect 1900 21400 1940 21440
rect 5068 21400 5108 21440
rect 12652 21400 12692 21440
rect 20332 21400 20372 21440
rect 21676 21400 21716 21440
rect 29836 21400 29876 21440
rect 31276 21400 31316 21440
rect 32140 21400 32180 21440
rect 36748 21400 36788 21440
rect 40108 21400 40148 21440
rect 44524 21400 44564 21440
rect 46732 21400 46772 21440
rect 49036 21400 49076 21440
rect 49708 21400 49748 21440
rect 4780 21316 4820 21356
rect 10444 21316 10484 21356
rect 12460 21316 12500 21356
rect 13132 21316 13172 21356
rect 40780 21316 40820 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4396 20980 4436 21020
rect 6028 20980 6068 21020
rect 14092 20980 14132 21020
rect 14668 20980 14708 21020
rect 15628 20980 15668 21020
rect 25516 20980 25556 21020
rect 32236 20980 32276 21020
rect 33100 20980 33140 21020
rect 42892 20980 42932 21020
rect 44236 20980 44276 21020
rect 10636 20896 10676 20936
rect 16492 20896 16532 20936
rect 17068 20896 17108 20936
rect 23596 20870 23636 20910
rect 23788 20896 23828 20936
rect 30028 20896 30068 20936
rect 6220 20812 6260 20852
rect 19948 20812 19988 20852
rect 30796 20812 30836 20852
rect 39340 20812 39380 20852
rect 4492 20728 4532 20768
rect 4684 20728 4724 20768
rect 4780 20728 4820 20768
rect 4876 20728 4916 20768
rect 4972 20728 5012 20768
rect 5548 20728 5588 20768
rect 5740 20728 5780 20768
rect 6412 20728 6452 20768
rect 6508 20728 6548 20768
rect 6604 20728 6644 20768
rect 6700 20728 6740 20768
rect 6892 20728 6932 20768
rect 7756 20728 7796 20768
rect 8812 20728 8852 20768
rect 8908 20728 8948 20768
rect 9100 20728 9140 20768
rect 9964 20728 10004 20768
rect 10348 20728 10388 20768
rect 10444 20728 10484 20768
rect 10636 20728 10676 20768
rect 10828 20728 10868 20768
rect 12076 20728 12116 20768
rect 12940 20728 12980 20768
rect 14572 20728 14612 20768
rect 15148 20728 15188 20768
rect 19852 20728 19892 20768
rect 20044 20728 20084 20768
rect 20524 20728 20564 20768
rect 20620 20728 20660 20768
rect 21388 20728 21428 20768
rect 21580 20742 21620 20782
rect 21680 20747 21720 20787
rect 21868 20728 21908 20768
rect 21964 20728 22004 20768
rect 22060 20728 22100 20768
rect 22540 20728 22580 20768
rect 22636 20728 22676 20768
rect 22732 20728 22772 20768
rect 22828 20728 22868 20768
rect 23020 20728 23060 20768
rect 23116 20728 23156 20768
rect 23212 20728 23252 20768
rect 23308 20728 23348 20768
rect 23596 20728 23636 20768
rect 24076 20728 24116 20768
rect 24172 20728 24212 20768
rect 24268 20728 24308 20768
rect 25036 20728 25076 20768
rect 25228 20728 25268 20768
rect 25324 20728 25364 20768
rect 25708 20728 25748 20768
rect 26092 20728 26132 20768
rect 26476 20728 26516 20768
rect 27436 20728 27476 20768
rect 31660 20728 31700 20768
rect 32332 20728 32372 20768
rect 32716 20728 32756 20768
rect 35596 20728 35636 20768
rect 35980 20728 36020 20768
rect 36844 20728 36884 20768
rect 38380 20742 38420 20782
rect 38860 20728 38900 20768
rect 39436 20728 39476 20768
rect 39820 20728 39860 20768
rect 39916 20728 39956 20768
rect 40492 20728 40532 20768
rect 40876 20728 40916 20768
rect 41740 20728 41780 20768
rect 43084 20728 43124 20768
rect 44044 20728 44084 20768
rect 44908 20728 44948 20768
rect 45388 20728 45428 20768
rect 46348 20728 46388 20768
rect 46540 20728 46580 20768
rect 49036 20728 49076 20768
rect 49900 20728 49940 20768
rect 50284 20728 50324 20768
rect 9004 20644 9044 20684
rect 11500 20644 11540 20684
rect 11692 20644 11732 20684
rect 26188 20644 26228 20684
rect 652 20560 692 20600
rect 5644 20560 5684 20600
rect 6028 20560 6068 20600
rect 9292 20560 9332 20600
rect 20812 20560 20852 20600
rect 21484 20560 21524 20600
rect 22156 20560 22196 20600
rect 23980 20560 24020 20600
rect 37996 20560 38036 20600
rect 38188 20560 38228 20600
rect 43756 20560 43796 20600
rect 43948 20560 43988 20600
rect 47212 20560 47252 20600
rect 47884 20560 47924 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 652 20224 692 20264
rect 4108 20224 4148 20264
rect 8044 20224 8084 20264
rect 14092 20224 14132 20264
rect 18988 20224 19028 20264
rect 25036 20224 25076 20264
rect 29068 20224 29108 20264
rect 41932 20224 41972 20264
rect 45196 20224 45236 20264
rect 8812 20140 8852 20180
rect 24460 20140 24500 20180
rect 24748 20140 24788 20180
rect 25516 20140 25556 20180
rect 27820 20140 27860 20180
rect 37804 20140 37844 20180
rect 38380 20140 38420 20180
rect 39244 20140 39284 20180
rect 44620 20140 44660 20180
rect 47596 20140 47636 20180
rect 4012 20056 4052 20096
rect 4876 20056 4916 20096
rect 5068 20056 5108 20096
rect 5644 20056 5684 20096
rect 6028 20056 6068 20096
rect 6892 20056 6932 20096
rect 8524 20056 8564 20096
rect 9196 20056 9236 20096
rect 10060 20056 10100 20096
rect 11404 20056 11444 20096
rect 11596 20056 11636 20096
rect 11692 20056 11732 20096
rect 12556 20056 12596 20096
rect 13132 20056 13172 20096
rect 13420 20056 13460 20096
rect 14284 20056 14324 20096
rect 15244 20056 15284 20096
rect 15628 20056 15668 20096
rect 17164 20056 17204 20096
rect 17260 20056 17300 20096
rect 17452 20056 17492 20096
rect 18316 20056 18356 20096
rect 19180 20056 19220 20096
rect 19276 20056 19316 20096
rect 19468 20056 19508 20096
rect 20332 20056 20372 20096
rect 21196 20056 21236 20096
rect 21292 20056 21332 20096
rect 21772 20056 21812 20096
rect 21964 20056 22004 20096
rect 22060 20056 22100 20096
rect 22540 20056 22580 20096
rect 22636 20056 22676 20096
rect 23308 20056 23348 20096
rect 23404 20056 23444 20096
rect 23884 20077 23924 20117
rect 24076 20056 24116 20096
rect 24268 20056 24308 20096
rect 24364 20056 24404 20096
rect 24556 20056 24596 20096
rect 24940 20056 24980 20096
rect 25036 20056 25076 20096
rect 25612 20056 25652 20096
rect 25996 20056 26036 20096
rect 26572 20056 26612 20096
rect 27532 20056 27572 20096
rect 28588 20056 28628 20096
rect 29164 20056 29204 20096
rect 29548 20056 29588 20096
rect 29932 20056 29972 20096
rect 30796 20056 30836 20096
rect 32044 20056 32084 20096
rect 36652 20056 36692 20096
rect 37516 20056 37556 20096
rect 37900 20056 37940 20096
rect 37996 20056 38036 20096
rect 38092 20056 38132 20096
rect 38284 20056 38324 20096
rect 38476 20056 38516 20096
rect 38572 20056 38612 20096
rect 38764 20056 38804 20096
rect 38956 20056 38996 20096
rect 39340 20056 39380 20096
rect 39628 20056 39668 20096
rect 40396 20056 40436 20096
rect 41260 20056 41300 20096
rect 41740 20056 41780 20096
rect 41836 20056 41876 20096
rect 42028 20056 42068 20096
rect 43372 20056 43412 20096
rect 44236 20056 44276 20096
rect 46348 20056 46388 20096
rect 47212 20056 47252 20096
rect 11212 19972 11252 20012
rect 13228 19972 13268 20012
rect 18796 19972 18836 20012
rect 19660 19972 19700 20012
rect 21004 19972 21044 20012
rect 22924 19972 22964 20012
rect 23692 19972 23732 20012
rect 36556 19972 36596 20012
rect 38860 19972 38900 20012
rect 42220 19972 42260 20012
rect 2380 19888 2420 19928
rect 5452 19888 5492 19928
rect 12748 19888 12788 19928
rect 16972 19888 17012 19928
rect 33004 19888 33044 19928
rect 33772 19888 33812 19928
rect 36076 19888 36116 19928
rect 3820 19804 3860 19844
rect 4876 19804 4916 19844
rect 8428 19804 8468 19844
rect 11404 19804 11444 19844
rect 11884 19804 11924 19844
rect 16300 19804 16340 19844
rect 17452 19804 17492 19844
rect 17644 19804 17684 19844
rect 19468 19804 19508 19844
rect 21772 19804 21812 19844
rect 23980 19804 24020 19844
rect 26860 19804 26900 19844
rect 28204 19804 28244 19844
rect 29356 19804 29396 19844
rect 36844 19804 36884 19844
rect 39532 19804 39572 19844
rect 40684 19804 40724 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 6508 19468 6548 19508
rect 14284 19468 14324 19508
rect 20908 19468 20948 19508
rect 25708 19468 25748 19508
rect 27148 19468 27188 19508
rect 30316 19468 30356 19508
rect 38188 19468 38228 19508
rect 43180 19468 43220 19508
rect 8524 19384 8564 19424
rect 9292 19384 9332 19424
rect 21484 19384 21524 19424
rect 32332 19384 32372 19424
rect 35212 19384 35252 19424
rect 39148 19384 39188 19424
rect 42892 19384 42932 19424
rect 45100 19384 45140 19424
rect 4300 19300 4340 19340
rect 8716 19300 8756 19340
rect 2284 19216 2324 19256
rect 3148 19216 3188 19256
rect 4684 19216 4724 19256
rect 5548 19216 5588 19256
rect 5740 19216 5780 19256
rect 5836 19216 5876 19256
rect 6028 19216 6068 19256
rect 6124 19216 6164 19256
rect 6220 19216 6260 19256
rect 6316 19216 6356 19256
rect 6508 19216 6548 19256
rect 6700 19216 6740 19256
rect 6796 19216 6836 19256
rect 6988 19216 7028 19256
rect 7180 19216 7220 19256
rect 7852 19216 7892 19256
rect 8044 19216 8084 19256
rect 10636 19216 10676 19256
rect 11020 19216 11060 19256
rect 11116 19216 11156 19256
rect 11212 19216 11252 19256
rect 11308 19216 11348 19256
rect 11884 19216 11924 19256
rect 12268 19216 12308 19256
rect 13132 19216 13172 19256
rect 14860 19216 14900 19256
rect 16108 19216 16148 19256
rect 17356 19216 17396 19256
rect 18220 19216 18260 19256
rect 19660 19216 19700 19256
rect 20812 19216 20852 19256
rect 21004 19216 21044 19256
rect 22156 19216 22196 19256
rect 22444 19216 22484 19256
rect 22636 19216 22676 19256
rect 22732 19216 22772 19256
rect 23212 19216 23252 19256
rect 23308 19216 23348 19256
rect 23404 19216 23444 19256
rect 23500 19216 23540 19256
rect 23692 19216 23732 19256
rect 23788 19216 23828 19256
rect 23884 19216 23924 19256
rect 23980 19216 24020 19256
rect 25228 19216 25268 19256
rect 25324 19216 25364 19256
rect 25420 19216 25460 19256
rect 25708 19216 25748 19256
rect 25900 19216 25940 19256
rect 25996 19216 26036 19256
rect 26956 19216 26996 19256
rect 28300 19216 28340 19256
rect 28588 19216 28628 19256
rect 28780 19216 28820 19256
rect 29164 19216 29204 19256
rect 29740 19216 29780 19256
rect 29836 19216 29876 19256
rect 30316 19216 30356 19256
rect 30508 19216 30548 19256
rect 32140 19216 32180 19256
rect 32332 19216 32372 19256
rect 32524 19216 32564 19256
rect 32908 19216 32948 19256
rect 33772 19216 33812 19256
rect 34924 19216 34964 19256
rect 35596 19216 35636 19256
rect 36556 19216 36596 19256
rect 36844 19216 36884 19256
rect 37804 19216 37844 19256
rect 38188 19216 38228 19256
rect 38380 19216 38420 19256
rect 38476 19216 38516 19256
rect 38764 19216 38804 19256
rect 38860 19216 38900 19256
rect 38956 19216 38996 19256
rect 39628 19216 39668 19256
rect 39916 19216 39956 19256
rect 40012 19216 40052 19256
rect 40108 19216 40148 19256
rect 41068 19216 41108 19256
rect 42220 19216 42260 19256
rect 42316 19216 42356 19256
rect 42412 19216 42452 19256
rect 42508 19216 42548 19256
rect 43852 19216 43892 19256
rect 44044 19216 44084 19256
rect 1900 19132 1940 19172
rect 7084 19132 7124 19172
rect 16972 19132 17012 19172
rect 20524 19132 20564 19172
rect 40396 19132 40436 19172
rect 652 19048 692 19088
rect 5356 19048 5396 19088
rect 5644 19048 5684 19088
rect 7948 19048 7988 19088
rect 9964 19048 10004 19088
rect 15244 19048 15284 19088
rect 16780 19048 16820 19088
rect 19372 19048 19412 19088
rect 22444 19048 22484 19088
rect 25516 19048 25556 19088
rect 27340 19048 27380 19088
rect 28108 19048 28148 19088
rect 29260 19048 29300 19088
rect 30124 19048 30164 19088
rect 38668 19048 38708 19088
rect 39724 19048 39764 19088
rect 40204 19048 40244 19088
rect 44716 19048 44756 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 652 18712 692 18752
rect 2860 18712 2900 18752
rect 3244 18712 3284 18752
rect 3532 18712 3572 18752
rect 9292 18712 9332 18752
rect 9964 18712 10004 18752
rect 14764 18712 14804 18752
rect 17356 18712 17396 18752
rect 22636 18754 22676 18794
rect 19084 18712 19124 18752
rect 20908 18712 20948 18752
rect 21388 18712 21428 18752
rect 27916 18712 27956 18752
rect 32908 18712 32948 18752
rect 40492 18712 40532 18752
rect 17164 18628 17204 18668
rect 21100 18628 21140 18668
rect 28204 18628 28244 18668
rect 32140 18628 32180 18668
rect 37900 18628 37940 18668
rect 2764 18544 2804 18584
rect 2956 18544 2996 18584
rect 3052 18544 3092 18584
rect 3436 18544 3476 18584
rect 3724 18544 3764 18584
rect 4588 18544 4628 18584
rect 5836 18544 5876 18584
rect 6220 18544 6260 18584
rect 6412 18544 6452 18584
rect 6508 18544 6548 18584
rect 6700 18544 6740 18584
rect 6796 18544 6836 18584
rect 6892 18544 6932 18584
rect 6988 18544 7028 18584
rect 7180 18544 7220 18584
rect 7852 18544 7892 18584
rect 8044 18544 8084 18584
rect 8236 18544 8276 18584
rect 8332 18544 8372 18584
rect 8812 18544 8852 18584
rect 10636 18544 10676 18584
rect 15916 18544 15956 18584
rect 16780 18544 16820 18584
rect 18028 18544 18068 18584
rect 18892 18544 18932 18584
rect 19084 18544 19124 18584
rect 19276 18544 19316 18584
rect 19372 18544 19412 18584
rect 19564 18544 19604 18584
rect 19756 18544 19796 18584
rect 20620 18544 20660 18584
rect 20716 18544 20756 18584
rect 21292 18544 21332 18584
rect 21388 18544 21428 18584
rect 22444 18544 22484 18584
rect 22623 18544 22663 18584
rect 24172 18544 24212 18584
rect 24364 18544 24404 18584
rect 24460 18544 24500 18584
rect 24652 18544 24692 18584
rect 24844 18544 24884 18584
rect 26092 18544 26132 18584
rect 28012 18544 28052 18584
rect 28684 18544 28724 18584
rect 28780 18544 28820 18584
rect 29356 18544 29396 18584
rect 29548 18544 29588 18584
rect 29644 18544 29684 18584
rect 29836 18544 29876 18584
rect 30028 18544 30068 18584
rect 30316 18544 30356 18584
rect 30508 18544 30548 18584
rect 32524 18544 32564 18584
rect 33004 18544 33044 18584
rect 33100 18544 33140 18584
rect 33196 18544 33236 18584
rect 33676 18544 33716 18584
rect 34348 18544 34388 18584
rect 34540 18544 34580 18584
rect 34924 18544 34964 18584
rect 35788 18544 35828 18584
rect 37036 18544 37076 18584
rect 38284 18544 38324 18584
rect 39148 18544 39188 18584
rect 41644 18544 41684 18584
rect 42508 18544 42548 18584
rect 42892 18544 42932 18584
rect 44236 18544 44276 18584
rect 45484 18544 45524 18584
rect 46348 18544 46388 18584
rect 46732 18544 46772 18584
rect 5644 18460 5684 18500
rect 24748 18460 24788 18500
rect 27532 18460 27572 18500
rect 37420 18460 37460 18500
rect 1708 18376 1748 18416
rect 6412 18376 6452 18416
rect 10828 18376 10868 18416
rect 12556 18376 12596 18416
rect 24460 18376 24500 18416
rect 27724 18376 27764 18416
rect 4396 18292 4436 18332
rect 5260 18292 5300 18332
rect 5836 18292 5876 18332
rect 8044 18292 8084 18332
rect 9292 18292 9332 18332
rect 18220 18292 18260 18332
rect 19660 18292 19700 18332
rect 25612 18292 25652 18332
rect 28492 18292 28532 18332
rect 29356 18292 29396 18332
rect 29932 18292 29972 18332
rect 30316 18292 30356 18332
rect 40300 18292 40340 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 5452 17956 5492 17996
rect 11116 17956 11156 17996
rect 14476 17956 14516 17996
rect 18988 17956 19028 17996
rect 1036 17872 1076 17912
rect 6604 17872 6644 17912
rect 21100 17872 21140 17912
rect 24844 17872 24884 17912
rect 28012 17872 28052 17912
rect 29356 17872 29396 17912
rect 30028 17872 30068 17912
rect 30988 17872 31028 17912
rect 32428 17872 32468 17912
rect 35980 17872 36020 17912
rect 40492 17872 40532 17912
rect 41740 17872 41780 17912
rect 3628 17788 3668 17828
rect 17164 17788 17204 17828
rect 20812 17788 20852 17828
rect 24748 17788 24788 17828
rect 24940 17788 24980 17828
rect 28972 17788 29012 17828
rect 1612 17704 1652 17744
rect 2476 17704 2516 17744
rect 3916 17704 3956 17744
rect 4780 17704 4820 17744
rect 5836 17704 5876 17744
rect 5932 17704 5972 17744
rect 6028 17704 6068 17744
rect 6124 17704 6164 17744
rect 6508 17704 6548 17744
rect 6700 17704 6740 17744
rect 6796 17704 6836 17744
rect 6988 17704 7028 17744
rect 7372 17704 7412 17744
rect 7852 17704 7892 17744
rect 9100 17704 9140 17744
rect 9964 17704 10004 17744
rect 12076 17704 12116 17744
rect 12460 17704 12500 17744
rect 13324 17704 13364 17744
rect 15148 17704 15188 17744
rect 16012 17704 16052 17744
rect 17356 17704 17396 17744
rect 17452 17704 17492 17744
rect 17548 17704 17588 17744
rect 17644 17704 17684 17744
rect 17836 17704 17876 17744
rect 18508 17704 18548 17744
rect 18700 17704 18740 17744
rect 18796 17704 18836 17744
rect 18988 17704 19028 17744
rect 19180 17704 19220 17744
rect 19276 17704 19316 17744
rect 19468 17704 19508 17744
rect 19756 17704 19796 17744
rect 20620 17704 20660 17744
rect 20716 17704 20756 17744
rect 20908 17704 20948 17744
rect 21292 17704 21332 17744
rect 21388 17704 21428 17744
rect 21484 17704 21524 17744
rect 21580 17704 21620 17744
rect 21964 17704 22004 17744
rect 22828 17704 22868 17744
rect 23788 17704 23828 17744
rect 24268 17704 24308 17744
rect 24652 17704 24692 17744
rect 25036 17704 25076 17744
rect 25420 17704 25460 17744
rect 26380 17704 26420 17744
rect 27532 17704 27572 17744
rect 28012 17704 28052 17744
rect 28684 17704 28724 17744
rect 28780 17704 28820 17744
rect 29356 17704 29396 17744
rect 29740 17704 29780 17744
rect 29836 17704 29876 17744
rect 30028 17704 30068 17744
rect 30508 17704 30548 17744
rect 30700 17704 30740 17744
rect 30796 17704 30836 17744
rect 30988 17704 31028 17744
rect 31180 17704 31220 17744
rect 31852 17704 31892 17744
rect 33100 17704 33140 17744
rect 33196 17704 33236 17744
rect 33292 17704 33332 17744
rect 34252 17704 34292 17744
rect 34444 17704 34484 17744
rect 35308 17704 35348 17744
rect 36844 17704 36884 17744
rect 37708 17704 37748 17744
rect 38860 17704 38900 17744
rect 39532 17704 39572 17744
rect 40204 17704 40244 17744
rect 40300 17704 40340 17744
rect 40492 17704 40532 17744
rect 40684 17704 40724 17744
rect 41356 17704 41396 17744
rect 1228 17620 1268 17660
rect 4588 17620 4628 17660
rect 7468 17620 7508 17660
rect 8524 17620 8564 17660
rect 8716 17620 8756 17660
rect 14764 17620 14804 17660
rect 24460 17620 24500 17660
rect 26668 17620 26708 17660
rect 33388 17620 33428 17660
rect 33580 17620 33620 17660
rect 5644 17536 5684 17576
rect 19372 17536 19412 17576
rect 19660 17536 19700 17576
rect 22156 17536 22196 17576
rect 22348 17536 22388 17576
rect 24172 17536 24212 17576
rect 28204 17536 28244 17576
rect 29548 17536 29588 17576
rect 30604 17536 30644 17576
rect 37324 17536 37364 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 6988 17258 7028 17298
rect 652 17200 692 17240
rect 3724 17200 3764 17240
rect 6220 17200 6260 17240
rect 16300 17200 16340 17240
rect 18316 17200 18356 17240
rect 18412 17200 18452 17240
rect 18700 17200 18740 17240
rect 21868 17200 21908 17240
rect 22540 17200 22580 17240
rect 24844 17200 24884 17240
rect 25228 17200 25268 17240
rect 26572 17200 26612 17240
rect 16012 17116 16052 17156
rect 18220 17116 18260 17156
rect 18796 17116 18836 17156
rect 22252 17116 22292 17156
rect 43276 17116 43316 17156
rect 1324 17032 1364 17072
rect 1708 17032 1748 17072
rect 2572 17032 2612 17072
rect 3916 17032 3956 17072
rect 4876 17032 4916 17072
rect 5932 17032 5972 17072
rect 6124 17032 6164 17072
rect 6412 17032 6452 17072
rect 6508 17032 6548 17072
rect 7180 17032 7220 17072
rect 7084 16990 7124 17030
rect 8332 17032 8372 17072
rect 8524 17032 8564 17072
rect 9196 17032 9236 17072
rect 9388 17032 9428 17072
rect 9772 17032 9812 17072
rect 10636 17032 10676 17072
rect 11788 17032 11828 17072
rect 13996 17032 14036 17072
rect 15916 17032 15956 17072
rect 16108 17032 16148 17072
rect 16972 17032 17012 17072
rect 17164 17032 17204 17072
rect 17836 17032 17876 17072
rect 18028 17032 18068 17072
rect 18124 17032 18164 17072
rect 18892 17032 18932 17072
rect 18988 17032 19028 17072
rect 19180 17032 19220 17072
rect 20044 17032 20084 17072
rect 21004 17032 21044 17072
rect 21196 17032 21236 17072
rect 21964 17032 22004 17072
rect 22156 17032 22196 17072
rect 22348 17032 22388 17072
rect 22636 17032 22676 17072
rect 24268 17032 24308 17072
rect 24748 17032 24788 17072
rect 24940 17032 24980 17072
rect 25132 17032 25172 17072
rect 25420 17032 25460 17072
rect 25612 17032 25652 17072
rect 25708 17032 25748 17072
rect 25804 17032 25844 17072
rect 25900 17032 25940 17072
rect 26380 17032 26420 17072
rect 26572 17032 26612 17072
rect 27532 17032 27572 17072
rect 27916 17032 27956 17072
rect 28108 17032 28148 17072
rect 28204 17032 28244 17072
rect 28300 17032 28340 17072
rect 28396 17032 28436 17072
rect 28588 17032 28628 17072
rect 28684 17032 28724 17072
rect 28780 17032 28820 17072
rect 28876 17032 28916 17072
rect 29068 17032 29108 17072
rect 29260 17032 29300 17072
rect 29356 17032 29396 17072
rect 29548 17032 29588 17072
rect 29932 17032 29972 17072
rect 30412 17032 30452 17072
rect 30508 17032 30548 17072
rect 30700 17032 30740 17072
rect 30892 17032 30932 17072
rect 30988 17032 31028 17072
rect 31084 17032 31124 17072
rect 31180 17032 31220 17072
rect 31372 17032 31412 17072
rect 31468 17032 31508 17072
rect 32620 17032 32660 17072
rect 33292 17032 33332 17072
rect 33676 17032 33716 17072
rect 34540 17032 34580 17072
rect 36652 17032 36692 17072
rect 37324 17032 37364 17072
rect 37708 17032 37748 17072
rect 38572 17032 38612 17072
rect 42892 17032 42932 17072
rect 44140 17032 44180 17072
rect 6604 16948 6644 16988
rect 24460 16948 24500 16988
rect 27628 16948 27668 16988
rect 27820 16948 27860 16988
rect 29644 16948 29684 16988
rect 29836 16948 29876 16988
rect 31564 16948 31604 16988
rect 35692 16948 35732 16988
rect 37036 16948 37076 16988
rect 39724 16948 39764 16988
rect 6700 16864 6740 16904
rect 6796 16864 6836 16904
rect 7468 16864 7508 16904
rect 12076 16864 12116 16904
rect 15244 16864 15284 16904
rect 27724 16864 27764 16904
rect 29068 16864 29108 16904
rect 29740 16864 29780 16904
rect 30700 16864 30740 16904
rect 31660 16864 31700 16904
rect 5260 16780 5300 16820
rect 7660 16780 7700 16820
rect 14668 16780 14708 16820
rect 18700 16780 18740 16820
rect 21100 16780 21140 16820
rect 22828 16780 22868 16820
rect 24268 16780 24308 16820
rect 31756 16780 31796 16820
rect 31948 16780 31988 16820
rect 35980 16780 36020 16820
rect 36844 16780 36884 16820
rect 42604 16780 42644 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 8332 16444 8372 16484
rect 29644 16444 29684 16484
rect 36940 16444 36980 16484
rect 940 16360 980 16400
rect 2092 16360 2132 16400
rect 10252 16360 10292 16400
rect 13612 16360 13652 16400
rect 16204 16360 16244 16400
rect 16588 16360 16628 16400
rect 17548 16360 17588 16400
rect 21772 16360 21812 16400
rect 27244 16360 27284 16400
rect 31180 16360 31220 16400
rect 32620 16360 32660 16400
rect 37804 16360 37844 16400
rect 38188 16360 38228 16400
rect 16396 16276 16436 16316
rect 21580 16276 21620 16316
rect 27148 16276 27188 16316
rect 27340 16276 27380 16316
rect 34156 16276 34196 16316
rect 35212 16276 35252 16316
rect 41644 16276 41684 16316
rect 1132 16192 1172 16232
rect 1324 16192 1364 16232
rect 1516 16192 1556 16232
rect 1612 16192 1652 16232
rect 1804 16192 1844 16232
rect 1996 16192 2036 16232
rect 2188 16192 2228 16232
rect 2284 16192 2324 16232
rect 3148 16192 3188 16232
rect 4012 16192 4052 16232
rect 4204 16192 4244 16232
rect 4876 16192 4916 16232
rect 5260 16192 5300 16232
rect 5356 16192 5396 16232
rect 6412 16192 6452 16232
rect 6604 16192 6644 16232
rect 7276 16192 7316 16232
rect 8140 16192 8180 16232
rect 8332 16192 8372 16232
rect 8620 16192 8660 16232
rect 9580 16192 9620 16232
rect 10924 16192 10964 16232
rect 11596 16192 11636 16232
rect 12460 16192 12500 16232
rect 14188 16192 14228 16232
rect 15052 16192 15092 16232
rect 16012 16192 16052 16232
rect 16204 16192 16244 16232
rect 16780 16192 16820 16232
rect 16876 16192 16916 16232
rect 16972 16192 17012 16232
rect 17068 16192 17108 16232
rect 17260 16192 17300 16232
rect 17356 16192 17396 16232
rect 17548 16192 17588 16232
rect 18700 16192 18740 16232
rect 20140 16192 20180 16232
rect 20236 16192 20276 16232
rect 20428 16192 20468 16232
rect 20620 16192 20660 16232
rect 20812 16192 20852 16232
rect 20908 16192 20948 16232
rect 21772 16192 21812 16232
rect 23884 16192 23924 16232
rect 24076 16192 24116 16232
rect 25228 16192 25268 16232
rect 25900 16192 25940 16232
rect 27052 16192 27092 16232
rect 27436 16192 27476 16232
rect 27916 16192 27956 16232
rect 28012 16192 28052 16232
rect 28108 16192 28148 16232
rect 29356 16192 29396 16232
rect 29452 16192 29492 16232
rect 29644 16192 29684 16232
rect 30412 16192 30452 16232
rect 30508 16192 30548 16232
rect 30700 16192 30740 16232
rect 31084 16192 31124 16232
rect 31276 16192 31316 16232
rect 32140 16192 32180 16232
rect 32332 16192 32372 16232
rect 32428 16192 32468 16232
rect 34060 16192 34100 16232
rect 34252 16192 34292 16232
rect 35980 16192 36020 16232
rect 36652 16192 36692 16232
rect 36940 16192 36980 16232
rect 37132 16171 37172 16211
rect 37228 16171 37268 16211
rect 37324 16192 37364 16232
rect 37996 16192 38036 16232
rect 38188 16192 38228 16232
rect 38380 16192 38420 16232
rect 39628 16192 39668 16232
rect 40492 16192 40532 16232
rect 41836 16192 41876 16232
rect 1228 16108 1268 16148
rect 5068 16108 5108 16148
rect 11212 16108 11252 16148
rect 32524 16108 32564 16148
rect 39052 16108 39092 16148
rect 39244 16108 39284 16148
rect 1708 16024 1748 16064
rect 2476 16024 2516 16064
rect 3340 16024 3380 16064
rect 5356 16024 5396 16064
rect 5740 16024 5780 16064
rect 7468 16024 7508 16064
rect 8908 16024 8948 16064
rect 18220 16024 18260 16064
rect 20428 16024 20468 16064
rect 20908 16024 20948 16064
rect 23980 16024 24020 16064
rect 24748 16024 24788 16064
rect 25516 16024 25556 16064
rect 25708 16024 25748 16064
rect 30700 16024 30740 16064
rect 31468 16024 31508 16064
rect 32620 16024 32660 16064
rect 37420 16024 37460 16064
rect 42508 16024 42548 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 748 15688 788 15728
rect 3916 15688 3956 15728
rect 7084 15688 7124 15728
rect 7660 15688 7700 15728
rect 10348 15688 10388 15728
rect 20140 15688 20180 15728
rect 21772 15692 21812 15732
rect 28492 15688 28532 15728
rect 29260 15688 29300 15728
rect 29932 15688 29972 15728
rect 33580 15688 33620 15728
rect 38092 15688 38132 15728
rect 7948 15604 7988 15644
rect 26092 15604 26132 15644
rect 27340 15604 27380 15644
rect 28588 15604 28628 15644
rect 29836 15604 29876 15644
rect 1132 15520 1172 15560
rect 1516 15520 1556 15560
rect 2380 15520 2420 15560
rect 3820 15520 3860 15560
rect 4012 15520 4052 15560
rect 4876 15520 4916 15560
rect 5164 15520 5204 15560
rect 5356 15520 5396 15560
rect 5452 15520 5492 15560
rect 5644 15520 5684 15560
rect 6508 15520 6548 15560
rect 6604 15520 6644 15560
rect 6700 15520 6740 15560
rect 6796 15520 6836 15560
rect 6988 15520 7028 15560
rect 7180 15520 7220 15560
rect 7276 15520 7316 15560
rect 7468 15520 7508 15560
rect 7564 15520 7604 15560
rect 7756 15520 7796 15560
rect 8332 15520 8372 15560
rect 9196 15520 9236 15560
rect 11980 15520 12020 15560
rect 12556 15520 12596 15560
rect 14380 15520 14420 15560
rect 15244 15520 15284 15560
rect 15628 15520 15668 15560
rect 15820 15520 15860 15560
rect 16492 15520 16532 15560
rect 17644 15520 17684 15560
rect 18412 15520 18452 15560
rect 18508 15520 18548 15560
rect 18604 15520 18644 15560
rect 18796 15520 18836 15560
rect 18892 15520 18932 15560
rect 18988 15520 19028 15560
rect 19084 15520 19124 15560
rect 19276 15520 19316 15560
rect 19468 15520 19508 15560
rect 19660 15520 19700 15560
rect 19756 15520 19796 15560
rect 19948 15520 19988 15560
rect 20140 15520 20180 15560
rect 20332 15520 20372 15560
rect 20428 15520 20468 15560
rect 20620 15520 20660 15560
rect 20716 15520 20756 15560
rect 20812 15520 20852 15560
rect 20908 15520 20948 15560
rect 21868 15520 21908 15560
rect 21964 15520 22004 15560
rect 25228 15520 25268 15560
rect 26860 15520 26900 15560
rect 27532 15520 27572 15560
rect 27820 15520 27860 15560
rect 28684 15520 28724 15560
rect 28780 15520 28820 15560
rect 28972 15520 29012 15560
rect 29068 15520 29108 15560
rect 29164 15520 29204 15560
rect 29644 15520 29684 15560
rect 29740 15520 29780 15560
rect 30316 15520 30356 15560
rect 31468 15520 31508 15560
rect 31564 15520 31604 15560
rect 31660 15520 31700 15560
rect 31756 15520 31796 15560
rect 32332 15520 32372 15560
rect 32524 15520 32564 15560
rect 32620 15520 32660 15560
rect 33100 15520 33140 15560
rect 33196 15520 33236 15560
rect 33388 15520 33428 15560
rect 33676 15520 33716 15560
rect 34060 15520 34100 15560
rect 34156 15520 34196 15560
rect 34252 15520 34292 15560
rect 34348 15520 34388 15560
rect 34540 15520 34580 15560
rect 35212 15520 35252 15560
rect 35404 15520 35444 15560
rect 35788 15520 35828 15560
rect 36652 15520 36692 15560
rect 38188 15520 38228 15560
rect 38284 15520 38324 15560
rect 38380 15520 38420 15560
rect 40972 15520 41012 15560
rect 41932 15520 41972 15560
rect 43948 15520 43988 15560
rect 5260 15436 5300 15476
rect 11212 15436 11252 15476
rect 23884 15436 23924 15476
rect 24364 15436 24404 15476
rect 19468 15352 19508 15392
rect 19660 15352 19700 15392
rect 28684 15352 28724 15392
rect 29932 15352 29972 15392
rect 32620 15352 32660 15392
rect 39724 15352 39764 15392
rect 3532 15268 3572 15308
rect 4204 15268 4244 15308
rect 6316 15268 6356 15308
rect 12652 15268 12692 15308
rect 13228 15268 13268 15308
rect 17068 15268 17108 15308
rect 22252 15268 22292 15308
rect 23692 15268 23732 15308
rect 26284 15268 26324 15308
rect 30604 15268 30644 15308
rect 33388 15268 33428 15308
rect 33868 15268 33908 15308
rect 37804 15268 37844 15308
rect 44428 15268 44468 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4780 14932 4820 14972
rect 5644 14932 5684 14972
rect 11116 14932 11156 14972
rect 11980 14932 12020 14972
rect 13804 14932 13844 14972
rect 24844 14932 24884 14972
rect 27244 14932 27284 14972
rect 30892 14932 30932 14972
rect 31468 14932 31508 14972
rect 32428 14932 32468 14972
rect 34444 14932 34484 14972
rect 1708 14848 1748 14888
rect 8236 14848 8276 14888
rect 8524 14848 8564 14888
rect 9868 14848 9908 14888
rect 16684 14848 16724 14888
rect 19084 14848 19124 14888
rect 10060 14764 10100 14804
rect 18988 14764 19028 14804
rect 19180 14806 19220 14846
rect 21004 14848 21044 14888
rect 22252 14848 22292 14888
rect 25132 14848 25172 14888
rect 31084 14848 31124 14888
rect 33292 14848 33332 14888
rect 37900 14848 37940 14888
rect 39052 14848 39092 14888
rect 41356 14848 41396 14888
rect 46924 14848 46964 14888
rect 20908 14764 20948 14804
rect 21100 14764 21140 14804
rect 22156 14764 22196 14804
rect 22348 14764 22388 14804
rect 26860 14764 26900 14804
rect 30700 14764 30740 14804
rect 33196 14764 33236 14804
rect 33388 14764 33428 14804
rect 2380 14680 2420 14720
rect 2764 14680 2804 14720
rect 3628 14680 3668 14720
rect 5164 14680 5204 14720
rect 5260 14680 5300 14720
rect 5356 14680 5396 14720
rect 5452 14680 5492 14720
rect 5836 14680 5876 14720
rect 6220 14680 6260 14720
rect 7084 14680 7124 14720
rect 8908 14680 8948 14720
rect 9100 14680 9140 14720
rect 10444 14680 10484 14720
rect 11308 14680 11348 14720
rect 12268 14680 12308 14720
rect 12652 14659 12692 14699
rect 12748 14659 12788 14699
rect 12844 14680 12884 14720
rect 13228 14680 13268 14720
rect 14956 14680 14996 14720
rect 15244 14680 15284 14720
rect 15340 14680 15380 14720
rect 15532 14680 15572 14720
rect 15724 14680 15764 14720
rect 16204 14680 16244 14720
rect 16300 14680 16340 14720
rect 16492 14680 16532 14720
rect 16684 14680 16724 14720
rect 16972 14680 17012 14720
rect 18124 14680 18164 14720
rect 18508 14680 18548 14720
rect 18892 14680 18932 14720
rect 19276 14680 19316 14720
rect 19756 14680 19796 14720
rect 19852 14680 19892 14720
rect 20044 14680 20084 14720
rect 20332 14680 20372 14720
rect 20428 14680 20468 14720
rect 20524 14680 20564 14720
rect 20620 14680 20660 14720
rect 20812 14680 20852 14720
rect 21196 14680 21236 14720
rect 21388 14680 21428 14720
rect 21484 14680 21524 14720
rect 21580 14680 21620 14720
rect 22060 14680 22100 14720
rect 22444 14680 22484 14720
rect 23596 14680 23636 14720
rect 23692 14680 23732 14720
rect 23788 14680 23828 14720
rect 23980 14680 24020 14720
rect 24076 14680 24116 14720
rect 24172 14680 24212 14720
rect 24364 14680 24404 14720
rect 24556 14680 24596 14720
rect 24652 14680 24692 14720
rect 25420 14680 25460 14720
rect 25516 14680 25556 14720
rect 25804 14680 25844 14720
rect 26188 14680 26228 14720
rect 26764 14680 26804 14720
rect 26956 14680 26996 14720
rect 27148 14680 27188 14720
rect 27340 14703 27380 14743
rect 27532 14680 27572 14720
rect 27724 14680 27764 14720
rect 28108 14680 28148 14720
rect 28204 14680 28244 14720
rect 28684 14680 28724 14720
rect 28780 14680 28820 14720
rect 28972 14680 29012 14720
rect 29164 14680 29204 14720
rect 29260 14680 29300 14720
rect 29356 14680 29396 14720
rect 29452 14680 29492 14720
rect 29644 14680 29684 14720
rect 29740 14680 29780 14720
rect 29932 14680 29972 14720
rect 31084 14680 31124 14720
rect 31276 14680 31316 14720
rect 31468 14680 31508 14720
rect 31756 14680 31796 14720
rect 31948 14680 31988 14720
rect 15436 14596 15476 14636
rect 15820 14596 15860 14636
rect 18604 14596 18644 14636
rect 27628 14596 27668 14636
rect 29836 14596 29876 14636
rect 31660 14638 31700 14678
rect 32044 14680 32084 14720
rect 32140 14680 32180 14720
rect 32236 14680 32276 14720
rect 32716 14680 32756 14720
rect 32812 14680 32852 14720
rect 33100 14680 33140 14720
rect 33484 14680 33524 14720
rect 33676 14680 33716 14720
rect 33772 14680 33812 14720
rect 33868 14680 33908 14720
rect 33964 14680 34004 14720
rect 34156 14680 34196 14720
rect 34252 14680 34292 14720
rect 34444 14680 34484 14720
rect 34636 14680 34676 14720
rect 34732 14680 34772 14720
rect 34828 14680 34868 14720
rect 37612 14680 37652 14720
rect 39724 14680 39764 14720
rect 40972 14680 41012 14720
rect 41068 14680 41108 14720
rect 41740 14680 41780 14720
rect 42124 14680 42164 14720
rect 42988 14680 43028 14720
rect 44140 14680 44180 14720
rect 44524 14680 44564 14720
rect 45676 14680 45716 14720
rect 46540 14680 46580 14720
rect 47596 14680 47636 14720
rect 652 14512 692 14552
rect 1036 14512 1076 14552
rect 9004 14512 9044 14552
rect 11788 14512 11828 14552
rect 12556 14512 12596 14552
rect 14284 14512 14324 14552
rect 17452 14512 17492 14552
rect 19948 14512 19988 14552
rect 23500 14512 23540 14552
rect 26092 14512 26132 14552
rect 26380 14512 26420 14552
rect 28492 14512 28532 14552
rect 28876 14512 28916 14552
rect 32908 14508 32948 14548
rect 40876 14508 40916 14548
rect 45004 14512 45044 14552
rect 46924 14512 46964 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 652 14176 692 14216
rect 4012 14176 4052 14216
rect 4300 14176 4340 14216
rect 5644 14176 5684 14216
rect 6316 14176 6356 14216
rect 6604 14176 6644 14216
rect 9772 14176 9812 14216
rect 15628 14176 15668 14216
rect 17164 14176 17204 14216
rect 18412 14176 18452 14216
rect 21100 14176 21140 14216
rect 22252 14176 22292 14216
rect 22444 14176 22484 14216
rect 23116 14176 23156 14216
rect 26092 14176 26132 14216
rect 35212 14176 35252 14216
rect 36172 14176 36212 14216
rect 37132 14176 37172 14216
rect 38380 14176 38420 14216
rect 41740 14176 41780 14216
rect 42028 14176 42068 14216
rect 20044 14092 20084 14132
rect 22924 14092 22964 14132
rect 27436 14092 27476 14132
rect 3244 14008 3284 14048
rect 3436 14008 3476 14048
rect 4204 13991 4244 14031
rect 4588 14008 4628 14048
rect 4684 14008 4724 14048
rect 4876 14008 4916 14048
rect 5068 14008 5108 14048
rect 5164 14008 5204 14048
rect 5356 14008 5396 14048
rect 5548 14008 5588 14048
rect 5740 14008 5780 14048
rect 5836 14008 5876 14048
rect 6028 14008 6068 14048
rect 6124 14008 6164 14048
rect 6316 14008 6356 14048
rect 6700 14008 6740 14048
rect 8044 14008 8084 14048
rect 10924 14008 10964 14048
rect 11788 14008 11828 14048
rect 12172 14008 12212 14048
rect 12460 14008 12500 14048
rect 13132 14008 13172 14048
rect 13804 14008 13844 14048
rect 14764 14008 14804 14048
rect 15724 14008 15764 14048
rect 15820 14008 15860 14048
rect 15916 14008 15956 14048
rect 17068 14008 17108 14048
rect 17452 14008 17492 14048
rect 18124 14008 18164 14048
rect 18604 14008 18644 14048
rect 18705 14017 18745 14057
rect 18892 14008 18932 14048
rect 18988 14008 19028 14048
rect 19084 14008 19124 14048
rect 19180 14008 19220 14048
rect 19660 14008 19700 14048
rect 19948 14008 19988 14048
rect 20620 14008 20660 14048
rect 20716 14008 20756 14048
rect 20908 14008 20948 14048
rect 21004 14008 21044 14048
rect 21105 14008 21145 14048
rect 21388 14008 21428 14048
rect 21772 14008 21812 14048
rect 21964 14008 22004 14048
rect 22636 14008 22676 14048
rect 24268 14008 24308 14048
rect 26476 14008 26516 14048
rect 27532 14008 27572 14048
rect 27820 14008 27860 14048
rect 28204 14008 28244 14048
rect 28300 14008 28340 14048
rect 28396 14008 28436 14048
rect 28492 14008 28532 14048
rect 30220 14008 30260 14048
rect 30316 14008 30356 14048
rect 30412 14008 30452 14048
rect 30508 14008 30548 14048
rect 31756 14008 31796 14048
rect 31948 14029 31988 14069
rect 32140 14008 32180 14048
rect 32524 14008 32564 14048
rect 32716 14008 32756 14048
rect 33100 14008 33140 14048
rect 33292 14008 33332 14048
rect 33676 14008 33716 14048
rect 33868 14008 33908 14048
rect 34156 14008 34196 14048
rect 34924 14008 34964 14048
rect 35020 14008 35060 14048
rect 35404 14008 35444 14048
rect 35692 14008 35732 14048
rect 35884 14008 35924 14048
rect 35980 14008 36020 14048
rect 36364 14008 36404 14048
rect 36556 14008 36596 14048
rect 36652 14008 36692 14048
rect 36844 14008 36884 14048
rect 36940 14008 36980 14048
rect 37324 14008 37364 14048
rect 37612 14008 37652 14048
rect 37996 14008 38036 14048
rect 38860 14008 38900 14048
rect 40684 14008 40724 14048
rect 41548 14008 41588 14048
rect 41932 14008 41972 14048
rect 42508 14008 42548 14048
rect 43468 14008 43508 14048
rect 44140 14008 44180 14048
rect 44524 14008 44564 14048
rect 45388 14008 45428 14048
rect 46636 14008 46676 14048
rect 17644 13924 17684 13964
rect 21484 13924 21524 13964
rect 21676 13924 21716 13964
rect 32236 13924 32276 13964
rect 32428 13924 32468 13964
rect 32812 13922 32852 13962
rect 33004 13924 33044 13964
rect 33388 13924 33428 13964
rect 33580 13924 33620 13964
rect 34060 13924 34100 13964
rect 3820 13840 3860 13880
rect 4876 13840 4916 13880
rect 5068 13840 5108 13880
rect 7372 13840 7412 13880
rect 8812 13840 8852 13880
rect 14092 13840 14132 13880
rect 15148 13840 15188 13880
rect 17548 13840 17588 13880
rect 21580 13840 21620 13880
rect 24556 13840 24596 13880
rect 24940 13840 24980 13880
rect 27148 13840 27188 13880
rect 32332 13840 32372 13880
rect 32908 13840 32948 13880
rect 33484 13840 33524 13880
rect 35692 13840 35732 13880
rect 39532 13840 39572 13880
rect 3436 13756 3476 13796
rect 14476 13756 14516 13796
rect 16876 13756 16916 13796
rect 18220 13756 18260 13796
rect 20332 13756 20372 13796
rect 25900 13756 25940 13796
rect 31852 13756 31892 13796
rect 36364 13756 36404 13796
rect 37612 13756 37652 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 23308 13420 23348 13460
rect 25804 13420 25844 13460
rect 30124 13420 30164 13460
rect 30604 13420 30644 13460
rect 31660 13420 31700 13460
rect 32908 13420 32948 13460
rect 3436 13336 3476 13376
rect 5356 13336 5396 13376
rect 12940 13336 12980 13376
rect 17836 13336 17876 13376
rect 19084 13336 19124 13376
rect 19852 13336 19892 13376
rect 20908 13336 20948 13376
rect 28684 13336 28724 13376
rect 29740 13336 29780 13376
rect 32236 13336 32276 13376
rect 42412 13336 42452 13376
rect 17740 13252 17780 13292
rect 17932 13252 17972 13292
rect 19756 13252 19796 13292
rect 19948 13252 19988 13292
rect 22348 13252 22388 13292
rect 32140 13252 32180 13292
rect 32332 13252 32372 13292
rect 42316 13252 42356 13292
rect 42508 13252 42548 13292
rect 3820 13168 3860 13208
rect 3916 13168 3956 13208
rect 4012 13168 4052 13208
rect 4972 13168 5012 13208
rect 5548 13168 5588 13208
rect 5644 13168 5684 13208
rect 5740 13168 5780 13208
rect 5836 13168 5876 13208
rect 6700 13168 6740 13208
rect 7852 13168 7892 13208
rect 9292 13168 9332 13208
rect 10156 13168 10196 13208
rect 11404 13168 11444 13208
rect 11884 13168 11924 13208
rect 11980 13168 12020 13208
rect 12172 13168 12212 13208
rect 12364 13168 12404 13208
rect 12460 13168 12500 13208
rect 12652 13168 12692 13208
rect 14092 13168 14132 13208
rect 14956 13168 14996 13208
rect 16204 13168 16244 13208
rect 17644 13168 17684 13208
rect 18028 13168 18068 13208
rect 18412 13168 18452 13208
rect 18700 13168 18740 13208
rect 18796 13168 18836 13208
rect 19276 13168 19316 13208
rect 19468 13168 19508 13208
rect 19660 13168 19700 13208
rect 20044 13168 20084 13208
rect 20428 13168 20468 13208
rect 20620 13153 20660 13193
rect 20716 13168 20756 13208
rect 20908 13168 20948 13208
rect 21100 13168 21140 13208
rect 21196 13168 21236 13208
rect 21292 13168 21332 13208
rect 21580 13168 21620 13208
rect 21772 13168 21812 13208
rect 22252 13168 22292 13208
rect 22444 13168 22484 13208
rect 22732 13168 22772 13208
rect 23308 13168 23348 13208
rect 23500 13168 23540 13208
rect 24652 13168 24692 13208
rect 25612 13168 25652 13208
rect 26188 13168 26228 13208
rect 26476 13168 26516 13208
rect 26764 13168 26804 13208
rect 26956 13168 26996 13208
rect 27724 13168 27764 13208
rect 27820 13168 27860 13208
rect 27916 13168 27956 13208
rect 28012 13168 28052 13208
rect 28300 13168 28340 13208
rect 28396 13168 28436 13208
rect 29068 13168 29108 13208
rect 29164 13168 29204 13208
rect 29260 13168 29300 13208
rect 29356 13168 29396 13208
rect 29740 13168 29780 13208
rect 30305 13168 30345 13208
rect 30412 13168 30452 13208
rect 30604 13168 30644 13208
rect 30796 13182 30836 13222
rect 30892 13168 30932 13208
rect 31564 13168 31604 13208
rect 31756 13168 31796 13208
rect 32044 13168 32084 13208
rect 32428 13168 32468 13208
rect 32812 13168 32852 13208
rect 33004 13168 33044 13208
rect 33580 13168 33620 13208
rect 33676 13168 33716 13208
rect 34060 13168 34100 13208
rect 34348 13168 34388 13208
rect 34924 13168 34964 13208
rect 35020 13168 35060 13208
rect 35404 13168 35444 13208
rect 35500 13168 35540 13208
rect 35692 13168 35732 13208
rect 35788 13168 35828 13208
rect 35889 13168 35929 13208
rect 36172 13168 36212 13208
rect 36460 13168 36500 13208
rect 37324 13168 37364 13208
rect 37420 13168 37460 13208
rect 37516 13168 37556 13208
rect 37612 13168 37652 13208
rect 37804 13168 37844 13208
rect 38764 13168 38804 13208
rect 39052 13168 39092 13208
rect 39436 13168 39476 13208
rect 40300 13168 40340 13208
rect 41452 13168 41492 13208
rect 41740 13168 41780 13208
rect 41932 13168 41972 13208
rect 42028 13168 42068 13208
rect 42220 13168 42260 13208
rect 42604 13168 42644 13208
rect 42796 13168 42836 13208
rect 43084 13168 43124 13208
rect 43564 13168 43604 13208
rect 44428 13168 44468 13208
rect 44812 13168 44852 13208
rect 45676 13168 45716 13208
rect 46828 13168 46868 13208
rect 47116 13168 47156 13208
rect 47308 13168 47348 13208
rect 47404 13168 47444 13208
rect 10540 13084 10580 13124
rect 10732 13084 10772 13124
rect 12556 13084 12596 13124
rect 15340 13084 15380 13124
rect 21676 13084 21716 13124
rect 22924 13084 22964 13124
rect 26092 13084 26132 13124
rect 30220 13084 30260 13124
rect 36364 13084 36404 13124
rect 43276 13084 43316 13124
rect 652 13000 692 13040
rect 4108 13000 4148 13040
rect 4300 13000 4340 13040
rect 6028 13000 6068 13040
rect 7372 13000 7412 13040
rect 8140 13000 8180 13040
rect 12076 13000 12116 13040
rect 15532 13000 15572 13040
rect 19372 13000 19412 13040
rect 20332 13000 20372 13040
rect 21388 13000 21428 13040
rect 22636 13000 22676 13040
rect 29548 13000 29588 13040
rect 30124 13000 30164 13040
rect 33868 13000 33908 13040
rect 34156 13000 34196 13040
rect 35212 13000 35252 13040
rect 35788 13000 35828 13040
rect 41740 13000 41780 13040
rect 44236 13000 44276 13040
rect 47116 13000 47156 13040
rect 28204 12942 28244 12982
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 652 12664 692 12704
rect 8812 12664 8852 12704
rect 27532 12664 27572 12704
rect 27820 12664 27860 12704
rect 28492 12664 28532 12704
rect 31852 12664 31892 12704
rect 35404 12664 35444 12704
rect 37996 12664 38036 12704
rect 38476 12664 38516 12704
rect 42124 12664 42164 12704
rect 10540 12580 10580 12620
rect 13612 12580 13652 12620
rect 16684 12580 16724 12620
rect 28972 12580 29012 12620
rect 32428 12580 32468 12620
rect 40684 12580 40724 12620
rect 42028 12580 42068 12620
rect 43852 12580 43892 12620
rect 2956 12496 2996 12536
rect 3340 12496 3380 12536
rect 4204 12496 4244 12536
rect 5452 12496 5492 12536
rect 5644 12496 5684 12536
rect 6028 12496 6068 12536
rect 6892 12496 6932 12536
rect 8044 12496 8084 12536
rect 8524 12496 8564 12536
rect 8620 12496 8660 12536
rect 9004 12496 9044 12536
rect 9676 12496 9716 12536
rect 9868 12496 9908 12536
rect 10732 12496 10772 12536
rect 11116 12496 11156 12536
rect 11212 12496 11252 12536
rect 11308 12496 11348 12536
rect 11404 12496 11444 12536
rect 11692 12496 11732 12536
rect 12940 12496 12980 12536
rect 14860 12496 14900 12536
rect 16588 12496 16628 12536
rect 16780 12496 16820 12536
rect 17068 12496 17108 12536
rect 17356 12523 17396 12563
rect 17452 12496 17492 12536
rect 17932 12496 17972 12536
rect 18316 12496 18356 12536
rect 18508 12496 18548 12536
rect 18604 12496 18644 12536
rect 18700 12496 18740 12536
rect 18796 12496 18836 12536
rect 19180 12496 19220 12536
rect 19564 12496 19604 12536
rect 19948 12496 19988 12536
rect 20044 12496 20084 12536
rect 20236 12496 20276 12536
rect 20428 12496 20468 12536
rect 20524 12496 20564 12536
rect 20716 12496 20756 12536
rect 20812 12496 20852 12536
rect 20913 12496 20953 12536
rect 21196 12496 21236 12536
rect 21388 12496 21428 12536
rect 21484 12496 21524 12536
rect 21676 12496 21716 12536
rect 21772 12496 21812 12536
rect 22252 12496 22292 12536
rect 22348 12496 22388 12536
rect 22636 12496 22676 12536
rect 26284 12496 26324 12536
rect 27244 12496 27284 12536
rect 27340 12496 27380 12536
rect 27916 12496 27956 12536
rect 28012 12496 28052 12536
rect 28108 12496 28148 12536
rect 28300 12496 28340 12536
rect 28396 12496 28436 12536
rect 28588 12496 28628 12536
rect 28780 12496 28820 12536
rect 28876 12496 28916 12536
rect 29068 12496 29108 12536
rect 29260 12496 29300 12536
rect 29452 12496 29492 12536
rect 30412 12496 30452 12536
rect 30796 12496 30836 12536
rect 30988 12496 31028 12536
rect 31372 12496 31412 12536
rect 31564 12496 31604 12536
rect 31660 12496 31700 12536
rect 31852 12496 31892 12536
rect 31948 12496 31988 12536
rect 32105 12481 32145 12521
rect 32332 12496 32372 12536
rect 32524 12496 32564 12536
rect 34060 12496 34100 12536
rect 34156 12496 34196 12536
rect 34348 12496 34388 12536
rect 34444 12496 34484 12536
rect 34599 12496 34639 12536
rect 34828 12496 34868 12536
rect 34924 12496 34964 12536
rect 35308 12496 35348 12536
rect 35596 12496 35636 12536
rect 37036 12496 37076 12536
rect 37228 12496 37268 12536
rect 37324 12496 37364 12536
rect 37516 12496 37556 12536
rect 37804 12496 37844 12536
rect 38188 12496 38228 12536
rect 38284 12496 38324 12536
rect 38668 12496 38708 12536
rect 38764 12496 38804 12536
rect 38956 12496 38996 12536
rect 39244 12496 39284 12536
rect 39628 12496 39668 12536
rect 41356 12496 41396 12536
rect 41836 12496 41876 12536
rect 41932 12496 41972 12536
rect 42604 12496 42644 12536
rect 42700 12496 42740 12536
rect 43180 12496 43220 12536
rect 44044 12496 44084 12536
rect 44428 12496 44468 12536
rect 45292 12496 45332 12536
rect 47596 12496 47636 12536
rect 48652 12496 48692 12536
rect 18028 12412 18068 12452
rect 18220 12412 18260 12452
rect 19276 12412 19316 12452
rect 19468 12412 19508 12452
rect 29356 12412 29396 12452
rect 30508 12412 30548 12452
rect 30700 12412 30740 12452
rect 31084 12412 31124 12452
rect 31276 12412 31316 12452
rect 37612 12412 37652 12452
rect 18124 12328 18164 12368
rect 19372 12328 19412 12368
rect 20236 12328 20276 12368
rect 21964 12328 22004 12368
rect 30604 12328 30644 12368
rect 31180 12328 31220 12368
rect 42124 12328 42164 12368
rect 42892 12328 42932 12368
rect 10828 12244 10868 12284
rect 12364 12244 12404 12284
rect 14668 12244 14708 12284
rect 17740 12244 17780 12284
rect 20428 12244 20468 12284
rect 21196 12244 21236 12284
rect 25612 12244 25652 12284
rect 34060 12244 34100 12284
rect 37036 12244 37076 12284
rect 38956 12244 38996 12284
rect 40204 12244 40244 12284
rect 41932 12244 41972 12284
rect 46444 12244 46484 12284
rect 46924 12244 46964 12284
rect 47980 12244 48020 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 6412 11908 6452 11948
rect 10156 11908 10196 11948
rect 12940 11908 12980 11948
rect 17740 11908 17780 11948
rect 27532 11908 27572 11948
rect 44716 11908 44756 11948
rect 45100 11908 45140 11948
rect 49324 11908 49364 11948
rect 4012 11824 4052 11864
rect 11404 11824 11444 11864
rect 14572 11824 14612 11864
rect 14956 11824 14996 11864
rect 16780 11824 16820 11864
rect 18988 11824 19028 11864
rect 31660 11824 31700 11864
rect 32044 11824 32084 11864
rect 6220 11740 6260 11780
rect 18892 11740 18932 11780
rect 19084 11740 19124 11780
rect 24844 11740 24884 11780
rect 26860 11740 26900 11780
rect 46732 11740 46772 11780
rect 3724 11656 3764 11696
rect 3820 11656 3860 11696
rect 4012 11656 4052 11696
rect 4204 11656 4244 11696
rect 4396 11656 4436 11696
rect 4492 11656 4532 11696
rect 4684 11656 4724 11696
rect 5548 11656 5588 11696
rect 6604 11656 6644 11696
rect 7948 11656 7988 11696
rect 8236 11656 8276 11696
rect 8428 11656 8468 11696
rect 8620 11656 8660 11696
rect 8716 11656 8756 11696
rect 8908 11656 8948 11696
rect 9004 11656 9044 11696
rect 9388 11656 9428 11696
rect 9580 11656 9620 11696
rect 9676 11656 9716 11696
rect 9868 11656 9908 11696
rect 9964 11656 10004 11696
rect 10156 11656 10196 11696
rect 11596 11656 11636 11696
rect 11692 11656 11732 11696
rect 11788 11656 11828 11696
rect 11884 11656 11924 11696
rect 12076 11656 12116 11696
rect 13036 11656 13076 11696
rect 13228 11656 13268 11696
rect 14092 11656 14132 11696
rect 14188 11656 14228 11696
rect 14284 11656 14324 11696
rect 14380 11656 14420 11696
rect 16108 11656 16148 11696
rect 16396 11656 16436 11696
rect 17068 11656 17108 11696
rect 17356 11656 17396 11696
rect 17452 11656 17492 11696
rect 18220 11656 18260 11696
rect 18316 11656 18356 11696
rect 18412 11656 18452 11696
rect 18796 11656 18836 11696
rect 19180 11656 19220 11696
rect 19852 11656 19892 11696
rect 19948 11656 19988 11696
rect 20044 11656 20084 11696
rect 20236 11656 20276 11696
rect 20332 11656 20372 11696
rect 20524 11671 20564 11711
rect 20620 11656 20660 11696
rect 20777 11671 20817 11711
rect 21100 11656 21140 11696
rect 21196 11656 21236 11696
rect 21388 11656 21428 11696
rect 21484 11656 21524 11696
rect 21641 11671 21681 11711
rect 23500 11656 23540 11696
rect 23596 11656 23636 11696
rect 23692 11656 23732 11696
rect 23980 11656 24020 11696
rect 26572 11656 26612 11696
rect 26668 11656 26708 11696
rect 27052 11656 27092 11696
rect 28012 11656 28052 11696
rect 28300 11656 28340 11696
rect 28492 11656 28532 11696
rect 28876 11656 28916 11696
rect 29068 11656 29108 11696
rect 29164 11656 29204 11696
rect 31468 11656 31508 11696
rect 31660 11656 31700 11696
rect 31948 11656 31988 11696
rect 32140 11656 32180 11696
rect 32236 11656 32276 11696
rect 32428 11656 32468 11696
rect 32524 11656 32564 11696
rect 32620 11656 32660 11696
rect 32908 11656 32948 11696
rect 33004 11656 33044 11696
rect 33772 11656 33812 11696
rect 33868 11656 33908 11696
rect 33964 11656 34004 11696
rect 34156 11656 34196 11696
rect 34252 11656 34292 11696
rect 34732 11656 34772 11696
rect 34828 11656 34868 11696
rect 34924 11656 34964 11696
rect 35212 11656 35252 11696
rect 36268 11656 36308 11696
rect 36556 11656 36596 11696
rect 36652 11656 36692 11696
rect 37420 11656 37460 11696
rect 38572 11656 38612 11696
rect 39244 11656 39284 11696
rect 39436 11656 39476 11696
rect 39532 11656 39572 11696
rect 40396 11656 40436 11696
rect 40492 11656 40532 11696
rect 41260 11656 41300 11696
rect 42124 11656 42164 11696
rect 43468 11656 43508 11696
rect 44332 11656 44372 11696
rect 44812 11656 44852 11696
rect 45772 11656 45812 11696
rect 46444 11656 46484 11696
rect 46540 11656 46580 11696
rect 46924 11656 46964 11696
rect 47308 11656 47348 11696
rect 48172 11656 48212 11696
rect 16492 11572 16532 11612
rect 32716 11572 32756 11612
rect 40876 11572 40916 11612
rect 652 11488 692 11528
rect 4300 11488 4340 11528
rect 5356 11488 5396 11528
rect 6700 11488 6740 11528
rect 8140 11488 8180 11528
rect 9196 11488 9236 11528
rect 9484 11488 9524 11528
rect 12748 11488 12788 11528
rect 13900 11488 13940 11528
rect 18124 11488 18164 11528
rect 19756 11488 19796 11528
rect 20428 11488 20468 11528
rect 21388 11488 21428 11528
rect 24460 11488 24500 11528
rect 28396 11488 28436 11528
rect 28972 11488 29012 11528
rect 33676 11488 33716 11528
rect 34444 11488 34484 11528
rect 34636 11488 34676 11528
rect 35308 11488 35348 11528
rect 36172 11488 36212 11528
rect 36844 11488 36884 11528
rect 37132 11488 37172 11528
rect 38092 11488 38132 11528
rect 39532 11488 39572 11528
rect 40684 11488 40724 11528
rect 43276 11488 43316 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 652 11152 692 11192
rect 3724 11152 3764 11192
rect 5548 11152 5588 11192
rect 9100 11152 9140 11192
rect 11308 11152 11348 11192
rect 16300 11152 16340 11192
rect 16780 11152 16820 11192
rect 17068 11152 17108 11192
rect 17260 11152 17300 11192
rect 27052 11152 27092 11192
rect 31756 11152 31796 11192
rect 35212 11152 35252 11192
rect 37516 11152 37556 11192
rect 40012 11152 40052 11192
rect 40876 11152 40916 11192
rect 42412 11152 42452 11192
rect 44236 11152 44276 11192
rect 45100 11152 45140 11192
rect 46636 11152 46676 11192
rect 48556 11152 48596 11192
rect 48844 11152 48884 11192
rect 10156 11068 10196 11108
rect 13708 11068 13748 11108
rect 29164 11068 29204 11108
rect 37804 11068 37844 11108
rect 42316 11068 42356 11108
rect 48460 11068 48500 11108
rect 2572 10984 2612 11024
rect 2668 10984 2708 11024
rect 2860 10984 2900 11024
rect 3628 10984 3668 11024
rect 4300 10984 4340 11024
rect 5260 10984 5300 11024
rect 5740 10984 5780 11024
rect 5836 10984 5876 11024
rect 5932 10984 5972 11024
rect 6028 10984 6068 11024
rect 6988 10984 7028 11024
rect 7660 10984 7700 11024
rect 7756 10984 7796 11024
rect 7852 10984 7892 11024
rect 7948 10984 7988 11024
rect 8140 10984 8180 11024
rect 8428 10984 8468 11024
rect 8620 10984 8660 11024
rect 8908 10984 8948 11024
rect 9292 10984 9332 11024
rect 9388 10984 9428 11024
rect 9676 10984 9716 11024
rect 9868 10984 9908 11024
rect 9484 10942 9524 10982
rect 9964 10984 10004 11024
rect 10060 10984 10100 11024
rect 12460 10984 12500 11024
rect 13324 10984 13364 11024
rect 13900 10984 13940 11024
rect 14284 10984 14324 11024
rect 15148 10984 15188 11024
rect 16876 10984 16916 11024
rect 17356 10984 17396 11024
rect 17452 10984 17492 11024
rect 17548 10984 17588 11024
rect 18412 10984 18452 11024
rect 18604 10984 18644 11024
rect 19468 10984 19508 11024
rect 19564 10984 19604 11024
rect 19756 10984 19796 11024
rect 20524 10984 20564 11024
rect 20908 10984 20948 11024
rect 23596 10984 23636 11024
rect 23692 10984 23732 11024
rect 23884 10984 23924 11024
rect 24076 10984 24116 11024
rect 24172 10984 24212 11024
rect 24268 10984 24308 11024
rect 24364 10984 24404 11024
rect 24748 10984 24788 11024
rect 24844 10984 24884 11024
rect 27340 10984 27380 11024
rect 27532 10984 27572 11024
rect 27724 10984 27764 11024
rect 28108 10984 28148 11024
rect 29260 10984 29300 11024
rect 29548 10984 29588 11024
rect 30796 10984 30836 11024
rect 31468 10984 31508 11024
rect 31564 10984 31604 11024
rect 31948 10984 31988 11024
rect 32332 10984 32372 11024
rect 32524 10984 32564 11024
rect 32908 10984 32948 11024
rect 17740 10900 17780 10940
rect 20620 10900 20660 10940
rect 20812 10900 20852 10940
rect 24940 10900 24980 10940
rect 32222 10942 32262 10982
rect 33100 10984 33140 11024
rect 33196 10984 33236 11024
rect 33292 10984 33332 11024
rect 33388 10984 33428 11024
rect 34924 10984 34964 11024
rect 35020 10984 35060 11024
rect 35500 10984 35540 11024
rect 35596 10984 35636 11024
rect 35692 10984 35732 11024
rect 35788 10984 35828 11024
rect 36172 10984 36212 11024
rect 36268 10984 36308 11024
rect 36364 10984 36404 11024
rect 36460 10984 36500 11024
rect 36652 10984 36692 11024
rect 37036 10984 37076 11024
rect 37228 10984 37268 11024
rect 37324 10984 37364 11024
rect 37708 10984 37748 11024
rect 37900 10984 37940 11024
rect 37996 10984 38036 11024
rect 38188 10984 38228 11024
rect 38380 10984 38420 11024
rect 38476 10984 38516 11024
rect 38668 10984 38708 11024
rect 38764 10984 38804 11024
rect 38956 10984 38996 11024
rect 39820 10984 39860 11024
rect 40684 10984 40724 11024
rect 41548 10984 41588 11024
rect 41740 10984 41780 11024
rect 41932 10984 41972 11024
rect 42124 10984 42164 11024
rect 42220 10984 42260 11024
rect 43660 10984 43700 11024
rect 43948 10984 43988 11024
rect 44908 10984 44948 11024
rect 45772 10984 45812 11024
rect 46156 10984 46196 11024
rect 47404 10984 47444 11024
rect 48268 10984 48308 11024
rect 48364 10984 48404 11024
rect 48940 10984 48980 11024
rect 32044 10900 32084 10940
rect 32620 10900 32660 10940
rect 32812 10900 32852 10940
rect 36748 10900 36788 10940
rect 36940 10900 36980 10940
rect 41836 10900 41876 10940
rect 1996 10816 2036 10856
rect 2572 10816 2612 10856
rect 4108 10816 4148 10856
rect 8428 10816 8468 10856
rect 20716 10816 20756 10856
rect 25036 10816 25076 10856
rect 28012 10816 28052 10856
rect 28876 10816 28916 10856
rect 30124 10816 30164 10856
rect 3436 10732 3476 10772
rect 4972 10732 5012 10772
rect 6316 10732 6356 10772
rect 8908 10732 8948 10772
rect 11308 10732 11348 10772
rect 19276 10732 19316 10772
rect 19756 10732 19796 10772
rect 23884 10732 23924 10772
rect 25132 10732 25172 10772
rect 32140 10774 32180 10814
rect 32716 10816 32756 10856
rect 36844 10816 36884 10856
rect 42988 10816 43028 10856
rect 48364 10816 48404 10856
rect 38188 10732 38228 10772
rect 38764 10732 38804 10772
rect 39148 10732 39188 10772
rect 40012 10732 40052 10772
rect 42412 10732 42452 10772
rect 44044 10732 44084 10772
rect 48076 10732 48116 10772
rect 49132 10732 49172 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4204 10396 4244 10436
rect 7468 10396 7508 10436
rect 9580 10396 9620 10436
rect 18220 10396 18260 10436
rect 23980 10396 24020 10436
rect 26284 10396 26324 10436
rect 29356 10396 29396 10436
rect 33484 10396 33524 10436
rect 39148 10396 39188 10436
rect 40204 10396 40244 10436
rect 42892 10396 42932 10436
rect 44236 10396 44276 10436
rect 46348 10396 46388 10436
rect 47020 10396 47060 10436
rect 8236 10312 8276 10352
rect 10252 10312 10292 10352
rect 14092 10312 14132 10352
rect 16012 10312 16052 10352
rect 21196 10312 21236 10352
rect 23020 10312 23060 10352
rect 31564 10312 31604 10352
rect 33100 10312 33140 10352
rect 45292 10312 45332 10352
rect 3916 10228 3956 10268
rect 8332 10228 8372 10268
rect 15436 10228 15476 10268
rect 25036 10228 25076 10268
rect 31468 10228 31508 10268
rect 31660 10228 31700 10268
rect 32812 10228 32852 10268
rect 37708 10228 37748 10268
rect 1516 10144 1556 10184
rect 1900 10144 1940 10184
rect 2764 10144 2804 10184
rect 4876 10144 4916 10184
rect 5068 10144 5108 10184
rect 5452 10144 5492 10184
rect 6316 10144 6356 10184
rect 8428 10144 8468 10184
rect 8524 10144 8564 10184
rect 9100 10144 9140 10184
rect 9196 10144 9236 10184
rect 9580 10144 9620 10184
rect 9868 10144 9908 10184
rect 10540 10144 10580 10184
rect 10636 10144 10676 10184
rect 10732 10144 10772 10184
rect 11596 10144 11636 10184
rect 11980 10144 12020 10184
rect 12172 10144 12212 10184
rect 12268 10144 12308 10184
rect 13132 10144 13172 10184
rect 13324 10144 13364 10184
rect 13420 10144 13460 10184
rect 16300 10144 16340 10184
rect 16588 10144 16628 10184
rect 17260 10144 17300 10184
rect 17740 10144 17780 10184
rect 17932 10144 17972 10184
rect 18028 10144 18068 10184
rect 18604 10144 18644 10184
rect 18892 10144 18932 10184
rect 19660 10144 19700 10184
rect 20236 10144 20276 10184
rect 20332 10144 20372 10184
rect 20428 10144 20468 10184
rect 20524 10144 20564 10184
rect 20716 10144 20756 10184
rect 20908 10144 20948 10184
rect 21004 10144 21044 10184
rect 21868 10144 21908 10184
rect 22060 10144 22100 10184
rect 22156 10144 22196 10184
rect 22252 10144 22292 10184
rect 22348 10144 22388 10184
rect 22732 10144 22772 10184
rect 22924 10144 22964 10184
rect 23020 10144 23060 10184
rect 23212 10144 23252 10184
rect 23308 10144 23348 10184
rect 23500 10144 23540 10184
rect 23596 10144 23636 10184
rect 23697 10144 23737 10184
rect 23980 10144 24020 10184
rect 24076 10144 24116 10184
rect 24268 10144 24308 10184
rect 24364 10144 24404 10184
rect 24521 10159 24561 10199
rect 24844 10144 24884 10184
rect 25132 10144 25172 10184
rect 25420 10144 25460 10184
rect 25516 10144 25556 10184
rect 25612 10144 25652 10184
rect 26668 10144 26708 10184
rect 26956 10144 26996 10184
rect 27724 10144 27764 10184
rect 28012 10144 28052 10184
rect 29452 10144 29492 10184
rect 29644 10144 29684 10184
rect 29836 10144 29876 10184
rect 30220 10144 30260 10184
rect 30412 10144 30452 10184
rect 30700 10144 30740 10184
rect 31372 10144 31412 10184
rect 31756 10144 31796 10184
rect 31982 10151 32022 10191
rect 32140 10144 32180 10184
rect 32236 10144 32276 10184
rect 32428 10144 32468 10184
rect 32524 10144 32564 10184
rect 32716 10144 32756 10184
rect 32908 10144 32948 10184
rect 33100 10144 33140 10184
rect 33292 10144 33332 10184
rect 33580 10144 33620 10184
rect 33868 10144 33908 10184
rect 34156 10144 34196 10184
rect 34348 10144 34388 10184
rect 34540 10144 34580 10184
rect 34636 10144 34676 10184
rect 34828 10144 34868 10184
rect 34924 10144 34964 10184
rect 35020 10144 35060 10184
rect 35308 10144 35348 10184
rect 35404 10144 35444 10184
rect 35596 10159 35636 10199
rect 35692 10144 35732 10184
rect 35793 10144 35833 10184
rect 36268 10144 36308 10184
rect 36364 10144 36404 10184
rect 36556 10144 36596 10184
rect 36748 10144 36788 10184
rect 36844 10144 36884 10184
rect 37132 10144 37172 10184
rect 37228 10144 37268 10184
rect 37324 10144 37364 10184
rect 37516 10144 37556 10184
rect 37804 10144 37844 10184
rect 37996 10144 38036 10184
rect 39820 10144 39860 10184
rect 41356 10144 41396 10184
rect 42220 10144 42260 10184
rect 42604 10144 42644 10184
rect 43180 10144 43220 10184
rect 43276 10144 43316 10184
rect 43564 10144 43604 10184
rect 44428 10144 44468 10184
rect 45292 10144 45332 10184
rect 45484 10144 45524 10184
rect 45676 10144 45716 10184
rect 46636 10144 46676 10184
rect 48172 10144 48212 10184
rect 49036 10144 49076 10184
rect 49420 10144 49460 10184
rect 12076 10060 12116 10100
rect 18508 10060 18548 10100
rect 19372 10060 19412 10100
rect 20812 10060 20852 10100
rect 25324 10060 25364 10100
rect 26572 10060 26612 10100
rect 28204 10060 28244 10100
rect 29740 10060 29780 10100
rect 30508 10060 30548 10100
rect 34060 10060 34100 10100
rect 38668 10060 38708 10100
rect 652 9976 692 10016
rect 8428 9976 8468 10016
rect 9388 9976 9428 10016
rect 10444 9976 10484 10016
rect 10924 9976 10964 10016
rect 12460 9976 12500 10016
rect 17836 9976 17876 10016
rect 19180 9976 19220 10016
rect 23404 9976 23444 10016
rect 29356 9976 29396 10016
rect 32044 9976 32084 10016
rect 35116 9976 35156 10016
rect 35596 9976 35636 10016
rect 36076 9976 36116 10016
rect 36652 9976 36692 10016
rect 37036 9976 37076 10016
rect 43372 9972 43412 10012
rect 45100 9976 45140 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 652 9640 692 9680
rect 5068 9640 5108 9680
rect 7084 9640 7124 9680
rect 9484 9640 9524 9680
rect 9772 9640 9812 9680
rect 12652 9640 12692 9680
rect 16012 9640 16052 9680
rect 16876 9640 16916 9680
rect 21964 9640 22004 9680
rect 24652 9640 24692 9680
rect 25132 9640 25172 9680
rect 27052 9640 27092 9680
rect 30796 9640 30836 9680
rect 37324 9640 37364 9680
rect 44716 9640 44756 9680
rect 48172 9640 48212 9680
rect 9388 9556 9428 9596
rect 10252 9556 10292 9596
rect 16492 9556 16532 9596
rect 23692 9556 23732 9596
rect 27916 9556 27956 9596
rect 29548 9556 29588 9596
rect 30220 9556 30260 9596
rect 1708 9472 1748 9512
rect 1900 9472 1940 9512
rect 2284 9472 2324 9512
rect 2380 9472 2420 9512
rect 3532 9472 3572 9512
rect 4204 9472 4244 9512
rect 4300 9472 4340 9512
rect 4588 9472 4628 9512
rect 4780 9472 4820 9512
rect 4876 9472 4916 9512
rect 5740 9472 5780 9512
rect 5932 9472 5972 9512
rect 6124 9472 6164 9512
rect 6988 9472 7028 9512
rect 7180 9472 7220 9512
rect 7276 9472 7316 9512
rect 7468 9472 7508 9512
rect 7564 9472 7604 9512
rect 8332 9472 8372 9512
rect 9004 9472 9044 9512
rect 9196 9472 9236 9512
rect 9292 9472 9332 9512
rect 9772 9472 9812 9512
rect 9964 9472 10004 9512
rect 10060 9472 10100 9512
rect 10636 9472 10676 9512
rect 11500 9472 11540 9512
rect 13612 9472 13652 9512
rect 13996 9472 14036 9512
rect 14860 9472 14900 9512
rect 16396 9472 16436 9512
rect 16588 9472 16628 9512
rect 16780 9472 16820 9512
rect 16972 9472 17012 9512
rect 17068 9472 17108 9512
rect 17260 9472 17300 9512
rect 17452 9472 17492 9512
rect 17548 9472 17588 9512
rect 17740 9472 17780 9512
rect 17836 9472 17876 9512
rect 18028 9472 18068 9512
rect 18316 9472 18356 9512
rect 19084 9472 19124 9512
rect 20332 9472 20372 9512
rect 20524 9472 20564 9512
rect 20716 9472 20756 9512
rect 20812 9472 20852 9512
rect 21004 9472 21044 9512
rect 21964 9472 22004 9512
rect 22060 9472 22100 9512
rect 22444 9472 22484 9512
rect 22540 9472 22580 9512
rect 22636 9472 22676 9512
rect 22732 9472 22772 9512
rect 23212 9472 23252 9512
rect 23596 9472 23636 9512
rect 23980 9472 24020 9512
rect 24172 9472 24212 9512
rect 24364 9472 24404 9512
rect 24460 9472 24500 9512
rect 24844 9472 24884 9512
rect 24940 9472 24980 9512
rect 25036 9472 25076 9512
rect 25324 9472 25364 9512
rect 25516 9472 25556 9512
rect 26956 9472 26996 9512
rect 27244 9472 27284 9512
rect 27436 9472 27476 9512
rect 27820 9472 27860 9512
rect 28492 9472 28532 9512
rect 28588 9472 28628 9512
rect 29644 9472 29684 9512
rect 29932 9472 29972 9512
rect 30316 9472 30356 9512
rect 30412 9472 30452 9512
rect 30508 9472 30548 9512
rect 30700 9472 30740 9512
rect 30892 9472 30932 9512
rect 31276 9472 31316 9512
rect 31660 9472 31700 9512
rect 31948 9472 31988 9512
rect 34156 9472 34196 9512
rect 34444 9472 34484 9512
rect 34828 9472 34868 9512
rect 34924 9472 34964 9512
rect 35404 9472 35444 9512
rect 35500 9472 35540 9512
rect 35596 9472 35636 9512
rect 35692 9472 35732 9512
rect 35884 9472 35924 9512
rect 36172 9472 36212 9512
rect 37420 9472 37460 9512
rect 38188 9472 38228 9512
rect 38284 9472 38324 9512
rect 38476 9472 38516 9512
rect 38860 9472 38900 9512
rect 39052 9472 39092 9512
rect 39436 9472 39476 9512
rect 40300 9472 40340 9512
rect 41452 9472 41492 9512
rect 42124 9472 42164 9512
rect 42988 9472 43028 9512
rect 43084 9472 43124 9512
rect 43276 9472 43316 9512
rect 44140 9472 44180 9512
rect 44428 9472 44468 9512
rect 44620 9472 44660 9512
rect 44908 9472 44948 9512
rect 45196 9472 45236 9512
rect 46060 9472 46100 9512
rect 47788 9472 47828 9512
rect 48844 9472 48884 9512
rect 2092 9388 2132 9428
rect 7660 9398 7700 9438
rect 21868 9388 21908 9428
rect 28396 9388 28436 9428
rect 31372 9388 31412 9428
rect 31564 9388 31604 9428
rect 35020 9388 35060 9428
rect 38572 9388 38612 9428
rect 38764 9388 38804 9428
rect 41740 9388 41780 9428
rect 47020 9388 47060 9428
rect 1516 9304 1556 9344
rect 4012 9304 4052 9344
rect 4876 9304 4916 9344
rect 7756 9304 7796 9344
rect 9292 9304 9332 9344
rect 18028 9304 18068 9344
rect 18892 9304 18932 9344
rect 21772 9304 21812 9344
rect 22252 9304 22292 9344
rect 28204 9304 28244 9344
rect 28300 9304 28340 9344
rect 29260 9304 29300 9344
rect 31468 9304 31508 9344
rect 32236 9304 32276 9344
rect 34444 9304 34484 9344
rect 35116 9304 35156 9344
rect 35884 9304 35924 9344
rect 38668 9304 38708 9344
rect 43180 9304 43220 9344
rect 1900 9220 1940 9260
rect 2860 9220 2900 9260
rect 5932 9220 5972 9260
rect 7852 9220 7892 9260
rect 17260 9220 17300 9260
rect 20332 9220 20372 9260
rect 21004 9220 21044 9260
rect 24172 9220 24212 9260
rect 25420 9220 25460 9260
rect 32428 9220 32468 9260
rect 35212 9220 35252 9260
rect 42796 9220 42836 9260
rect 43468 9220 43508 9260
rect 45868 9220 45908 9260
rect 46732 9220 46772 9260
rect 48172 9220 48212 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 8908 8884 8948 8924
rect 17164 8884 17204 8924
rect 18316 8884 18356 8924
rect 22828 8884 22868 8924
rect 24940 8884 24980 8924
rect 49036 8884 49076 8924
rect 3724 8800 3764 8840
rect 11404 8800 11444 8840
rect 12172 8800 12212 8840
rect 16492 8800 16532 8840
rect 20428 8800 20468 8840
rect 21964 8800 22004 8840
rect 29260 8800 29300 8840
rect 31564 8800 31604 8840
rect 32236 8800 32276 8840
rect 34060 8800 34100 8840
rect 37900 8800 37940 8840
rect 41068 8800 41108 8840
rect 44332 8800 44372 8840
rect 45772 8800 45812 8840
rect 15628 8716 15668 8756
rect 20332 8716 20372 8756
rect 20524 8716 20564 8756
rect 28492 8716 28532 8756
rect 33772 8716 33812 8756
rect 1036 8632 1076 8672
rect 1420 8632 1460 8672
rect 2284 8632 2324 8672
rect 3436 8632 3476 8672
rect 3724 8632 3764 8672
rect 3916 8632 3956 8672
rect 4108 8632 4148 8672
rect 4492 8632 4532 8672
rect 5356 8632 5396 8672
rect 6604 8632 6644 8672
rect 7468 8632 7508 8672
rect 7660 8632 7700 8672
rect 7756 8632 7796 8672
rect 7948 8632 7988 8672
rect 8236 8632 8276 8672
rect 9676 8632 9716 8672
rect 9868 8632 9908 8672
rect 10444 8632 10484 8672
rect 10540 8632 10580 8672
rect 10636 8632 10676 8672
rect 11404 8632 11444 8672
rect 11596 8632 11636 8672
rect 11692 8632 11732 8672
rect 11980 8632 12020 8672
rect 13420 8632 13460 8672
rect 14380 8632 14420 8672
rect 15532 8632 15572 8672
rect 15724 8632 15764 8672
rect 16012 8632 16052 8672
rect 17164 8632 17204 8672
rect 17356 8632 17396 8672
rect 17548 8632 17588 8672
rect 17740 8632 17780 8672
rect 17836 8632 17876 8672
rect 18316 8632 18356 8672
rect 18508 8632 18548 8672
rect 18700 8632 18740 8672
rect 19756 8632 19796 8672
rect 19852 8632 19892 8672
rect 19948 8632 19988 8672
rect 20044 8632 20084 8672
rect 20236 8632 20276 8672
rect 20620 8632 20660 8672
rect 20908 8632 20948 8672
rect 21004 8632 21044 8672
rect 21100 8632 21140 8672
rect 21388 8632 21428 8672
rect 21484 8632 21524 8672
rect 21580 8632 21620 8672
rect 21868 8632 21908 8672
rect 22060 8632 22100 8672
rect 22732 8632 22772 8672
rect 22919 8611 22959 8651
rect 23116 8632 23156 8672
rect 23308 8632 23348 8672
rect 23404 8632 23444 8672
rect 23788 8632 23828 8672
rect 23884 8632 23924 8672
rect 24076 8632 24116 8672
rect 24172 8632 24212 8672
rect 24268 8632 24308 8672
rect 24364 8632 24404 8672
rect 24556 8632 24596 8672
rect 24748 8632 24788 8672
rect 25036 8632 25076 8672
rect 25708 8632 25748 8672
rect 26284 8632 26324 8672
rect 26380 8632 26420 8672
rect 26476 8632 26516 8672
rect 27239 8632 27279 8672
rect 27340 8632 27380 8672
rect 27436 8632 27476 8672
rect 27628 8632 27668 8672
rect 27724 8632 27764 8672
rect 27916 8628 27956 8668
rect 28012 8632 28052 8672
rect 28115 8628 28155 8668
rect 28211 8637 28251 8677
rect 28396 8632 28436 8672
rect 28588 8632 28628 8672
rect 28972 8632 29012 8672
rect 29164 8632 29204 8672
rect 29356 8632 29396 8672
rect 29548 8632 29588 8672
rect 29644 8632 29684 8672
rect 29740 8632 29780 8672
rect 29836 8632 29876 8672
rect 30065 8632 30105 8672
rect 30220 8632 30260 8672
rect 30316 8632 30356 8672
rect 30508 8632 30548 8672
rect 30604 8632 30644 8672
rect 31660 8632 31700 8672
rect 31948 8632 31988 8672
rect 33580 8632 33620 8672
rect 33868 8632 33908 8672
rect 34348 8632 34388 8672
rect 34444 8632 34484 8672
rect 34732 8632 34772 8672
rect 35020 8632 35060 8672
rect 35596 8632 35636 8672
rect 35692 8632 35732 8672
rect 35788 8632 35828 8672
rect 35980 8632 36020 8672
rect 36076 8632 36116 8672
rect 37612 8632 37652 8672
rect 37900 8632 37940 8672
rect 38764 8632 38804 8672
rect 38956 8632 38996 8672
rect 39820 8632 39860 8672
rect 40012 8632 40052 8672
rect 40876 8632 40916 8672
rect 41164 8632 41204 8672
rect 41644 8632 41684 8672
rect 41740 8632 41780 8672
rect 42604 8632 42644 8672
rect 42796 8632 42836 8672
rect 43660 8632 43700 8672
rect 45196 8632 45236 8672
rect 45484 8632 45524 8672
rect 46444 8632 46484 8672
rect 46636 8632 46676 8672
rect 47020 8632 47060 8672
rect 47884 8632 47924 8672
rect 9100 8548 9140 8588
rect 9772 8548 9812 8588
rect 11884 8548 11924 8588
rect 17644 8548 17684 8588
rect 21676 8548 21716 8588
rect 23212 8548 23252 8588
rect 41548 8548 41588 8588
rect 652 8464 692 8504
rect 6796 8464 6836 8504
rect 7948 8464 7988 8504
rect 10732 8464 10772 8504
rect 18796 8464 18836 8504
rect 21196 8464 21236 8504
rect 23596 8464 23636 8504
rect 24652 8464 24692 8504
rect 25804 8464 25844 8504
rect 26188 8464 26228 8504
rect 27532 8464 27572 8504
rect 28876 8464 28916 8504
rect 30412 8464 30452 8504
rect 34540 8460 34580 8500
rect 35212 8464 35252 8504
rect 35500 8464 35540 8504
rect 36268 8464 36308 8504
rect 38092 8464 38132 8504
rect 39628 8464 39668 8504
rect 39916 8464 39956 8504
rect 40204 8464 40244 8504
rect 41356 8464 41396 8504
rect 41452 8464 41492 8504
rect 41932 8464 41972 8504
rect 43468 8464 43508 8504
rect 44524 8464 44564 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 1516 8128 1556 8168
rect 3724 8128 3764 8168
rect 4876 8128 4916 8168
rect 5548 8128 5588 8168
rect 8140 8128 8180 8168
rect 8236 8128 8276 8168
rect 10828 8128 10868 8168
rect 15916 8128 15956 8168
rect 17356 8128 17396 8168
rect 21196 8128 21236 8168
rect 23500 8128 23540 8168
rect 25228 8128 25268 8168
rect 34924 8128 34964 8168
rect 36364 8128 36404 8168
rect 37804 8128 37844 8168
rect 8044 8044 8084 8084
rect 11116 8044 11156 8084
rect 11692 8044 11732 8084
rect 21580 8044 21620 8084
rect 844 7960 884 8000
rect 1036 7960 1076 8000
rect 1132 7960 1172 8000
rect 1324 7960 1364 8000
rect 1420 7960 1460 8000
rect 1612 7960 1652 8000
rect 2476 7960 2516 8000
rect 3532 7960 3572 8000
rect 4396 7960 4436 8000
rect 4684 7960 4724 8000
rect 5068 7960 5108 8000
rect 5356 7960 5396 8000
rect 5836 7960 5876 8000
rect 6028 7960 6068 8000
rect 7564 7960 7604 8000
rect 7852 7960 7892 8000
rect 7948 7960 7988 8000
rect 9100 7960 9140 8000
rect 9484 7960 9524 8000
rect 9580 7960 9620 8000
rect 9676 7960 9716 8000
rect 9772 7960 9812 8000
rect 9964 7960 10004 8000
rect 10156 7960 10196 8000
rect 10252 7960 10292 8000
rect 10828 7960 10868 8000
rect 10924 7960 10964 8000
rect 12076 7960 12116 8000
rect 12940 7960 12980 8000
rect 15820 7960 15860 8000
rect 16876 7960 16916 8000
rect 17068 7960 17108 8000
rect 17164 7960 17204 8000
rect 17260 7960 17300 8000
rect 17836 7960 17876 8000
rect 17932 7960 17972 8000
rect 20332 7960 20372 8000
rect 20716 7960 20756 8000
rect 20812 7960 20852 8000
rect 21004 7960 21044 8000
rect 21100 7960 21140 8000
rect 21257 7945 21297 7985
rect 21484 7960 21524 8000
rect 21676 7960 21716 8000
rect 22348 7960 22388 8000
rect 22444 7960 22484 8000
rect 22540 7960 22580 8000
rect 22732 7960 22772 8000
rect 22924 7960 22964 8000
rect 23020 7960 23060 8000
rect 23212 7960 23252 8000
rect 23308 7960 23348 8000
rect 23692 7960 23732 8000
rect 23788 7960 23828 8000
rect 23884 7960 23924 8000
rect 23980 7960 24020 8000
rect 24460 7960 24500 8000
rect 24556 7960 24596 8000
rect 24652 7960 24692 8000
rect 24748 7960 24788 8000
rect 24940 7960 24980 8000
rect 25036 7960 25076 8000
rect 25420 7960 25460 8000
rect 25612 7960 25652 8000
rect 25708 7960 25748 8000
rect 25991 7960 26031 8000
rect 26092 7960 26132 8000
rect 26188 7960 26228 8000
rect 26380 7960 26420 8000
rect 26476 7960 26516 8000
rect 27052 7960 27092 8000
rect 27148 7960 27188 8000
rect 27244 7960 27284 8000
rect 27340 7960 27380 8000
rect 27532 7960 27572 8000
rect 29836 7960 29876 8000
rect 29932 7960 29972 8000
rect 30028 7960 30068 8000
rect 30124 7960 30164 8000
rect 31276 7960 31316 8000
rect 31468 7960 31508 8000
rect 31852 7960 31892 8000
rect 32236 7960 32276 8000
rect 34060 7960 34100 8000
rect 34252 7960 34292 8000
rect 34348 7960 34388 8000
rect 34574 7945 34614 7985
rect 34732 7960 34772 8000
rect 34828 7960 34868 8000
rect 35020 7960 35060 8000
rect 35116 7960 35156 8000
rect 35308 7973 35348 8013
rect 35500 7960 35540 8000
rect 35692 7960 35732 8000
rect 35788 7960 35828 8000
rect 35884 7981 35924 8021
rect 35980 7960 36020 8000
rect 36212 7960 36252 8000
rect 36364 7960 36404 8000
rect 36460 7960 36500 8000
rect 36652 7960 36692 8000
rect 36748 7960 36788 8000
rect 36940 7960 36980 8000
rect 37036 7960 37076 8000
rect 37228 7960 37268 8000
rect 37708 7960 37748 8000
rect 37996 7960 38036 8000
rect 38092 7960 38132 8000
rect 38284 7960 38324 8000
rect 38572 7960 38612 8000
rect 38764 7960 38804 8000
rect 38956 7960 38996 8000
rect 40204 7960 40244 8000
rect 41068 7960 41108 8000
rect 41452 7960 41492 8000
rect 41932 7960 41972 8000
rect 43084 7960 43124 8000
rect 43948 7960 43988 8000
rect 44332 7960 44372 8000
rect 44812 7960 44852 8000
rect 46060 7960 46100 8000
rect 46924 7960 46964 8000
rect 47308 7960 47348 8000
rect 17548 7876 17588 7916
rect 18892 7876 18932 7916
rect 31948 7876 31988 7916
rect 32140 7876 32180 7916
rect 1132 7792 1172 7832
rect 4684 7792 4724 7832
rect 6412 7792 6452 7832
rect 10444 7792 10484 7832
rect 14860 7792 14900 7832
rect 20428 7792 20468 7832
rect 23020 7792 23060 7832
rect 25708 7792 25748 7832
rect 31468 7792 31508 7832
rect 32044 7792 32084 7832
rect 34348 7792 34388 7832
rect 36940 7792 36980 7832
rect 38284 7792 38324 7832
rect 1804 7708 1844 7748
rect 2860 7708 2900 7748
rect 3724 7708 3764 7748
rect 5932 7708 5972 7748
rect 7084 7708 7124 7748
rect 8428 7708 8468 7748
rect 14092 7708 14132 7748
rect 16204 7708 16244 7748
rect 19084 7708 19124 7748
rect 26476 7708 26516 7748
rect 27820 7708 27860 7748
rect 35404 7708 35444 7748
rect 37516 7708 37556 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 8812 7372 8852 7412
rect 23596 7372 23636 7412
rect 25036 7372 25076 7412
rect 25228 7372 25268 7412
rect 26380 7372 26420 7412
rect 27724 7372 27764 7412
rect 34252 7372 34292 7412
rect 34444 7372 34484 7412
rect 37612 7372 37652 7412
rect 40108 7372 40148 7412
rect 43276 7372 43316 7412
rect 4012 7288 4052 7328
rect 9388 7288 9428 7328
rect 10252 7288 10292 7328
rect 21196 7288 21236 7328
rect 23212 7288 23252 7328
rect 29644 7288 29684 7328
rect 30220 7288 30260 7328
rect 31372 7288 31412 7328
rect 32428 7288 32468 7328
rect 33004 7288 33044 7328
rect 35116 7288 35156 7328
rect 42892 7288 42932 7328
rect 23116 7204 23156 7244
rect 23308 7204 23348 7244
rect 27340 7204 27380 7244
rect 29548 7204 29588 7244
rect 29740 7204 29780 7244
rect 30124 7204 30164 7244
rect 30316 7204 30356 7244
rect 32332 7204 32372 7244
rect 844 7120 884 7160
rect 1228 7120 1268 7160
rect 2092 7120 2132 7160
rect 3340 7120 3380 7160
rect 3724 7120 3764 7160
rect 3820 7120 3860 7160
rect 4876 7120 4916 7160
rect 5068 7120 5108 7160
rect 6316 7120 6356 7160
rect 7180 7120 7220 7160
rect 8620 7120 8660 7160
rect 8812 7120 8852 7160
rect 9004 7120 9044 7160
rect 9196 7120 9236 7160
rect 9388 7120 9428 7160
rect 9580 7120 9620 7160
rect 9676 7120 9716 7160
rect 11116 7120 11156 7160
rect 12076 7120 12116 7160
rect 13132 7120 13172 7160
rect 13996 7120 14036 7160
rect 14380 7120 14420 7160
rect 14764 7120 14804 7160
rect 15628 7120 15668 7160
rect 16876 7120 16916 7160
rect 17356 7120 17396 7160
rect 17644 7120 17684 7160
rect 18508 7120 18548 7160
rect 18700 7120 18740 7160
rect 18796 7120 18836 7160
rect 18988 7120 19028 7160
rect 20428 7120 20468 7160
rect 20620 7120 20660 7160
rect 20812 7120 20852 7160
rect 21004 7120 21044 7160
rect 21484 7120 21524 7160
rect 21580 7120 21620 7160
rect 22252 7120 22292 7160
rect 22348 7120 22388 7160
rect 22540 7120 22580 7160
rect 22636 7120 22676 7160
rect 23020 7120 23060 7160
rect 23404 7120 23444 7160
rect 23596 7120 23636 7160
rect 23692 7120 23732 7160
rect 23884 7120 23924 7160
rect 23980 7120 24020 7160
rect 24081 7120 24121 7160
rect 24364 7120 24404 7160
rect 24460 7120 24500 7160
rect 24556 7120 24596 7160
rect 24652 7120 24692 7160
rect 24844 7120 24884 7160
rect 25036 7120 25076 7160
rect 25324 7120 25364 7160
rect 26380 7120 26420 7160
rect 26572 7120 26612 7160
rect 27148 7120 27188 7160
rect 27436 7120 27476 7160
rect 27628 7120 27668 7160
rect 27820 7120 27860 7160
rect 29068 7120 29108 7160
rect 29260 7120 29300 7160
rect 29452 7120 29492 7160
rect 29836 7120 29876 7160
rect 30028 7120 30068 7160
rect 30412 7120 30452 7160
rect 30700 7162 30740 7202
rect 32524 7204 32564 7244
rect 32908 7204 32948 7244
rect 33100 7204 33140 7244
rect 35020 7204 35060 7244
rect 35212 7204 35252 7244
rect 35692 7204 35732 7244
rect 40588 7204 40628 7244
rect 30604 7120 30644 7160
rect 30796 7120 30836 7160
rect 30892 7120 30932 7160
rect 31660 7120 31700 7160
rect 31756 7120 31796 7160
rect 32236 7120 32276 7160
rect 32620 7120 32660 7160
rect 32812 7120 32852 7160
rect 33196 7120 33236 7160
rect 34156 7120 34196 7160
rect 34444 7120 34484 7160
rect 34636 7120 34676 7160
rect 34924 7120 34964 7160
rect 35308 7120 35348 7160
rect 35884 7120 35924 7160
rect 36844 7120 36884 7160
rect 37324 7120 37364 7160
rect 37420 7120 37460 7160
rect 37612 7120 37652 7160
rect 37804 7120 37844 7160
rect 37996 7120 38036 7160
rect 38092 7120 38132 7160
rect 38476 7120 38516 7160
rect 39436 7120 39476 7160
rect 40396 7120 40436 7160
rect 41260 7120 41300 7160
rect 41452 7120 41492 7160
rect 41836 7120 41876 7160
rect 42220 7120 42260 7160
rect 43180 7120 43220 7160
rect 43276 7120 43316 7160
rect 43756 7120 43796 7160
rect 44620 7120 44660 7160
rect 46252 7120 46292 7160
rect 46636 7120 46676 7160
rect 47020 7120 47060 7160
rect 5932 7036 5972 7076
rect 9100 7036 9140 7076
rect 41932 7036 41972 7076
rect 43372 7036 43412 7076
rect 46540 7036 46580 7076
rect 3724 6952 3764 6992
rect 4204 6952 4244 6992
rect 5740 6952 5780 6992
rect 8332 6952 8372 6992
rect 10444 6952 10484 6992
rect 11404 6952 11444 6992
rect 17164 6952 17204 6992
rect 17836 6952 17876 6992
rect 18892 6952 18932 6992
rect 20524 6952 20564 6992
rect 21676 6948 21716 6988
rect 22828 6952 22868 6992
rect 31852 6948 31892 6988
rect 36364 6952 36404 6992
rect 37612 6952 37652 6992
rect 38092 6952 38132 6992
rect 39148 6952 39188 6992
rect 43468 6952 43508 6992
rect 44428 6952 44468 6992
rect 45292 6952 45332 6992
rect 45580 6952 45620 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 652 6616 692 6656
rect 7756 6616 7796 6656
rect 8332 6616 8372 6656
rect 9484 6616 9524 6656
rect 10156 6616 10196 6656
rect 12844 6616 12884 6656
rect 18220 6616 18260 6656
rect 30124 6616 30164 6656
rect 33196 6616 33236 6656
rect 34060 6616 34100 6656
rect 34636 6616 34676 6656
rect 35308 6616 35348 6656
rect 36076 6616 36116 6656
rect 10444 6532 10484 6572
rect 18124 6532 18164 6572
rect 2188 6448 2228 6488
rect 2380 6448 2420 6488
rect 2764 6448 2804 6488
rect 2860 6448 2900 6488
rect 3628 6448 3668 6488
rect 4492 6448 4532 6488
rect 5164 6448 5204 6488
rect 5452 6448 5492 6488
rect 5548 6448 5588 6488
rect 5740 6448 5780 6488
rect 6604 6448 6644 6488
rect 6796 6448 6836 6488
rect 7084 6448 7124 6488
rect 7276 6448 7316 6488
rect 7468 6448 7508 6488
rect 7564 6448 7604 6488
rect 8236 6448 8276 6488
rect 8428 6448 8468 6488
rect 8620 6448 8660 6488
rect 8812 6448 8852 6488
rect 9004 6448 9044 6488
rect 9196 6448 9236 6488
rect 9388 6448 9428 6488
rect 9772 6448 9812 6488
rect 9964 6448 10004 6488
rect 10060 6448 10100 6488
rect 10252 6448 10292 6488
rect 10828 6448 10868 6488
rect 11692 6448 11732 6488
rect 13612 6448 13652 6488
rect 13900 6448 13940 6488
rect 15532 6448 15572 6488
rect 16396 6448 16436 6488
rect 16780 6448 16820 6488
rect 17452 6448 17492 6488
rect 17932 6448 17972 6488
rect 18892 6490 18932 6530
rect 18028 6448 18068 6488
rect 18796 6448 18836 6488
rect 19084 6448 19124 6488
rect 19276 6448 19316 6488
rect 19372 6448 19412 6488
rect 19468 6448 19508 6488
rect 19564 6448 19604 6488
rect 19756 6448 19796 6488
rect 19852 6448 19892 6488
rect 19948 6448 19988 6488
rect 22924 6490 22964 6530
rect 31372 6532 31412 6572
rect 35596 6532 35636 6572
rect 38764 6532 38804 6572
rect 20044 6448 20084 6488
rect 22540 6448 22580 6488
rect 23116 6448 23156 6488
rect 23500 6448 23540 6488
rect 23692 6448 23732 6488
rect 24076 6448 24116 6488
rect 24268 6448 24308 6488
rect 24460 6448 24500 6488
rect 27244 6448 27284 6488
rect 27628 6448 27668 6488
rect 28204 6448 28244 6488
rect 28396 6448 28436 6488
rect 28588 6448 28628 6488
rect 28780 6448 28820 6488
rect 28972 6448 29012 6488
rect 29164 6448 29204 6488
rect 29260 6448 29300 6488
rect 29452 6448 29492 6488
rect 29644 6448 29684 6488
rect 29836 6448 29876 6488
rect 29932 6448 29972 6488
rect 31276 6448 31316 6488
rect 31468 6448 31508 6488
rect 31660 6448 31700 6488
rect 31852 6448 31892 6488
rect 32044 6448 32084 6488
rect 32428 6448 32468 6488
rect 32716 6448 32756 6488
rect 33868 6448 33908 6488
rect 34156 6448 34196 6488
rect 34348 6448 34388 6488
rect 35020 6448 35060 6488
rect 35116 6448 35156 6488
rect 35404 6448 35444 6488
rect 35788 6448 35828 6488
rect 35884 6448 35924 6488
rect 36076 6448 36116 6488
rect 36268 6448 36308 6488
rect 37132 6448 37172 6488
rect 37708 6448 37748 6488
rect 37804 6448 37844 6488
rect 37900 6448 37940 6488
rect 37996 6448 38036 6488
rect 38284 6448 38324 6488
rect 38572 6448 38612 6488
rect 39244 6448 39284 6488
rect 39628 6448 39668 6488
rect 40492 6448 40532 6488
rect 41644 6448 41684 6488
rect 43180 6448 43220 6488
rect 44044 6448 44084 6488
rect 44428 6448 44468 6488
rect 44716 6448 44756 6488
rect 45868 6448 45908 6488
rect 46732 6448 46772 6488
rect 47116 6448 47156 6488
rect 2284 6364 2324 6404
rect 2572 6364 2612 6404
rect 22636 6364 22676 6404
rect 22828 6364 22868 6404
rect 23212 6364 23252 6404
rect 23404 6364 23444 6404
rect 23788 6364 23828 6404
rect 23980 6364 24020 6404
rect 27340 6364 27380 6404
rect 27532 6364 27572 6404
rect 29548 6364 29588 6404
rect 32140 6364 32180 6404
rect 32332 6364 32372 6404
rect 42028 6364 42068 6404
rect 1324 6280 1364 6320
rect 5740 6280 5780 6320
rect 8812 6280 8852 6320
rect 9100 6280 9140 6320
rect 9676 6280 9716 6320
rect 14092 6280 14132 6320
rect 16204 6280 16244 6320
rect 19084 6280 19124 6320
rect 22732 6280 22772 6320
rect 23308 6280 23348 6320
rect 23884 6280 23924 6320
rect 27436 6280 27476 6320
rect 4300 6196 4340 6236
rect 5932 6196 5972 6236
rect 7180 6196 7220 6236
rect 13612 6196 13652 6236
rect 18220 6196 18260 6236
rect 24268 6196 24308 6236
rect 28204 6196 28244 6236
rect 28588 6196 28628 6236
rect 28972 6196 29012 6236
rect 31756 6196 31796 6236
rect 32236 6238 32276 6278
rect 36940 6196 36980 6236
rect 37228 6196 37268 6236
rect 37516 6196 37556 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 6796 5860 6836 5900
rect 8908 5860 8948 5900
rect 15820 5860 15860 5900
rect 17068 5860 17108 5900
rect 22060 5860 22100 5900
rect 27148 5860 27188 5900
rect 34540 5860 34580 5900
rect 2284 5776 2324 5816
rect 21388 5776 21428 5816
rect 31564 5776 31604 5816
rect 32236 5776 32276 5816
rect 36364 5776 36404 5816
rect 37132 5776 37172 5816
rect 3628 5692 3668 5732
rect 24844 5692 24884 5732
rect 35788 5692 35828 5732
rect 37036 5692 37076 5732
rect 37228 5692 37268 5732
rect 3532 5608 3572 5648
rect 3724 5608 3764 5648
rect 3916 5608 3956 5648
rect 4012 5608 4052 5648
rect 4204 5608 4244 5648
rect 4396 5608 4436 5648
rect 4780 5608 4820 5648
rect 5644 5608 5684 5648
rect 7372 5608 7412 5648
rect 7468 5608 7508 5648
rect 7660 5608 7700 5648
rect 7756 5608 7796 5648
rect 8140 5608 8180 5648
rect 8236 5608 8276 5648
rect 8908 5608 8948 5648
rect 9004 5608 9044 5648
rect 9196 5608 9236 5648
rect 9292 5608 9332 5648
rect 9393 5608 9433 5648
rect 9676 5608 9716 5648
rect 9868 5608 9908 5648
rect 11884 5608 11924 5648
rect 11980 5608 12020 5648
rect 12076 5608 12116 5648
rect 12172 5608 12212 5648
rect 12940 5608 12980 5648
rect 13036 5608 13076 5648
rect 13132 5608 13172 5648
rect 13228 5608 13268 5648
rect 13420 5608 13460 5648
rect 13804 5608 13844 5648
rect 14668 5608 14708 5648
rect 16108 5608 16148 5648
rect 16204 5608 16244 5648
rect 16396 5608 16436 5648
rect 16588 5608 16628 5648
rect 16684 5608 16724 5648
rect 16780 5608 16820 5648
rect 16876 5608 16916 5648
rect 17068 5608 17108 5648
rect 17260 5608 17300 5648
rect 17356 5608 17396 5648
rect 17836 5608 17876 5648
rect 17932 5608 17972 5648
rect 18796 5608 18836 5648
rect 18892 5608 18932 5648
rect 19372 5608 19412 5648
rect 19660 5608 19700 5648
rect 19948 5608 19988 5648
rect 20140 5608 20180 5648
rect 20716 5608 20756 5648
rect 20812 5608 20852 5648
rect 21292 5608 21332 5648
rect 21484 5608 21524 5648
rect 22348 5608 22388 5648
rect 22444 5608 22484 5648
rect 23020 5608 23060 5648
rect 23212 5608 23252 5648
rect 23308 5608 23348 5648
rect 23500 5608 23540 5648
rect 23596 5608 23636 5648
rect 23788 5608 23828 5648
rect 23980 5608 24020 5648
rect 24076 5608 24116 5648
rect 24172 5608 24212 5648
rect 24364 5608 24404 5648
rect 24556 5608 24596 5648
rect 24748 5608 24788 5648
rect 24940 5608 24980 5648
rect 26285 5593 26325 5633
rect 26380 5594 26420 5634
rect 26572 5608 26612 5648
rect 26860 5608 26900 5648
rect 27820 5608 27860 5648
rect 28204 5608 28244 5648
rect 28396 5608 28436 5648
rect 28492 5608 28532 5648
rect 28876 5608 28916 5648
rect 28972 5608 29012 5648
rect 29644 5608 29684 5648
rect 29740 5608 29780 5648
rect 29836 5608 29876 5648
rect 31084 5608 31124 5648
rect 31372 5608 31412 5648
rect 31852 5608 31892 5648
rect 31948 5608 31988 5648
rect 32524 5608 32564 5648
rect 32620 5608 32660 5648
rect 32908 5608 32948 5648
rect 33004 5608 33044 5648
rect 33100 5608 33140 5648
rect 33292 5608 33332 5648
rect 33484 5608 33524 5648
rect 34444 5608 34484 5648
rect 34732 5608 34772 5648
rect 34828 5608 34868 5648
rect 34924 5608 34964 5648
rect 35404 5608 35444 5648
rect 35500 5608 35540 5648
rect 36652 5608 36692 5648
rect 36940 5608 36980 5648
rect 37324 5608 37364 5648
rect 37612 5608 37652 5648
rect 38572 5608 38612 5648
rect 38668 5608 38708 5648
rect 39532 5608 39572 5648
rect 40492 5608 40532 5648
rect 40684 5608 40724 5648
rect 40876 5608 40916 5648
rect 40972 5608 41012 5648
rect 42220 5608 42260 5648
rect 42412 5608 42452 5648
rect 42604 5608 42644 5648
rect 42700 5608 42740 5648
rect 42892 5608 42932 5648
rect 43948 5608 43988 5648
rect 44236 5608 44276 5648
rect 44716 5608 44756 5648
rect 44908 5608 44948 5648
rect 45004 5608 45044 5648
rect 8332 5524 8372 5564
rect 16300 5524 16340 5564
rect 18700 5524 18740 5564
rect 19180 5524 19220 5564
rect 20524 5524 20564 5564
rect 38860 5524 38900 5564
rect 40780 5524 40820 5564
rect 42796 5524 42836 5564
rect 44428 5524 44468 5564
rect 44812 5524 44852 5564
rect 652 5440 692 5480
rect 1036 5440 1076 5480
rect 4204 5440 4244 5480
rect 7180 5440 7220 5480
rect 7948 5440 7988 5480
rect 8428 5440 8468 5480
rect 8524 5440 8564 5480
rect 9772 5440 9812 5480
rect 17548 5440 17588 5480
rect 18508 5440 18548 5480
rect 18604 5440 18644 5480
rect 20812 5440 20852 5480
rect 22540 5436 22580 5476
rect 23116 5440 23156 5480
rect 23692 5440 23732 5480
rect 24460 5440 24500 5480
rect 26476 5440 26516 5480
rect 28300 5440 28340 5480
rect 29260 5440 29300 5480
rect 29932 5440 29972 5480
rect 31276 5440 31316 5480
rect 32044 5436 32084 5476
rect 32716 5436 32756 5476
rect 33388 5440 33428 5480
rect 35020 5440 35060 5480
rect 35212 5440 35252 5480
rect 38284 5440 38324 5480
rect 39820 5440 39860 5480
rect 42316 5440 42356 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 652 5104 692 5144
rect 7948 5104 7988 5144
rect 8716 5104 8756 5144
rect 9676 5108 9716 5148
rect 12076 5104 12116 5144
rect 21484 5104 21524 5144
rect 24268 5104 24308 5144
rect 27052 5104 27092 5144
rect 29260 5104 29300 5144
rect 30220 5104 30260 5144
rect 30316 5104 30356 5144
rect 30892 5104 30932 5144
rect 4780 5020 4820 5060
rect 5164 5020 5204 5060
rect 16012 5020 16052 5060
rect 16396 5020 16436 5060
rect 21580 5020 21620 5060
rect 23884 5020 23924 5060
rect 24364 5020 24404 5060
rect 28780 5020 28820 5060
rect 30412 5020 30452 5060
rect 30988 5020 31028 5060
rect 1708 4936 1748 4976
rect 2092 4936 2132 4976
rect 2956 4936 2996 4976
rect 4204 4936 4244 4976
rect 4588 4936 4628 4976
rect 4684 4936 4724 4976
rect 4876 4936 4916 4976
rect 5068 4936 5108 4976
rect 5260 4936 5300 4976
rect 6604 4936 6644 4976
rect 7468 4936 7508 4976
rect 7660 4936 7700 4976
rect 7756 4936 7796 4976
rect 8620 4936 8660 4976
rect 8716 4936 8756 4976
rect 9484 4936 9524 4976
rect 9580 4936 9620 4976
rect 9868 4936 9908 4976
rect 10060 4936 10100 4976
rect 10156 4936 10196 4976
rect 10348 4936 10388 4976
rect 10540 4936 10580 4976
rect 11596 4936 11636 4976
rect 14668 4936 14708 4976
rect 15916 4936 15956 4976
rect 16108 4936 16148 4976
rect 17260 4936 17300 4976
rect 17548 4936 17588 4976
rect 17740 4936 17780 4976
rect 17836 4936 17876 4976
rect 18028 4936 18068 4976
rect 19084 4936 19124 4976
rect 19180 4936 19220 4976
rect 19276 4936 19316 4976
rect 19372 4936 19412 4976
rect 20044 4936 20084 4976
rect 20236 4936 20276 4976
rect 20428 4936 20468 4976
rect 20524 4936 20564 4976
rect 20620 4936 20660 4976
rect 20716 4936 20756 4976
rect 21676 4936 21716 4976
rect 21772 4936 21812 4976
rect 22732 4936 22772 4976
rect 22924 4936 22964 4976
rect 23116 4936 23156 4976
rect 23308 4936 23348 4976
rect 23404 4936 23444 4976
rect 23692 4936 23732 4976
rect 23788 4936 23828 4976
rect 23980 4936 24020 4976
rect 24460 4936 24500 4976
rect 24556 4936 24596 4976
rect 24748 4936 24788 4976
rect 25036 4936 25076 4976
rect 26092 4936 26132 4976
rect 26188 4936 26228 4976
rect 26284 4936 26324 4976
rect 26380 4936 26420 4976
rect 26572 4936 26612 4976
rect 26668 4936 26708 4976
rect 26764 4936 26804 4976
rect 26860 4936 26900 4976
rect 27244 4936 27284 4976
rect 27340 4936 27380 4976
rect 27532 4936 27572 4976
rect 27916 4936 27956 4976
rect 28684 4936 28724 4976
rect 28876 4936 28916 4976
rect 28972 4936 29012 4976
rect 29164 4936 29204 4976
rect 29356 4936 29396 4976
rect 29452 4936 29492 4976
rect 29644 4936 29684 4976
rect 29740 4936 29780 4976
rect 29836 4936 29876 4976
rect 29932 4936 29972 4976
rect 30508 4936 30548 4976
rect 30604 4936 30644 4976
rect 31084 4936 31124 4976
rect 31180 4936 31220 4976
rect 31564 4936 31604 4976
rect 32620 4936 32660 4976
rect 32716 4936 32756 4976
rect 32908 4936 32948 4976
rect 34252 4936 34292 4976
rect 35116 4936 35156 4976
rect 35308 4936 35348 4976
rect 36556 4936 36596 4976
rect 37420 4936 37460 4976
rect 37804 4936 37844 4976
rect 38188 4936 38228 4976
rect 38380 4936 38420 4976
rect 39244 4936 39284 4976
rect 39628 4936 39668 4976
rect 40492 4936 40532 4976
rect 41644 4936 41684 4976
rect 8812 4852 8852 4892
rect 10444 4852 10484 4892
rect 8908 4810 8948 4850
rect 20140 4852 20180 4892
rect 28108 4852 28148 4892
rect 33868 4852 33908 4892
rect 5452 4768 5492 4808
rect 9196 4768 9236 4808
rect 12748 4768 12788 4808
rect 15052 4768 15092 4808
rect 24460 4768 24500 4808
rect 27628 4768 27668 4808
rect 33676 4768 33716 4808
rect 5932 4684 5972 4724
rect 6796 4684 6836 4724
rect 9868 4684 9908 4724
rect 11884 4684 11924 4724
rect 13996 4684 14036 4724
rect 17548 4684 17588 4724
rect 18700 4684 18740 4724
rect 21676 4684 21716 4724
rect 22732 4684 22772 4724
rect 23116 4684 23156 4724
rect 25036 4684 25076 4724
rect 31084 4684 31124 4724
rect 31948 4684 31988 4724
rect 32908 4684 32948 4724
rect 34444 4684 34484 4724
rect 38092 4684 38132 4724
rect 39052 4684 39092 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 14188 4348 14228 4388
rect 23500 4348 23540 4388
rect 24556 4348 24596 4388
rect 26380 4348 26420 4388
rect 34252 4348 34292 4388
rect 40780 4348 40820 4388
rect 9196 4264 9236 4304
rect 13132 4264 13172 4304
rect 22252 4264 22292 4304
rect 26668 4264 26708 4304
rect 27628 4264 27668 4304
rect 28300 4264 28340 4304
rect 9580 4180 9620 4220
rect 18316 4180 18356 4220
rect 22924 4180 22964 4220
rect 34540 4180 34580 4220
rect 4300 4096 4340 4136
rect 4684 4096 4724 4136
rect 5548 4096 5588 4136
rect 7660 4096 7700 4136
rect 7948 4096 7988 4136
rect 8140 4096 8180 4136
rect 8812 4096 8852 4136
rect 9388 4096 9428 4136
rect 9676 4096 9716 4136
rect 9868 4096 9908 4136
rect 9964 4096 10004 4136
rect 10156 4096 10196 4136
rect 10348 4096 10388 4136
rect 10444 4096 10484 4136
rect 10540 4096 10580 4136
rect 10636 4096 10676 4136
rect 10924 4096 10964 4136
rect 11020 4096 11060 4136
rect 11116 4096 11156 4136
rect 11404 4096 11444 4136
rect 11500 4096 11540 4136
rect 11596 4096 11636 4136
rect 11788 4096 11828 4136
rect 11884 4096 11924 4136
rect 11980 4096 12020 4136
rect 12076 4096 12116 4136
rect 12940 4096 12980 4136
rect 13132 4096 13172 4136
rect 13324 4096 13364 4136
rect 13420 4096 13460 4136
rect 13612 4096 13652 4136
rect 13804 4096 13844 4136
rect 15340 4096 15380 4136
rect 16204 4096 16244 4136
rect 16588 4096 16628 4136
rect 16972 4096 17012 4136
rect 17068 4096 17108 4136
rect 17164 4096 17204 4136
rect 17260 4096 17300 4136
rect 17644 4096 17684 4136
rect 17740 4096 17780 4136
rect 17932 4096 17972 4136
rect 18124 4096 18164 4136
rect 18412 4096 18452 4136
rect 18604 4096 18644 4136
rect 18700 4096 18740 4136
rect 18796 4096 18836 4136
rect 18892 4096 18932 4136
rect 19372 4096 19412 4136
rect 20332 4096 20372 4136
rect 20812 4096 20852 4136
rect 20908 4096 20948 4136
rect 23788 4096 23828 4136
rect 24172 4096 24212 4136
rect 24268 4096 24308 4136
rect 25132 4096 25172 4136
rect 25228 4096 25268 4136
rect 25324 4096 25364 4136
rect 25420 4096 25460 4136
rect 25612 4096 25652 4136
rect 25804 4096 25844 4136
rect 25900 4096 25940 4136
rect 26092 4096 26132 4136
rect 26188 4096 26228 4136
rect 26380 4096 26420 4136
rect 26764 4096 26804 4136
rect 26860 4096 26900 4136
rect 27340 4096 27380 4136
rect 27532 4096 27572 4136
rect 27628 4096 27668 4136
rect 27820 4096 27860 4136
rect 27916 4096 27956 4136
rect 28108 4096 28148 4136
rect 28588 4096 28628 4136
rect 28684 4096 28724 4136
rect 29260 4096 29300 4136
rect 29548 4096 29588 4136
rect 31372 4096 31412 4136
rect 31468 4096 31508 4136
rect 31564 4096 31604 4136
rect 31660 4096 31700 4136
rect 31852 4096 31892 4136
rect 32236 4096 32276 4136
rect 33100 4096 33140 4136
rect 35308 4096 35348 4136
rect 35884 4096 35924 4136
rect 36268 4096 36308 4136
rect 36652 4096 36692 4136
rect 37324 4096 37364 4136
rect 37516 4096 37556 4136
rect 38188 4096 38228 4136
rect 38380 4096 38420 4136
rect 38764 4096 38804 4136
rect 39628 4096 39668 4136
rect 28012 4012 28052 4052
rect 36364 4012 36404 4052
rect 652 3928 692 3968
rect 6700 3928 6740 3968
rect 6988 3928 7028 3968
rect 7852 3928 7892 3968
rect 10060 3928 10100 3968
rect 10828 3928 10868 3968
rect 11308 3928 11348 3968
rect 12268 3928 12308 3968
rect 17836 3928 17876 3968
rect 20620 3928 20660 3968
rect 24076 3924 24116 3964
rect 25708 3928 25748 3968
rect 29068 3928 29108 3968
rect 34252 3928 34292 3968
rect 28780 3870 28820 3910
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 652 3592 692 3632
rect 7756 3592 7796 3632
rect 8140 3592 8180 3632
rect 8812 3592 8852 3632
rect 10156 3592 10196 3632
rect 14092 3592 14132 3632
rect 15820 3592 15860 3632
rect 16780 3592 16820 3632
rect 17548 3592 17588 3632
rect 17740 3592 17780 3632
rect 20620 3592 20660 3632
rect 23788 3592 23828 3632
rect 23980 3592 24020 3632
rect 25516 3592 25556 3632
rect 28588 3592 28628 3632
rect 28876 3592 28916 3632
rect 29164 3592 29204 3632
rect 32908 3592 32948 3632
rect 35020 3592 35060 3632
rect 5356 3508 5396 3548
rect 11692 3508 11732 3548
rect 17068 3508 17108 3548
rect 19756 3508 19796 3548
rect 29260 3508 29300 3548
rect 29740 3508 29780 3548
rect 35308 3508 35348 3548
rect 5740 3424 5780 3464
rect 6604 3424 6644 3464
rect 7948 3424 7988 3464
rect 8044 3424 8084 3464
rect 8236 3424 8276 3464
rect 8716 3424 8756 3464
rect 8908 3424 8948 3464
rect 9004 3424 9044 3464
rect 9196 3424 9236 3464
rect 9868 3424 9908 3464
rect 10060 3424 10100 3464
rect 11308 3424 11348 3464
rect 12076 3424 12116 3464
rect 12940 3424 12980 3464
rect 15916 3424 15956 3464
rect 16300 3424 16340 3464
rect 16396 3424 16436 3464
rect 16492 3424 16532 3464
rect 16588 3424 16628 3464
rect 16876 3424 16916 3464
rect 17260 3424 17300 3464
rect 17356 3424 17396 3464
rect 17452 3424 17492 3464
rect 17836 3424 17876 3464
rect 17932 3424 17972 3464
rect 18028 3424 18068 3464
rect 19276 3424 19316 3464
rect 19564 3424 19604 3464
rect 20332 3424 20372 3464
rect 20428 3424 20468 3464
rect 20524 3424 20564 3464
rect 20812 3424 20852 3464
rect 20908 3424 20948 3464
rect 21004 3424 21044 3464
rect 21100 3424 21140 3464
rect 21292 3424 21332 3464
rect 21388 3424 21428 3464
rect 21484 3424 21524 3464
rect 21580 3424 21620 3464
rect 22444 3424 22484 3464
rect 22636 3424 22676 3464
rect 22732 3424 22772 3464
rect 22924 3424 22964 3464
rect 23500 3424 23540 3464
rect 23596 3424 23636 3464
rect 23692 3424 23732 3464
rect 24076 3424 24116 3464
rect 24172 3424 24212 3464
rect 24268 3424 24308 3464
rect 24460 3424 24500 3464
rect 26380 3424 26420 3464
rect 26764 3424 26804 3464
rect 27436 3424 27476 3464
rect 27628 3424 27668 3464
rect 27820 3424 27860 3464
rect 27916 3424 27956 3464
rect 28108 3424 28148 3464
rect 28204 3424 28244 3464
rect 28300 3424 28340 3464
rect 28396 3424 28436 3464
rect 28684 3424 28724 3464
rect 29356 3424 29396 3464
rect 29452 3424 29492 3464
rect 29644 3424 29684 3464
rect 29836 3424 29876 3464
rect 31276 3424 31316 3464
rect 31372 3424 31412 3464
rect 31468 3424 31508 3464
rect 31564 3424 31604 3464
rect 31756 3424 31796 3464
rect 32044 3424 32084 3464
rect 33580 3424 33620 3464
rect 34348 3424 34388 3464
rect 36172 3424 36212 3464
rect 37228 3424 37268 3464
rect 38380 3424 38420 3464
rect 39244 3424 39284 3464
rect 39628 3424 39668 3464
rect 25324 3340 25364 3380
rect 4780 3256 4820 3296
rect 32332 3256 32372 3296
rect 33772 3256 33812 3296
rect 10636 3172 10676 3212
rect 16108 3172 16148 3212
rect 21772 3172 21812 3212
rect 22924 3172 22964 3212
rect 25132 3172 25172 3212
rect 25708 3172 25748 3212
rect 27628 3172 27668 3212
rect 29164 3172 29204 3212
rect 32044 3172 32084 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 7372 2836 7412 2876
rect 8236 2836 8276 2876
rect 16300 2836 16340 2876
rect 16780 2836 16820 2876
rect 20428 2836 20468 2876
rect 24172 2836 24212 2876
rect 25132 2836 25172 2876
rect 26572 2836 26612 2876
rect 27052 2836 27092 2876
rect 35692 2836 35732 2876
rect 36652 2836 36692 2876
rect 37996 2836 38036 2876
rect 5836 2752 5876 2792
rect 32428 2752 32468 2792
rect 844 2668 884 2708
rect 20620 2668 20660 2708
rect 7084 2584 7124 2624
rect 7180 2584 7220 2624
rect 7372 2584 7412 2624
rect 7564 2584 7604 2624
rect 7660 2584 7700 2624
rect 9388 2584 9428 2624
rect 10252 2584 10292 2624
rect 10636 2584 10676 2624
rect 15820 2584 15860 2624
rect 15916 2584 15956 2624
rect 16012 2584 16052 2624
rect 16108 2584 16148 2624
rect 16300 2584 16340 2624
rect 16492 2584 16532 2624
rect 16588 2584 16628 2624
rect 16972 2584 17012 2624
rect 17068 2584 17108 2624
rect 17164 2586 17204 2626
rect 17356 2584 17396 2624
rect 17548 2584 17588 2624
rect 17836 2584 17876 2624
rect 18316 2584 18356 2624
rect 18412 2584 18452 2624
rect 18508 2584 18548 2624
rect 19276 2584 19316 2624
rect 19372 2584 19412 2624
rect 19468 2584 19508 2624
rect 19852 2584 19892 2624
rect 19948 2584 19988 2624
rect 20140 2584 20180 2624
rect 20236 2584 20276 2624
rect 20428 2584 20468 2624
rect 21292 2584 21332 2624
rect 21772 2584 21812 2624
rect 22156 2584 22196 2624
rect 23020 2584 23060 2624
rect 25324 2584 25364 2624
rect 25900 2584 25940 2624
rect 27148 2584 27188 2624
rect 27532 2584 27572 2624
rect 27916 2584 27956 2624
rect 28108 2584 28148 2624
rect 28492 2584 28532 2624
rect 29164 2584 29204 2624
rect 29356 2584 29396 2624
rect 29452 2584 29492 2624
rect 29644 2584 29684 2624
rect 29740 2584 29780 2624
rect 29836 2584 29876 2624
rect 29932 2584 29972 2624
rect 30316 2584 30356 2624
rect 31276 2584 31316 2624
rect 31564 2584 31604 2624
rect 32236 2551 32276 2591
rect 33292 2584 33332 2624
rect 33676 2584 33716 2624
rect 34540 2584 34580 2624
rect 35980 2584 36020 2624
rect 37516 2584 37556 2624
rect 37612 2584 37652 2624
rect 37804 2584 37844 2624
rect 37996 2584 38036 2624
rect 38188 2584 38228 2624
rect 38284 2584 38324 2624
rect 18028 2500 18068 2540
rect 18604 2500 18644 2540
rect 27436 2500 27476 2540
rect 28588 2500 28628 2540
rect 37708 2500 37748 2540
rect 652 2416 692 2456
rect 19180 2416 19220 2456
rect 19660 2416 19700 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 17452 2080 17492 2120
rect 21772 2080 21812 2120
rect 22540 1996 22580 2036
rect 22924 1996 22964 2036
rect 16300 1912 16340 1952
rect 16492 1912 16532 1952
rect 16876 1912 16916 1952
rect 16972 1922 17012 1962
rect 17548 1912 17588 1952
rect 17644 1912 17684 1952
rect 17740 1912 17780 1952
rect 17932 1912 17972 1952
rect 18028 1912 18068 1952
rect 18220 1912 18260 1952
rect 18988 1912 19028 1952
rect 19372 1912 19412 1952
rect 20236 1912 20276 1952
rect 21484 1912 21524 1952
rect 21676 1912 21716 1952
rect 21964 1912 22004 1952
rect 22444 1912 22484 1952
rect 22636 1912 22676 1952
rect 23308 1912 23348 1952
rect 24172 1912 24212 1952
rect 25612 1912 25652 1952
rect 25996 1912 26036 1952
rect 26860 1912 26900 1952
rect 28012 1912 28052 1952
rect 28876 1912 28916 1952
rect 29260 1912 29300 1952
rect 30124 1912 30164 1952
rect 31276 1912 31316 1952
rect 31564 1912 31604 1952
rect 31948 1912 31988 1952
rect 32812 1912 32852 1952
rect 34060 1912 34100 1952
rect 17164 1744 17204 1784
rect 18220 1744 18260 1784
rect 18796 1744 18836 1784
rect 16492 1660 16532 1700
rect 25324 1660 25364 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 23404 1240 23444 1280
rect 26092 1240 26132 1280
rect 29644 1240 29684 1280
rect 17356 1156 17396 1196
rect 17260 1072 17300 1112
rect 17452 1072 17492 1112
rect 19276 1072 19316 1112
rect 19468 1072 19508 1112
rect 19564 1072 19604 1112
rect 26668 1072 26708 1112
rect 26860 1072 26900 1112
rect 19372 904 19412 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 9676 38417 9716 38502
rect 9675 38408 9717 38417
rect 9675 38368 9676 38408
rect 9716 38368 9717 38408
rect 9675 38359 9717 38368
rect 11883 38408 11925 38417
rect 11883 38368 11884 38408
rect 11924 38368 11925 38408
rect 11883 38359 11925 38368
rect 9580 38240 9620 38249
rect 9868 38240 9908 38249
rect 9484 38200 9580 38240
rect 9620 38200 9868 38240
rect 8044 38072 8084 38081
rect 3112 37820 3480 37829
rect 8044 37820 8084 38032
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 7852 37780 8084 37820
rect 267 37568 309 37577
rect 267 37528 268 37568
rect 308 37528 309 37568
rect 267 37519 309 37528
rect 268 20945 308 37519
rect 7084 37400 7124 37409
rect 7852 37400 7892 37780
rect 7124 37360 7316 37400
rect 7084 37351 7124 37360
rect 6988 37232 7028 37241
rect 6700 37192 6988 37232
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 6508 36728 6548 36737
rect 4300 36560 4340 36569
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 4300 35888 4340 36520
rect 4684 36560 4724 36569
rect 4724 36520 4820 36560
rect 4684 36511 4724 36520
rect 4300 35839 4340 35848
rect 3435 35804 3477 35813
rect 3435 35764 3436 35804
rect 3476 35764 3477 35804
rect 3435 35755 3477 35764
rect 3915 35804 3957 35813
rect 3915 35764 3916 35804
rect 3956 35764 3957 35804
rect 3915 35755 3957 35764
rect 3436 35300 3476 35755
rect 3916 35670 3956 35755
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3436 35251 3476 35260
rect 3244 35216 3284 35225
rect 1996 35048 2036 35057
rect 1324 34544 1364 34553
rect 1228 33704 1268 33713
rect 1324 33704 1364 34504
rect 1900 34376 1940 34385
rect 1996 34376 2036 35008
rect 3244 34973 3284 35176
rect 3339 35216 3381 35225
rect 3339 35176 3340 35216
rect 3380 35176 3381 35216
rect 3339 35167 3381 35176
rect 3532 35216 3572 35225
rect 3340 35082 3380 35167
rect 3243 34964 3285 34973
rect 3243 34924 3244 34964
rect 3284 34924 3285 34964
rect 3243 34915 3285 34924
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 3532 34385 3572 35176
rect 3723 35216 3765 35225
rect 3723 35176 3724 35216
rect 3764 35176 3765 35216
rect 3723 35167 3765 35176
rect 3820 35216 3860 35225
rect 3627 34964 3669 34973
rect 3627 34924 3628 34964
rect 3668 34924 3669 34964
rect 3627 34915 3669 34924
rect 1940 34336 2036 34376
rect 2764 34376 2804 34385
rect 3531 34376 3573 34385
rect 2804 34336 2900 34376
rect 1900 34327 1940 34336
rect 2764 34327 2804 34336
rect 1516 34292 1556 34301
rect 1556 34252 1748 34292
rect 1516 34243 1556 34252
rect 1612 33704 1652 33713
rect 1324 33664 1612 33704
rect 1131 33452 1173 33461
rect 1131 33412 1132 33452
rect 1172 33412 1173 33452
rect 1131 33403 1173 33412
rect 1132 32276 1172 33403
rect 1228 33377 1268 33664
rect 1612 33655 1652 33664
rect 1227 33368 1269 33377
rect 1227 33328 1228 33368
rect 1268 33328 1269 33368
rect 1227 33319 1269 33328
rect 1708 33125 1748 34252
rect 2476 33704 2516 33713
rect 2860 33704 2900 34336
rect 3531 34336 3532 34376
rect 3572 34336 3573 34376
rect 3531 34327 3573 34336
rect 3628 34301 3668 34915
rect 3627 34292 3669 34301
rect 3627 34252 3628 34292
rect 3668 34252 3669 34292
rect 3627 34243 3669 34252
rect 3724 33797 3764 35167
rect 3820 34805 3860 35176
rect 3916 35216 3956 35225
rect 3819 34796 3861 34805
rect 3819 34756 3820 34796
rect 3860 34756 3861 34796
rect 3819 34747 3861 34756
rect 3916 34721 3956 35176
rect 4012 35216 4052 35225
rect 3915 34712 3957 34721
rect 3915 34672 3916 34712
rect 3956 34672 3957 34712
rect 3915 34663 3957 34672
rect 3915 34208 3957 34217
rect 3915 34168 3916 34208
rect 3956 34168 3957 34208
rect 3915 34159 3957 34168
rect 3916 34074 3956 34159
rect 4012 33965 4052 35176
rect 4204 35216 4244 35225
rect 4204 34637 4244 35176
rect 4588 35216 4628 35225
rect 4780 35216 4820 36520
rect 5164 35888 5204 35897
rect 5204 35848 5396 35888
rect 5164 35839 5204 35848
rect 4628 35176 4820 35216
rect 4588 35167 4628 35176
rect 4683 34964 4725 34973
rect 4683 34924 4684 34964
rect 4724 34924 4725 34964
rect 4683 34915 4725 34924
rect 4203 34628 4245 34637
rect 4203 34588 4204 34628
rect 4244 34588 4245 34628
rect 4203 34579 4245 34588
rect 4491 34376 4533 34385
rect 4491 34336 4492 34376
rect 4532 34336 4533 34376
rect 4491 34327 4533 34336
rect 4588 34376 4628 34385
rect 4492 34242 4532 34327
rect 4588 34208 4628 34336
rect 4684 34376 4724 34915
rect 5067 34712 5109 34721
rect 5067 34672 5068 34712
rect 5108 34672 5109 34712
rect 5067 34663 5109 34672
rect 4779 34460 4821 34469
rect 4779 34420 4780 34460
rect 4820 34420 4821 34460
rect 4779 34411 4821 34420
rect 4684 34327 4724 34336
rect 4780 34376 4820 34411
rect 5068 34376 5108 34663
rect 5259 34544 5301 34553
rect 5259 34504 5260 34544
rect 5300 34504 5301 34544
rect 5259 34495 5301 34504
rect 5260 34421 5300 34495
rect 4780 34325 4820 34336
rect 4876 34336 5068 34376
rect 4876 34208 4916 34336
rect 5068 34327 5108 34336
rect 5164 34376 5204 34385
rect 5260 34372 5300 34381
rect 5164 34292 5204 34336
rect 5164 34252 5300 34292
rect 4588 34168 4916 34208
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 4011 33956 4053 33965
rect 4011 33916 4012 33956
rect 4052 33916 4053 33956
rect 4011 33907 4053 33916
rect 3531 33788 3573 33797
rect 3531 33748 3532 33788
rect 3572 33748 3573 33788
rect 3531 33739 3573 33748
rect 3723 33788 3765 33797
rect 3723 33748 3724 33788
rect 3764 33748 3765 33788
rect 3723 33739 3765 33748
rect 4011 33788 4053 33797
rect 4011 33748 4012 33788
rect 4052 33748 4053 33788
rect 4011 33739 4053 33748
rect 2516 33664 2900 33704
rect 2476 33655 2516 33664
rect 2475 33200 2517 33209
rect 2380 33160 2476 33200
rect 2516 33160 2517 33200
rect 1707 33116 1749 33125
rect 1707 33076 1708 33116
rect 1748 33076 1749 33116
rect 1707 33067 1749 33076
rect 2380 33116 2420 33160
rect 2475 33151 2517 33160
rect 2380 33067 2420 33076
rect 1612 33032 1652 33041
rect 1612 32780 1652 32992
rect 1995 33032 2037 33041
rect 1995 32992 1996 33032
rect 2036 32992 2037 33032
rect 1995 32983 2037 32992
rect 1132 32227 1172 32236
rect 1516 32740 1652 32780
rect 1516 32192 1556 32740
rect 1516 32143 1556 32152
rect 1324 31520 1364 31529
rect 1364 31480 1652 31520
rect 1324 31471 1364 31480
rect 1612 31352 1652 31480
rect 1900 31352 1940 31361
rect 1612 31312 1900 31352
rect 1900 31303 1940 31312
rect 1516 31268 1556 31277
rect 1516 31184 1556 31228
rect 1996 31184 2036 32983
rect 2476 32864 2516 32873
rect 2476 32369 2516 32824
rect 2667 32864 2709 32873
rect 2667 32824 2668 32864
rect 2708 32824 2709 32864
rect 2667 32815 2709 32824
rect 2764 32864 2804 32873
rect 2668 32730 2708 32815
rect 2475 32360 2517 32369
rect 2475 32320 2476 32360
rect 2516 32320 2517 32360
rect 2475 32311 2517 32320
rect 2379 32192 2421 32201
rect 2379 32152 2380 32192
rect 2420 32152 2421 32192
rect 2379 32143 2421 32152
rect 2380 32058 2420 32143
rect 2764 31613 2804 32824
rect 2860 32789 2900 33664
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 3243 33116 3285 33125
rect 3243 33076 3244 33116
rect 3284 33076 3285 33116
rect 3243 33067 3285 33076
rect 3244 32982 3284 33067
rect 3532 32957 3572 33739
rect 3819 33704 3861 33713
rect 3819 33664 3820 33704
rect 3860 33664 3861 33704
rect 3819 33655 3861 33664
rect 4012 33704 4052 33739
rect 3627 33620 3669 33629
rect 3627 33580 3628 33620
rect 3668 33580 3669 33620
rect 3627 33571 3669 33580
rect 3628 33486 3668 33571
rect 3820 33570 3860 33655
rect 4012 33653 4052 33664
rect 4108 33704 4148 33713
rect 4300 33704 4340 33713
rect 3819 33452 3861 33461
rect 3819 33412 3820 33452
rect 3860 33412 3861 33452
rect 3819 33403 3861 33412
rect 3820 33318 3860 33403
rect 3723 33116 3765 33125
rect 3723 33076 3724 33116
rect 3764 33076 3765 33116
rect 3723 33067 3765 33076
rect 3051 32948 3093 32957
rect 3051 32908 3052 32948
rect 3092 32908 3093 32948
rect 3051 32899 3093 32908
rect 3531 32948 3573 32957
rect 3531 32908 3532 32948
rect 3572 32908 3573 32948
rect 3531 32899 3573 32908
rect 2955 32864 2997 32873
rect 2955 32824 2956 32864
rect 2996 32824 2997 32864
rect 2955 32815 2997 32824
rect 3052 32864 3092 32899
rect 2859 32780 2901 32789
rect 2859 32740 2860 32780
rect 2900 32740 2901 32780
rect 2859 32731 2901 32740
rect 2860 32201 2900 32731
rect 2956 32730 2996 32815
rect 3052 32813 3092 32824
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3532 32864 3572 32899
rect 3244 32730 3284 32815
rect 3532 32814 3572 32824
rect 3724 32864 3764 33067
rect 4108 32957 4148 33664
rect 4204 33664 4300 33704
rect 4107 32948 4149 32957
rect 4107 32908 4108 32948
rect 4148 32908 4149 32948
rect 4107 32899 4149 32908
rect 3724 32815 3764 32824
rect 3916 32864 3956 32873
rect 3723 32360 3765 32369
rect 3723 32320 3724 32360
rect 3764 32320 3765 32360
rect 3723 32311 3765 32320
rect 3724 32226 3764 32311
rect 2859 32192 2901 32201
rect 2859 32152 2860 32192
rect 2900 32152 2901 32192
rect 2859 32143 2901 32152
rect 2763 31604 2805 31613
rect 2763 31564 2764 31604
rect 2804 31564 2805 31604
rect 2763 31555 2805 31564
rect 2764 31352 2804 31361
rect 2860 31352 2900 32143
rect 3916 31949 3956 32824
rect 3531 31940 3573 31949
rect 3531 31900 3532 31940
rect 3572 31900 3573 31940
rect 3531 31891 3573 31900
rect 3915 31940 3957 31949
rect 3915 31900 3916 31940
rect 3956 31900 3957 31940
rect 3915 31891 3957 31900
rect 3532 31806 3572 31891
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3915 31688 3957 31697
rect 3915 31648 3916 31688
rect 3956 31648 3957 31688
rect 3915 31639 3957 31648
rect 3819 31604 3861 31613
rect 3819 31564 3820 31604
rect 3860 31564 3861 31604
rect 3819 31555 3861 31564
rect 1516 31144 2036 31184
rect 2572 31312 2764 31352
rect 2804 31312 2900 31352
rect 1804 30512 1844 30521
rect 1323 30428 1365 30437
rect 1323 30388 1324 30428
rect 1364 30388 1365 30428
rect 1323 30379 1365 30388
rect 1324 29840 1364 30379
rect 1324 29791 1364 29800
rect 1708 29840 1748 29849
rect 1804 29840 1844 30472
rect 1748 29800 1844 29840
rect 2572 29840 2612 31312
rect 2764 31303 2804 31312
rect 3820 30848 3860 31555
rect 3916 31520 3956 31639
rect 3916 31471 3956 31480
rect 4011 31436 4053 31445
rect 4011 31396 4012 31436
rect 4052 31396 4053 31436
rect 4011 31387 4053 31396
rect 3916 30848 3956 30857
rect 3820 30808 3916 30848
rect 3916 30799 3956 30808
rect 3724 30680 3764 30689
rect 3052 30437 3092 30522
rect 3051 30428 3093 30437
rect 3051 30388 3052 30428
rect 3092 30388 3093 30428
rect 3051 30379 3093 30388
rect 3724 30269 3764 30640
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3723 30260 3765 30269
rect 3723 30220 3724 30260
rect 3764 30220 3765 30260
rect 3723 30211 3765 30220
rect 3819 30176 3861 30185
rect 3819 30136 3820 30176
rect 3860 30136 3861 30176
rect 3819 30127 3861 30136
rect 3723 30092 3765 30101
rect 3723 30052 3724 30092
rect 3764 30052 3765 30092
rect 3723 30043 3765 30052
rect 3724 29958 3764 30043
rect 1708 29791 1748 29800
rect 2572 29791 2612 29800
rect 2667 29840 2709 29849
rect 2667 29800 2668 29840
rect 2708 29800 2709 29840
rect 2667 29791 2709 29800
rect 1323 29252 1365 29261
rect 1323 29212 1324 29252
rect 1364 29212 1365 29252
rect 1323 29203 1365 29212
rect 1324 29118 1364 29203
rect 1708 29168 1748 29177
rect 1708 29009 1748 29128
rect 2571 29168 2613 29177
rect 2571 29128 2572 29168
rect 2612 29128 2613 29168
rect 2571 29119 2613 29128
rect 2572 29034 2612 29119
rect 1131 29000 1173 29009
rect 1131 28960 1132 29000
rect 1172 28960 1173 29000
rect 1131 28951 1173 28960
rect 1707 29000 1749 29009
rect 1707 28960 1708 29000
rect 1748 28960 1749 29000
rect 1707 28951 1749 28960
rect 1132 28866 1172 28951
rect 2572 28580 2612 28589
rect 2668 28580 2708 29791
rect 3723 29756 3765 29765
rect 3723 29716 3724 29756
rect 3764 29716 3765 29756
rect 3723 29707 3765 29716
rect 3724 29336 3764 29707
rect 3724 29287 3764 29296
rect 3531 29168 3573 29177
rect 3531 29128 3532 29168
rect 3572 29128 3573 29168
rect 3531 29119 3573 29128
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 2763 28664 2805 28673
rect 2763 28624 2764 28664
rect 2804 28624 2805 28664
rect 2763 28615 2805 28624
rect 2612 28540 2708 28580
rect 2572 28531 2612 28540
rect 1708 28496 1748 28505
rect 1612 28456 1708 28496
rect 1228 27656 1268 27665
rect 1228 26909 1268 27616
rect 1612 27656 1652 28456
rect 1708 28447 1748 28456
rect 2668 28328 2708 28337
rect 2764 28328 2804 28615
rect 3532 28580 3572 29119
rect 3820 29000 3860 30127
rect 4012 29765 4052 31387
rect 4204 30848 4244 33664
rect 4300 33655 4340 33664
rect 4492 33704 4532 33713
rect 4300 33452 4340 33461
rect 4300 33041 4340 33412
rect 4492 33125 4532 33664
rect 4588 33704 4628 33713
rect 4779 33704 4821 33713
rect 4628 33664 4724 33704
rect 4588 33655 4628 33664
rect 4491 33116 4533 33125
rect 4491 33076 4492 33116
rect 4532 33076 4533 33116
rect 4491 33067 4533 33076
rect 4299 33032 4341 33041
rect 4299 32992 4300 33032
rect 4340 32992 4341 33032
rect 4684 33032 4724 33664
rect 4779 33664 4780 33704
rect 4820 33664 4821 33704
rect 4779 33655 4821 33664
rect 4876 33704 4916 34168
rect 4972 34208 5012 34217
rect 5012 34168 5204 34208
rect 4972 34159 5012 34168
rect 4780 33570 4820 33655
rect 4876 33293 4916 33664
rect 4972 33704 5012 33713
rect 4875 33284 4917 33293
rect 4875 33244 4876 33284
rect 4916 33244 4917 33284
rect 4875 33235 4917 33244
rect 4684 32992 4916 33032
rect 4299 32983 4341 32992
rect 4780 32864 4820 32873
rect 4588 32780 4628 32791
rect 4588 32705 4628 32740
rect 4587 32696 4629 32705
rect 4587 32656 4588 32696
rect 4628 32656 4629 32696
rect 4587 32647 4629 32656
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4683 32360 4725 32369
rect 4683 32320 4684 32360
rect 4724 32320 4725 32360
rect 4683 32311 4725 32320
rect 4396 32192 4436 32201
rect 4300 32152 4396 32192
rect 4300 31445 4340 32152
rect 4396 32143 4436 32152
rect 4491 31940 4533 31949
rect 4491 31900 4492 31940
rect 4532 31900 4533 31940
rect 4491 31891 4533 31900
rect 4395 31520 4437 31529
rect 4395 31480 4396 31520
rect 4436 31480 4437 31520
rect 4395 31471 4437 31480
rect 4299 31436 4341 31445
rect 4299 31396 4300 31436
rect 4340 31396 4341 31436
rect 4299 31387 4341 31396
rect 4396 31352 4436 31471
rect 4396 31303 4436 31312
rect 4492 31352 4532 31891
rect 4492 31303 4532 31312
rect 4684 31268 4724 32311
rect 4780 31697 4820 32824
rect 4779 31688 4821 31697
rect 4779 31648 4780 31688
rect 4820 31648 4821 31688
rect 4779 31639 4821 31648
rect 4780 31352 4820 31639
rect 4876 31613 4916 32992
rect 4972 32705 5012 33664
rect 5067 33704 5109 33713
rect 5067 33664 5068 33704
rect 5108 33664 5109 33704
rect 5067 33655 5109 33664
rect 5068 33570 5108 33655
rect 5067 33116 5109 33125
rect 5067 33076 5068 33116
rect 5108 33076 5109 33116
rect 5067 33067 5109 33076
rect 4971 32696 5013 32705
rect 4971 32656 4972 32696
rect 5012 32656 5013 32696
rect 4971 32647 5013 32656
rect 4875 31604 4917 31613
rect 4875 31564 4876 31604
rect 4916 31564 4917 31604
rect 4875 31555 4917 31564
rect 4876 31436 4916 31445
rect 4876 31352 4916 31396
rect 4780 31312 4916 31352
rect 4972 31352 5012 31361
rect 4684 31228 4916 31268
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4780 30848 4820 30857
rect 4204 30808 4780 30848
rect 4780 30799 4820 30808
rect 4587 30680 4629 30689
rect 4587 30640 4588 30680
rect 4628 30640 4629 30680
rect 4587 30631 4629 30640
rect 4876 30680 4916 31228
rect 4972 30857 5012 31312
rect 4971 30848 5013 30857
rect 4971 30808 4972 30848
rect 5012 30808 5013 30848
rect 4971 30799 5013 30808
rect 4876 30631 4916 30640
rect 4971 30680 5013 30689
rect 4971 30640 4972 30680
rect 5012 30640 5013 30680
rect 4971 30631 5013 30640
rect 5068 30680 5108 33067
rect 5164 32873 5204 34168
rect 5260 33881 5300 34252
rect 5259 33872 5301 33881
rect 5259 33832 5260 33872
rect 5300 33832 5301 33872
rect 5259 33823 5301 33832
rect 5163 32864 5205 32873
rect 5163 32824 5164 32864
rect 5204 32824 5205 32864
rect 5163 32815 5205 32824
rect 5356 32789 5396 35848
rect 6315 35720 6357 35729
rect 6315 35680 6316 35720
rect 6356 35680 6357 35720
rect 6315 35671 6357 35680
rect 6316 35586 6356 35671
rect 6411 35636 6453 35645
rect 6508 35636 6548 36688
rect 6603 36644 6645 36653
rect 6603 36604 6604 36644
rect 6644 36604 6645 36644
rect 6603 36595 6645 36604
rect 6604 36510 6644 36595
rect 6700 36308 6740 37192
rect 6988 37183 7028 37192
rect 7180 36728 7220 36737
rect 6987 36560 7029 36569
rect 6987 36520 6988 36560
rect 7028 36520 7029 36560
rect 6987 36511 7029 36520
rect 6988 36426 7028 36511
rect 6604 36268 6740 36308
rect 6604 35888 6644 36268
rect 6892 36140 6932 36149
rect 7180 36140 7220 36688
rect 6932 36100 7220 36140
rect 6892 36091 6932 36100
rect 6700 35897 6740 35982
rect 6604 35839 6644 35848
rect 6699 35888 6741 35897
rect 6699 35848 6700 35888
rect 6740 35848 6741 35888
rect 6699 35839 6741 35848
rect 6891 35888 6933 35897
rect 6891 35848 6892 35888
rect 6932 35848 6933 35888
rect 6891 35839 6933 35848
rect 6892 35754 6932 35839
rect 6795 35720 6837 35729
rect 6795 35680 6796 35720
rect 6836 35680 6837 35720
rect 6795 35671 6837 35680
rect 7084 35720 7124 35731
rect 6411 35596 6412 35636
rect 6452 35596 6548 35636
rect 6411 35587 6453 35596
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5452 35082 5492 35167
rect 5451 34796 5493 34805
rect 5451 34756 5452 34796
rect 5492 34756 5493 34796
rect 5451 34747 5493 34756
rect 5452 34628 5492 34747
rect 5452 34579 5492 34588
rect 5643 34544 5685 34553
rect 5643 34504 5644 34544
rect 5684 34504 5685 34544
rect 5643 34495 5685 34504
rect 5451 34040 5493 34049
rect 5451 34000 5452 34040
rect 5492 34000 5493 34040
rect 5451 33991 5493 34000
rect 5452 33704 5492 33991
rect 5547 33956 5589 33965
rect 5547 33916 5548 33956
rect 5588 33916 5589 33956
rect 5547 33907 5589 33916
rect 5452 33655 5492 33664
rect 5548 32864 5588 33907
rect 5644 33713 5684 34495
rect 6315 34460 6357 34469
rect 6315 34420 6316 34460
rect 6356 34420 6357 34460
rect 6315 34411 6357 34420
rect 6124 34376 6164 34385
rect 6028 34336 6124 34376
rect 5643 33704 5685 33713
rect 5643 33664 5644 33704
rect 5684 33664 5685 33704
rect 5643 33655 5685 33664
rect 5835 33704 5877 33713
rect 5835 33664 5836 33704
rect 5876 33664 5877 33704
rect 5835 33655 5877 33664
rect 5643 33368 5685 33377
rect 5643 33328 5644 33368
rect 5684 33328 5685 33368
rect 5643 33319 5685 33328
rect 5644 33116 5684 33319
rect 5644 33067 5684 33076
rect 5644 32864 5684 32873
rect 5548 32824 5644 32864
rect 5644 32815 5684 32824
rect 5836 32864 5876 33655
rect 6028 33629 6068 34336
rect 6124 34327 6164 34336
rect 6219 34376 6261 34385
rect 6219 34336 6220 34376
rect 6260 34336 6261 34376
rect 6219 34327 6261 34336
rect 6316 34376 6356 34411
rect 6123 33872 6165 33881
rect 6123 33832 6124 33872
rect 6164 33832 6165 33872
rect 6123 33823 6165 33832
rect 6124 33738 6164 33823
rect 6027 33620 6069 33629
rect 6027 33580 6028 33620
rect 6068 33580 6069 33620
rect 6027 33571 6069 33580
rect 6123 33452 6165 33461
rect 6123 33412 6124 33452
rect 6164 33412 6165 33452
rect 6123 33403 6165 33412
rect 6124 33318 6164 33403
rect 5931 33200 5973 33209
rect 5931 33160 5932 33200
rect 5972 33160 5973 33200
rect 5931 33151 5973 33160
rect 5836 32815 5876 32824
rect 5932 32864 5972 33151
rect 6220 33116 6260 34327
rect 6316 34325 6356 34336
rect 6412 34376 6452 35587
rect 6796 35216 6836 35671
rect 7084 35645 7124 35680
rect 7083 35636 7125 35645
rect 7083 35596 7084 35636
rect 7124 35596 7125 35636
rect 7083 35587 7125 35596
rect 6603 35132 6645 35141
rect 6603 35092 6604 35132
rect 6644 35092 6645 35132
rect 6603 35083 6645 35092
rect 6604 34998 6644 35083
rect 6796 35057 6836 35176
rect 6891 35132 6933 35141
rect 6891 35092 6892 35132
rect 6932 35092 6933 35132
rect 6891 35083 6933 35092
rect 6795 35048 6837 35057
rect 6795 35008 6796 35048
rect 6836 35008 6837 35048
rect 6795 34999 6837 35008
rect 6507 34712 6549 34721
rect 6507 34672 6508 34712
rect 6548 34672 6549 34712
rect 6507 34663 6549 34672
rect 6412 34327 6452 34336
rect 6508 34376 6548 34663
rect 6796 34637 6836 34722
rect 6795 34628 6837 34637
rect 6795 34588 6796 34628
rect 6836 34588 6837 34628
rect 6795 34579 6837 34588
rect 6508 34301 6548 34336
rect 6604 34376 6644 34385
rect 6796 34376 6836 34385
rect 6644 34336 6796 34376
rect 6604 34327 6644 34336
rect 6796 34327 6836 34336
rect 6507 34292 6549 34301
rect 6507 34252 6508 34292
rect 6548 34252 6549 34292
rect 6507 34243 6549 34252
rect 6315 34208 6357 34217
rect 6315 34168 6316 34208
rect 6356 34168 6357 34208
rect 6315 34159 6357 34168
rect 6316 33536 6356 34159
rect 6507 34124 6549 34133
rect 6507 34084 6508 34124
rect 6548 34084 6549 34124
rect 6507 34075 6549 34084
rect 6508 33724 6548 34075
rect 6412 33704 6452 33713
rect 6508 33675 6548 33684
rect 6892 33704 6932 35083
rect 7276 34973 7316 37360
rect 7852 37351 7892 37360
rect 8716 37400 8756 37409
rect 7467 37316 7509 37325
rect 7467 37276 7468 37316
rect 7508 37276 7509 37316
rect 7467 37267 7509 37276
rect 8331 37316 8373 37325
rect 8331 37276 8332 37316
rect 8372 37276 8373 37316
rect 8331 37267 8373 37276
rect 7468 37182 7508 37267
rect 7564 36728 7604 36737
rect 7564 36569 7604 36688
rect 8043 36644 8085 36653
rect 8043 36604 8044 36644
rect 8084 36604 8085 36644
rect 8043 36595 8085 36604
rect 7563 36560 7605 36569
rect 7563 36520 7564 36560
rect 7604 36520 7605 36560
rect 7563 36511 7605 36520
rect 7756 35888 7796 35897
rect 7660 35216 7700 35225
rect 7371 35048 7413 35057
rect 7371 35008 7372 35048
rect 7412 35008 7413 35048
rect 7371 34999 7413 35008
rect 7275 34964 7317 34973
rect 7275 34924 7276 34964
rect 7316 34924 7317 34964
rect 7275 34915 7317 34924
rect 6987 34544 7029 34553
rect 6987 34504 6988 34544
rect 7028 34504 7029 34544
rect 6987 34495 7029 34504
rect 6988 34376 7028 34495
rect 7372 34469 7412 34999
rect 7467 34964 7509 34973
rect 7467 34924 7468 34964
rect 7508 34924 7509 34964
rect 7467 34915 7509 34924
rect 7468 34830 7508 34915
rect 7660 34805 7700 35176
rect 7756 35141 7796 35848
rect 8044 35888 8084 36595
rect 8332 36140 8372 37267
rect 8332 36091 8372 36100
rect 8428 36728 8468 36737
rect 8716 36728 8756 37360
rect 8468 36688 8756 36728
rect 8139 35972 8181 35981
rect 8139 35932 8140 35972
rect 8180 35932 8181 35972
rect 8139 35923 8181 35932
rect 8044 35839 8084 35848
rect 8140 35888 8180 35923
rect 8140 35837 8180 35848
rect 8331 35888 8373 35897
rect 8331 35848 8332 35888
rect 8372 35848 8373 35888
rect 8331 35839 8373 35848
rect 8332 35754 8372 35839
rect 8139 35720 8181 35729
rect 8139 35680 8140 35720
rect 8180 35680 8181 35720
rect 8139 35671 8181 35680
rect 8044 35216 8084 35225
rect 7852 35176 8044 35216
rect 7755 35132 7797 35141
rect 7755 35092 7756 35132
rect 7796 35092 7797 35132
rect 7755 35083 7797 35092
rect 7756 34964 7796 34973
rect 7659 34796 7701 34805
rect 7659 34756 7660 34796
rect 7700 34756 7701 34796
rect 7659 34747 7701 34756
rect 7756 34628 7796 34924
rect 7660 34588 7796 34628
rect 7371 34460 7413 34469
rect 7371 34420 7372 34460
rect 7412 34420 7413 34460
rect 7371 34411 7413 34420
rect 6988 34327 7028 34336
rect 7083 34376 7125 34385
rect 7276 34376 7316 34385
rect 7083 34336 7084 34376
rect 7124 34336 7125 34376
rect 7083 34327 7125 34336
rect 7180 34336 7276 34376
rect 7084 34242 7124 34327
rect 6987 34040 7029 34049
rect 6987 34000 6988 34040
rect 7028 34000 7029 34040
rect 6987 33991 7029 34000
rect 6412 33620 6452 33664
rect 6892 33655 6932 33664
rect 6988 33704 7028 33991
rect 6988 33655 7028 33664
rect 6412 33580 6556 33620
rect 6516 33536 6556 33580
rect 6316 33496 6452 33536
rect 6220 33067 6260 33076
rect 6219 32948 6261 32957
rect 6219 32908 6220 32948
rect 6260 32908 6261 32948
rect 6219 32899 6261 32908
rect 6124 32864 6164 32873
rect 5932 32815 5972 32824
rect 6028 32824 6124 32864
rect 5355 32780 5397 32789
rect 5355 32740 5356 32780
rect 5396 32740 5397 32780
rect 5355 32731 5397 32740
rect 5452 32780 5492 32789
rect 5260 32360 5300 32369
rect 5356 32360 5396 32731
rect 5300 32320 5396 32360
rect 5452 32528 5492 32740
rect 6028 32528 6068 32824
rect 6124 32815 6164 32824
rect 5452 32488 6068 32528
rect 5260 32311 5300 32320
rect 5452 32108 5492 32488
rect 6123 32444 6165 32453
rect 6123 32404 6124 32444
rect 6164 32404 6165 32444
rect 6123 32395 6165 32404
rect 5356 32068 5492 32108
rect 5740 32192 5780 32201
rect 5356 30689 5396 32068
rect 5740 32033 5780 32152
rect 6124 32192 6164 32395
rect 6124 32143 6164 32152
rect 5739 32024 5781 32033
rect 5739 31984 5740 32024
rect 5780 31984 5781 32024
rect 5739 31975 5781 31984
rect 6028 32024 6068 32033
rect 6220 32024 6260 32899
rect 6315 32696 6357 32705
rect 6315 32656 6316 32696
rect 6356 32656 6357 32696
rect 6315 32647 6357 32656
rect 6316 32192 6356 32647
rect 6412 32360 6452 33496
rect 6508 33496 6556 33536
rect 6508 32873 6548 33496
rect 6603 33452 6645 33461
rect 6603 33412 6604 33452
rect 6644 33412 6645 33452
rect 6603 33403 6645 33412
rect 6507 32864 6549 32873
rect 6507 32824 6508 32864
rect 6548 32824 6549 32864
rect 6507 32815 6549 32824
rect 6412 32311 6452 32320
rect 6316 32143 6356 32152
rect 6068 31984 6260 32024
rect 6028 31975 6068 31984
rect 6315 31604 6357 31613
rect 6315 31564 6316 31604
rect 6356 31564 6357 31604
rect 6315 31555 6357 31564
rect 6316 31520 6356 31555
rect 6508 31529 6548 32815
rect 6604 32192 6644 33403
rect 6699 33032 6741 33041
rect 6699 32992 6700 33032
rect 6740 32992 6741 33032
rect 6699 32983 6741 32992
rect 6700 32898 6740 32983
rect 7180 32948 7220 34336
rect 7276 34327 7316 34336
rect 7372 34376 7412 34411
rect 7275 33032 7317 33041
rect 7275 32992 7276 33032
rect 7316 32992 7317 33032
rect 7275 32983 7317 32992
rect 6796 32908 7220 32948
rect 6796 32360 6836 32908
rect 7276 32864 7316 32983
rect 7276 32815 7316 32824
rect 6892 32780 6932 32789
rect 6932 32740 7220 32780
rect 6892 32731 6932 32740
rect 7180 32360 7220 32740
rect 7276 32360 7316 32369
rect 7180 32320 7276 32360
rect 6796 32311 6836 32320
rect 7276 32311 7316 32320
rect 7372 32285 7412 34336
rect 7563 34376 7605 34385
rect 7563 34336 7564 34376
rect 7604 34336 7605 34376
rect 7563 34327 7605 34336
rect 7564 34242 7604 34327
rect 7467 34208 7509 34217
rect 7467 34168 7468 34208
rect 7508 34168 7509 34208
rect 7467 34159 7509 34168
rect 7468 34074 7508 34159
rect 7468 33713 7508 33798
rect 7467 33704 7509 33713
rect 7467 33664 7468 33704
rect 7508 33664 7509 33704
rect 7467 33655 7509 33664
rect 7660 33536 7700 34588
rect 7756 34292 7796 34303
rect 7756 34217 7796 34252
rect 7755 34208 7797 34217
rect 7755 34168 7756 34208
rect 7796 34168 7797 34208
rect 7755 34159 7797 34168
rect 7468 33496 7700 33536
rect 7371 32276 7413 32285
rect 7371 32236 7372 32276
rect 7412 32236 7413 32276
rect 7371 32227 7413 32236
rect 6700 32192 6740 32201
rect 6604 32152 6700 32192
rect 6700 32143 6740 32152
rect 7179 32192 7221 32201
rect 7179 32152 7180 32192
rect 7220 32152 7221 32192
rect 7179 32143 7221 32152
rect 7372 32192 7412 32227
rect 7180 32058 7220 32143
rect 7372 32142 7412 32152
rect 7468 32192 7508 33496
rect 7468 32143 7508 32152
rect 7852 32024 7892 35176
rect 8044 35167 8084 35176
rect 8140 34376 8180 35671
rect 8428 35384 8468 36688
rect 9099 36476 9141 36485
rect 9099 36436 9100 36476
rect 9140 36436 9141 36476
rect 9099 36427 9141 36436
rect 8524 36056 8564 36065
rect 8524 35729 8564 36016
rect 9004 35888 9044 35897
rect 8907 35804 8949 35813
rect 8907 35764 8908 35804
rect 8948 35764 8949 35804
rect 8907 35755 8949 35764
rect 8523 35720 8565 35729
rect 8523 35680 8524 35720
rect 8564 35680 8565 35720
rect 8523 35671 8565 35680
rect 8908 35670 8948 35755
rect 8524 35384 8564 35393
rect 8428 35344 8524 35384
rect 9004 35384 9044 35848
rect 9100 35888 9140 36427
rect 9484 36308 9524 38200
rect 9580 38191 9620 38200
rect 9868 38191 9908 38200
rect 10540 38240 10580 38249
rect 9771 37736 9813 37745
rect 9771 37696 9772 37736
rect 9812 37696 9813 37736
rect 9771 37687 9813 37696
rect 9579 36644 9621 36653
rect 9579 36604 9580 36644
rect 9620 36604 9621 36644
rect 9579 36595 9621 36604
rect 9580 36510 9620 36595
rect 9484 36268 9620 36308
rect 9195 35972 9237 35981
rect 9195 35932 9196 35972
rect 9236 35932 9237 35972
rect 9195 35923 9237 35932
rect 9100 35839 9140 35848
rect 9196 35888 9236 35923
rect 9196 35837 9236 35848
rect 9387 35888 9429 35897
rect 9387 35848 9388 35888
rect 9428 35848 9429 35888
rect 9387 35839 9429 35848
rect 9484 35888 9524 35897
rect 9388 35754 9428 35839
rect 9196 35384 9236 35393
rect 9484 35384 9524 35848
rect 9580 35888 9620 36268
rect 9675 35972 9717 35981
rect 9675 35932 9676 35972
rect 9716 35932 9717 35972
rect 9675 35923 9717 35932
rect 9580 35839 9620 35848
rect 9676 35888 9716 35923
rect 9772 35888 9812 37687
rect 10540 37661 10580 38200
rect 10732 38240 10772 38249
rect 11596 38240 11636 38249
rect 11788 38240 11828 38249
rect 10732 38081 10772 38200
rect 11500 38200 11596 38240
rect 10731 38072 10773 38081
rect 10731 38032 10732 38072
rect 10772 38032 10773 38072
rect 10731 38023 10773 38032
rect 11403 37988 11445 37997
rect 11403 37948 11404 37988
rect 11444 37948 11445 37988
rect 11403 37939 11445 37948
rect 11404 37854 11444 37939
rect 11500 37829 11540 38200
rect 11596 38191 11636 38200
rect 11692 38200 11788 38240
rect 11595 38072 11637 38081
rect 11595 38032 11596 38072
rect 11636 38032 11637 38072
rect 11595 38023 11637 38032
rect 11596 37938 11636 38023
rect 11499 37820 11541 37829
rect 11499 37780 11500 37820
rect 11540 37780 11541 37820
rect 11499 37771 11541 37780
rect 9867 37652 9909 37661
rect 9867 37612 9868 37652
rect 9908 37612 9909 37652
rect 9867 37603 9909 37612
rect 10539 37652 10581 37661
rect 10539 37612 10540 37652
rect 10580 37612 10581 37652
rect 10539 37603 10581 37612
rect 9868 37518 9908 37603
rect 11692 37568 11732 38200
rect 11788 38191 11828 38200
rect 11884 38240 11924 38359
rect 11884 38191 11924 38200
rect 12268 38072 12308 38081
rect 12268 37820 12308 38032
rect 12843 37988 12885 37997
rect 12843 37948 12844 37988
rect 12884 37948 12885 37988
rect 12843 37939 12885 37948
rect 12268 37780 12500 37820
rect 11212 37528 11732 37568
rect 10060 37400 10100 37409
rect 9964 37360 10060 37400
rect 9868 37232 9908 37241
rect 9868 36821 9908 37192
rect 9964 36896 10004 37360
rect 10060 37351 10100 37360
rect 10059 37232 10101 37241
rect 10059 37192 10060 37232
rect 10100 37192 10101 37232
rect 10059 37183 10101 37192
rect 10156 37232 10196 37241
rect 10443 37232 10485 37241
rect 10196 37192 10388 37232
rect 10156 37183 10196 37192
rect 9964 36847 10004 36856
rect 9867 36812 9909 36821
rect 9867 36772 9868 36812
rect 9908 36772 9909 36812
rect 9867 36763 9909 36772
rect 9963 36476 10005 36485
rect 9963 36436 9964 36476
rect 10004 36436 10005 36476
rect 9963 36427 10005 36436
rect 9964 36342 10004 36427
rect 9868 35888 9908 35897
rect 9772 35848 9868 35888
rect 9676 35837 9716 35848
rect 9868 35839 9908 35848
rect 9964 35888 10004 35897
rect 9964 35384 10004 35848
rect 10060 35888 10100 37183
rect 10348 36980 10388 37192
rect 10443 37192 10444 37232
rect 10484 37192 10485 37232
rect 10443 37183 10485 37192
rect 10444 37098 10484 37183
rect 10348 36940 11156 36980
rect 10827 36812 10869 36821
rect 10827 36772 10828 36812
rect 10868 36772 10869 36812
rect 10827 36763 10869 36772
rect 10636 36728 10676 36739
rect 10636 36653 10676 36688
rect 10635 36644 10677 36653
rect 10635 36604 10636 36644
rect 10676 36604 10772 36644
rect 10635 36595 10677 36604
rect 10155 35972 10197 35981
rect 10155 35932 10156 35972
rect 10196 35932 10197 35972
rect 10155 35923 10197 35932
rect 10060 35839 10100 35848
rect 10156 35888 10196 35923
rect 10156 35813 10196 35848
rect 10444 35888 10484 35897
rect 10155 35804 10197 35813
rect 10155 35764 10156 35804
rect 10196 35764 10197 35804
rect 10155 35755 10197 35764
rect 10156 35724 10196 35755
rect 9004 35344 9196 35384
rect 9236 35344 10004 35384
rect 8428 35225 8468 35344
rect 8524 35335 8564 35344
rect 9196 35335 9236 35344
rect 8427 35216 8469 35225
rect 8427 35176 8428 35216
rect 8468 35176 8469 35216
rect 8427 35167 8469 35176
rect 9580 35216 9620 35225
rect 9388 35132 9428 35141
rect 8140 34327 8180 34336
rect 8716 34964 8756 34973
rect 8716 34376 8756 34924
rect 9388 34553 9428 35092
rect 9387 34544 9429 34553
rect 9387 34504 9388 34544
rect 9428 34504 9429 34544
rect 9387 34495 9429 34504
rect 9580 34469 9620 35176
rect 9676 35216 9716 35344
rect 9676 35167 9716 35176
rect 9772 35216 9812 35225
rect 9772 34964 9812 35176
rect 9867 35216 9909 35225
rect 9867 35176 9868 35216
rect 9908 35176 9909 35216
rect 9867 35167 9909 35176
rect 9868 35082 9908 35167
rect 10060 34964 10100 34973
rect 9772 34924 10060 34964
rect 9579 34460 9621 34469
rect 9579 34420 9580 34460
rect 9620 34420 9621 34460
rect 9579 34411 9621 34420
rect 9004 34376 9044 34385
rect 8716 34336 9004 34376
rect 8043 34292 8085 34301
rect 8043 34252 8044 34292
rect 8084 34252 8085 34292
rect 8043 34243 8085 34252
rect 7948 33690 7988 33699
rect 7948 32789 7988 33650
rect 7947 32780 7989 32789
rect 7947 32740 7948 32780
rect 7988 32740 7989 32780
rect 7947 32731 7989 32740
rect 7948 32201 7988 32286
rect 7947 32192 7989 32201
rect 7947 32152 7948 32192
rect 7988 32152 7989 32192
rect 7947 32143 7989 32152
rect 8044 32192 8084 34243
rect 8139 33788 8181 33797
rect 8139 33748 8140 33788
rect 8180 33748 8181 33788
rect 8139 33739 8181 33748
rect 8427 33788 8469 33797
rect 8427 33748 8428 33788
rect 8468 33748 8469 33788
rect 8427 33739 8469 33748
rect 8140 33654 8180 33739
rect 8140 32864 8180 32873
rect 8140 32705 8180 32824
rect 8139 32696 8181 32705
rect 8139 32656 8140 32696
rect 8180 32656 8181 32696
rect 8139 32647 8181 32656
rect 8235 32276 8277 32285
rect 8235 32236 8236 32276
rect 8276 32236 8277 32276
rect 8235 32227 8277 32236
rect 8044 32143 8084 32152
rect 8139 32192 8181 32201
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8236 32192 8276 32227
rect 8140 32058 8180 32143
rect 8236 32141 8276 32152
rect 7947 32024 7989 32033
rect 7852 31984 7948 32024
rect 7988 31984 7989 32024
rect 7947 31975 7989 31984
rect 6892 31529 6932 31614
rect 6316 31469 6356 31480
rect 6507 31520 6549 31529
rect 6507 31480 6508 31520
rect 6548 31480 6549 31520
rect 6507 31471 6549 31480
rect 6891 31520 6933 31529
rect 6891 31480 6892 31520
rect 6932 31480 6933 31520
rect 6891 31471 6933 31480
rect 5451 31436 5493 31445
rect 5451 31396 5452 31436
rect 5492 31396 5493 31436
rect 5451 31387 5493 31396
rect 5452 31352 5492 31387
rect 5452 31301 5492 31312
rect 5932 31357 5972 31366
rect 5932 31277 5972 31317
rect 6412 31352 6452 31361
rect 7084 31352 7124 31361
rect 6452 31312 7084 31352
rect 6412 31303 6452 31312
rect 7084 31303 7124 31312
rect 7756 31352 7796 31361
rect 5931 31268 5973 31277
rect 5931 31228 5932 31268
rect 5972 31228 5973 31268
rect 5931 31219 5973 31228
rect 6123 31184 6165 31193
rect 6123 31144 6124 31184
rect 6164 31144 6165 31184
rect 6123 31135 6165 31144
rect 7659 31184 7701 31193
rect 7659 31144 7660 31184
rect 7700 31144 7701 31184
rect 7659 31135 7701 31144
rect 6124 31050 6164 31135
rect 7563 31100 7605 31109
rect 7563 31060 7564 31100
rect 7604 31060 7605 31100
rect 7563 31051 7605 31060
rect 7564 30848 7604 31051
rect 7564 30799 7604 30808
rect 4395 30176 4437 30185
rect 4395 30136 4396 30176
rect 4436 30136 4437 30176
rect 4395 30127 4437 30136
rect 4203 29924 4245 29933
rect 4203 29884 4204 29924
rect 4244 29884 4245 29924
rect 4203 29875 4245 29884
rect 4204 29840 4244 29875
rect 4204 29789 4244 29800
rect 4300 29840 4340 29851
rect 4300 29765 4340 29800
rect 4396 29840 4436 30127
rect 4588 30101 4628 30631
rect 4972 30546 5012 30631
rect 5068 30269 5108 30640
rect 5355 30680 5397 30689
rect 5355 30640 5356 30680
rect 5396 30640 5397 30680
rect 5355 30631 5397 30640
rect 5547 30680 5589 30689
rect 5547 30640 5548 30680
rect 5588 30640 5589 30680
rect 5547 30631 5589 30640
rect 5836 30680 5876 30689
rect 5356 30512 5396 30521
rect 5396 30472 5492 30512
rect 5356 30463 5396 30472
rect 4875 30260 4917 30269
rect 4875 30220 4876 30260
rect 4916 30220 4917 30260
rect 4875 30211 4917 30220
rect 5067 30260 5109 30269
rect 5067 30220 5068 30260
rect 5108 30220 5109 30260
rect 5067 30211 5109 30220
rect 5355 30260 5397 30269
rect 5355 30220 5356 30260
rect 5396 30220 5397 30260
rect 5355 30211 5397 30220
rect 4683 30176 4725 30185
rect 4683 30136 4684 30176
rect 4724 30136 4725 30176
rect 4683 30127 4725 30136
rect 4587 30092 4629 30101
rect 4587 30052 4588 30092
rect 4628 30052 4629 30092
rect 4587 30043 4629 30052
rect 4396 29791 4436 29800
rect 4587 29840 4629 29849
rect 4587 29800 4588 29840
rect 4628 29800 4629 29840
rect 4587 29791 4629 29800
rect 4684 29840 4724 30127
rect 4876 30092 4916 30211
rect 4876 30043 4916 30052
rect 5259 30092 5301 30101
rect 5259 30052 5260 30092
rect 5300 30052 5301 30092
rect 5259 30043 5301 30052
rect 5163 29924 5205 29933
rect 5163 29884 5164 29924
rect 5204 29884 5205 29924
rect 5163 29875 5205 29884
rect 4684 29791 4724 29800
rect 4876 29840 4916 29849
rect 5068 29840 5108 29849
rect 4916 29800 5068 29840
rect 4876 29791 4916 29800
rect 5068 29791 5108 29800
rect 5164 29840 5204 29875
rect 4011 29756 4053 29765
rect 4011 29716 4012 29756
rect 4052 29716 4053 29756
rect 4011 29707 4053 29716
rect 4299 29756 4341 29765
rect 4299 29716 4300 29756
rect 4340 29716 4341 29756
rect 4299 29707 4341 29716
rect 4588 29706 4628 29791
rect 5164 29789 5204 29800
rect 5260 29840 5300 30043
rect 5260 29791 5300 29800
rect 5356 29840 5396 30211
rect 5356 29791 5396 29800
rect 4108 29672 4148 29681
rect 3915 29252 3957 29261
rect 3915 29212 3916 29252
rect 3956 29212 3957 29252
rect 3915 29203 3957 29212
rect 3916 29118 3956 29203
rect 4108 29000 4148 29632
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 4875 29252 4917 29261
rect 4875 29212 4876 29252
rect 4916 29212 4917 29252
rect 4875 29203 4917 29212
rect 4588 29168 4628 29177
rect 4588 29000 4628 29128
rect 4876 29118 4916 29203
rect 5260 29168 5300 29177
rect 5452 29168 5492 30472
rect 5300 29128 5492 29168
rect 5260 29119 5300 29128
rect 5548 29000 5588 30631
rect 5836 30269 5876 30640
rect 6028 30680 6068 30691
rect 6220 30680 6260 30689
rect 6028 30605 6068 30640
rect 6124 30640 6220 30680
rect 6027 30596 6069 30605
rect 6027 30556 6028 30596
rect 6068 30556 6069 30596
rect 6027 30547 6069 30556
rect 5835 30260 5877 30269
rect 5835 30220 5836 30260
rect 5876 30220 5877 30260
rect 5835 30211 5877 30220
rect 6124 29840 6164 30640
rect 6220 30631 6260 30640
rect 6315 30680 6357 30689
rect 6315 30640 6316 30680
rect 6356 30640 6357 30680
rect 6315 30631 6357 30640
rect 6412 30680 6452 30689
rect 6316 30546 6356 30631
rect 6412 30092 6452 30640
rect 6508 30680 6548 30689
rect 6508 30605 6548 30640
rect 7563 30680 7605 30689
rect 7563 30640 7564 30680
rect 7604 30640 7605 30680
rect 7563 30631 7605 30640
rect 6507 30596 6549 30605
rect 6507 30556 6508 30596
rect 6548 30556 6549 30596
rect 6507 30547 6549 30556
rect 6508 30260 6548 30547
rect 6508 30220 6644 30260
rect 6604 30101 6644 30220
rect 6508 30092 6548 30101
rect 6412 30052 6508 30092
rect 6508 30043 6548 30052
rect 6603 30092 6645 30101
rect 6603 30052 6604 30092
rect 6644 30052 6645 30092
rect 6603 30043 6645 30052
rect 6316 29840 6356 29849
rect 6604 29840 6644 30043
rect 6028 29800 6164 29840
rect 6220 29800 6316 29840
rect 5644 29672 5684 29681
rect 5644 29261 5684 29632
rect 5643 29252 5685 29261
rect 5643 29212 5644 29252
rect 5684 29212 5685 29252
rect 5643 29203 5685 29212
rect 3820 28960 3956 29000
rect 3532 28531 3572 28540
rect 2708 28288 2804 28328
rect 2860 28328 2900 28337
rect 2668 28279 2708 28288
rect 2860 27665 2900 28288
rect 3819 28328 3861 28337
rect 3819 28288 3820 28328
rect 3860 28288 3861 28328
rect 3819 28279 3861 28288
rect 3820 28194 3860 28279
rect 2955 27740 2997 27749
rect 2955 27700 2956 27740
rect 2996 27700 2997 27740
rect 2955 27691 2997 27700
rect 1612 27607 1652 27616
rect 2475 27656 2517 27665
rect 2475 27616 2476 27656
rect 2516 27616 2517 27656
rect 2475 27607 2517 27616
rect 2571 27656 2613 27665
rect 2571 27616 2572 27656
rect 2612 27616 2613 27656
rect 2571 27607 2613 27616
rect 2859 27656 2901 27665
rect 2859 27616 2860 27656
rect 2900 27616 2901 27656
rect 2859 27607 2901 27616
rect 2476 27522 2516 27607
rect 2188 26984 2228 26993
rect 1227 26900 1269 26909
rect 1227 26860 1228 26900
rect 1268 26860 1269 26900
rect 1227 26851 1269 26860
rect 1899 26732 1941 26741
rect 1899 26692 1900 26732
rect 1940 26692 1941 26732
rect 1899 26683 1941 26692
rect 1707 26648 1749 26657
rect 1707 26608 1708 26648
rect 1748 26608 1749 26648
rect 1707 26599 1749 26608
rect 843 26396 885 26405
rect 843 26356 844 26396
rect 884 26356 885 26396
rect 843 26347 885 26356
rect 844 24800 884 26347
rect 1708 26228 1748 26599
rect 1708 26179 1748 26188
rect 1516 25976 1556 25985
rect 1420 25304 1460 25313
rect 1516 25304 1556 25936
rect 1460 25264 1556 25304
rect 1420 25255 1460 25264
rect 1036 25220 1076 25229
rect 1036 24809 1076 25180
rect 844 24751 884 24760
rect 1035 24800 1077 24809
rect 1035 24760 1036 24800
rect 1076 24760 1077 24800
rect 1035 24751 1077 24760
rect 939 24716 981 24725
rect 939 24676 940 24716
rect 980 24676 981 24716
rect 939 24667 981 24676
rect 940 24632 980 24667
rect 940 24581 980 24592
rect 1900 24632 1940 26683
rect 2092 26144 2132 26153
rect 2188 26144 2228 26944
rect 2572 26489 2612 27607
rect 2763 27068 2805 27077
rect 2763 27028 2764 27068
rect 2804 27028 2805 27068
rect 2763 27019 2805 27028
rect 2764 26934 2804 27019
rect 2860 26816 2900 26825
rect 2956 26816 2996 27691
rect 3820 27656 3860 27665
rect 3627 27572 3669 27581
rect 3627 27532 3628 27572
rect 3668 27532 3669 27572
rect 3627 27523 3669 27532
rect 3628 27438 3668 27523
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3820 27077 3860 27616
rect 3916 27656 3956 28960
rect 4012 28960 4148 29000
rect 4204 28960 4628 29000
rect 5164 28960 5588 29000
rect 4012 27656 4052 28960
rect 4108 28160 4148 28169
rect 4108 27833 4148 28120
rect 4107 27824 4149 27833
rect 4107 27784 4108 27824
rect 4148 27784 4149 27824
rect 4107 27775 4149 27784
rect 4108 27656 4148 27665
rect 4012 27616 4108 27656
rect 3916 27607 3956 27616
rect 4108 27607 4148 27616
rect 4108 27488 4148 27497
rect 4204 27488 4244 28960
rect 4875 28496 4917 28505
rect 4875 28456 4876 28496
rect 4916 28456 4917 28496
rect 4875 28447 4917 28456
rect 4780 28328 4820 28337
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4148 27448 4244 27488
rect 4492 27656 4532 27665
rect 4108 27439 4148 27448
rect 3915 27404 3957 27413
rect 3915 27364 3916 27404
rect 3956 27364 3957 27404
rect 3915 27355 3957 27364
rect 3819 27068 3861 27077
rect 3819 27028 3820 27068
rect 3860 27028 3861 27068
rect 3819 27019 3861 27028
rect 2900 26776 2996 26816
rect 3148 26816 3188 26825
rect 2860 26767 2900 26776
rect 3052 26648 3092 26657
rect 2283 26480 2325 26489
rect 2283 26440 2284 26480
rect 2324 26440 2325 26480
rect 2283 26431 2325 26440
rect 2571 26480 2613 26489
rect 2571 26440 2572 26480
rect 2612 26440 2613 26480
rect 2571 26431 2613 26440
rect 2955 26480 2997 26489
rect 2955 26440 2956 26480
rect 2996 26440 2997 26480
rect 2955 26431 2997 26440
rect 2132 26104 2228 26144
rect 2092 26095 2132 26104
rect 2187 25892 2229 25901
rect 2187 25852 2188 25892
rect 2228 25852 2229 25892
rect 2187 25843 2229 25852
rect 1995 24800 2037 24809
rect 1995 24760 1996 24800
rect 2036 24760 2037 24800
rect 1995 24751 2037 24760
rect 1996 24666 2036 24751
rect 1900 24583 1940 24592
rect 2091 24632 2133 24641
rect 2091 24592 2092 24632
rect 2132 24592 2133 24632
rect 2091 24583 2133 24592
rect 2188 24632 2228 25843
rect 2188 24583 2228 24592
rect 2284 25304 2324 26431
rect 2956 26144 2996 26431
rect 2956 26095 2996 26104
rect 3052 25901 3092 26608
rect 3148 26489 3188 26776
rect 3340 26816 3380 26825
rect 3147 26480 3189 26489
rect 3147 26440 3148 26480
rect 3188 26440 3189 26480
rect 3147 26431 3189 26440
rect 3340 26405 3380 26776
rect 3436 26816 3476 26825
rect 3436 26573 3476 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 3916 26816 3956 27355
rect 4492 27329 4532 27616
rect 4780 27581 4820 28288
rect 4779 27572 4821 27581
rect 4779 27532 4780 27572
rect 4820 27532 4821 27572
rect 4779 27523 4821 27532
rect 4683 27404 4725 27413
rect 4683 27364 4684 27404
rect 4724 27364 4725 27404
rect 4683 27355 4725 27364
rect 4491 27320 4533 27329
rect 4491 27280 4492 27320
rect 4532 27280 4533 27320
rect 4491 27271 4533 27280
rect 3916 26767 3956 26776
rect 4012 26944 4244 26984
rect 4012 26816 4052 26944
rect 4012 26767 4052 26776
rect 4108 26816 4148 26825
rect 3628 26682 3668 26767
rect 3819 26732 3861 26741
rect 3819 26692 3820 26732
rect 3860 26692 3861 26732
rect 3819 26683 3861 26692
rect 3531 26648 3573 26657
rect 3531 26608 3532 26648
rect 3572 26608 3573 26648
rect 3531 26599 3573 26608
rect 3435 26564 3477 26573
rect 3435 26524 3436 26564
rect 3476 26524 3477 26564
rect 3435 26515 3477 26524
rect 3532 26514 3572 26599
rect 3820 26598 3860 26683
rect 3627 26480 3669 26489
rect 3627 26440 3628 26480
rect 3668 26440 3669 26480
rect 3627 26431 3669 26440
rect 3339 26396 3381 26405
rect 3339 26356 3340 26396
rect 3380 26356 3381 26396
rect 3339 26347 3381 26356
rect 3051 25892 3093 25901
rect 3051 25852 3052 25892
rect 3092 25852 3093 25892
rect 3051 25843 3093 25852
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3435 25556 3477 25565
rect 3435 25516 3436 25556
rect 3476 25516 3477 25556
rect 3435 25507 3477 25516
rect 3436 25422 3476 25507
rect 2092 24498 2132 24583
rect 1324 24464 1364 24473
rect 1324 23960 1364 24424
rect 1708 24464 1748 24473
rect 1611 24380 1653 24389
rect 1611 24340 1612 24380
rect 1652 24340 1653 24380
rect 1611 24331 1653 24340
rect 1324 23920 1556 23960
rect 1516 23792 1556 23920
rect 1516 23743 1556 23752
rect 1131 23708 1173 23717
rect 1131 23668 1132 23708
rect 1172 23668 1173 23708
rect 1131 23659 1173 23668
rect 1132 23574 1172 23659
rect 1420 23204 1460 23213
rect 1612 23204 1652 24331
rect 1708 23960 1748 24424
rect 2284 23960 2324 25264
rect 3628 25229 3668 26431
rect 4108 26228 4148 26776
rect 4012 26188 4148 26228
rect 2475 25220 2517 25229
rect 2475 25180 2476 25220
rect 2516 25180 2517 25220
rect 2475 25171 2517 25180
rect 3627 25220 3669 25229
rect 3627 25180 3628 25220
rect 3668 25180 3669 25220
rect 3627 25171 3669 25180
rect 3915 25220 3957 25229
rect 3915 25180 3916 25220
rect 3956 25180 3957 25220
rect 3915 25171 3957 25180
rect 2379 24632 2421 24641
rect 2379 24592 2380 24632
rect 2420 24592 2421 24632
rect 2379 24583 2421 24592
rect 2476 24632 2516 25171
rect 3628 25086 3668 25171
rect 2476 24583 2516 24592
rect 2572 24632 2612 24643
rect 2380 24137 2420 24583
rect 2572 24557 2612 24592
rect 2667 24632 2709 24641
rect 2667 24592 2668 24632
rect 2708 24592 2709 24632
rect 2667 24583 2709 24592
rect 3532 24632 3572 24641
rect 3916 24632 3956 25171
rect 4012 25145 4052 26188
rect 4204 26144 4244 26944
rect 4395 26816 4437 26825
rect 4395 26776 4396 26816
rect 4436 26776 4437 26816
rect 4395 26767 4437 26776
rect 4492 26816 4532 27271
rect 4684 27270 4724 27355
rect 4876 27068 4916 28447
rect 4492 26767 4532 26776
rect 4588 27028 4876 27068
rect 4588 26816 4628 27028
rect 4876 27019 4916 27028
rect 4972 28328 5012 28337
rect 4588 26767 4628 26776
rect 4684 26816 4724 26827
rect 4396 26682 4436 26767
rect 4684 26741 4724 26776
rect 4972 26741 5012 28288
rect 5068 28328 5108 28337
rect 5068 27749 5108 28288
rect 5164 28328 5204 28960
rect 5931 28916 5973 28925
rect 5931 28876 5932 28916
rect 5972 28876 5973 28916
rect 5931 28867 5973 28876
rect 5451 28496 5493 28505
rect 5451 28456 5452 28496
rect 5492 28456 5493 28496
rect 5451 28447 5493 28456
rect 5067 27740 5109 27749
rect 5067 27700 5068 27740
rect 5108 27700 5109 27740
rect 5164 27740 5204 28288
rect 5452 28328 5492 28447
rect 5835 28412 5877 28421
rect 5835 28372 5836 28412
rect 5876 28372 5877 28412
rect 5835 28363 5877 28372
rect 5452 28279 5492 28288
rect 5836 28328 5876 28363
rect 5836 28277 5876 28288
rect 5260 28160 5300 28169
rect 5260 27917 5300 28120
rect 5548 28160 5588 28169
rect 5259 27908 5301 27917
rect 5259 27868 5260 27908
rect 5300 27868 5301 27908
rect 5259 27859 5301 27868
rect 5548 27749 5588 28120
rect 5740 28160 5780 28169
rect 5780 28120 5876 28160
rect 5740 28111 5780 28120
rect 5739 27908 5781 27917
rect 5739 27868 5740 27908
rect 5780 27868 5781 27908
rect 5739 27859 5781 27868
rect 5260 27740 5300 27749
rect 5164 27700 5260 27740
rect 5067 27691 5109 27700
rect 4683 26732 4725 26741
rect 4683 26692 4684 26732
rect 4724 26692 4725 26732
rect 4683 26683 4725 26692
rect 4971 26732 5013 26741
rect 4971 26692 4972 26732
rect 5012 26692 5013 26732
rect 4971 26683 5013 26692
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4396 26144 4436 26153
rect 4684 26144 4724 26153
rect 4204 26104 4396 26144
rect 4436 26104 4684 26144
rect 4396 26095 4436 26104
rect 4684 26095 4724 26104
rect 4107 26060 4149 26069
rect 4107 26020 4108 26060
rect 4148 26020 4149 26060
rect 4107 26011 4149 26020
rect 4108 25926 4148 26011
rect 4492 25892 4532 25901
rect 4203 25304 4245 25313
rect 4203 25264 4204 25304
rect 4244 25264 4245 25304
rect 4203 25255 4245 25264
rect 4300 25304 4340 25315
rect 4011 25136 4053 25145
rect 4011 25096 4012 25136
rect 4052 25096 4053 25136
rect 4011 25087 4053 25096
rect 4011 24800 4053 24809
rect 4011 24760 4012 24800
rect 4052 24760 4053 24800
rect 4011 24751 4053 24760
rect 4204 24800 4244 25255
rect 4300 25229 4340 25264
rect 4299 25220 4341 25229
rect 4299 25180 4300 25220
rect 4340 25180 4341 25220
rect 4299 25171 4341 25180
rect 4492 25145 4532 25852
rect 4588 25304 4628 25315
rect 4588 25229 4628 25264
rect 4587 25220 4629 25229
rect 4587 25180 4588 25220
rect 4628 25180 4629 25220
rect 4587 25171 4629 25180
rect 4779 25220 4821 25229
rect 4779 25180 4780 25220
rect 4820 25180 4821 25220
rect 4779 25171 4821 25180
rect 4491 25136 4533 25145
rect 4491 25096 4492 25136
rect 4532 25096 4533 25136
rect 4491 25087 4533 25096
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4204 24751 4244 24760
rect 2571 24548 2613 24557
rect 2571 24508 2572 24548
rect 2612 24508 2613 24548
rect 2571 24499 2613 24508
rect 2668 24498 2708 24583
rect 2859 24380 2901 24389
rect 2859 24340 2860 24380
rect 2900 24340 2901 24380
rect 2859 24331 2901 24340
rect 2860 24246 2900 24331
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 2379 24128 2421 24137
rect 2379 24088 2380 24128
rect 2420 24088 2421 24128
rect 2379 24079 2421 24088
rect 3532 24053 3572 24592
rect 3628 24592 3916 24632
rect 3531 24044 3573 24053
rect 3531 24004 3532 24044
rect 3572 24004 3573 24044
rect 3531 23995 3573 24004
rect 2667 23960 2709 23969
rect 1708 23920 1844 23960
rect 2284 23920 2420 23960
rect 1460 23164 1652 23204
rect 1420 23155 1460 23164
rect 1804 23120 1844 23920
rect 2380 23792 2420 23920
rect 2667 23920 2668 23960
rect 2708 23920 2709 23960
rect 2667 23911 2709 23920
rect 2380 23743 2420 23752
rect 1804 23071 1844 23080
rect 2668 23120 2708 23911
rect 3532 23876 3572 23885
rect 3628 23876 3668 24592
rect 3916 24583 3956 24592
rect 4012 24632 4052 24751
rect 4395 24716 4437 24725
rect 4395 24676 4396 24716
rect 4436 24676 4437 24716
rect 4395 24667 4437 24676
rect 4012 24583 4052 24592
rect 4108 24632 4148 24641
rect 4108 24221 4148 24592
rect 4396 24582 4436 24667
rect 4587 24632 4629 24641
rect 4587 24592 4588 24632
rect 4628 24592 4629 24632
rect 4587 24583 4629 24592
rect 4107 24212 4149 24221
rect 4107 24172 4108 24212
rect 4148 24172 4149 24212
rect 4107 24163 4149 24172
rect 4011 24044 4053 24053
rect 4011 24004 4012 24044
rect 4052 24004 4053 24044
rect 4011 23995 4053 24004
rect 4203 24044 4245 24053
rect 4203 24004 4204 24044
rect 4244 24004 4245 24044
rect 4203 23995 4245 24004
rect 4012 23960 4052 23995
rect 4012 23909 4052 23920
rect 3572 23836 3668 23876
rect 3532 23827 3572 23836
rect 3723 23792 3765 23801
rect 3723 23752 3724 23792
rect 3764 23752 3765 23792
rect 3723 23743 3765 23752
rect 3820 23792 3860 23801
rect 3724 23658 3764 23743
rect 3820 23549 3860 23752
rect 4012 23792 4052 23801
rect 3819 23540 3861 23549
rect 3819 23500 3820 23540
rect 3860 23500 3861 23540
rect 3819 23491 3861 23500
rect 3819 23288 3861 23297
rect 3819 23248 3820 23288
rect 3860 23248 3861 23288
rect 3819 23239 3861 23248
rect 3820 23154 3860 23239
rect 2708 23080 2996 23120
rect 2668 23071 2708 23080
rect 652 23036 692 23045
rect 652 22457 692 22996
rect 844 22868 884 22877
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 652 22112 692 22121
rect 652 21617 692 22072
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 267 20936 309 20945
rect 267 20896 268 20936
rect 308 20896 309 20936
rect 267 20887 309 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 652 20600 692 20719
rect 652 20551 692 20560
rect 652 20264 692 20273
rect 652 19937 692 20224
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18954 692 19039
rect 844 18845 884 22828
rect 1516 22448 1556 22457
rect 1556 22408 2420 22448
rect 1516 22399 1556 22408
rect 2092 22280 2132 22289
rect 1900 22240 2092 22280
rect 1707 22196 1749 22205
rect 1707 22156 1708 22196
rect 1748 22156 1749 22196
rect 1707 22147 1749 22156
rect 1708 22062 1748 22147
rect 1900 21440 1940 22240
rect 2092 22231 2132 22240
rect 2092 21608 2132 21617
rect 2380 21608 2420 22408
rect 2956 22280 2996 23080
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4012 22289 4052 23752
rect 4204 23792 4244 23995
rect 4204 23743 4244 23752
rect 4300 23792 4340 23801
rect 4300 23624 4340 23752
rect 4588 23792 4628 24583
rect 4780 24473 4820 25171
rect 5163 25052 5205 25061
rect 5163 25012 5164 25052
rect 5204 25012 5205 25052
rect 5163 25003 5205 25012
rect 5164 24809 5204 25003
rect 5163 24800 5205 24809
rect 5163 24760 5164 24800
rect 5204 24760 5205 24800
rect 5163 24751 5205 24760
rect 5068 24632 5108 24641
rect 4779 24464 4821 24473
rect 4779 24424 4780 24464
rect 4820 24424 4821 24464
rect 4779 24415 4821 24424
rect 4780 24053 4820 24415
rect 4779 24044 4821 24053
rect 4779 24004 4780 24044
rect 4820 24004 4821 24044
rect 4779 23995 4821 24004
rect 4588 23743 4628 23752
rect 4684 23717 4724 23802
rect 4780 23792 4820 23995
rect 4683 23708 4725 23717
rect 4683 23668 4684 23708
rect 4724 23668 4725 23708
rect 4683 23659 4725 23668
rect 4204 23584 4340 23624
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4108 22532 4148 23071
rect 4108 22483 4148 22492
rect 4011 22280 4053 22289
rect 2996 22240 3380 22280
rect 2956 22231 2996 22240
rect 2476 21608 2516 21617
rect 2380 21568 2476 21608
rect 2092 21449 2132 21568
rect 2476 21559 2516 21568
rect 3340 21608 3380 22240
rect 4011 22240 4012 22280
rect 4052 22240 4053 22280
rect 4011 22231 4053 22240
rect 3340 21559 3380 21568
rect 1900 21391 1940 21400
rect 2091 21440 2133 21449
rect 2091 21400 2092 21440
rect 2132 21400 2133 21440
rect 2091 21391 2133 21400
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4204 21020 4244 23584
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 4491 23288 4533 23297
rect 4780 23288 4820 23752
rect 4875 23792 4917 23801
rect 4875 23752 4876 23792
rect 4916 23752 4917 23792
rect 4875 23743 4917 23752
rect 4876 23658 4916 23743
rect 5068 23297 5108 24592
rect 5164 24212 5204 24751
rect 5260 24557 5300 27700
rect 5547 27740 5589 27749
rect 5547 27700 5548 27740
rect 5588 27700 5589 27740
rect 5547 27691 5589 27700
rect 5644 27656 5684 27665
rect 5548 26816 5588 26825
rect 5451 26732 5493 26741
rect 5451 26692 5452 26732
rect 5492 26692 5493 26732
rect 5451 26683 5493 26692
rect 5355 26144 5397 26153
rect 5355 26104 5356 26144
rect 5396 26104 5397 26144
rect 5355 26095 5397 26104
rect 5356 25565 5396 26095
rect 5355 25556 5397 25565
rect 5355 25516 5356 25556
rect 5396 25516 5397 25556
rect 5355 25507 5397 25516
rect 5452 25304 5492 26683
rect 5548 26069 5588 26776
rect 5644 26144 5684 27616
rect 5740 26816 5780 27859
rect 5836 27488 5876 28120
rect 5932 27656 5972 28867
rect 6028 28328 6068 29800
rect 6123 29168 6165 29177
rect 6123 29128 6124 29168
rect 6164 29128 6165 29168
rect 6123 29119 6165 29128
rect 6124 29034 6164 29119
rect 6124 28580 6164 28589
rect 6220 28580 6260 29800
rect 6316 29791 6356 29800
rect 6412 29800 6644 29840
rect 7180 29840 7220 29849
rect 7468 29840 7508 29849
rect 7220 29800 7316 29840
rect 6412 29000 6452 29800
rect 7180 29791 7220 29800
rect 6164 28540 6260 28580
rect 6316 28960 6452 29000
rect 6508 29672 6548 29681
rect 6124 28531 6164 28540
rect 6124 28328 6164 28337
rect 6028 28288 6124 28328
rect 6124 28279 6164 28288
rect 6316 28328 6356 28960
rect 6508 28673 6548 29632
rect 7276 29093 7316 29800
rect 7372 29672 7412 29681
rect 7275 29084 7317 29093
rect 7275 29044 7276 29084
rect 7316 29044 7317 29084
rect 7275 29035 7317 29044
rect 6507 28664 6549 28673
rect 7372 28664 7412 29632
rect 7468 29345 7508 29800
rect 7467 29336 7509 29345
rect 7467 29296 7468 29336
rect 7508 29296 7509 29336
rect 7467 29287 7509 29296
rect 7564 29177 7604 30631
rect 7563 29168 7605 29177
rect 7563 29128 7564 29168
rect 7604 29128 7605 29168
rect 7563 29119 7605 29128
rect 6507 28624 6508 28664
rect 6548 28624 6549 28664
rect 6507 28615 6549 28624
rect 6604 28624 7412 28664
rect 6316 28279 6356 28288
rect 6412 28328 6452 28337
rect 6604 28328 6644 28624
rect 7564 28496 7604 29119
rect 7468 28456 7604 28496
rect 6700 28337 6740 28368
rect 6452 28288 6644 28328
rect 6699 28328 6741 28337
rect 6699 28288 6700 28328
rect 6740 28288 6741 28328
rect 6412 28279 6452 28288
rect 6699 28279 6741 28288
rect 6700 28244 6740 28279
rect 6603 28160 6645 28169
rect 6603 28120 6604 28160
rect 6644 28120 6645 28160
rect 6603 28111 6645 28120
rect 6028 27665 6068 27750
rect 5932 27607 5972 27616
rect 6027 27656 6069 27665
rect 6027 27616 6028 27656
rect 6068 27616 6069 27656
rect 6027 27607 6069 27616
rect 6604 27656 6644 28111
rect 6604 27607 6644 27616
rect 5836 27448 6068 27488
rect 5835 26900 5877 26909
rect 5835 26860 5836 26900
rect 5876 26860 5877 26900
rect 5835 26851 5877 26860
rect 5740 26767 5780 26776
rect 5836 26732 5876 26851
rect 5932 26816 5972 26827
rect 5932 26741 5972 26776
rect 6028 26816 6068 27448
rect 6316 27404 6356 27413
rect 6028 26767 6068 26776
rect 6220 27364 6316 27404
rect 6220 26816 6260 27364
rect 6316 27355 6356 27364
rect 6508 27404 6548 27413
rect 6412 26909 6452 26940
rect 6411 26900 6453 26909
rect 6411 26860 6412 26900
rect 6452 26860 6453 26900
rect 6411 26851 6453 26860
rect 6220 26767 6260 26776
rect 6412 26816 6452 26851
rect 6508 26825 6548 27364
rect 6700 26900 6740 28204
rect 6796 27656 6836 27665
rect 6796 27161 6836 27616
rect 6892 27656 6932 27665
rect 6892 27413 6932 27616
rect 6988 27656 7028 27665
rect 6891 27404 6933 27413
rect 6891 27364 6892 27404
rect 6932 27364 6933 27404
rect 6891 27355 6933 27364
rect 6988 27329 7028 27616
rect 7083 27656 7125 27665
rect 7083 27616 7084 27656
rect 7124 27616 7125 27656
rect 7083 27607 7125 27616
rect 7084 27522 7124 27607
rect 7275 27404 7317 27413
rect 7275 27364 7276 27404
rect 7316 27364 7317 27404
rect 7275 27355 7317 27364
rect 6987 27320 7029 27329
rect 6987 27280 6988 27320
rect 7028 27280 7029 27320
rect 6987 27271 7029 27280
rect 7276 27270 7316 27355
rect 6795 27152 6837 27161
rect 6795 27112 6796 27152
rect 6836 27112 6837 27152
rect 6795 27103 6837 27112
rect 7468 26909 7508 28456
rect 7563 28328 7605 28337
rect 7563 28288 7564 28328
rect 7604 28288 7605 28328
rect 7563 28279 7605 28288
rect 7564 28194 7604 28279
rect 7563 27152 7605 27161
rect 7563 27112 7564 27152
rect 7604 27112 7605 27152
rect 7563 27103 7605 27112
rect 7467 26900 7509 26909
rect 6700 26860 6836 26900
rect 5836 26683 5876 26692
rect 5931 26732 5973 26741
rect 5931 26692 5932 26732
rect 5972 26692 5973 26732
rect 5931 26683 5973 26692
rect 6316 26732 6356 26741
rect 6316 26573 6356 26692
rect 6315 26564 6357 26573
rect 6315 26524 6316 26564
rect 6356 26524 6357 26564
rect 6315 26515 6357 26524
rect 5931 26396 5973 26405
rect 5931 26356 5932 26396
rect 5972 26356 5973 26396
rect 5931 26347 5973 26356
rect 5836 26144 5876 26153
rect 5644 26104 5836 26144
rect 5547 26060 5589 26069
rect 5547 26020 5548 26060
rect 5588 26020 5589 26060
rect 5547 26011 5589 26020
rect 5452 25255 5492 25264
rect 5836 25078 5876 26104
rect 5932 25304 5972 26347
rect 6123 26144 6165 26153
rect 6123 26104 6124 26144
rect 6164 26104 6165 26144
rect 6123 26095 6165 26104
rect 6220 26144 6260 26155
rect 6124 26010 6164 26095
rect 6220 26069 6260 26104
rect 6219 26060 6261 26069
rect 6219 26020 6220 26060
rect 6260 26020 6261 26060
rect 6219 26011 6261 26020
rect 6315 25556 6357 25565
rect 6315 25516 6316 25556
rect 6356 25516 6357 25556
rect 6315 25507 6357 25516
rect 6316 25422 6356 25507
rect 5932 25255 5972 25264
rect 6027 25304 6069 25313
rect 6412 25304 6452 26776
rect 6507 26816 6549 26825
rect 6507 26776 6508 26816
rect 6548 26776 6549 26816
rect 6507 26767 6549 26776
rect 6699 26732 6741 26741
rect 6699 26692 6700 26732
rect 6740 26692 6741 26732
rect 6699 26683 6741 26692
rect 6507 26648 6549 26657
rect 6507 26608 6508 26648
rect 6548 26608 6549 26648
rect 6507 26599 6549 26608
rect 6508 25976 6548 26599
rect 6700 26598 6740 26683
rect 6603 26312 6645 26321
rect 6603 26272 6604 26312
rect 6644 26272 6645 26312
rect 6603 26263 6645 26272
rect 6508 25927 6548 25936
rect 6027 25264 6028 25304
rect 6068 25264 6069 25304
rect 6027 25255 6069 25264
rect 6316 25264 6452 25304
rect 6028 25170 6068 25255
rect 5931 25136 5973 25145
rect 5931 25096 5932 25136
rect 5972 25096 5973 25136
rect 5931 25087 5973 25096
rect 6219 25136 6261 25145
rect 6219 25096 6220 25136
rect 6260 25096 6261 25136
rect 6219 25087 6261 25096
rect 5835 25012 5836 25061
rect 5876 25012 5877 25061
rect 5835 25003 5877 25012
rect 5452 24760 5876 24800
rect 5452 24632 5492 24760
rect 5452 24583 5492 24592
rect 5548 24632 5588 24641
rect 5259 24548 5301 24557
rect 5259 24508 5260 24548
rect 5300 24508 5301 24548
rect 5259 24499 5301 24508
rect 5260 24389 5300 24499
rect 5259 24380 5301 24389
rect 5259 24340 5260 24380
rect 5300 24340 5301 24380
rect 5259 24331 5301 24340
rect 5355 24212 5397 24221
rect 5164 24172 5300 24212
rect 5164 23792 5204 23801
rect 4491 23248 4492 23288
rect 4532 23248 4533 23288
rect 4491 23239 4533 23248
rect 4588 23248 4820 23288
rect 5067 23288 5109 23297
rect 5067 23248 5068 23288
rect 5108 23248 5109 23288
rect 4395 22364 4437 22373
rect 4395 22324 4396 22364
rect 4436 22324 4437 22364
rect 4395 22315 4437 22324
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4396 22280 4436 22315
rect 4300 22146 4340 22231
rect 4396 22229 4436 22240
rect 4492 22280 4532 23239
rect 4492 22231 4532 22240
rect 4588 22280 4628 23248
rect 5067 23239 5109 23248
rect 4972 23120 5012 23129
rect 5164 23120 5204 23752
rect 5012 23080 5204 23120
rect 5260 23792 5300 24172
rect 5355 24172 5356 24212
rect 5396 24172 5397 24212
rect 5355 24163 5397 24172
rect 4779 22868 4821 22877
rect 4779 22828 4780 22868
rect 4820 22828 4821 22868
rect 4779 22819 4821 22828
rect 4780 22734 4820 22819
rect 4972 22709 5012 23080
rect 5260 22793 5300 23752
rect 5356 23792 5396 24163
rect 5356 23743 5396 23752
rect 5452 23792 5492 23801
rect 5548 23792 5588 24592
rect 5644 24632 5684 24643
rect 5644 24557 5684 24592
rect 5739 24632 5781 24641
rect 5739 24592 5740 24632
rect 5780 24592 5781 24632
rect 5739 24583 5781 24592
rect 5643 24548 5685 24557
rect 5643 24508 5644 24548
rect 5684 24508 5685 24548
rect 5643 24499 5685 24508
rect 5740 24498 5780 24583
rect 5643 24380 5685 24389
rect 5643 24340 5644 24380
rect 5684 24340 5685 24380
rect 5643 24331 5685 24340
rect 5492 23752 5588 23792
rect 5452 23743 5492 23752
rect 5644 23708 5684 24331
rect 5548 23668 5684 23708
rect 5548 22868 5588 23668
rect 5643 23540 5685 23549
rect 5643 23500 5644 23540
rect 5684 23500 5685 23540
rect 5643 23491 5685 23500
rect 5644 23288 5684 23491
rect 5836 23288 5876 24760
rect 5932 24632 5972 25087
rect 6123 24716 6165 24725
rect 6123 24676 6124 24716
rect 6164 24676 6165 24716
rect 6123 24667 6165 24676
rect 5932 24583 5972 24592
rect 6028 24632 6068 24641
rect 6028 24473 6068 24592
rect 6124 24582 6164 24667
rect 6220 24632 6260 25087
rect 6220 24583 6260 24592
rect 6027 24464 6069 24473
rect 6027 24424 6028 24464
rect 6068 24424 6069 24464
rect 6027 24415 6069 24424
rect 6316 24221 6356 25264
rect 6507 25052 6549 25061
rect 6507 25012 6508 25052
rect 6548 25012 6549 25052
rect 6507 25003 6549 25012
rect 6508 24641 6548 25003
rect 6604 24800 6644 26263
rect 6700 25136 6740 25147
rect 6700 25061 6740 25096
rect 6699 25052 6741 25061
rect 6699 25012 6700 25052
rect 6740 25012 6741 25052
rect 6699 25003 6741 25012
rect 6700 24800 6740 24809
rect 6604 24760 6700 24800
rect 6700 24751 6740 24760
rect 6412 24632 6452 24641
rect 6412 24473 6452 24592
rect 6507 24632 6549 24641
rect 6507 24592 6508 24632
rect 6548 24592 6549 24632
rect 6507 24583 6549 24592
rect 6604 24632 6644 24641
rect 6508 24498 6548 24583
rect 6411 24464 6453 24473
rect 6411 24424 6412 24464
rect 6452 24424 6453 24464
rect 6411 24415 6453 24424
rect 6604 24389 6644 24592
rect 6603 24380 6645 24389
rect 6603 24340 6604 24380
rect 6644 24340 6645 24380
rect 6603 24331 6645 24340
rect 6315 24212 6357 24221
rect 6315 24172 6316 24212
rect 6356 24172 6357 24212
rect 6315 24163 6357 24172
rect 6123 23960 6165 23969
rect 6123 23920 6124 23960
rect 6164 23920 6165 23960
rect 6123 23911 6165 23920
rect 6124 23826 6164 23911
rect 6604 23792 6644 23801
rect 6796 23792 6836 26860
rect 7467 26860 7468 26900
rect 7508 26860 7509 26900
rect 7467 26851 7509 26860
rect 7564 26816 7604 27103
rect 7564 26767 7604 26776
rect 7084 26648 7124 26657
rect 7084 26489 7124 26608
rect 7083 26480 7125 26489
rect 7083 26440 7084 26480
rect 7124 26440 7125 26480
rect 7083 26431 7125 26440
rect 6892 26144 6932 26153
rect 6892 25985 6932 26104
rect 6891 25976 6933 25985
rect 6891 25936 6892 25976
rect 6932 25936 6933 25976
rect 6891 25927 6933 25936
rect 7564 25892 7604 25901
rect 7564 25313 7604 25852
rect 7563 25304 7605 25313
rect 7563 25264 7564 25304
rect 7604 25264 7605 25304
rect 7563 25255 7605 25264
rect 7563 24716 7605 24725
rect 7563 24676 7564 24716
rect 7604 24676 7605 24716
rect 7563 24667 7605 24676
rect 7564 24632 7604 24667
rect 7660 24632 7700 31135
rect 7756 31109 7796 31312
rect 7755 31100 7797 31109
rect 7755 31060 7756 31100
rect 7796 31060 7797 31100
rect 7755 31051 7797 31060
rect 7852 30008 7892 30017
rect 7755 29924 7797 29933
rect 7755 29884 7756 29924
rect 7796 29884 7797 29924
rect 7755 29875 7797 29884
rect 7756 27908 7796 29875
rect 7852 29000 7892 29968
rect 7948 29336 7988 31975
rect 8043 31268 8085 31277
rect 8043 31228 8044 31268
rect 8084 31228 8085 31268
rect 8043 31219 8085 31228
rect 8044 30689 8084 31219
rect 8043 30680 8085 30689
rect 8043 30640 8044 30680
rect 8084 30640 8085 30680
rect 8043 30631 8085 30640
rect 8043 30092 8085 30101
rect 8043 30052 8044 30092
rect 8084 30052 8085 30092
rect 8043 30043 8085 30052
rect 8044 29840 8084 30043
rect 8235 29924 8277 29933
rect 8235 29884 8236 29924
rect 8276 29884 8277 29924
rect 8235 29875 8277 29884
rect 8044 29791 8084 29800
rect 8140 29840 8180 29849
rect 7948 29287 7988 29296
rect 7852 28960 7988 29000
rect 7851 28412 7893 28421
rect 7851 28372 7852 28412
rect 7892 28372 7893 28412
rect 7851 28363 7893 28372
rect 7852 28278 7892 28363
rect 7756 27868 7892 27908
rect 7755 27740 7797 27749
rect 7755 27700 7756 27740
rect 7796 27700 7797 27740
rect 7755 27691 7797 27700
rect 7756 26564 7796 27691
rect 7852 27329 7892 27868
rect 7948 27497 7988 28960
rect 8140 28169 8180 29800
rect 8236 29840 8276 29875
rect 8236 29789 8276 29800
rect 8331 29840 8373 29849
rect 8331 29800 8332 29840
rect 8372 29800 8373 29840
rect 8331 29791 8373 29800
rect 8332 29706 8372 29791
rect 8428 29504 8468 33739
rect 8716 32705 8756 34336
rect 9004 34327 9044 34336
rect 9387 34376 9429 34385
rect 9387 34336 9388 34376
rect 9428 34336 9429 34376
rect 9387 34327 9429 34336
rect 9388 33872 9428 34327
rect 9388 33823 9428 33832
rect 9484 33704 9524 33713
rect 9772 33704 9812 34924
rect 10060 34915 10100 34924
rect 10155 34712 10197 34721
rect 10155 34672 10156 34712
rect 10196 34672 10197 34712
rect 10155 34663 10197 34672
rect 10156 34628 10196 34663
rect 10156 34577 10196 34588
rect 10059 34544 10101 34553
rect 10444 34544 10484 35848
rect 10732 35888 10772 36604
rect 10732 35839 10772 35848
rect 10828 35888 10868 36763
rect 11116 36728 11156 36940
rect 11116 36679 11156 36688
rect 11212 36728 11252 37528
rect 11596 37400 11636 37409
rect 12460 37400 12500 37780
rect 11636 37360 11732 37400
rect 11596 37351 11636 37360
rect 11115 36056 11157 36065
rect 11115 36016 11116 36056
rect 11156 36016 11157 36056
rect 11115 36007 11157 36016
rect 11116 35922 11156 36007
rect 10828 35839 10868 35848
rect 11212 35813 11252 36688
rect 11404 36728 11444 36737
rect 11444 36688 11540 36728
rect 11404 36679 11444 36688
rect 11403 36560 11445 36569
rect 11403 36520 11404 36560
rect 11444 36520 11445 36560
rect 11403 36511 11445 36520
rect 11404 36426 11444 36511
rect 11211 35804 11253 35813
rect 11211 35764 11212 35804
rect 11252 35764 11253 35804
rect 11211 35755 11253 35764
rect 11115 35720 11157 35729
rect 11115 35680 11116 35720
rect 11156 35680 11157 35720
rect 11115 35671 11157 35680
rect 10923 35300 10965 35309
rect 10923 35260 10924 35300
rect 10964 35260 10965 35300
rect 10923 35251 10965 35260
rect 10732 35216 10772 35225
rect 10539 35048 10581 35057
rect 10539 35008 10540 35048
rect 10580 35008 10581 35048
rect 10539 34999 10581 35008
rect 10059 34504 10060 34544
rect 10100 34504 10101 34544
rect 10059 34495 10101 34504
rect 10348 34504 10484 34544
rect 10060 34133 10100 34495
rect 10156 34208 10196 34217
rect 10196 34168 10292 34208
rect 10156 34159 10196 34168
rect 10059 34124 10101 34133
rect 10059 34084 10060 34124
rect 10100 34084 10101 34124
rect 10059 34075 10101 34084
rect 9524 33664 9812 33704
rect 10060 33704 10100 34075
rect 10156 33704 10196 33713
rect 10060 33664 10156 33704
rect 9484 33655 9524 33664
rect 10156 33655 10196 33664
rect 9867 33536 9909 33545
rect 9867 33496 9868 33536
rect 9908 33496 9909 33536
rect 9867 33487 9909 33496
rect 9868 33402 9908 33487
rect 9963 33200 10005 33209
rect 9963 33160 9964 33200
rect 10004 33160 10005 33200
rect 9963 33151 10005 33160
rect 9291 32948 9333 32957
rect 9291 32908 9292 32948
rect 9332 32908 9333 32948
rect 9291 32899 9333 32908
rect 9292 32814 9332 32899
rect 9964 32873 10004 33151
rect 9963 32864 10005 32873
rect 9963 32824 9964 32864
rect 10004 32824 10005 32864
rect 9963 32815 10005 32824
rect 10252 32864 10292 34168
rect 10348 33209 10388 34504
rect 10443 34376 10485 34385
rect 10443 34336 10444 34376
rect 10484 34336 10485 34376
rect 10443 34327 10485 34336
rect 10540 34376 10580 34999
rect 10732 34721 10772 35176
rect 10924 35166 10964 35251
rect 11020 35216 11060 35225
rect 10731 34712 10773 34721
rect 10731 34672 10732 34712
rect 10772 34672 10773 34712
rect 10731 34663 10773 34672
rect 10732 34544 10772 34553
rect 10772 34504 10964 34544
rect 10732 34495 10772 34504
rect 10540 34327 10580 34336
rect 10732 34376 10772 34385
rect 10444 34242 10484 34327
rect 10732 34049 10772 34336
rect 10924 34376 10964 34504
rect 10924 34327 10964 34336
rect 11020 34301 11060 35176
rect 11116 35216 11156 35671
rect 11500 35309 11540 36688
rect 11595 35888 11637 35897
rect 11595 35848 11596 35888
rect 11636 35848 11637 35888
rect 11595 35839 11637 35848
rect 11596 35754 11636 35839
rect 11692 35720 11732 37360
rect 12460 37351 12500 37360
rect 12844 37400 12884 37939
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 12844 37351 12884 37360
rect 13996 37400 14036 37409
rect 13996 37241 14036 37360
rect 16396 37400 16436 37409
rect 13995 37232 14037 37241
rect 13995 37192 13996 37232
rect 14036 37192 14037 37232
rect 13995 37183 14037 37192
rect 14668 37232 14708 37241
rect 15724 37232 15764 37241
rect 14708 37192 14900 37232
rect 14668 37183 14708 37192
rect 11788 36728 11828 36737
rect 11788 36569 11828 36688
rect 13996 36569 14036 37183
rect 14860 36728 14900 37192
rect 15531 36896 15573 36905
rect 15531 36856 15532 36896
rect 15572 36856 15573 36896
rect 15531 36847 15573 36856
rect 15532 36762 15572 36847
rect 14860 36679 14900 36688
rect 14955 36728 14997 36737
rect 14955 36688 14956 36728
rect 14996 36688 14997 36728
rect 14955 36679 14997 36688
rect 15339 36728 15381 36737
rect 15339 36688 15340 36728
rect 15380 36688 15381 36728
rect 15339 36679 15381 36688
rect 15436 36728 15476 36737
rect 14956 36594 14996 36679
rect 15340 36594 15380 36679
rect 11787 36560 11829 36569
rect 12652 36560 12692 36569
rect 11787 36520 11788 36560
rect 11828 36520 11829 36560
rect 11787 36511 11829 36520
rect 12556 36520 12652 36560
rect 12460 36476 12500 36485
rect 11980 36436 12460 36476
rect 11788 35888 11828 35897
rect 11980 35888 12020 36436
rect 12460 36427 12500 36436
rect 11828 35848 11924 35888
rect 11788 35839 11828 35848
rect 11692 35680 11828 35720
rect 11499 35300 11541 35309
rect 11499 35260 11500 35300
rect 11540 35260 11541 35300
rect 11499 35251 11541 35260
rect 11116 35167 11156 35176
rect 11211 35216 11253 35225
rect 11404 35216 11444 35225
rect 11211 35176 11212 35216
rect 11252 35176 11404 35216
rect 11211 35167 11253 35176
rect 11404 35167 11444 35176
rect 11212 35082 11252 35167
rect 11019 34292 11061 34301
rect 11019 34252 11020 34292
rect 11060 34252 11061 34292
rect 11019 34243 11061 34252
rect 10731 34040 10773 34049
rect 10731 34000 10732 34040
rect 10772 34000 10773 34040
rect 10731 33991 10773 34000
rect 11020 33788 11060 34243
rect 11596 34208 11636 34217
rect 11020 33739 11060 33748
rect 11308 34168 11596 34208
rect 11308 33788 11348 34168
rect 11596 34159 11636 34168
rect 11308 33739 11348 33748
rect 11788 33713 11828 35680
rect 11884 35225 11924 35848
rect 11980 35839 12020 35848
rect 12364 35888 12404 35897
rect 12556 35888 12596 36520
rect 12652 36511 12692 36520
rect 13995 36560 14037 36569
rect 13995 36520 13996 36560
rect 14036 36520 14037 36560
rect 13995 36511 14037 36520
rect 14859 36560 14901 36569
rect 14859 36520 14860 36560
rect 14900 36520 14901 36560
rect 14859 36511 14901 36520
rect 14572 36056 14612 36065
rect 13900 36016 14572 36056
rect 12843 35972 12885 35981
rect 12843 35932 12844 35972
rect 12884 35932 12885 35972
rect 12843 35923 12885 35932
rect 12404 35848 12596 35888
rect 12364 35839 12404 35848
rect 11883 35216 11925 35225
rect 11883 35176 11884 35216
rect 11924 35176 11925 35216
rect 11883 35167 11925 35176
rect 12363 35216 12405 35225
rect 12363 35176 12364 35216
rect 12404 35176 12405 35216
rect 12363 35167 12405 35176
rect 12364 35082 12404 35167
rect 11980 34376 12020 34385
rect 11980 34133 12020 34336
rect 12364 34208 12404 34219
rect 12364 34133 12404 34168
rect 11979 34124 12021 34133
rect 11979 34084 11980 34124
rect 12020 34084 12021 34124
rect 11979 34075 12021 34084
rect 12363 34124 12405 34133
rect 12363 34084 12364 34124
rect 12404 34084 12405 34124
rect 12363 34075 12405 34084
rect 11883 34040 11925 34049
rect 11883 34000 11884 34040
rect 11924 34000 11925 34040
rect 11883 33991 11925 34000
rect 11692 33704 11732 33713
rect 11692 33545 11732 33664
rect 11787 33704 11829 33713
rect 11787 33664 11788 33704
rect 11828 33664 11829 33704
rect 11787 33655 11829 33664
rect 11691 33536 11733 33545
rect 11691 33496 11692 33536
rect 11732 33496 11733 33536
rect 11691 33487 11733 33496
rect 10347 33200 10389 33209
rect 10347 33160 10348 33200
rect 10388 33160 10389 33200
rect 10347 33151 10389 33160
rect 10635 33032 10677 33041
rect 10635 32992 10636 33032
rect 10676 32992 10677 33032
rect 10635 32983 10677 32992
rect 10347 32948 10389 32957
rect 10347 32908 10348 32948
rect 10388 32908 10389 32948
rect 10347 32899 10389 32908
rect 10252 32815 10292 32824
rect 10348 32864 10388 32899
rect 10636 32898 10676 32983
rect 11691 32948 11733 32957
rect 11691 32908 11692 32948
rect 11732 32908 11733 32948
rect 11691 32899 11733 32908
rect 8811 32780 8853 32789
rect 8811 32740 8812 32780
rect 8852 32740 8853 32780
rect 8811 32731 8853 32740
rect 8715 32696 8757 32705
rect 8715 32656 8716 32696
rect 8756 32656 8757 32696
rect 8715 32647 8757 32656
rect 8716 30680 8756 32647
rect 8812 32621 8852 32731
rect 9964 32730 10004 32815
rect 8811 32612 8853 32621
rect 8811 32572 8812 32612
rect 8852 32572 8853 32612
rect 8811 32563 8853 32572
rect 8812 31352 8852 32563
rect 9579 32192 9621 32201
rect 9579 32152 9580 32192
rect 9620 32152 9621 32192
rect 9579 32143 9621 32152
rect 10252 32192 10292 32201
rect 10348 32192 10388 32824
rect 10292 32152 10388 32192
rect 10828 32864 10868 32873
rect 10252 32143 10292 32152
rect 9387 32024 9429 32033
rect 9387 31984 9388 32024
rect 9428 31984 9429 32024
rect 9387 31975 9429 31984
rect 9388 31890 9428 31975
rect 9483 31520 9525 31529
rect 9483 31480 9484 31520
rect 9524 31480 9525 31520
rect 9483 31471 9525 31480
rect 8812 31303 8852 31312
rect 9484 30680 9524 31471
rect 9580 31352 9620 32143
rect 10347 32024 10389 32033
rect 10347 31984 10348 32024
rect 10388 31984 10389 32024
rect 10347 31975 10389 31984
rect 10059 31940 10101 31949
rect 10059 31900 10060 31940
rect 10100 31900 10101 31940
rect 10059 31891 10101 31900
rect 9963 31604 10005 31613
rect 9963 31564 9964 31604
rect 10004 31564 10005 31604
rect 9963 31555 10005 31564
rect 9771 31520 9813 31529
rect 9771 31480 9772 31520
rect 9812 31480 9813 31520
rect 9771 31471 9813 31480
rect 9772 31386 9812 31471
rect 9676 31352 9716 31361
rect 9580 31312 9676 31352
rect 9676 31303 9716 31312
rect 9964 31352 10004 31555
rect 9964 31303 10004 31312
rect 9964 30764 10004 30773
rect 10060 30764 10100 31891
rect 10348 31352 10388 31975
rect 10443 31940 10485 31949
rect 10443 31900 10444 31940
rect 10484 31900 10485 31940
rect 10443 31891 10485 31900
rect 10444 31806 10484 31891
rect 10828 31529 10868 32824
rect 10923 32864 10965 32873
rect 10923 32824 10924 32864
rect 10964 32824 10965 32864
rect 10923 32815 10965 32824
rect 11116 32864 11156 32873
rect 11404 32864 11444 32873
rect 11156 32824 11404 32864
rect 11116 32815 11156 32824
rect 11404 32815 11444 32824
rect 11500 32864 11540 32873
rect 10924 32730 10964 32815
rect 11019 32780 11061 32789
rect 11019 32740 11020 32780
rect 11060 32740 11061 32780
rect 11019 32731 11061 32740
rect 11020 32646 11060 32731
rect 11500 32705 11540 32824
rect 11596 32864 11636 32873
rect 11499 32696 11541 32705
rect 11499 32656 11500 32696
rect 11540 32656 11541 32696
rect 11499 32647 11541 32656
rect 11116 32192 11156 32201
rect 10924 32152 11116 32192
rect 10827 31520 10869 31529
rect 10827 31480 10828 31520
rect 10868 31480 10869 31520
rect 10827 31471 10869 31480
rect 10348 31303 10388 31312
rect 10924 30848 10964 32152
rect 11116 32143 11156 32152
rect 11308 31940 11348 31949
rect 11308 31613 11348 31900
rect 11307 31604 11349 31613
rect 11307 31564 11308 31604
rect 11348 31564 11349 31604
rect 11307 31555 11349 31564
rect 11211 31520 11253 31529
rect 11211 31480 11212 31520
rect 11252 31480 11253 31520
rect 11211 31471 11253 31480
rect 11212 31352 11252 31471
rect 11019 31184 11061 31193
rect 11019 31144 11020 31184
rect 11060 31144 11061 31184
rect 11019 31135 11061 31144
rect 10924 30799 10964 30808
rect 10004 30724 10100 30764
rect 9964 30715 10004 30724
rect 9580 30680 9620 30689
rect 9484 30640 9580 30680
rect 8716 30631 8756 30640
rect 9580 30631 9620 30640
rect 10731 30680 10773 30689
rect 10731 30640 10732 30680
rect 10772 30640 10773 30680
rect 10731 30631 10773 30640
rect 10828 30680 10868 30689
rect 10732 30546 10772 30631
rect 9963 30512 10005 30521
rect 9963 30472 9964 30512
rect 10004 30472 10005 30512
rect 9963 30463 10005 30472
rect 8715 30092 8757 30101
rect 8715 30052 8716 30092
rect 8756 30052 8757 30092
rect 8715 30043 8757 30052
rect 8523 29840 8565 29849
rect 8523 29800 8524 29840
rect 8564 29800 8565 29840
rect 8523 29791 8565 29800
rect 8716 29840 8756 30043
rect 9868 30008 9908 30017
rect 8812 29849 8852 29934
rect 8716 29791 8756 29800
rect 8811 29840 8853 29849
rect 8811 29800 8812 29840
rect 8852 29800 8853 29840
rect 8811 29791 8853 29800
rect 9676 29840 9716 29851
rect 8524 29706 8564 29791
rect 9676 29765 9716 29800
rect 8619 29756 8661 29765
rect 8619 29716 8620 29756
rect 8660 29716 8661 29756
rect 8619 29707 8661 29716
rect 9675 29756 9717 29765
rect 9675 29716 9676 29756
rect 9716 29716 9717 29756
rect 9675 29707 9717 29716
rect 8620 29622 8660 29707
rect 9004 29672 9044 29681
rect 8716 29632 9004 29672
rect 8428 29464 8660 29504
rect 8428 29168 8468 29177
rect 8428 28337 8468 29128
rect 8620 28496 8660 29464
rect 8716 29252 8756 29632
rect 9004 29623 9044 29632
rect 8716 29203 8756 29212
rect 9100 29168 9140 29177
rect 9868 29168 9908 29968
rect 9140 29128 9908 29168
rect 9964 29168 10004 30463
rect 10828 30101 10868 30640
rect 11020 30680 11060 31135
rect 11020 30631 11060 30640
rect 11212 30521 11252 31312
rect 11211 30512 11253 30521
rect 11211 30472 11212 30512
rect 11252 30472 11253 30512
rect 11211 30463 11253 30472
rect 11500 30512 11540 32647
rect 11596 31613 11636 32824
rect 11692 32864 11732 32899
rect 11692 32813 11732 32824
rect 11787 32864 11829 32873
rect 11787 32824 11788 32864
rect 11828 32824 11829 32864
rect 11787 32815 11829 32824
rect 11884 32864 11924 33991
rect 11884 32815 11924 32824
rect 11980 32864 12020 34075
rect 12556 33704 12596 33713
rect 12651 33704 12693 33713
rect 12596 33664 12652 33704
rect 12692 33664 12693 33704
rect 12556 33655 12596 33664
rect 12651 33655 12693 33664
rect 12267 33032 12309 33041
rect 12267 32992 12268 33032
rect 12308 32992 12309 33032
rect 12267 32983 12309 32992
rect 12171 32948 12213 32957
rect 12171 32908 12172 32948
rect 12212 32908 12213 32948
rect 12171 32899 12213 32908
rect 11788 32192 11828 32815
rect 11980 32705 12020 32824
rect 12076 32864 12116 32875
rect 12076 32789 12116 32824
rect 12172 32864 12212 32899
rect 12075 32780 12117 32789
rect 12075 32740 12076 32780
rect 12116 32740 12117 32780
rect 12075 32731 12117 32740
rect 11979 32696 12021 32705
rect 11979 32656 11980 32696
rect 12020 32656 12021 32696
rect 11979 32647 12021 32656
rect 12172 32360 12212 32824
rect 12076 32320 12212 32360
rect 11980 32192 12020 32201
rect 11788 32152 11980 32192
rect 11980 32143 12020 32152
rect 11595 31604 11637 31613
rect 11595 31564 11596 31604
rect 11636 31564 11637 31604
rect 11595 31555 11637 31564
rect 12076 31277 12116 32320
rect 12172 32192 12212 32201
rect 12268 32192 12308 32983
rect 12556 32873 12596 32958
rect 12652 32948 12692 33655
rect 12748 32948 12788 32957
rect 12652 32908 12748 32948
rect 12555 32864 12597 32873
rect 12555 32824 12556 32864
rect 12596 32824 12597 32864
rect 12555 32815 12597 32824
rect 12460 32696 12500 32705
rect 12652 32696 12692 32908
rect 12748 32899 12788 32908
rect 12363 32612 12405 32621
rect 12363 32572 12364 32612
rect 12404 32572 12405 32612
rect 12363 32563 12405 32572
rect 12364 32285 12404 32563
rect 12363 32276 12405 32285
rect 12363 32236 12364 32276
rect 12404 32236 12405 32276
rect 12363 32227 12405 32236
rect 12212 32152 12308 32192
rect 12364 32192 12404 32227
rect 12172 32143 12212 32152
rect 12364 32141 12404 32152
rect 12267 31940 12309 31949
rect 12267 31900 12268 31940
rect 12308 31900 12309 31940
rect 12267 31891 12309 31900
rect 12268 31806 12308 31891
rect 12363 31604 12405 31613
rect 12363 31564 12364 31604
rect 12404 31564 12405 31604
rect 12363 31555 12405 31564
rect 12364 31520 12404 31555
rect 12364 31469 12404 31480
rect 12460 31445 12500 32656
rect 12556 32656 12692 32696
rect 12556 31529 12596 32656
rect 12747 32192 12789 32201
rect 12747 32152 12748 32192
rect 12788 32152 12789 32192
rect 12747 32143 12789 32152
rect 12748 31781 12788 32143
rect 12747 31772 12789 31781
rect 12747 31732 12748 31772
rect 12788 31732 12789 31772
rect 12747 31723 12789 31732
rect 12555 31520 12597 31529
rect 12555 31480 12556 31520
rect 12596 31480 12597 31520
rect 12555 31471 12597 31480
rect 12459 31436 12501 31445
rect 12459 31396 12460 31436
rect 12500 31396 12501 31436
rect 12459 31387 12501 31396
rect 12844 31361 12884 35923
rect 13228 35888 13268 35897
rect 13268 35848 13364 35888
rect 13228 35839 13268 35848
rect 13227 35048 13269 35057
rect 13227 35008 13228 35048
rect 13268 35008 13269 35048
rect 13227 34999 13269 35008
rect 13228 34914 13268 34999
rect 13324 34628 13364 35848
rect 13324 34579 13364 34588
rect 13420 35216 13460 35225
rect 13036 34376 13076 34385
rect 13036 33713 13076 34336
rect 13131 33872 13173 33881
rect 13131 33832 13132 33872
rect 13172 33832 13173 33872
rect 13131 33823 13173 33832
rect 13035 33704 13077 33713
rect 13035 33664 13036 33704
rect 13076 33664 13077 33704
rect 13035 33655 13077 33664
rect 13132 33452 13172 33823
rect 13036 33412 13172 33452
rect 12939 33200 12981 33209
rect 12939 33160 12940 33200
rect 12980 33160 12981 33200
rect 12939 33151 12981 33160
rect 12940 32201 12980 33151
rect 13036 32789 13076 33412
rect 13035 32780 13077 32789
rect 13035 32740 13036 32780
rect 13076 32740 13077 32780
rect 13035 32731 13077 32740
rect 12939 32192 12981 32201
rect 12939 32152 12940 32192
rect 12980 32152 12981 32192
rect 12939 32143 12981 32152
rect 13036 32192 13076 32731
rect 13132 32696 13172 32705
rect 13132 32453 13172 32656
rect 13131 32444 13173 32453
rect 13131 32404 13132 32444
rect 13172 32404 13173 32444
rect 13131 32395 13173 32404
rect 13036 32143 13076 32152
rect 13132 32192 13172 32201
rect 13132 32117 13172 32152
rect 13131 32108 13173 32117
rect 13420 32108 13460 35176
rect 13611 35216 13653 35225
rect 13611 35176 13612 35216
rect 13652 35176 13653 35216
rect 13611 35167 13653 35176
rect 13612 35082 13652 35167
rect 13707 33872 13749 33881
rect 13707 33832 13708 33872
rect 13748 33832 13749 33872
rect 13707 33823 13749 33832
rect 13708 33738 13748 33823
rect 13611 32864 13653 32873
rect 13611 32824 13612 32864
rect 13652 32824 13653 32864
rect 13611 32815 13653 32824
rect 13804 32864 13844 32873
rect 13612 32360 13652 32815
rect 13804 32453 13844 32824
rect 13900 32528 13940 36016
rect 14572 36007 14612 36016
rect 14860 35888 14900 36511
rect 14860 35839 14900 35848
rect 14956 35888 14996 35897
rect 14956 35729 14996 35848
rect 15244 35888 15284 35897
rect 14379 35720 14421 35729
rect 14379 35680 14380 35720
rect 14420 35680 14421 35720
rect 14379 35671 14421 35680
rect 14955 35720 14997 35729
rect 14955 35680 14956 35720
rect 14996 35680 14997 35720
rect 14955 35671 14997 35680
rect 14380 35586 14420 35671
rect 14092 35216 14132 35225
rect 13996 34376 14036 34385
rect 13996 34049 14036 34336
rect 13995 34040 14037 34049
rect 13995 34000 13996 34040
rect 14036 34000 14037 34040
rect 13995 33991 14037 34000
rect 14092 33881 14132 35176
rect 14955 35048 14997 35057
rect 14955 35008 14956 35048
rect 14996 35008 14997 35048
rect 14955 34999 14997 35008
rect 14764 34964 14804 34973
rect 14380 34924 14764 34964
rect 14380 34376 14420 34924
rect 14764 34915 14804 34924
rect 14380 34327 14420 34336
rect 14956 34376 14996 34999
rect 14956 34327 14996 34336
rect 14572 34292 14612 34301
rect 14612 34252 14804 34292
rect 14572 34243 14612 34252
rect 14284 34208 14324 34217
rect 14091 33872 14133 33881
rect 14091 33832 14092 33872
rect 14132 33832 14133 33872
rect 14091 33823 14133 33832
rect 14092 33452 14132 33461
rect 13996 32864 14036 32873
rect 14092 32864 14132 33412
rect 14036 32824 14132 32864
rect 13996 32815 14036 32824
rect 14284 32537 14324 34168
rect 14571 34124 14613 34133
rect 14571 34084 14572 34124
rect 14612 34084 14613 34124
rect 14571 34075 14613 34084
rect 14572 33125 14612 34075
rect 14764 33872 14804 34252
rect 14956 33872 14996 33881
rect 14764 33832 14956 33872
rect 14956 33823 14996 33832
rect 14764 33704 14804 33713
rect 14571 33116 14613 33125
rect 14571 33076 14572 33116
rect 14612 33076 14613 33116
rect 14571 33067 14613 33076
rect 14379 32864 14421 32873
rect 14379 32824 14380 32864
rect 14420 32824 14421 32864
rect 14379 32815 14421 32824
rect 14380 32730 14420 32815
rect 14283 32528 14325 32537
rect 13900 32488 14132 32528
rect 13803 32444 13845 32453
rect 13803 32404 13804 32444
rect 13844 32404 13845 32444
rect 13803 32395 13845 32404
rect 13612 32311 13652 32320
rect 13707 32360 13749 32369
rect 13707 32320 13708 32360
rect 13748 32320 13749 32360
rect 13707 32311 13749 32320
rect 13131 32068 13132 32108
rect 13172 32068 13173 32108
rect 13131 32059 13173 32068
rect 13228 32068 13460 32108
rect 12939 31940 12981 31949
rect 12939 31900 12940 31940
rect 12980 31900 12981 31940
rect 12939 31891 12981 31900
rect 12556 31352 12596 31361
rect 12075 31268 12117 31277
rect 12075 31228 12076 31268
rect 12116 31228 12117 31268
rect 12075 31219 12117 31228
rect 12076 30680 12116 30689
rect 12556 30680 12596 31312
rect 12652 31352 12692 31361
rect 12652 31109 12692 31312
rect 12748 31352 12788 31361
rect 12651 31100 12693 31109
rect 12651 31060 12652 31100
rect 12692 31060 12693 31100
rect 12651 31051 12693 31060
rect 12748 30941 12788 31312
rect 12843 31352 12885 31361
rect 12843 31312 12844 31352
rect 12884 31312 12885 31352
rect 12843 31303 12885 31312
rect 12843 31184 12885 31193
rect 12843 31144 12844 31184
rect 12884 31144 12885 31184
rect 12843 31135 12885 31144
rect 12844 31050 12884 31135
rect 12747 30932 12789 30941
rect 12747 30892 12748 30932
rect 12788 30892 12789 30932
rect 12747 30883 12789 30892
rect 11500 30463 11540 30472
rect 11884 30640 12076 30680
rect 10827 30092 10869 30101
rect 10827 30052 10828 30092
rect 10868 30052 10869 30092
rect 10827 30043 10869 30052
rect 10827 29924 10869 29933
rect 10827 29884 10828 29924
rect 10868 29884 10964 29924
rect 10827 29875 10869 29884
rect 10924 29840 10964 29884
rect 10924 29791 10964 29800
rect 11884 29840 11924 30640
rect 12076 30631 12116 30640
rect 12460 30640 12556 30680
rect 12460 30092 12500 30640
rect 12556 30631 12596 30640
rect 12652 30680 12692 30689
rect 12652 30269 12692 30640
rect 12748 30680 12788 30883
rect 12843 30848 12885 30857
rect 12843 30808 12844 30848
rect 12884 30808 12885 30848
rect 12843 30799 12885 30808
rect 12844 30714 12884 30799
rect 12748 30631 12788 30640
rect 12843 30596 12885 30605
rect 12843 30556 12844 30596
rect 12884 30556 12885 30596
rect 12843 30547 12885 30556
rect 12651 30260 12693 30269
rect 12460 30043 12500 30052
rect 12556 30220 12652 30260
rect 12692 30220 12693 30260
rect 12171 29924 12213 29933
rect 12171 29884 12172 29924
rect 12212 29884 12213 29924
rect 12171 29875 12213 29884
rect 11787 29336 11829 29345
rect 11787 29296 11788 29336
rect 11828 29296 11829 29336
rect 11787 29287 11829 29296
rect 11788 29202 11828 29287
rect 9100 29119 9140 29128
rect 9964 29119 10004 29128
rect 11691 29000 11733 29009
rect 11691 28960 11692 29000
rect 11732 28960 11733 29000
rect 11884 29000 11924 29800
rect 12172 29840 12212 29875
rect 12172 29789 12212 29800
rect 12460 29168 12500 29177
rect 12556 29168 12596 30220
rect 12651 30211 12693 30220
rect 12500 29128 12596 29168
rect 12460 29119 12500 29128
rect 11884 28960 12020 29000
rect 11691 28951 11733 28960
rect 10347 28916 10389 28925
rect 10347 28876 10348 28916
rect 10388 28876 10389 28916
rect 10347 28867 10389 28876
rect 11115 28916 11157 28925
rect 11115 28876 11116 28916
rect 11156 28876 11157 28916
rect 11115 28867 11157 28876
rect 11499 28916 11541 28925
rect 11499 28876 11500 28916
rect 11540 28876 11541 28916
rect 11499 28867 11541 28876
rect 8620 28456 8852 28496
rect 8427 28328 8469 28337
rect 8427 28288 8428 28328
rect 8468 28288 8469 28328
rect 8427 28279 8469 28288
rect 8524 28328 8564 28337
rect 8716 28328 8756 28337
rect 8139 28160 8181 28169
rect 8139 28120 8140 28160
rect 8180 28120 8181 28160
rect 8139 28111 8181 28120
rect 8139 27656 8181 27665
rect 8139 27616 8140 27656
rect 8180 27616 8181 27656
rect 8139 27607 8181 27616
rect 8427 27656 8469 27665
rect 8427 27616 8428 27656
rect 8468 27616 8469 27656
rect 8427 27607 8469 27616
rect 7947 27488 7989 27497
rect 7947 27448 7948 27488
rect 7988 27448 7989 27488
rect 7947 27439 7989 27448
rect 7851 27320 7893 27329
rect 7851 27280 7852 27320
rect 7892 27280 7893 27320
rect 7851 27271 7893 27280
rect 7947 27152 7989 27161
rect 7947 27112 7948 27152
rect 7988 27112 7989 27152
rect 7947 27103 7989 27112
rect 7851 26816 7893 26825
rect 7851 26776 7852 26816
rect 7892 26776 7893 26816
rect 7851 26767 7893 26776
rect 7948 26816 7988 27103
rect 7948 26767 7988 26776
rect 8140 26816 8180 27607
rect 8428 27522 8468 27607
rect 8524 27413 8564 28288
rect 8620 28288 8716 28328
rect 8523 27404 8565 27413
rect 8523 27364 8524 27404
rect 8564 27364 8565 27404
rect 8523 27355 8565 27364
rect 8620 27236 8660 28288
rect 8716 28279 8756 28288
rect 8812 28160 8852 28456
rect 10348 28328 10388 28867
rect 11116 28782 11156 28867
rect 10348 28279 10388 28288
rect 8140 26767 8180 26776
rect 8236 27196 8660 27236
rect 8716 28120 8852 28160
rect 9388 28160 9428 28169
rect 9675 28160 9717 28169
rect 9428 28120 9524 28160
rect 7852 26682 7892 26767
rect 8044 26732 8084 26741
rect 8044 26648 8084 26692
rect 8236 26648 8276 27196
rect 8427 27068 8469 27077
rect 8427 27028 8428 27068
rect 8468 27028 8469 27068
rect 8427 27019 8469 27028
rect 8428 26934 8468 27019
rect 8523 26900 8565 26909
rect 8523 26860 8524 26900
rect 8564 26860 8565 26900
rect 8523 26851 8565 26860
rect 8332 26816 8372 26825
rect 8332 26657 8372 26776
rect 8524 26816 8564 26851
rect 8524 26765 8564 26776
rect 8044 26608 8276 26648
rect 8331 26648 8373 26657
rect 8331 26608 8332 26648
rect 8372 26608 8373 26648
rect 8331 26599 8373 26608
rect 7756 26524 8084 26564
rect 7947 26396 7989 26405
rect 7947 26356 7948 26396
rect 7988 26356 7989 26396
rect 7947 26347 7989 26356
rect 7755 26312 7797 26321
rect 7755 26272 7756 26312
rect 7796 26272 7797 26312
rect 7755 26263 7797 26272
rect 7756 26144 7796 26263
rect 7756 26095 7796 26104
rect 7851 26144 7893 26153
rect 7851 26104 7852 26144
rect 7892 26104 7893 26144
rect 7851 26095 7893 26104
rect 7948 26144 7988 26347
rect 7948 26095 7988 26104
rect 8044 26144 8084 26524
rect 8716 26405 8756 28120
rect 9388 28111 9428 28120
rect 9484 27740 9524 28120
rect 9675 28120 9676 28160
rect 9716 28120 9717 28160
rect 9675 28111 9717 28120
rect 10540 28160 10580 28169
rect 9676 28026 9716 28111
rect 10059 27908 10101 27917
rect 10059 27868 10060 27908
rect 10100 27868 10101 27908
rect 10059 27859 10101 27868
rect 9676 27740 9716 27749
rect 9484 27700 9676 27740
rect 9676 27691 9716 27700
rect 9292 27656 9332 27665
rect 9292 27497 9332 27616
rect 9291 27488 9333 27497
rect 9291 27448 9292 27488
rect 9332 27448 9333 27488
rect 9291 27439 9333 27448
rect 10060 27488 10100 27859
rect 10540 27749 10580 28120
rect 10539 27740 10581 27749
rect 10539 27700 10540 27740
rect 10580 27700 10581 27740
rect 10539 27691 10581 27700
rect 10923 27740 10965 27749
rect 10923 27700 10924 27740
rect 10964 27700 10965 27740
rect 10923 27691 10965 27700
rect 10924 27656 10964 27691
rect 11212 27656 11252 27665
rect 10924 27605 10964 27616
rect 11020 27616 11212 27656
rect 10060 27439 10100 27448
rect 10252 27404 10292 27413
rect 9963 27320 10005 27329
rect 9963 27280 9964 27320
rect 10004 27280 10005 27320
rect 9963 27271 10005 27280
rect 9483 27152 9525 27161
rect 8812 27112 9332 27152
rect 8715 26396 8757 26405
rect 8715 26356 8716 26396
rect 8756 26356 8757 26396
rect 8715 26347 8757 26356
rect 8812 26228 8852 27112
rect 9292 27068 9332 27112
rect 9483 27112 9484 27152
rect 9524 27112 9525 27152
rect 9483 27103 9525 27112
rect 9771 27152 9813 27161
rect 9771 27112 9772 27152
rect 9812 27112 9813 27152
rect 9771 27103 9813 27112
rect 9292 27019 9332 27028
rect 9100 26984 9140 26993
rect 8907 26900 8949 26909
rect 8907 26860 8908 26900
rect 8948 26860 8949 26900
rect 8907 26851 8949 26860
rect 8812 26179 8852 26188
rect 8044 26095 8084 26104
rect 7755 25976 7797 25985
rect 7755 25936 7756 25976
rect 7796 25936 7797 25976
rect 7755 25927 7797 25936
rect 7756 25842 7796 25927
rect 7852 25304 7892 26095
rect 8428 25976 8468 25985
rect 8468 25936 8756 25976
rect 8428 25927 8468 25936
rect 8716 25304 8756 25936
rect 8908 25817 8948 26851
rect 9100 26144 9140 26944
rect 9291 26816 9333 26825
rect 9291 26776 9292 26816
rect 9332 26776 9333 26816
rect 9291 26767 9333 26776
rect 9484 26816 9524 27103
rect 9484 26767 9524 26776
rect 9580 26816 9620 26825
rect 9292 26682 9332 26767
rect 9580 26732 9620 26776
rect 9772 26816 9812 27103
rect 9867 26900 9909 26909
rect 9867 26860 9868 26900
rect 9908 26860 9909 26900
rect 9867 26851 9909 26860
rect 9772 26767 9812 26776
rect 9868 26816 9908 26851
rect 9868 26765 9908 26776
rect 9964 26816 10004 27271
rect 10252 26993 10292 27364
rect 10539 27152 10581 27161
rect 10539 27112 10540 27152
rect 10580 27112 10581 27152
rect 10539 27103 10581 27112
rect 10251 26984 10293 26993
rect 10251 26944 10252 26984
rect 10292 26944 10293 26984
rect 10251 26935 10293 26944
rect 10251 26816 10293 26825
rect 10004 26776 10196 26816
rect 9964 26767 10004 26776
rect 9675 26732 9717 26741
rect 9580 26692 9676 26732
rect 9716 26692 9717 26732
rect 9675 26683 9717 26692
rect 10059 26648 10101 26657
rect 10059 26608 10060 26648
rect 10100 26608 10101 26648
rect 10059 26599 10101 26608
rect 10060 26514 10100 26599
rect 10156 26564 10196 26776
rect 10251 26776 10252 26816
rect 10292 26776 10293 26816
rect 10251 26767 10293 26776
rect 10348 26816 10388 26825
rect 10252 26682 10292 26767
rect 10348 26564 10388 26776
rect 10156 26524 10388 26564
rect 10444 26816 10484 26825
rect 10444 26489 10484 26776
rect 10540 26816 10580 27103
rect 10443 26480 10485 26489
rect 10443 26440 10444 26480
rect 10484 26440 10485 26480
rect 10443 26431 10485 26440
rect 9196 26144 9236 26153
rect 9100 26104 9196 26144
rect 9196 26095 9236 26104
rect 10059 26144 10101 26153
rect 10059 26104 10060 26144
rect 10100 26104 10101 26144
rect 10059 26095 10101 26104
rect 10060 26010 10100 26095
rect 8907 25808 8949 25817
rect 8907 25768 8908 25808
rect 8948 25768 8949 25808
rect 8907 25759 8949 25768
rect 7892 25264 8084 25304
rect 7852 25255 7892 25264
rect 7947 24884 7989 24893
rect 7947 24844 7948 24884
rect 7988 24844 7989 24884
rect 7947 24835 7989 24844
rect 7756 24632 7796 24641
rect 7660 24592 7756 24632
rect 7564 24581 7604 24592
rect 7756 24583 7796 24592
rect 7948 24632 7988 24835
rect 7948 24557 7988 24592
rect 7852 24548 7892 24557
rect 7275 24464 7317 24473
rect 7275 24424 7276 24464
rect 7316 24424 7317 24464
rect 7275 24415 7317 24424
rect 6644 23752 6836 23792
rect 6892 24380 6932 24389
rect 6892 23792 6932 24340
rect 6604 23743 6644 23752
rect 6892 23743 6932 23752
rect 7276 23792 7316 24415
rect 7852 24305 7892 24508
rect 7947 24548 7989 24557
rect 7947 24508 7948 24548
rect 7988 24508 7989 24548
rect 7947 24499 7989 24508
rect 7948 24468 7988 24499
rect 7851 24296 7893 24305
rect 7851 24256 7852 24296
rect 7892 24256 7893 24296
rect 7851 24247 7893 24256
rect 8044 23969 8084 25264
rect 8716 25255 8756 25264
rect 8620 24632 8660 24641
rect 8524 24592 8620 24632
rect 8139 24464 8181 24473
rect 8139 24424 8140 24464
rect 8180 24424 8181 24464
rect 8139 24415 8181 24424
rect 8140 24330 8180 24415
rect 8043 23960 8085 23969
rect 8043 23920 8044 23960
rect 8084 23920 8085 23960
rect 8043 23911 8085 23920
rect 8044 23792 8084 23911
rect 8140 23792 8180 23801
rect 8044 23752 8140 23792
rect 7276 23743 7316 23752
rect 8140 23743 8180 23752
rect 5932 23288 5972 23297
rect 5836 23248 5932 23288
rect 5644 23239 5684 23248
rect 5932 23239 5972 23248
rect 5835 23120 5877 23129
rect 5835 23080 5836 23120
rect 5876 23080 5877 23120
rect 5835 23071 5877 23080
rect 6124 23120 6164 23129
rect 7180 23120 7220 23129
rect 5836 22986 5876 23071
rect 5452 22828 5588 22868
rect 5644 22868 5684 22877
rect 6027 22868 6069 22877
rect 5684 22828 5780 22868
rect 5259 22784 5301 22793
rect 5259 22744 5260 22784
rect 5300 22744 5301 22784
rect 5259 22735 5301 22744
rect 4971 22700 5013 22709
rect 4971 22660 4972 22700
rect 5012 22660 5013 22700
rect 4971 22651 5013 22660
rect 5452 22373 5492 22828
rect 5644 22819 5684 22828
rect 5547 22700 5589 22709
rect 5547 22660 5548 22700
rect 5588 22660 5589 22700
rect 5547 22651 5589 22660
rect 5451 22364 5493 22373
rect 5451 22324 5452 22364
rect 5492 22324 5493 22364
rect 5451 22315 5493 22324
rect 4588 22231 4628 22240
rect 4780 22280 4820 22289
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4491 21776 4533 21785
rect 4491 21736 4492 21776
rect 4532 21736 4533 21776
rect 4491 21727 4533 21736
rect 4492 21642 4532 21727
rect 4780 21524 4820 22240
rect 4972 22280 5012 22289
rect 4875 22196 4917 22205
rect 4875 22156 4876 22196
rect 4916 22156 4917 22196
rect 4875 22147 4917 22156
rect 4876 22062 4916 22147
rect 4875 21692 4917 21701
rect 4875 21652 4876 21692
rect 4916 21652 4917 21692
rect 4875 21643 4917 21652
rect 4876 21608 4916 21643
rect 4876 21557 4916 21568
rect 4684 21484 4820 21524
rect 4396 21020 4436 21029
rect 4204 20980 4396 21020
rect 4396 20971 4436 20980
rect 4491 20768 4533 20777
rect 4491 20728 4492 20768
rect 4532 20728 4533 20768
rect 4491 20719 4533 20728
rect 4684 20768 4724 21484
rect 4972 21440 5012 22240
rect 5068 22280 5108 22289
rect 5068 21785 5108 22240
rect 5548 22280 5588 22651
rect 5643 22364 5685 22373
rect 5643 22324 5644 22364
rect 5684 22324 5685 22364
rect 5643 22315 5685 22324
rect 5548 22231 5588 22240
rect 5452 22112 5492 22121
rect 5163 21944 5205 21953
rect 5163 21904 5164 21944
rect 5204 21904 5205 21944
rect 5163 21895 5205 21904
rect 5067 21776 5109 21785
rect 5067 21736 5068 21776
rect 5108 21736 5109 21776
rect 5067 21727 5109 21736
rect 5068 21608 5108 21617
rect 5164 21608 5204 21895
rect 5260 21617 5300 21702
rect 5452 21692 5492 22072
rect 5547 21944 5589 21953
rect 5547 21904 5548 21944
rect 5588 21904 5589 21944
rect 5547 21895 5589 21904
rect 5548 21776 5588 21895
rect 5548 21727 5588 21736
rect 5356 21652 5492 21692
rect 5108 21568 5204 21608
rect 5259 21608 5301 21617
rect 5259 21568 5260 21608
rect 5300 21568 5301 21608
rect 5068 21559 5108 21568
rect 5259 21559 5301 21568
rect 5356 21608 5396 21652
rect 5356 21559 5396 21568
rect 5644 21608 5684 22315
rect 4780 21400 5012 21440
rect 5067 21440 5109 21449
rect 5067 21400 5068 21440
rect 5108 21400 5109 21440
rect 4780 21356 4820 21400
rect 5067 21391 5109 21400
rect 4780 21307 4820 21316
rect 5068 21306 5108 21391
rect 4971 21272 5013 21281
rect 4971 21232 4972 21272
rect 5012 21232 5013 21272
rect 4971 21223 5013 21232
rect 4779 21188 4821 21197
rect 4779 21148 4780 21188
rect 4820 21148 4821 21188
rect 4779 21139 4821 21148
rect 4684 20719 4724 20728
rect 4780 20768 4820 21139
rect 4780 20719 4820 20728
rect 4875 20768 4917 20777
rect 4875 20728 4876 20768
rect 4916 20728 4917 20768
rect 4875 20719 4917 20728
rect 4972 20768 5012 21223
rect 5644 21197 5684 21568
rect 5740 21608 5780 22828
rect 6027 22828 6028 22868
rect 6068 22828 6069 22868
rect 6027 22819 6069 22828
rect 5932 22448 5972 22457
rect 5932 21617 5972 22408
rect 6028 21692 6068 22819
rect 6124 22793 6164 23080
rect 6412 23080 7180 23120
rect 6123 22784 6165 22793
rect 6123 22744 6124 22784
rect 6164 22744 6165 22784
rect 6123 22735 6165 22744
rect 6412 22532 6452 23080
rect 7180 23071 7220 23080
rect 8044 23120 8084 23129
rect 8084 23080 8180 23120
rect 8044 23071 8084 23080
rect 6507 22868 6549 22877
rect 6507 22828 6508 22868
rect 6548 22828 6549 22868
rect 6507 22819 6549 22828
rect 7372 22868 7412 22877
rect 6508 22734 6548 22819
rect 7372 22709 7412 22828
rect 7851 22784 7893 22793
rect 7851 22744 7852 22784
rect 7892 22744 7893 22784
rect 7851 22735 7893 22744
rect 7371 22700 7413 22709
rect 7371 22660 7372 22700
rect 7412 22660 7413 22700
rect 7371 22651 7413 22660
rect 6412 22483 6452 22492
rect 7563 22364 7605 22373
rect 7563 22324 7564 22364
rect 7604 22324 7605 22364
rect 7563 22315 7605 22324
rect 6123 22280 6165 22289
rect 6123 22240 6124 22280
rect 6164 22240 6165 22280
rect 6123 22231 6165 22240
rect 6220 22280 6260 22289
rect 6124 22146 6164 22231
rect 6124 21692 6164 21701
rect 6028 21652 6124 21692
rect 6124 21643 6164 21652
rect 5740 21559 5780 21568
rect 5836 21608 5876 21617
rect 5836 21449 5876 21568
rect 5931 21608 5973 21617
rect 5931 21568 5932 21608
rect 5972 21568 5973 21608
rect 5931 21559 5973 21568
rect 6220 21449 6260 22240
rect 6412 22280 6452 22289
rect 7276 22280 7316 22291
rect 6452 22240 6740 22280
rect 6412 22231 6452 22240
rect 6604 22112 6644 22121
rect 6604 21701 6644 22072
rect 6603 21692 6645 21701
rect 6603 21652 6604 21692
rect 6644 21652 6645 21692
rect 6603 21643 6645 21652
rect 6507 21608 6549 21617
rect 6507 21568 6508 21608
rect 6548 21568 6549 21608
rect 6507 21559 6549 21568
rect 6508 21474 6548 21559
rect 6603 21524 6645 21533
rect 6603 21484 6604 21524
rect 6644 21484 6645 21524
rect 6603 21475 6645 21484
rect 5835 21440 5877 21449
rect 5835 21400 5836 21440
rect 5876 21400 5877 21440
rect 5835 21391 5877 21400
rect 6219 21440 6261 21449
rect 6219 21400 6220 21440
rect 6260 21400 6261 21440
rect 6219 21391 6261 21400
rect 5643 21188 5685 21197
rect 5643 21148 5644 21188
rect 5684 21148 5685 21188
rect 5643 21139 5685 21148
rect 5836 21020 5876 21391
rect 6604 21356 6644 21475
rect 6508 21316 6644 21356
rect 6028 21020 6068 21029
rect 5836 20980 6028 21020
rect 6028 20971 6068 20980
rect 6219 20852 6261 20861
rect 6219 20812 6220 20852
rect 6260 20812 6261 20852
rect 6219 20803 6261 20812
rect 4492 20634 4532 20719
rect 4876 20634 4916 20719
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4108 20273 4148 20358
rect 4972 20357 5012 20728
rect 5163 20768 5205 20777
rect 5163 20728 5164 20768
rect 5204 20728 5205 20768
rect 5163 20719 5205 20728
rect 5548 20768 5588 20777
rect 4971 20348 5013 20357
rect 4971 20308 4972 20348
rect 5012 20308 5013 20348
rect 4971 20299 5013 20308
rect 4107 20264 4149 20273
rect 4107 20224 4108 20264
rect 4148 20224 4149 20264
rect 4107 20215 4149 20224
rect 3531 20096 3573 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 4012 20096 4052 20107
rect 2380 19928 2420 19937
rect 2284 19888 2380 19928
rect 2284 19256 2324 19888
rect 2380 19879 2420 19888
rect 2955 19844 2997 19853
rect 2955 19804 2956 19844
rect 2996 19804 2997 19844
rect 2955 19795 2997 19804
rect 2284 19207 2324 19216
rect 1900 19172 1940 19181
rect 843 18836 885 18845
rect 843 18796 844 18836
rect 884 18796 885 18836
rect 843 18787 885 18796
rect 1900 18761 1940 19132
rect 2283 19088 2325 19097
rect 2283 19048 2284 19088
rect 2324 19048 2325 19088
rect 2283 19039 2325 19048
rect 652 18752 692 18761
rect 652 18257 692 18712
rect 1899 18752 1941 18761
rect 1899 18712 1900 18752
rect 1940 18712 1941 18752
rect 1899 18703 1941 18712
rect 1995 18584 2037 18593
rect 1995 18544 1996 18584
rect 2036 18544 2037 18584
rect 1995 18535 2037 18544
rect 1708 18416 1748 18425
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 1036 17912 1076 17921
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 17240 692 17359
rect 652 17191 692 17200
rect 1036 17081 1076 17872
rect 1612 17744 1652 17753
rect 1708 17744 1748 18376
rect 1652 17704 1748 17744
rect 1612 17695 1652 17704
rect 1228 17660 1268 17669
rect 1035 17072 1077 17081
rect 1035 17032 1036 17072
rect 1076 17032 1077 17072
rect 1035 17023 1077 17032
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 14552 692 16519
rect 1228 16409 1268 17620
rect 1324 17072 1364 17081
rect 1707 17072 1749 17081
rect 1364 17032 1460 17072
rect 1324 17023 1364 17032
rect 940 16400 980 16409
rect 747 15728 789 15737
rect 747 15688 748 15728
rect 788 15688 789 15728
rect 747 15679 789 15688
rect 748 15594 788 15679
rect 940 14729 980 16360
rect 1227 16400 1269 16409
rect 1227 16360 1228 16400
rect 1268 16360 1269 16400
rect 1227 16351 1269 16360
rect 1132 16232 1172 16241
rect 1132 15989 1172 16192
rect 1324 16232 1364 16241
rect 1227 16148 1269 16157
rect 1227 16108 1228 16148
rect 1268 16108 1269 16148
rect 1227 16099 1269 16108
rect 1228 16014 1268 16099
rect 1131 15980 1173 15989
rect 1131 15940 1132 15980
rect 1172 15940 1173 15980
rect 1131 15931 1173 15940
rect 1131 15560 1173 15569
rect 1131 15520 1132 15560
rect 1172 15520 1173 15560
rect 1131 15511 1173 15520
rect 1132 15426 1172 15511
rect 1035 14888 1077 14897
rect 1035 14848 1036 14888
rect 1076 14848 1077 14888
rect 1035 14839 1077 14848
rect 939 14720 981 14729
rect 939 14680 940 14720
rect 980 14680 981 14720
rect 939 14671 981 14680
rect 652 14503 692 14512
rect 1036 14552 1076 14839
rect 1036 14503 1076 14512
rect 652 14216 692 14225
rect 652 14057 692 14176
rect 1324 14141 1364 16192
rect 1420 16073 1460 17032
rect 1707 17032 1708 17072
rect 1748 17032 1749 17072
rect 1707 17023 1749 17032
rect 1708 16938 1748 17023
rect 1516 16232 1556 16241
rect 1419 16064 1461 16073
rect 1419 16024 1420 16064
rect 1460 16024 1461 16064
rect 1419 16015 1461 16024
rect 1516 15728 1556 16192
rect 1611 16232 1653 16241
rect 1611 16192 1612 16232
rect 1652 16192 1653 16232
rect 1611 16183 1653 16192
rect 1804 16232 1844 16241
rect 1996 16232 2036 18535
rect 2091 16400 2133 16409
rect 2091 16360 2092 16400
rect 2132 16360 2133 16400
rect 2091 16351 2133 16360
rect 2092 16266 2132 16351
rect 2187 16316 2229 16325
rect 2187 16276 2188 16316
rect 2228 16276 2229 16316
rect 2187 16267 2229 16276
rect 1844 16192 1996 16232
rect 1804 16183 1844 16192
rect 1996 16183 2036 16192
rect 2188 16232 2228 16267
rect 1612 16098 1652 16183
rect 2188 16181 2228 16192
rect 2284 16232 2324 19039
rect 2571 18920 2613 18929
rect 2571 18880 2572 18920
rect 2612 18880 2613 18920
rect 2571 18871 2613 18880
rect 2476 17744 2516 17753
rect 2572 17744 2612 18871
rect 2859 18752 2901 18761
rect 2859 18712 2860 18752
rect 2900 18712 2901 18752
rect 2859 18703 2901 18712
rect 2860 18618 2900 18703
rect 2763 18584 2805 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 2956 18584 2996 19795
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3532 19508 3572 20047
rect 4012 20021 4052 20056
rect 4875 20096 4917 20105
rect 4972 20096 5012 20299
rect 5164 20273 5204 20719
rect 5259 20600 5301 20609
rect 5259 20560 5260 20600
rect 5300 20560 5301 20600
rect 5259 20551 5301 20560
rect 5163 20264 5205 20273
rect 5163 20224 5164 20264
rect 5204 20224 5205 20264
rect 5163 20215 5205 20224
rect 4875 20056 4876 20096
rect 4916 20056 5012 20096
rect 5068 20096 5108 20105
rect 4875 20047 4917 20056
rect 4011 20012 4053 20021
rect 4011 19972 4012 20012
rect 4052 19972 4053 20012
rect 4011 19963 4053 19972
rect 3436 19468 3572 19508
rect 3820 19844 3860 19853
rect 3148 19256 3188 19265
rect 3148 18929 3188 19216
rect 3243 19004 3285 19013
rect 3243 18964 3244 19004
rect 3284 18964 3285 19004
rect 3243 18955 3285 18964
rect 3147 18920 3189 18929
rect 3147 18880 3148 18920
rect 3188 18880 3189 18920
rect 3147 18871 3189 18880
rect 3244 18752 3284 18955
rect 2956 18535 2996 18544
rect 3052 18712 3244 18752
rect 3052 18584 3092 18712
rect 3244 18703 3284 18712
rect 3052 18535 3092 18544
rect 3436 18584 3476 19468
rect 3820 19265 3860 19804
rect 3819 19256 3861 19265
rect 3819 19216 3820 19256
rect 3860 19216 3861 19256
rect 3819 19207 3861 19216
rect 3820 19097 3860 19207
rect 3819 19088 3861 19097
rect 3819 19048 3820 19088
rect 3860 19048 3861 19088
rect 3819 19039 3861 19048
rect 4012 19013 4052 19963
rect 4876 19962 4916 20047
rect 4875 19844 4917 19853
rect 4875 19804 4876 19844
rect 4916 19804 4917 19844
rect 4875 19795 4917 19804
rect 4876 19710 4916 19795
rect 4300 19340 4340 19349
rect 4340 19300 4724 19340
rect 4300 19291 4340 19300
rect 4684 19256 4724 19300
rect 4724 19216 4820 19256
rect 4684 19207 4724 19216
rect 4011 19004 4053 19013
rect 4011 18964 4012 19004
rect 4052 18964 4053 19004
rect 4011 18955 4053 18964
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3531 18752 3573 18761
rect 3531 18712 3532 18752
rect 3572 18712 3573 18752
rect 3531 18703 3573 18712
rect 4107 18752 4149 18761
rect 4107 18712 4108 18752
rect 4148 18712 4149 18752
rect 4107 18703 4149 18712
rect 3532 18618 3572 18703
rect 3724 18584 3764 18593
rect 3436 18535 3476 18544
rect 3628 18544 3724 18584
rect 2764 18257 2804 18535
rect 2763 18248 2805 18257
rect 2763 18208 2764 18248
rect 2804 18208 2805 18248
rect 2763 18199 2805 18208
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3628 17837 3668 18544
rect 3724 18535 3764 18544
rect 3627 17828 3669 17837
rect 3627 17788 3628 17828
rect 3668 17788 3669 17828
rect 3627 17779 3669 17788
rect 2516 17704 2612 17744
rect 2476 17695 2516 17704
rect 2572 17081 2612 17704
rect 3628 17694 3668 17779
rect 3916 17744 3956 17753
rect 3724 17704 3916 17744
rect 3724 17240 3764 17704
rect 3916 17695 3956 17704
rect 3724 17191 3764 17200
rect 2571 17072 2613 17081
rect 2571 17032 2572 17072
rect 2612 17032 2613 17072
rect 2571 17023 2613 17032
rect 3627 17072 3669 17081
rect 3916 17072 3956 17081
rect 3627 17032 3628 17072
rect 3668 17032 3916 17072
rect 3627 17023 3669 17032
rect 3916 17023 3956 17032
rect 2572 16938 2612 17023
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 2284 16183 2324 16192
rect 3148 16232 3188 16241
rect 1708 16064 1748 16073
rect 1516 15688 1652 15728
rect 1516 15560 1556 15569
rect 1516 14888 1556 15520
rect 1612 15233 1652 15688
rect 1708 15569 1748 16024
rect 2476 16064 2516 16075
rect 2476 15989 2516 16024
rect 2475 15980 2517 15989
rect 2475 15940 2476 15980
rect 2516 15940 2517 15980
rect 2475 15931 2517 15940
rect 2476 15653 2516 15931
rect 2475 15644 2517 15653
rect 2475 15604 2476 15644
rect 2516 15604 2517 15644
rect 2475 15595 2517 15604
rect 1707 15560 1749 15569
rect 1707 15520 1708 15560
rect 1748 15520 1749 15560
rect 1707 15511 1749 15520
rect 2379 15560 2421 15569
rect 2379 15520 2380 15560
rect 2420 15520 2421 15560
rect 2379 15511 2421 15520
rect 2380 15426 2420 15511
rect 2379 15308 2421 15317
rect 2379 15268 2380 15308
rect 2420 15268 2421 15308
rect 3148 15308 3188 16192
rect 3339 16064 3381 16073
rect 3339 16024 3340 16064
rect 3380 16024 3381 16064
rect 3339 16015 3381 16024
rect 3340 15930 3380 16015
rect 3628 15569 3668 17023
rect 4012 16232 4052 16241
rect 3915 15980 3957 15989
rect 3915 15940 3916 15980
rect 3956 15940 3957 15980
rect 3915 15931 3957 15940
rect 3916 15728 3956 15931
rect 4012 15737 4052 16192
rect 4108 15980 4148 18703
rect 4588 18584 4628 18593
rect 4780 18584 4820 19216
rect 5068 18761 5108 20056
rect 5067 18752 5109 18761
rect 5067 18712 5068 18752
rect 5108 18712 5109 18752
rect 5067 18703 5109 18712
rect 4628 18544 4820 18584
rect 4588 18535 4628 18544
rect 5067 18500 5109 18509
rect 5067 18460 5068 18500
rect 5108 18460 5109 18500
rect 5067 18451 5109 18460
rect 4396 18332 4436 18341
rect 4396 17753 4436 18292
rect 4780 17837 4820 17868
rect 4779 17828 4821 17837
rect 4779 17788 4780 17828
rect 4820 17788 4821 17828
rect 4779 17779 4821 17788
rect 4971 17828 5013 17837
rect 4971 17788 4972 17828
rect 5012 17788 5013 17828
rect 4971 17779 5013 17788
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4588 17669 4628 17754
rect 4780 17744 4820 17779
rect 4587 17660 4629 17669
rect 4587 17620 4588 17660
rect 4628 17620 4629 17660
rect 4587 17611 4629 17620
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4203 16232 4245 16241
rect 4203 16192 4204 16232
rect 4244 16192 4245 16232
rect 4203 16183 4245 16192
rect 4204 16098 4244 16183
rect 4108 15940 4244 15980
rect 4107 15812 4149 15821
rect 4107 15772 4108 15812
rect 4148 15772 4149 15812
rect 4107 15763 4149 15772
rect 3916 15679 3956 15688
rect 4011 15728 4053 15737
rect 4011 15688 4012 15728
rect 4052 15688 4053 15728
rect 4011 15679 4053 15688
rect 3627 15560 3669 15569
rect 3627 15520 3628 15560
rect 3668 15520 3669 15560
rect 3627 15511 3669 15520
rect 3820 15560 3860 15569
rect 3532 15308 3572 15317
rect 3148 15268 3532 15308
rect 2379 15259 2421 15268
rect 1611 15224 1653 15233
rect 1611 15184 1612 15224
rect 1652 15184 1653 15224
rect 1611 15175 1653 15184
rect 1708 14888 1748 14897
rect 1516 14848 1708 14888
rect 1708 14839 1748 14848
rect 2380 14720 2420 15259
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3532 14981 3572 15268
rect 3531 14972 3573 14981
rect 3531 14932 3532 14972
rect 3572 14932 3573 14972
rect 3531 14923 3573 14932
rect 3628 14729 3668 15511
rect 3820 15233 3860 15520
rect 4012 15560 4052 15569
rect 4108 15560 4148 15763
rect 4052 15520 4148 15560
rect 4012 15511 4052 15520
rect 4204 15476 4244 15940
rect 4780 15905 4820 17704
rect 4972 17669 5012 17779
rect 4971 17660 5013 17669
rect 4971 17620 4972 17660
rect 5012 17620 5013 17660
rect 4971 17611 5013 17620
rect 4875 17072 4917 17081
rect 4875 17032 4876 17072
rect 4916 17032 4917 17072
rect 4875 17023 4917 17032
rect 4876 16938 4916 17023
rect 4875 16232 4917 16241
rect 4875 16192 4876 16232
rect 4916 16192 4917 16232
rect 4875 16183 4917 16192
rect 4876 16098 4916 16183
rect 4972 15980 5012 17611
rect 5068 16409 5108 18451
rect 5164 17996 5204 20215
rect 5260 18509 5300 20551
rect 5548 20189 5588 20728
rect 5739 20768 5781 20777
rect 5739 20728 5740 20768
rect 5780 20728 5781 20768
rect 5739 20719 5781 20728
rect 5740 20634 5780 20719
rect 6220 20718 6260 20803
rect 6412 20768 6452 20777
rect 5643 20600 5685 20609
rect 5643 20560 5644 20600
rect 5684 20560 5685 20600
rect 5643 20551 5685 20560
rect 6028 20600 6068 20609
rect 6412 20600 6452 20728
rect 6508 20768 6548 21316
rect 6508 20719 6548 20728
rect 6604 20768 6644 20777
rect 6068 20560 6452 20600
rect 6028 20551 6068 20560
rect 5644 20466 5684 20551
rect 5547 20180 5589 20189
rect 5547 20140 5548 20180
rect 5588 20140 5589 20180
rect 5547 20131 5589 20140
rect 5643 20096 5685 20105
rect 6028 20096 6068 20105
rect 5643 20056 5644 20096
rect 5684 20056 5685 20096
rect 5643 20047 5685 20056
rect 5740 20056 6028 20096
rect 5644 19962 5684 20047
rect 5452 19928 5492 19937
rect 5452 19844 5492 19888
rect 5740 19844 5780 20056
rect 6028 20047 6068 20056
rect 6027 19928 6069 19937
rect 6027 19888 6028 19928
rect 6068 19888 6069 19928
rect 6027 19879 6069 19888
rect 5452 19804 5780 19844
rect 5548 19265 5588 19350
rect 5931 19340 5973 19349
rect 5931 19300 5932 19340
rect 5972 19300 5973 19340
rect 5931 19291 5973 19300
rect 5547 19256 5589 19265
rect 5547 19216 5548 19256
rect 5588 19216 5589 19256
rect 5547 19207 5589 19216
rect 5740 19256 5780 19265
rect 5356 19088 5396 19097
rect 5644 19088 5684 19097
rect 5356 18761 5396 19048
rect 5548 19048 5644 19088
rect 5355 18752 5397 18761
rect 5355 18712 5356 18752
rect 5396 18712 5397 18752
rect 5355 18703 5397 18712
rect 5259 18500 5301 18509
rect 5259 18460 5260 18500
rect 5300 18460 5301 18500
rect 5259 18451 5301 18460
rect 5259 18332 5301 18341
rect 5259 18292 5260 18332
rect 5300 18292 5301 18332
rect 5259 18283 5301 18292
rect 5260 18198 5300 18283
rect 5452 17996 5492 18005
rect 5164 17956 5452 17996
rect 5452 17947 5492 17956
rect 5355 17576 5397 17585
rect 5355 17536 5356 17576
rect 5396 17536 5397 17576
rect 5355 17527 5397 17536
rect 5260 16820 5300 16829
rect 5164 16780 5260 16820
rect 5067 16400 5109 16409
rect 5067 16360 5068 16400
rect 5108 16360 5109 16400
rect 5067 16351 5109 16360
rect 4876 15940 5012 15980
rect 5068 16148 5108 16157
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4779 15896 4821 15905
rect 4779 15856 4780 15896
rect 4820 15856 4821 15896
rect 4779 15847 4821 15856
rect 4876 15728 4916 15940
rect 5068 15905 5108 16108
rect 5067 15896 5109 15905
rect 5067 15856 5068 15896
rect 5108 15856 5109 15896
rect 5067 15847 5109 15856
rect 4780 15688 4916 15728
rect 4971 15728 5013 15737
rect 5164 15728 5204 16780
rect 5260 16771 5300 16780
rect 5356 16484 5396 17527
rect 5548 17072 5588 19048
rect 5644 19039 5684 19048
rect 5643 18584 5685 18593
rect 5643 18544 5644 18584
rect 5684 18544 5685 18584
rect 5643 18535 5685 18544
rect 5644 18500 5684 18535
rect 5644 18449 5684 18460
rect 5740 17837 5780 19216
rect 5836 19256 5876 19265
rect 5836 18677 5876 19216
rect 5835 18668 5877 18677
rect 5835 18628 5836 18668
rect 5876 18628 5877 18668
rect 5835 18619 5877 18628
rect 5836 18584 5876 18619
rect 5932 18593 5972 19291
rect 6028 19256 6068 19879
rect 6028 19207 6068 19216
rect 6124 19256 6164 20560
rect 6507 20096 6549 20105
rect 6507 20056 6508 20096
rect 6548 20056 6549 20096
rect 6507 20047 6549 20056
rect 6508 19508 6548 20047
rect 6604 20021 6644 20728
rect 6700 20768 6740 22240
rect 7276 22205 7316 22240
rect 7467 22280 7509 22289
rect 7467 22240 7468 22280
rect 7508 22240 7509 22280
rect 7467 22231 7509 22240
rect 7564 22280 7604 22315
rect 7275 22196 7317 22205
rect 7275 22156 7276 22196
rect 7316 22156 7317 22196
rect 7275 22147 7317 22156
rect 7468 22146 7508 22231
rect 7564 22229 7604 22240
rect 7852 22280 7892 22735
rect 7852 22231 7892 22240
rect 8140 22280 8180 23080
rect 8524 22532 8564 24592
rect 8620 24583 8660 24592
rect 8812 24632 8852 24641
rect 8908 24632 8948 25759
rect 9963 25640 10005 25649
rect 9963 25600 9964 25640
rect 10004 25600 10005 25640
rect 9963 25591 10005 25600
rect 9291 25388 9333 25397
rect 9291 25348 9292 25388
rect 9332 25348 9333 25388
rect 9291 25339 9333 25348
rect 9099 25304 9141 25313
rect 9099 25264 9100 25304
rect 9140 25264 9141 25304
rect 9099 25255 9141 25264
rect 9100 25170 9140 25255
rect 9292 25254 9332 25339
rect 9387 25304 9429 25313
rect 9387 25264 9388 25304
rect 9428 25264 9429 25304
rect 9387 25255 9429 25264
rect 9676 25304 9716 25313
rect 9388 25170 9428 25255
rect 9580 25136 9620 25145
rect 9291 24968 9333 24977
rect 9291 24928 9292 24968
rect 9332 24928 9333 24968
rect 9291 24919 9333 24928
rect 9003 24716 9045 24725
rect 9003 24676 9004 24716
rect 9044 24676 9045 24716
rect 9003 24667 9045 24676
rect 8852 24592 8948 24632
rect 9004 24632 9044 24667
rect 8812 24583 8852 24592
rect 9004 24581 9044 24592
rect 8715 24464 8757 24473
rect 8715 24424 8716 24464
rect 8756 24424 8757 24464
rect 8715 24415 8757 24424
rect 8716 24330 8756 24415
rect 8715 23960 8757 23969
rect 8715 23920 8716 23960
rect 8756 23920 8757 23960
rect 8715 23911 8757 23920
rect 9292 23960 9332 24919
rect 9580 23969 9620 25096
rect 9676 24800 9716 25264
rect 9964 25304 10004 25591
rect 10444 25313 10484 26431
rect 10540 25733 10580 26776
rect 10828 26816 10868 26825
rect 11020 26816 11060 27616
rect 11212 27497 11252 27616
rect 11500 27656 11540 28867
rect 11692 28328 11732 28951
rect 11595 27740 11637 27749
rect 11595 27700 11596 27740
rect 11636 27700 11637 27740
rect 11595 27691 11637 27700
rect 11500 27607 11540 27616
rect 11596 27606 11636 27691
rect 11692 27665 11732 28288
rect 11691 27656 11733 27665
rect 11691 27616 11692 27656
rect 11732 27616 11733 27656
rect 11691 27607 11733 27616
rect 11211 27488 11253 27497
rect 11211 27448 11212 27488
rect 11252 27448 11253 27488
rect 11211 27439 11253 27448
rect 11115 27404 11157 27413
rect 11115 27364 11116 27404
rect 11156 27364 11157 27404
rect 11115 27355 11157 27364
rect 11884 27404 11924 27413
rect 10868 26776 11060 26816
rect 11116 26816 11156 27355
rect 10828 26767 10868 26776
rect 11116 26767 11156 26776
rect 11500 26984 11540 26993
rect 11212 26732 11252 26741
rect 11212 26312 11252 26692
rect 11403 26480 11445 26489
rect 11403 26440 11404 26480
rect 11444 26440 11445 26480
rect 11403 26431 11445 26440
rect 11212 26153 11252 26272
rect 11404 26312 11444 26431
rect 11404 26263 11444 26272
rect 11211 26144 11253 26153
rect 11211 26104 11212 26144
rect 11252 26104 11253 26144
rect 11211 26095 11253 26104
rect 11500 26069 11540 26944
rect 11884 26825 11924 27364
rect 11691 26816 11733 26825
rect 11691 26776 11692 26816
rect 11732 26776 11733 26816
rect 11691 26767 11733 26776
rect 11883 26816 11925 26825
rect 11883 26776 11884 26816
rect 11924 26776 11925 26816
rect 11883 26767 11925 26776
rect 11692 26682 11732 26767
rect 11787 26732 11829 26741
rect 11787 26692 11788 26732
rect 11828 26692 11829 26732
rect 11787 26683 11829 26692
rect 11788 26598 11828 26683
rect 11499 26060 11541 26069
rect 11499 26020 11500 26060
rect 11540 26020 11541 26060
rect 11499 26011 11541 26020
rect 10539 25724 10581 25733
rect 10539 25684 10540 25724
rect 10580 25684 10581 25724
rect 10539 25675 10581 25684
rect 9867 25136 9909 25145
rect 9867 25096 9868 25136
rect 9908 25096 9909 25136
rect 9867 25087 9909 25096
rect 9868 25002 9908 25087
rect 9964 24800 10004 25264
rect 10060 25304 10100 25313
rect 10060 24977 10100 25264
rect 10156 25304 10196 25313
rect 10059 24968 10101 24977
rect 10059 24928 10060 24968
rect 10100 24928 10101 24968
rect 10059 24919 10101 24928
rect 9676 24751 9716 24760
rect 9868 24760 10004 24800
rect 8716 23120 8756 23911
rect 9003 23288 9045 23297
rect 9003 23248 9004 23288
rect 9044 23248 9045 23288
rect 9003 23239 9045 23248
rect 8716 23071 8756 23080
rect 8811 23120 8853 23129
rect 8811 23080 8812 23120
rect 8852 23080 8853 23120
rect 8811 23071 8853 23080
rect 9004 23120 9044 23239
rect 9004 23071 9044 23080
rect 8812 22986 8852 23071
rect 9292 23045 9332 23920
rect 9579 23960 9621 23969
rect 9579 23920 9580 23960
rect 9620 23920 9621 23960
rect 9579 23911 9621 23920
rect 9676 23960 9716 23969
rect 9716 23920 9812 23960
rect 9676 23911 9716 23920
rect 9291 23036 9333 23045
rect 9291 22996 9292 23036
rect 9332 22996 9333 23036
rect 9291 22987 9333 22996
rect 9003 22952 9045 22961
rect 9003 22912 9004 22952
rect 9044 22912 9045 22952
rect 9003 22903 9045 22912
rect 9004 22818 9044 22903
rect 9196 22868 9236 22877
rect 8524 22483 8564 22492
rect 9196 22280 9236 22828
rect 9579 22868 9621 22877
rect 9579 22828 9580 22868
rect 9620 22828 9621 22868
rect 9579 22819 9621 22828
rect 9292 22280 9332 22289
rect 9196 22240 9292 22280
rect 7372 21608 7412 21617
rect 6892 20768 6932 20777
rect 6700 20719 6740 20728
rect 6796 20728 6892 20768
rect 6796 20357 6836 20728
rect 6892 20719 6932 20728
rect 6795 20348 6837 20357
rect 6795 20308 6796 20348
rect 6836 20308 6837 20348
rect 6795 20299 6837 20308
rect 6603 20012 6645 20021
rect 6603 19972 6604 20012
rect 6644 19972 6645 20012
rect 6603 19963 6645 19972
rect 6508 19459 6548 19468
rect 6604 19433 6644 19963
rect 6603 19424 6645 19433
rect 6603 19384 6604 19424
rect 6644 19384 6645 19424
rect 6603 19375 6645 19384
rect 6219 19340 6261 19349
rect 6219 19300 6220 19340
rect 6260 19300 6261 19340
rect 6219 19291 6261 19300
rect 6124 19207 6164 19216
rect 6220 19256 6260 19291
rect 6220 19205 6260 19216
rect 6316 19256 6356 19265
rect 6508 19256 6548 19265
rect 6700 19256 6740 19265
rect 6356 19216 6508 19256
rect 6316 19207 6356 19216
rect 6508 19207 6548 19216
rect 6604 19216 6700 19256
rect 6219 19088 6261 19097
rect 6219 19048 6220 19088
rect 6260 19048 6261 19088
rect 6219 19039 6261 19048
rect 6220 18845 6260 19039
rect 6219 18836 6261 18845
rect 6604 18836 6644 19216
rect 6700 19207 6740 19216
rect 6796 19256 6836 20299
rect 7372 20105 7412 21568
rect 8140 21533 8180 22240
rect 9292 22231 9332 22240
rect 9580 22280 9620 22819
rect 9772 22280 9812 23920
rect 9868 23792 9908 24760
rect 9963 24632 10005 24641
rect 9963 24592 9964 24632
rect 10004 24592 10005 24632
rect 9963 24583 10005 24592
rect 9964 24498 10004 24583
rect 10156 23960 10196 25264
rect 10443 25304 10485 25313
rect 10443 25264 10444 25304
rect 10484 25264 10485 25304
rect 10443 25255 10485 25264
rect 10540 25304 10580 25675
rect 11980 25649 12020 28960
rect 12556 28328 12596 28337
rect 12459 28244 12501 28253
rect 12459 28204 12460 28244
rect 12500 28204 12501 28244
rect 12459 28195 12501 28204
rect 12075 27656 12117 27665
rect 12075 27616 12076 27656
rect 12116 27616 12117 27656
rect 12075 27607 12117 27616
rect 12076 27522 12116 27607
rect 12364 27404 12404 27413
rect 12075 26144 12117 26153
rect 12075 26104 12076 26144
rect 12116 26104 12117 26144
rect 12075 26095 12117 26104
rect 12076 26010 12116 26095
rect 12075 25724 12117 25733
rect 12075 25684 12076 25724
rect 12116 25684 12117 25724
rect 12075 25675 12117 25684
rect 10731 25640 10773 25649
rect 10731 25600 10732 25640
rect 10772 25600 10773 25640
rect 10731 25591 10773 25600
rect 11979 25640 12021 25649
rect 11979 25600 11980 25640
rect 12020 25600 12021 25640
rect 11979 25591 12021 25600
rect 10636 25313 10676 25398
rect 10540 25136 10580 25264
rect 10635 25304 10677 25313
rect 10635 25264 10636 25304
rect 10676 25264 10677 25304
rect 10635 25255 10677 25264
rect 10732 25304 10772 25591
rect 11884 25481 11924 25566
rect 11019 25472 11061 25481
rect 11019 25432 11020 25472
rect 11060 25432 11061 25472
rect 11019 25423 11061 25432
rect 11883 25472 11925 25481
rect 11883 25432 11884 25472
rect 11924 25432 11925 25472
rect 11883 25423 11925 25432
rect 10732 25255 10772 25264
rect 10827 25304 10869 25313
rect 10827 25264 10828 25304
rect 10868 25264 10869 25304
rect 10827 25255 10869 25264
rect 11020 25304 11060 25423
rect 11020 25255 11060 25264
rect 11883 25304 11925 25313
rect 11883 25264 11884 25304
rect 11924 25264 11925 25304
rect 11883 25255 11925 25264
rect 12076 25304 12116 25675
rect 12076 25255 12116 25264
rect 12171 25304 12213 25313
rect 12171 25264 12172 25304
rect 12212 25264 12213 25304
rect 12171 25255 12213 25264
rect 10828 25170 10868 25255
rect 11884 25170 11924 25255
rect 12172 25170 12212 25255
rect 10444 25096 10580 25136
rect 10635 25136 10677 25145
rect 10635 25096 10636 25136
rect 10676 25096 10677 25136
rect 10251 24968 10293 24977
rect 10251 24928 10252 24968
rect 10292 24928 10293 24968
rect 10251 24919 10293 24928
rect 10252 24632 10292 24919
rect 10347 24716 10389 24725
rect 10347 24676 10348 24716
rect 10388 24676 10389 24716
rect 10347 24667 10389 24676
rect 10252 24583 10292 24592
rect 10348 24582 10388 24667
rect 10156 23920 10292 23960
rect 9964 23792 10004 23801
rect 9868 23752 9964 23792
rect 9964 23743 10004 23752
rect 10059 23792 10101 23801
rect 10059 23752 10060 23792
rect 10100 23752 10101 23792
rect 10059 23743 10101 23752
rect 10156 23792 10196 23801
rect 10060 23658 10100 23743
rect 9868 23624 9908 23633
rect 9868 23297 9908 23584
rect 9867 23288 9909 23297
rect 10156 23288 10196 23752
rect 9867 23248 9868 23288
rect 9908 23248 9909 23288
rect 9867 23239 9909 23248
rect 10060 23248 10196 23288
rect 9868 23120 9908 23131
rect 9868 23045 9908 23080
rect 9867 23036 9909 23045
rect 10060 23036 10100 23248
rect 10155 23120 10197 23129
rect 10252 23120 10292 23920
rect 10444 23876 10484 25096
rect 10635 25087 10677 25096
rect 11692 25136 11732 25145
rect 10636 24464 10676 25087
rect 10827 25052 10869 25061
rect 10827 25012 10828 25052
rect 10868 25012 10869 25052
rect 10827 25003 10869 25012
rect 10828 24800 10868 25003
rect 11307 24968 11349 24977
rect 11307 24928 11308 24968
rect 11348 24928 11349 24968
rect 11307 24919 11349 24928
rect 10828 24751 10868 24760
rect 11308 24473 11348 24919
rect 11692 24725 11732 25096
rect 11691 24716 11733 24725
rect 11691 24676 11692 24716
rect 11732 24676 11733 24716
rect 11691 24667 11733 24676
rect 12364 24641 12404 27364
rect 12460 27068 12500 28195
rect 12556 27917 12596 28288
rect 12555 27908 12597 27917
rect 12555 27868 12556 27908
rect 12596 27868 12597 27908
rect 12555 27859 12597 27868
rect 12747 27740 12789 27749
rect 12747 27700 12748 27740
rect 12788 27700 12789 27740
rect 12747 27691 12789 27700
rect 12460 27019 12500 27028
rect 12460 26816 12500 26825
rect 12460 26657 12500 26776
rect 12652 26816 12692 26825
rect 12459 26648 12501 26657
rect 12459 26608 12460 26648
rect 12500 26608 12501 26648
rect 12459 26599 12501 26608
rect 12460 25976 12500 25985
rect 12652 25976 12692 26776
rect 12748 26816 12788 27691
rect 12844 26816 12884 30547
rect 12940 30185 12980 31891
rect 13132 31697 13172 32059
rect 13131 31688 13173 31697
rect 13131 31648 13132 31688
rect 13172 31648 13173 31688
rect 13131 31639 13173 31648
rect 13228 31520 13268 32068
rect 13420 31940 13460 31949
rect 13036 31480 13268 31520
rect 13323 31520 13365 31529
rect 13323 31480 13324 31520
rect 13364 31480 13365 31520
rect 12939 30176 12981 30185
rect 12939 30136 12940 30176
rect 12980 30136 12981 30176
rect 12939 30127 12981 30136
rect 13036 29840 13076 31480
rect 13323 31471 13365 31480
rect 13227 31352 13269 31361
rect 13227 31312 13228 31352
rect 13268 31312 13269 31352
rect 13227 31303 13269 31312
rect 13324 31352 13364 31471
rect 13324 31303 13364 31312
rect 13228 31218 13268 31303
rect 13420 30848 13460 31900
rect 13515 31436 13557 31445
rect 13515 31396 13516 31436
rect 13556 31396 13557 31436
rect 13515 31387 13557 31396
rect 13516 31352 13556 31387
rect 13516 31301 13556 31312
rect 13612 31352 13652 31363
rect 13612 31277 13652 31312
rect 13611 31268 13653 31277
rect 13611 31228 13612 31268
rect 13652 31228 13653 31268
rect 13611 31219 13653 31228
rect 13708 31268 13748 32311
rect 13803 32192 13845 32201
rect 13803 32152 13804 32192
rect 13844 32152 13845 32192
rect 13803 32143 13845 32152
rect 13804 31352 13844 32143
rect 13995 31604 14037 31613
rect 13995 31564 13996 31604
rect 14036 31564 14037 31604
rect 13995 31555 14037 31564
rect 13996 31470 14036 31555
rect 13996 31352 14036 31361
rect 13804 31303 13844 31312
rect 13900 31312 13996 31352
rect 13708 31219 13748 31228
rect 13515 31100 13557 31109
rect 13515 31060 13516 31100
rect 13556 31060 13557 31100
rect 13515 31051 13557 31060
rect 13324 30808 13460 30848
rect 13131 30680 13173 30689
rect 13131 30640 13132 30680
rect 13172 30640 13173 30680
rect 13131 30631 13173 30640
rect 13132 30546 13172 30631
rect 13036 29000 13076 29800
rect 13324 29168 13364 30808
rect 13516 30764 13556 31051
rect 13611 31016 13653 31025
rect 13611 30976 13612 31016
rect 13652 30976 13653 31016
rect 13611 30967 13653 30976
rect 13516 30715 13556 30724
rect 13420 30680 13460 30689
rect 13420 30596 13460 30640
rect 13612 30596 13652 30967
rect 13900 30857 13940 31312
rect 13996 31303 14036 31312
rect 14092 31184 14132 32488
rect 14283 32488 14284 32528
rect 14324 32488 14325 32528
rect 14283 32479 14325 32488
rect 14284 32192 14324 32203
rect 14476 32201 14516 32286
rect 14284 32117 14324 32152
rect 14475 32192 14517 32201
rect 14475 32152 14476 32192
rect 14516 32152 14517 32192
rect 14475 32143 14517 32152
rect 14572 32192 14612 33067
rect 14764 32369 14804 33664
rect 15244 33032 15284 35848
rect 15339 35216 15381 35225
rect 15436 35216 15476 36688
rect 15627 36728 15669 36737
rect 15627 36688 15628 36728
rect 15668 36688 15669 36728
rect 15627 36679 15669 36688
rect 15628 36594 15668 36679
rect 15628 35888 15668 35897
rect 15724 35888 15764 37192
rect 16396 36905 16436 37360
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 16395 36896 16437 36905
rect 16395 36856 16396 36896
rect 16436 36856 16437 36896
rect 16395 36847 16437 36856
rect 16491 36812 16533 36821
rect 16491 36772 16492 36812
rect 16532 36772 16533 36812
rect 16491 36763 16533 36772
rect 17547 36812 17589 36821
rect 17547 36772 17548 36812
rect 17588 36772 17589 36812
rect 17547 36763 17589 36772
rect 15668 35848 15764 35888
rect 15820 36728 15860 36737
rect 15628 35839 15668 35848
rect 15820 35729 15860 36688
rect 16492 36678 16532 36763
rect 16683 36728 16725 36737
rect 16683 36688 16684 36728
rect 16724 36688 16725 36728
rect 16683 36679 16725 36688
rect 16780 36728 16820 36737
rect 16684 36594 16724 36679
rect 16011 36560 16053 36569
rect 16011 36520 16012 36560
rect 16052 36520 16053 36560
rect 16011 36511 16053 36520
rect 16012 35888 16052 36511
rect 16012 35839 16052 35848
rect 15819 35720 15861 35729
rect 15819 35680 15820 35720
rect 15860 35680 15861 35720
rect 15819 35671 15861 35680
rect 15339 35176 15340 35216
rect 15380 35176 15476 35216
rect 16203 35216 16245 35225
rect 16203 35176 16204 35216
rect 16244 35176 16245 35216
rect 15339 35167 15381 35176
rect 16203 35167 16245 35176
rect 16587 35216 16629 35225
rect 16587 35176 16588 35216
rect 16628 35176 16629 35216
rect 16587 35167 16629 35176
rect 16684 35216 16724 35225
rect 15340 35082 15380 35167
rect 16204 35082 16244 35167
rect 16491 35048 16533 35057
rect 16491 35008 16492 35048
rect 16532 35008 16533 35048
rect 16491 34999 16533 35008
rect 15820 34376 15860 34385
rect 15820 33713 15860 34336
rect 16108 33788 16148 33797
rect 15628 33704 15668 33713
rect 15531 33116 15573 33125
rect 15531 33076 15532 33116
rect 15572 33076 15573 33116
rect 15531 33067 15573 33076
rect 15244 32992 15476 33032
rect 14955 32864 14997 32873
rect 14955 32824 14956 32864
rect 14996 32824 14997 32864
rect 14955 32815 14997 32824
rect 15244 32864 15284 32873
rect 14859 32528 14901 32537
rect 14859 32488 14860 32528
rect 14900 32488 14901 32528
rect 14859 32479 14901 32488
rect 14763 32360 14805 32369
rect 14763 32320 14764 32360
rect 14804 32320 14805 32360
rect 14763 32311 14805 32320
rect 14668 32201 14708 32286
rect 14572 32143 14612 32152
rect 14667 32192 14709 32201
rect 14667 32152 14668 32192
rect 14708 32152 14709 32192
rect 14667 32143 14709 32152
rect 14764 32192 14804 32201
rect 14283 32108 14325 32117
rect 14283 32068 14284 32108
rect 14324 32068 14325 32108
rect 14283 32059 14325 32068
rect 14764 31445 14804 32152
rect 14187 31436 14229 31445
rect 14187 31396 14188 31436
rect 14228 31396 14229 31436
rect 14187 31387 14229 31396
rect 14763 31436 14805 31445
rect 14763 31396 14764 31436
rect 14804 31396 14805 31436
rect 14763 31387 14805 31396
rect 14188 31352 14228 31387
rect 14188 31301 14228 31312
rect 14283 31352 14325 31361
rect 14283 31312 14284 31352
rect 14324 31312 14325 31352
rect 14283 31303 14325 31312
rect 14667 31352 14709 31361
rect 14667 31312 14668 31352
rect 14708 31312 14709 31352
rect 14667 31303 14709 31312
rect 14284 31218 14324 31303
rect 14668 31218 14708 31303
rect 14764 31277 14804 31387
rect 14860 31352 14900 32479
rect 14956 32024 14996 32815
rect 15147 32696 15189 32705
rect 15147 32656 15148 32696
rect 15188 32656 15189 32696
rect 15147 32647 15189 32656
rect 14956 31975 14996 31984
rect 14955 31856 14997 31865
rect 14955 31816 14956 31856
rect 14996 31816 14997 31856
rect 14955 31807 14997 31816
rect 14860 31303 14900 31312
rect 14956 31352 14996 31807
rect 15148 31772 15188 32647
rect 15052 31732 15188 31772
rect 15052 31352 15092 31732
rect 15147 31604 15189 31613
rect 15147 31564 15148 31604
rect 15188 31564 15189 31604
rect 15147 31555 15189 31564
rect 15148 31470 15188 31555
rect 15148 31352 15188 31361
rect 15052 31312 15148 31352
rect 14956 31303 14996 31312
rect 15148 31303 15188 31312
rect 14763 31268 14805 31277
rect 14763 31228 14764 31268
rect 14804 31228 14805 31268
rect 14763 31219 14805 31228
rect 14572 31184 14612 31193
rect 14092 31144 14228 31184
rect 13995 31016 14037 31025
rect 14188 31016 14228 31144
rect 13995 30976 13996 31016
rect 14036 30976 14037 31016
rect 13995 30967 14037 30976
rect 14092 30976 14228 31016
rect 13899 30848 13941 30857
rect 13899 30808 13900 30848
rect 13940 30808 13941 30848
rect 13899 30799 13941 30808
rect 13996 30680 14036 30967
rect 13996 30631 14036 30640
rect 13420 30556 13652 30596
rect 13803 30428 13845 30437
rect 13803 30388 13804 30428
rect 13844 30388 13845 30428
rect 13803 30379 13845 30388
rect 13804 30294 13844 30379
rect 13419 30260 13461 30269
rect 13419 30220 13420 30260
rect 13460 30220 13461 30260
rect 13419 30211 13461 30220
rect 13420 30092 13460 30211
rect 13803 30176 13845 30185
rect 13803 30136 13804 30176
rect 13844 30136 13845 30176
rect 13803 30127 13845 30136
rect 13420 30043 13460 30052
rect 13708 29177 13748 29262
rect 13516 29168 13556 29177
rect 13324 29128 13516 29168
rect 13516 29119 13556 29128
rect 13707 29168 13749 29177
rect 13707 29128 13708 29168
rect 13748 29128 13749 29168
rect 13707 29119 13749 29128
rect 13804 29000 13844 30127
rect 13036 28960 13172 29000
rect 12939 28244 12981 28253
rect 12939 28204 12940 28244
rect 12980 28204 12981 28244
rect 12939 28195 12981 28204
rect 12940 28110 12980 28195
rect 13035 27656 13077 27665
rect 13035 27616 13036 27656
rect 13076 27616 13077 27656
rect 13035 27607 13077 27616
rect 13036 27522 13076 27607
rect 12940 26816 12980 26825
rect 12844 26776 12940 26816
rect 12748 26767 12788 26776
rect 12940 26767 12980 26776
rect 13036 26816 13076 26825
rect 13036 26657 13076 26776
rect 13132 26741 13172 28960
rect 13708 28960 13844 29000
rect 13611 28916 13653 28925
rect 13611 28876 13612 28916
rect 13652 28876 13653 28916
rect 13611 28867 13653 28876
rect 13612 28782 13652 28867
rect 13612 28496 13652 28505
rect 13324 27656 13364 27665
rect 13324 27497 13364 27616
rect 13323 27488 13365 27497
rect 13323 27448 13324 27488
rect 13364 27448 13365 27488
rect 13323 27439 13365 27448
rect 13228 26984 13268 26993
rect 13268 26944 13556 26984
rect 13228 26935 13268 26944
rect 13228 26816 13268 26825
rect 13131 26732 13173 26741
rect 13131 26692 13132 26732
rect 13172 26692 13173 26732
rect 13131 26683 13173 26692
rect 13035 26648 13077 26657
rect 13035 26608 13036 26648
rect 13076 26608 13077 26648
rect 13035 26599 13077 26608
rect 13131 26564 13173 26573
rect 13131 26524 13132 26564
rect 13172 26524 13173 26564
rect 13131 26515 13173 26524
rect 13035 26144 13077 26153
rect 13035 26104 13036 26144
rect 13076 26104 13077 26144
rect 13035 26095 13077 26104
rect 12652 25936 12884 25976
rect 12460 24893 12500 25936
rect 12747 25808 12789 25817
rect 12747 25768 12748 25808
rect 12788 25768 12789 25808
rect 12747 25759 12789 25768
rect 12651 25388 12693 25397
rect 12651 25348 12652 25388
rect 12692 25348 12693 25388
rect 12651 25339 12693 25348
rect 12555 25304 12597 25313
rect 12555 25264 12556 25304
rect 12596 25264 12597 25304
rect 12555 25255 12597 25264
rect 12556 25170 12596 25255
rect 12652 25254 12692 25339
rect 12748 25327 12788 25759
rect 12748 25278 12788 25287
rect 12844 25220 12884 25936
rect 12939 25640 12981 25649
rect 12939 25600 12940 25640
rect 12980 25600 12981 25640
rect 12939 25591 12981 25600
rect 12759 25180 12884 25220
rect 12759 25136 12799 25180
rect 12748 25096 12799 25136
rect 12459 24884 12501 24893
rect 12459 24844 12460 24884
rect 12500 24844 12501 24884
rect 12459 24835 12501 24844
rect 11979 24632 12021 24641
rect 11979 24592 11980 24632
rect 12020 24592 12021 24632
rect 11979 24583 12021 24592
rect 12363 24632 12405 24641
rect 12363 24592 12364 24632
rect 12404 24592 12405 24632
rect 12363 24583 12405 24592
rect 11980 24498 12020 24583
rect 12651 24548 12693 24557
rect 12651 24508 12652 24548
rect 12692 24508 12693 24548
rect 12651 24499 12693 24508
rect 10636 24415 10676 24424
rect 11307 24464 11349 24473
rect 11307 24424 11308 24464
rect 11348 24424 11349 24464
rect 11307 24415 11349 24424
rect 10444 23827 10484 23836
rect 11212 23792 11252 23801
rect 11212 23717 11252 23752
rect 11883 23792 11925 23801
rect 11883 23752 11884 23792
rect 11924 23752 11925 23792
rect 11883 23743 11925 23752
rect 11211 23708 11253 23717
rect 11211 23668 11212 23708
rect 11252 23668 11253 23708
rect 11211 23659 11253 23668
rect 11691 23708 11733 23717
rect 11691 23668 11692 23708
rect 11732 23668 11733 23708
rect 11691 23659 11733 23668
rect 11212 23129 11252 23659
rect 10155 23080 10156 23120
rect 10196 23080 10292 23120
rect 10732 23120 10772 23129
rect 10155 23071 10197 23080
rect 9867 22996 9868 23036
rect 9908 22996 9909 23036
rect 9867 22987 9909 22996
rect 9964 22996 10100 23036
rect 9964 22616 10004 22996
rect 10059 22868 10101 22877
rect 10059 22828 10060 22868
rect 10100 22828 10101 22868
rect 10059 22819 10101 22828
rect 10060 22734 10100 22819
rect 9964 22576 10100 22616
rect 9964 22280 10004 22289
rect 9772 22240 9964 22280
rect 9580 22231 9620 22240
rect 9964 22231 10004 22240
rect 8235 22196 8277 22205
rect 8235 22156 8236 22196
rect 8276 22156 8277 22196
rect 8235 22147 8277 22156
rect 8139 21524 8181 21533
rect 8139 21484 8140 21524
rect 8180 21484 8181 21524
rect 8139 21475 8181 21484
rect 7755 20852 7797 20861
rect 7755 20812 7756 20852
rect 7796 20812 7797 20852
rect 7755 20803 7797 20812
rect 7756 20768 7796 20803
rect 7756 20717 7796 20728
rect 8044 20264 8084 20273
rect 8236 20264 8276 22147
rect 9388 22112 9428 22121
rect 8812 22072 9388 22112
rect 8523 21524 8565 21533
rect 8523 21484 8524 21524
rect 8564 21484 8565 21524
rect 8523 21475 8565 21484
rect 8524 21390 8564 21475
rect 8812 20768 8852 22072
rect 9388 22063 9428 22072
rect 9580 21608 9620 21617
rect 9100 21568 9580 21608
rect 8907 20852 8949 20861
rect 8907 20812 8908 20852
rect 8948 20812 8949 20852
rect 8907 20803 8949 20812
rect 8812 20719 8852 20728
rect 8908 20768 8948 20803
rect 8908 20717 8948 20728
rect 9100 20768 9140 21568
rect 9580 21559 9620 21568
rect 9676 21608 9716 21617
rect 9100 20719 9140 20728
rect 9003 20684 9045 20693
rect 9003 20644 9004 20684
rect 9044 20644 9045 20684
rect 9003 20635 9045 20644
rect 9004 20550 9044 20635
rect 9292 20600 9332 20609
rect 9100 20560 9292 20600
rect 8084 20224 8276 20264
rect 8044 20215 8084 20224
rect 8812 20180 8852 20189
rect 9100 20180 9140 20560
rect 9292 20551 9332 20560
rect 8852 20140 9140 20180
rect 8812 20131 8852 20140
rect 6891 20096 6933 20105
rect 6891 20056 6892 20096
rect 6932 20056 6933 20096
rect 6891 20047 6933 20056
rect 7371 20096 7413 20105
rect 7371 20056 7372 20096
rect 7412 20056 7413 20096
rect 7371 20047 7413 20056
rect 8524 20096 8564 20105
rect 8715 20096 8757 20105
rect 8564 20056 8660 20096
rect 8524 20047 8564 20056
rect 6892 19962 6932 20047
rect 8428 19844 8468 19853
rect 8236 19804 8428 19844
rect 6988 19384 7316 19424
rect 6988 19256 7028 19384
rect 6836 19216 6988 19256
rect 6796 19207 6836 19216
rect 6988 19207 7028 19216
rect 7180 19256 7220 19265
rect 6219 18796 6220 18836
rect 6260 18796 6261 18836
rect 6219 18787 6261 18796
rect 6316 18796 6644 18836
rect 7084 19172 7124 19181
rect 5836 18533 5876 18544
rect 5931 18584 5973 18593
rect 5931 18544 5932 18584
rect 5972 18544 5973 18584
rect 5931 18535 5973 18544
rect 6220 18584 6260 18787
rect 5836 18332 5876 18341
rect 5836 18173 5876 18292
rect 5931 18332 5973 18341
rect 5931 18292 5932 18332
rect 5972 18292 5973 18332
rect 5931 18283 5973 18292
rect 5835 18164 5877 18173
rect 5835 18124 5836 18164
rect 5876 18124 5877 18164
rect 5835 18115 5877 18124
rect 5739 17828 5781 17837
rect 5739 17788 5740 17828
rect 5780 17788 5781 17828
rect 5739 17779 5781 17788
rect 5836 17744 5876 17753
rect 5739 17660 5781 17669
rect 5836 17660 5876 17704
rect 5932 17744 5972 18283
rect 6123 17828 6165 17837
rect 6123 17788 6124 17828
rect 6164 17788 6165 17828
rect 6123 17779 6165 17788
rect 5932 17695 5972 17704
rect 6027 17744 6069 17753
rect 6027 17704 6028 17744
rect 6068 17704 6069 17744
rect 6027 17695 6069 17704
rect 6124 17744 6164 17779
rect 5739 17620 5740 17660
rect 5780 17620 5876 17660
rect 5739 17611 5781 17620
rect 6028 17610 6068 17695
rect 6124 17693 6164 17704
rect 5643 17576 5685 17585
rect 6220 17576 6260 18544
rect 5643 17536 5644 17576
rect 5684 17536 5685 17576
rect 5643 17527 5685 17536
rect 6124 17536 6260 17576
rect 6316 17744 6356 18796
rect 7084 18752 7124 19132
rect 7180 18929 7220 19216
rect 7179 18920 7221 18929
rect 7179 18880 7180 18920
rect 7220 18880 7221 18920
rect 7179 18871 7221 18880
rect 6892 18712 7124 18752
rect 6412 18593 6452 18678
rect 6411 18584 6453 18593
rect 6411 18544 6412 18584
rect 6452 18544 6453 18584
rect 6411 18535 6453 18544
rect 6508 18584 6548 18595
rect 6508 18509 6548 18544
rect 6603 18584 6645 18593
rect 6603 18544 6604 18584
rect 6644 18544 6645 18584
rect 6603 18535 6645 18544
rect 6700 18584 6740 18593
rect 6507 18500 6549 18509
rect 6507 18460 6508 18500
rect 6548 18460 6549 18500
rect 6507 18451 6549 18460
rect 6411 18416 6453 18425
rect 6411 18376 6412 18416
rect 6452 18376 6453 18416
rect 6411 18367 6453 18376
rect 6412 18282 6452 18367
rect 6604 17912 6644 18535
rect 6700 17921 6740 18544
rect 6796 18584 6836 18593
rect 6796 18425 6836 18544
rect 6892 18584 6932 18712
rect 6795 18416 6837 18425
rect 6795 18376 6796 18416
rect 6836 18376 6837 18416
rect 6795 18367 6837 18376
rect 6604 17863 6644 17872
rect 6699 17912 6741 17921
rect 6699 17872 6700 17912
rect 6740 17872 6741 17912
rect 6699 17863 6741 17872
rect 6508 17744 6548 17753
rect 6316 17704 6508 17744
rect 5644 17442 5684 17527
rect 5932 17072 5972 17081
rect 5548 17032 5932 17072
rect 5932 17023 5972 17032
rect 6124 17072 6164 17536
rect 6220 17240 6260 17249
rect 6316 17240 6356 17704
rect 6508 17695 6548 17704
rect 6603 17744 6645 17753
rect 6700 17744 6740 17753
rect 6603 17704 6604 17744
rect 6644 17704 6700 17744
rect 6603 17695 6645 17704
rect 6700 17695 6740 17704
rect 6795 17744 6837 17753
rect 6795 17704 6796 17744
rect 6836 17704 6837 17744
rect 6795 17695 6837 17704
rect 6796 17610 6836 17695
rect 6892 17492 6932 18544
rect 6988 18584 7028 18593
rect 7180 18584 7220 18593
rect 7028 18544 7180 18584
rect 6988 18535 7028 18544
rect 7180 18535 7220 18544
rect 6988 17753 7028 17838
rect 6987 17744 7029 17753
rect 7276 17744 7316 19384
rect 8044 19265 8084 19350
rect 7852 19256 7892 19265
rect 7371 18920 7413 18929
rect 7371 18880 7372 18920
rect 7412 18880 7413 18920
rect 7371 18871 7413 18880
rect 7372 18509 7412 18871
rect 7852 18752 7892 19216
rect 8043 19256 8085 19265
rect 8043 19216 8044 19256
rect 8084 19216 8085 19256
rect 8043 19207 8085 19216
rect 7948 19088 7988 19097
rect 7988 19048 8180 19088
rect 7948 19039 7988 19048
rect 7852 18712 7988 18752
rect 7467 18668 7509 18677
rect 7467 18628 7468 18668
rect 7508 18628 7509 18668
rect 7467 18619 7509 18628
rect 7371 18500 7413 18509
rect 7371 18460 7372 18500
rect 7412 18460 7413 18500
rect 7371 18451 7413 18460
rect 6987 17704 6988 17744
rect 7028 17704 7316 17744
rect 7372 17744 7412 18451
rect 6987 17695 7029 17704
rect 7372 17695 7412 17704
rect 7468 17660 7508 18619
rect 7852 18584 7892 18593
rect 6987 17576 7029 17585
rect 7468 17576 7508 17620
rect 6987 17536 6988 17576
rect 7028 17536 7029 17576
rect 6987 17527 7029 17536
rect 7276 17536 7508 17576
rect 7564 18544 7852 18584
rect 6260 17200 6356 17240
rect 6700 17452 6932 17492
rect 6220 17191 6260 17200
rect 6124 17023 6164 17032
rect 6412 17072 6452 17081
rect 6315 16988 6357 16997
rect 6315 16948 6316 16988
rect 6356 16948 6357 16988
rect 6315 16939 6357 16948
rect 5260 16444 5588 16484
rect 5260 16232 5300 16444
rect 5260 16183 5300 16192
rect 5356 16232 5396 16241
rect 5396 16192 5492 16232
rect 5356 16183 5396 16192
rect 5356 16064 5404 16073
rect 5403 16024 5404 16064
rect 5356 16015 5404 16024
rect 5363 15936 5403 16015
rect 5452 15821 5492 16192
rect 5451 15812 5493 15821
rect 5451 15772 5452 15812
rect 5492 15772 5493 15812
rect 5451 15763 5493 15772
rect 4971 15688 4972 15728
rect 5012 15688 5013 15728
rect 4299 15644 4341 15653
rect 4299 15604 4300 15644
rect 4340 15604 4341 15644
rect 4299 15595 4341 15604
rect 4108 15436 4244 15476
rect 3819 15224 3861 15233
rect 3819 15184 3820 15224
rect 3860 15184 3861 15224
rect 3819 15175 3861 15184
rect 4011 15140 4053 15149
rect 4011 15100 4012 15140
rect 4052 15100 4053 15140
rect 4011 15091 4053 15100
rect 2380 14671 2420 14680
rect 2763 14720 2805 14729
rect 2763 14680 2764 14720
rect 2804 14680 2805 14720
rect 2763 14671 2805 14680
rect 3627 14720 3669 14729
rect 3627 14680 3628 14720
rect 3668 14680 3669 14720
rect 3627 14671 3669 14680
rect 2764 14586 2804 14671
rect 3628 14586 3668 14671
rect 4012 14309 4052 15091
rect 4011 14300 4053 14309
rect 4011 14260 4012 14300
rect 4052 14260 4053 14300
rect 4011 14251 4053 14260
rect 4012 14216 4052 14251
rect 4108 14225 4148 15436
rect 4203 15308 4245 15317
rect 4203 15268 4204 15308
rect 4244 15268 4245 15308
rect 4203 15259 4245 15268
rect 4204 15174 4244 15259
rect 4300 14552 4340 15595
rect 4780 15308 4820 15688
rect 4971 15679 5013 15688
rect 5068 15688 5204 15728
rect 5355 15728 5397 15737
rect 5355 15688 5356 15728
rect 5396 15688 5397 15728
rect 4876 15560 4916 15569
rect 4876 15485 4916 15520
rect 4875 15476 4917 15485
rect 4875 15436 4876 15476
rect 4916 15436 4917 15476
rect 4875 15427 4917 15436
rect 4876 15425 4916 15427
rect 4780 15268 4916 15308
rect 4779 15140 4821 15149
rect 4779 15100 4780 15140
rect 4820 15100 4821 15140
rect 4779 15091 4821 15100
rect 4780 14972 4820 15091
rect 4780 14923 4820 14932
rect 4204 14512 4340 14552
rect 3244 14176 3764 14216
rect 1323 14132 1365 14141
rect 1323 14092 1324 14132
rect 1364 14092 1365 14132
rect 1323 14083 1365 14092
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 3244 14048 3284 14176
rect 3244 13999 3284 14008
rect 3436 14048 3476 14057
rect 3476 14008 3668 14048
rect 3436 13999 3476 14008
rect 3436 13796 3476 13805
rect 3476 13756 3572 13796
rect 3436 13747 3476 13756
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3436 13376 3476 13385
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 2955 13040 2997 13049
rect 2955 13000 2956 13040
rect 2996 13000 2997 13040
rect 2955 12991 2997 13000
rect 652 12704 692 12713
rect 652 12377 692 12664
rect 2956 12536 2996 12991
rect 2956 12487 2996 12496
rect 3340 12536 3380 12545
rect 3436 12536 3476 13336
rect 3532 12629 3572 13756
rect 3628 13217 3668 14008
rect 3724 13628 3764 14176
rect 4012 14165 4052 14176
rect 4107 14216 4149 14225
rect 4107 14176 4108 14216
rect 4148 14176 4149 14216
rect 4204 14216 4244 14512
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4300 14216 4340 14225
rect 4204 14176 4300 14216
rect 4107 14167 4149 14176
rect 4300 14167 4340 14176
rect 4491 14216 4533 14225
rect 4491 14176 4492 14216
rect 4532 14176 4533 14216
rect 4491 14167 4533 14176
rect 4683 14216 4725 14225
rect 4683 14176 4684 14216
rect 4724 14176 4725 14216
rect 4876 14216 4916 15268
rect 4876 14176 4917 14216
rect 4683 14167 4725 14176
rect 4204 14031 4244 14059
rect 4492 14048 4532 14167
rect 4588 14048 4628 14057
rect 4492 14008 4588 14048
rect 4588 13999 4628 14008
rect 4684 14048 4724 14167
rect 4877 14132 4917 14176
rect 4684 13999 4724 14008
rect 4876 14092 4917 14132
rect 4876 14048 4916 14092
rect 4876 13999 4916 14008
rect 4204 13973 4244 13991
rect 4203 13964 4245 13973
rect 4203 13924 4204 13964
rect 4244 13924 4245 13964
rect 4203 13915 4245 13924
rect 3819 13880 3861 13889
rect 3819 13840 3820 13880
rect 3860 13840 3861 13880
rect 3819 13831 3861 13840
rect 4876 13880 4916 13889
rect 4972 13880 5012 15679
rect 5068 14552 5108 15688
rect 5355 15679 5397 15688
rect 5164 15560 5204 15569
rect 5164 15401 5204 15520
rect 5356 15560 5396 15679
rect 5356 15511 5396 15520
rect 5451 15560 5493 15569
rect 5451 15520 5452 15560
rect 5492 15520 5493 15560
rect 5451 15511 5493 15520
rect 5259 15476 5301 15485
rect 5259 15436 5260 15476
rect 5300 15436 5301 15476
rect 5259 15427 5301 15436
rect 5163 15392 5205 15401
rect 5163 15352 5164 15392
rect 5204 15352 5205 15392
rect 5163 15343 5205 15352
rect 5260 15342 5300 15427
rect 5163 15224 5205 15233
rect 5163 15184 5164 15224
rect 5204 15184 5205 15224
rect 5163 15175 5205 15184
rect 5164 14720 5204 15175
rect 5452 15065 5492 15511
rect 5451 15056 5493 15065
rect 5451 15016 5452 15056
rect 5492 15016 5493 15056
rect 5451 15007 5493 15016
rect 5355 14972 5397 14981
rect 5355 14932 5356 14972
rect 5396 14932 5397 14972
rect 5355 14923 5397 14932
rect 5259 14888 5301 14897
rect 5259 14848 5260 14888
rect 5300 14848 5301 14888
rect 5259 14839 5301 14848
rect 5164 14671 5204 14680
rect 5260 14720 5300 14839
rect 5260 14671 5300 14680
rect 5356 14720 5396 14923
rect 5356 14671 5396 14680
rect 5452 14720 5492 14729
rect 5548 14720 5588 16444
rect 5740 16064 5780 16073
rect 5644 16024 5740 16064
rect 5644 15737 5684 16024
rect 5740 16015 5780 16024
rect 5931 15896 5973 15905
rect 5931 15856 5932 15896
rect 5972 15856 5973 15896
rect 5931 15847 5973 15856
rect 6219 15896 6261 15905
rect 6219 15856 6220 15896
rect 6260 15856 6261 15896
rect 6219 15847 6261 15856
rect 5643 15728 5685 15737
rect 5643 15688 5644 15728
rect 5684 15688 5685 15728
rect 5643 15679 5685 15688
rect 5644 15560 5684 15569
rect 5644 15149 5684 15520
rect 5643 15140 5685 15149
rect 5643 15100 5644 15140
rect 5684 15100 5685 15140
rect 5643 15091 5685 15100
rect 5643 14972 5685 14981
rect 5643 14932 5644 14972
rect 5684 14932 5685 14972
rect 5643 14923 5685 14932
rect 5644 14838 5684 14923
rect 5492 14680 5588 14720
rect 5836 14720 5876 14729
rect 5068 14512 5204 14552
rect 5068 14057 5108 14142
rect 5067 14048 5109 14057
rect 5067 14008 5068 14048
rect 5108 14008 5109 14048
rect 5067 13999 5109 14008
rect 5164 14048 5204 14512
rect 5355 14384 5397 14393
rect 5355 14344 5356 14384
rect 5396 14344 5397 14384
rect 5355 14335 5397 14344
rect 5164 13999 5204 14008
rect 5356 14048 5396 14335
rect 5452 14057 5492 14680
rect 5547 14552 5589 14561
rect 5547 14512 5548 14552
rect 5588 14512 5589 14552
rect 5547 14503 5589 14512
rect 5356 13999 5396 14008
rect 5451 14048 5493 14057
rect 5451 14008 5452 14048
rect 5492 14008 5493 14048
rect 5451 13999 5493 14008
rect 5548 14048 5588 14503
rect 5644 14216 5684 14225
rect 5836 14216 5876 14680
rect 5684 14176 5876 14216
rect 5644 14167 5684 14176
rect 5548 13999 5588 14008
rect 5739 14048 5781 14057
rect 5739 14008 5740 14048
rect 5780 14008 5781 14048
rect 5739 13999 5781 14008
rect 5836 14048 5876 14057
rect 5932 14048 5972 15847
rect 6027 15812 6069 15821
rect 6027 15772 6028 15812
rect 6068 15772 6069 15812
rect 6027 15763 6069 15772
rect 5876 14008 5972 14048
rect 6028 14048 6068 15763
rect 6220 15485 6260 15847
rect 6316 15560 6356 16939
rect 6412 16409 6452 17032
rect 6508 17072 6548 17081
rect 6411 16400 6453 16409
rect 6411 16360 6412 16400
rect 6452 16360 6453 16400
rect 6411 16351 6453 16360
rect 6412 16232 6452 16241
rect 6412 15989 6452 16192
rect 6411 15980 6453 15989
rect 6411 15940 6412 15980
rect 6452 15940 6453 15980
rect 6411 15931 6453 15940
rect 6508 15905 6548 17032
rect 6603 16988 6645 16997
rect 6603 16948 6604 16988
rect 6644 16948 6645 16988
rect 6603 16939 6645 16948
rect 6604 16854 6644 16939
rect 6700 16904 6740 17452
rect 6988 17298 7028 17527
rect 6988 17249 7028 17258
rect 6987 17156 7029 17165
rect 6987 17116 6988 17156
rect 7028 17116 7029 17156
rect 6987 17107 7029 17116
rect 6988 16988 7028 17107
rect 7180 17072 7220 17083
rect 7084 17030 7124 17039
rect 7180 16997 7220 17032
rect 7084 16988 7124 16990
rect 6892 16948 7124 16988
rect 7179 16988 7221 16997
rect 7179 16948 7180 16988
rect 7220 16948 7221 16988
rect 6700 16855 6740 16864
rect 6795 16904 6837 16913
rect 6795 16864 6796 16904
rect 6836 16864 6837 16904
rect 6795 16855 6837 16864
rect 6796 16770 6836 16855
rect 6699 16736 6741 16745
rect 6699 16696 6700 16736
rect 6740 16696 6741 16736
rect 6699 16687 6741 16696
rect 6604 16232 6644 16241
rect 6507 15896 6549 15905
rect 6507 15856 6508 15896
rect 6548 15856 6549 15896
rect 6507 15847 6549 15856
rect 6604 15737 6644 16192
rect 6603 15728 6645 15737
rect 6603 15688 6604 15728
rect 6644 15688 6645 15728
rect 6603 15679 6645 15688
rect 6508 15560 6548 15569
rect 6316 15520 6508 15560
rect 6219 15476 6261 15485
rect 6219 15436 6220 15476
rect 6260 15436 6261 15476
rect 6219 15427 6261 15436
rect 6123 15224 6165 15233
rect 6123 15184 6124 15224
rect 6164 15184 6165 15224
rect 6123 15175 6165 15184
rect 5836 13999 5876 14008
rect 6028 13999 6068 14008
rect 6124 14048 6164 15175
rect 6220 14888 6260 15427
rect 6316 15317 6356 15402
rect 6315 15308 6357 15317
rect 6315 15268 6316 15308
rect 6356 15268 6357 15308
rect 6315 15259 6357 15268
rect 6411 14972 6453 14981
rect 6411 14932 6412 14972
rect 6452 14932 6453 14972
rect 6411 14923 6453 14932
rect 6220 14848 6356 14888
rect 6124 13999 6164 14008
rect 6220 14720 6260 14729
rect 5259 13964 5301 13973
rect 5259 13924 5260 13964
rect 5300 13924 5301 13964
rect 5259 13915 5301 13924
rect 5068 13880 5108 13889
rect 4972 13840 5068 13880
rect 3820 13746 3860 13831
rect 4876 13712 4916 13840
rect 5068 13831 5108 13840
rect 5260 13712 5300 13915
rect 5740 13914 5780 13999
rect 6123 13880 6165 13889
rect 6123 13840 6124 13880
rect 6164 13840 6165 13880
rect 6123 13831 6165 13840
rect 4876 13672 5300 13712
rect 3724 13588 3956 13628
rect 3627 13208 3669 13217
rect 3627 13168 3628 13208
rect 3668 13168 3669 13208
rect 3627 13159 3669 13168
rect 3820 13208 3860 13217
rect 3531 12620 3573 12629
rect 3531 12580 3532 12620
rect 3572 12580 3573 12620
rect 3531 12571 3573 12580
rect 3380 12496 3476 12536
rect 3340 12487 3380 12496
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3723 11948 3765 11957
rect 3723 11908 3724 11948
rect 3764 11908 3765 11948
rect 3723 11899 3765 11908
rect 3724 11696 3764 11899
rect 3820 11705 3860 13168
rect 3916 13208 3956 13588
rect 5355 13376 5397 13385
rect 5355 13336 5356 13376
rect 5396 13336 5397 13376
rect 5355 13327 5397 13336
rect 5356 13242 5396 13327
rect 5835 13292 5877 13301
rect 5835 13252 5836 13292
rect 5876 13252 5877 13292
rect 5835 13243 5877 13252
rect 3916 11957 3956 13168
rect 4012 13208 4052 13217
rect 4972 13208 5012 13217
rect 4012 12965 4052 13168
rect 4780 13168 4972 13208
rect 4300 13049 4340 13134
rect 4108 13040 4148 13049
rect 4299 13040 4341 13049
rect 4148 13000 4244 13040
rect 4108 12991 4148 13000
rect 4011 12956 4053 12965
rect 4011 12916 4012 12956
rect 4052 12916 4053 12956
rect 4011 12907 4053 12916
rect 4204 12704 4244 13000
rect 4299 13000 4300 13040
rect 4340 13000 4341 13040
rect 4299 12991 4341 13000
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4204 12664 4340 12704
rect 4204 12536 4244 12545
rect 4108 12496 4204 12536
rect 3915 11948 3957 11957
rect 3915 11908 3916 11948
rect 3956 11908 3957 11948
rect 3915 11899 3957 11908
rect 4012 11873 4052 11958
rect 4011 11864 4053 11873
rect 4011 11824 4012 11864
rect 4052 11824 4053 11864
rect 4011 11815 4053 11824
rect 3724 11647 3764 11656
rect 3819 11696 3861 11705
rect 3819 11656 3820 11696
rect 3860 11656 3861 11696
rect 3819 11647 3861 11656
rect 4012 11696 4052 11705
rect 3820 11562 3860 11647
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 652 11192 692 11201
rect 652 10697 692 11152
rect 3627 11192 3669 11201
rect 3627 11152 3628 11192
rect 3668 11152 3669 11192
rect 3627 11143 3669 11152
rect 3724 11192 3764 11201
rect 2572 11033 2612 11118
rect 2571 11024 2613 11033
rect 2571 10984 2572 11024
rect 2612 10984 2613 11024
rect 2571 10975 2613 10984
rect 2668 11024 2708 11033
rect 1515 10856 1557 10865
rect 1996 10856 2036 10865
rect 1515 10816 1516 10856
rect 1556 10816 1557 10856
rect 1515 10807 1557 10816
rect 1900 10816 1996 10856
rect 651 10688 693 10697
rect 651 10648 652 10688
rect 692 10648 693 10688
rect 651 10639 693 10648
rect 1516 10184 1556 10807
rect 1516 10135 1556 10144
rect 1900 10184 1940 10816
rect 1996 10807 2036 10816
rect 2571 10856 2613 10865
rect 2571 10816 2572 10856
rect 2612 10816 2613 10856
rect 2571 10807 2613 10816
rect 2572 10722 2612 10807
rect 2571 10184 2613 10193
rect 1900 10135 1940 10144
rect 2476 10144 2572 10184
rect 2612 10144 2613 10184
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9689
rect 652 9017 692 9640
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1708 9512 1748 9521
rect 1516 9344 1556 9353
rect 1035 9260 1077 9269
rect 1035 9220 1036 9260
rect 1076 9220 1077 9260
rect 1035 9211 1077 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 1036 8672 1076 9211
rect 1323 8924 1365 8933
rect 1323 8884 1324 8924
rect 1364 8884 1365 8924
rect 1323 8875 1365 8884
rect 1036 8623 1076 8632
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 1035 8168 1077 8177
rect 1035 8128 1036 8168
rect 1076 8128 1077 8168
rect 1035 8119 1077 8128
rect 844 8000 884 8011
rect 844 7925 884 7960
rect 1036 8000 1076 8119
rect 1036 7951 1076 7960
rect 1132 8000 1172 8009
rect 1324 8000 1364 8875
rect 1420 8672 1460 8681
rect 1516 8672 1556 9304
rect 1460 8632 1556 8672
rect 1420 8623 1460 8632
rect 1516 8168 1556 8177
rect 1612 8168 1652 9463
rect 1708 9353 1748 9472
rect 1900 9512 1940 9521
rect 1900 9428 1940 9472
rect 2284 9512 2324 9521
rect 2092 9428 2132 9437
rect 1900 9388 2092 9428
rect 2092 9379 2132 9388
rect 1707 9344 1749 9353
rect 1707 9304 1708 9344
rect 1748 9304 1749 9344
rect 1707 9295 1749 9304
rect 1556 8128 1652 8168
rect 1516 8119 1556 8128
rect 1419 8084 1461 8093
rect 1419 8044 1420 8084
rect 1460 8044 1461 8084
rect 1419 8035 1461 8044
rect 1172 7960 1268 8000
rect 1132 7951 1172 7960
rect 843 7916 885 7925
rect 843 7876 844 7916
rect 884 7876 885 7916
rect 843 7867 885 7876
rect 1131 7832 1173 7841
rect 1131 7792 1132 7832
rect 1172 7792 1173 7832
rect 1131 7783 1173 7792
rect 843 7748 885 7757
rect 843 7708 844 7748
rect 884 7708 885 7748
rect 843 7699 885 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 652 6656 692 7279
rect 844 7160 884 7699
rect 1132 7698 1172 7783
rect 1228 7337 1268 7960
rect 1324 7951 1364 7960
rect 1420 8000 1460 8035
rect 1420 7949 1460 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 1612 7866 1652 7951
rect 1708 7925 1748 9295
rect 1899 9260 1941 9269
rect 1899 9220 1900 9260
rect 1940 9220 1941 9260
rect 1899 9211 1941 9220
rect 1900 9126 1940 9211
rect 2284 8933 2324 9472
rect 2380 9512 2420 9521
rect 2283 8924 2325 8933
rect 2283 8884 2284 8924
rect 2324 8884 2325 8924
rect 2283 8875 2325 8884
rect 2380 8849 2420 9472
rect 2379 8840 2421 8849
rect 2379 8800 2380 8840
rect 2420 8800 2421 8840
rect 2379 8791 2421 8800
rect 2284 8672 2324 8681
rect 2476 8672 2516 10144
rect 2571 10135 2613 10144
rect 2572 10116 2612 10135
rect 2668 8849 2708 10984
rect 2860 11024 2900 11033
rect 2763 10184 2805 10193
rect 2763 10144 2764 10184
rect 2804 10144 2805 10184
rect 2763 10135 2805 10144
rect 2764 10050 2804 10135
rect 2860 9437 2900 10984
rect 3435 11024 3477 11033
rect 3435 10984 3436 11024
rect 3476 10984 3477 11024
rect 3435 10975 3477 10984
rect 3628 11024 3668 11143
rect 3436 10772 3476 10975
rect 3476 10732 3572 10772
rect 3436 10723 3476 10732
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3532 10025 3572 10732
rect 3531 10016 3573 10025
rect 3531 9976 3532 10016
rect 3572 9976 3573 10016
rect 3531 9967 3573 9976
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 2859 9428 2901 9437
rect 2859 9388 2860 9428
rect 2900 9388 2901 9428
rect 2859 9379 2901 9388
rect 3532 9378 3572 9463
rect 2860 9260 2900 9269
rect 2667 8840 2709 8849
rect 2667 8800 2668 8840
rect 2708 8800 2709 8840
rect 2667 8791 2709 8800
rect 2324 8632 2516 8672
rect 1707 7916 1749 7925
rect 1707 7876 1708 7916
rect 1748 7876 1749 7916
rect 1707 7867 1749 7876
rect 1995 7916 2037 7925
rect 1995 7876 1996 7916
rect 2036 7876 2037 7916
rect 1995 7867 2037 7876
rect 1803 7748 1845 7757
rect 1803 7708 1804 7748
rect 1844 7708 1845 7748
rect 1803 7699 1845 7708
rect 1804 7614 1844 7699
rect 1227 7328 1269 7337
rect 1227 7288 1228 7328
rect 1268 7288 1269 7328
rect 1227 7279 1269 7288
rect 844 7111 884 7120
rect 1228 7160 1268 7169
rect 1268 7120 1364 7160
rect 1228 7111 1268 7120
rect 652 6607 692 6616
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 652 5480 692 6439
rect 1324 6320 1364 7120
rect 1996 6488 2036 7867
rect 2092 7160 2132 7169
rect 2284 7160 2324 8632
rect 2860 8177 2900 9220
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3628 8924 3668 10984
rect 3724 10445 3764 11152
rect 4012 11117 4052 11656
rect 4011 11108 4053 11117
rect 4011 11068 4012 11108
rect 4052 11068 4053 11108
rect 4011 11059 4053 11068
rect 4108 11024 4148 12496
rect 4204 12487 4244 12496
rect 4204 11696 4244 11705
rect 4300 11696 4340 12664
rect 4491 11948 4533 11957
rect 4491 11908 4492 11948
rect 4532 11908 4533 11948
rect 4491 11899 4533 11908
rect 4396 11705 4436 11790
rect 4244 11656 4340 11696
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4204 11647 4244 11656
rect 4395 11647 4437 11656
rect 4492 11696 4532 11899
rect 4683 11864 4725 11873
rect 4683 11824 4684 11864
rect 4724 11824 4725 11864
rect 4683 11815 4725 11824
rect 4492 11647 4532 11656
rect 4684 11696 4724 11815
rect 4684 11647 4724 11656
rect 4300 11528 4340 11537
rect 4780 11528 4820 13168
rect 4972 13159 5012 13168
rect 5547 13208 5589 13217
rect 5547 13168 5548 13208
rect 5588 13168 5589 13208
rect 5547 13159 5589 13168
rect 5644 13208 5684 13217
rect 5548 13074 5588 13159
rect 5644 12965 5684 13168
rect 5740 13208 5780 13217
rect 5740 13040 5780 13168
rect 5836 13208 5876 13243
rect 5836 13157 5876 13168
rect 6028 13040 6068 13049
rect 5740 13000 6028 13040
rect 5643 12956 5685 12965
rect 5643 12916 5644 12956
rect 5684 12916 5685 12956
rect 5643 12907 5685 12916
rect 5643 12620 5685 12629
rect 5643 12580 5644 12620
rect 5684 12580 5685 12620
rect 5643 12571 5685 12580
rect 5452 12536 5492 12545
rect 5644 12536 5684 12571
rect 5492 12496 5588 12536
rect 5452 12487 5492 12496
rect 5548 11696 5588 12496
rect 5644 12485 5684 12496
rect 5740 11705 5780 13000
rect 6028 12991 6068 13000
rect 6028 12536 6068 12545
rect 6124 12536 6164 13831
rect 6220 13385 6260 14680
rect 6316 14216 6356 14848
rect 6316 14167 6356 14176
rect 6316 14048 6356 14057
rect 6412 14048 6452 14923
rect 6356 14008 6452 14048
rect 6316 13999 6356 14008
rect 6508 13973 6548 15520
rect 6604 15560 6644 15571
rect 6604 15485 6644 15520
rect 6700 15560 6740 16687
rect 6795 15896 6837 15905
rect 6795 15856 6796 15896
rect 6836 15856 6837 15896
rect 6795 15847 6837 15856
rect 6700 15511 6740 15520
rect 6796 15560 6836 15847
rect 6796 15511 6836 15520
rect 6603 15476 6645 15485
rect 6603 15436 6604 15476
rect 6644 15436 6645 15476
rect 6603 15427 6645 15436
rect 6699 15392 6741 15401
rect 6699 15352 6700 15392
rect 6740 15352 6741 15392
rect 6699 15343 6741 15352
rect 6603 14384 6645 14393
rect 6603 14344 6604 14384
rect 6644 14344 6645 14384
rect 6603 14335 6645 14344
rect 6604 14216 6644 14335
rect 6604 14167 6644 14176
rect 6700 14048 6740 15343
rect 6700 13999 6740 14008
rect 6507 13964 6549 13973
rect 6507 13924 6508 13964
rect 6548 13924 6549 13964
rect 6507 13915 6549 13924
rect 6219 13376 6261 13385
rect 6219 13336 6220 13376
rect 6260 13336 6261 13376
rect 6219 13327 6261 13336
rect 6892 13301 6932 16948
rect 7179 16939 7221 16948
rect 7276 16820 7316 17536
rect 7371 17072 7413 17081
rect 7371 17032 7372 17072
rect 7412 17032 7413 17072
rect 7371 17023 7413 17032
rect 7180 16780 7316 16820
rect 7180 15980 7220 16780
rect 7275 16232 7317 16241
rect 7275 16192 7276 16232
rect 7316 16192 7317 16232
rect 7275 16183 7317 16192
rect 7276 16098 7316 16183
rect 7180 15940 7316 15980
rect 7083 15728 7125 15737
rect 7083 15688 7084 15728
rect 7124 15688 7125 15728
rect 7083 15679 7125 15688
rect 7084 15594 7124 15679
rect 7179 15644 7221 15653
rect 7179 15604 7180 15644
rect 7220 15604 7221 15644
rect 7179 15595 7221 15604
rect 6987 15560 7029 15569
rect 6987 15520 6988 15560
rect 7028 15520 7029 15560
rect 6987 15511 7029 15520
rect 7180 15560 7220 15595
rect 6988 15426 7028 15511
rect 7180 15149 7220 15520
rect 7276 15560 7316 15940
rect 7276 15511 7316 15520
rect 7179 15140 7221 15149
rect 7179 15100 7180 15140
rect 7220 15100 7221 15140
rect 7179 15091 7221 15100
rect 7083 14720 7125 14729
rect 7083 14680 7084 14720
rect 7124 14680 7125 14720
rect 7083 14671 7125 14680
rect 7084 14586 7124 14671
rect 7372 13880 7412 17023
rect 7467 16904 7509 16913
rect 7467 16864 7468 16904
rect 7508 16864 7509 16904
rect 7467 16855 7509 16864
rect 7468 16770 7508 16855
rect 7564 16745 7604 18544
rect 7852 18535 7892 18544
rect 7948 18416 7988 18712
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 8044 18450 8084 18535
rect 7756 18376 7988 18416
rect 8140 18416 8180 19048
rect 8236 18584 8276 19804
rect 8428 19795 8468 19804
rect 8523 19424 8565 19433
rect 8523 19384 8524 19424
rect 8564 19384 8565 19424
rect 8523 19375 8565 19384
rect 8524 19290 8564 19375
rect 8620 18929 8660 20056
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 8715 20047 8757 20056
rect 9196 20096 9236 20105
rect 8716 19340 8756 20047
rect 9099 19424 9141 19433
rect 9099 19384 9100 19424
rect 9140 19384 9141 19424
rect 9196 19424 9236 20056
rect 9676 20021 9716 21568
rect 9771 21608 9813 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 9868 21608 9908 21617
rect 10060 21608 10100 22576
rect 9908 21568 10100 21608
rect 10156 21608 10196 23071
rect 10732 22961 10772 23080
rect 11211 23120 11253 23129
rect 11596 23120 11636 23129
rect 11211 23080 11212 23120
rect 11252 23080 11253 23120
rect 11211 23071 11253 23080
rect 11500 23080 11596 23120
rect 10731 22952 10773 22961
rect 10731 22912 10732 22952
rect 10772 22912 10773 22952
rect 10731 22903 10773 22912
rect 10924 22868 10964 22877
rect 10924 22373 10964 22828
rect 10923 22364 10965 22373
rect 10923 22324 10924 22364
rect 10964 22324 10965 22364
rect 10923 22315 10965 22324
rect 10828 22280 10868 22289
rect 9772 21474 9812 21559
rect 9868 20861 9908 21568
rect 10156 21559 10196 21568
rect 10252 22240 10828 22280
rect 9867 20852 9909 20861
rect 9867 20812 9868 20852
rect 9908 20812 9909 20852
rect 9867 20803 9909 20812
rect 9964 20768 10004 20779
rect 9964 20693 10004 20728
rect 9963 20684 10005 20693
rect 9963 20644 9964 20684
rect 10004 20644 10005 20684
rect 9963 20635 10005 20644
rect 10252 20180 10292 22240
rect 10828 22231 10868 22240
rect 11211 21692 11253 21701
rect 11211 21652 11212 21692
rect 11252 21652 11253 21692
rect 11211 21643 11253 21652
rect 10347 21356 10389 21365
rect 10347 21316 10348 21356
rect 10388 21316 10389 21356
rect 10347 21307 10389 21316
rect 10444 21356 10484 21365
rect 10348 20768 10388 21307
rect 10444 20861 10484 21316
rect 10636 20936 10676 20945
rect 10676 20896 10868 20936
rect 10636 20887 10676 20896
rect 10443 20852 10485 20861
rect 10443 20812 10444 20852
rect 10484 20812 10485 20852
rect 10443 20803 10485 20812
rect 10348 20719 10388 20728
rect 10444 20768 10484 20803
rect 10444 20525 10484 20728
rect 10635 20768 10677 20777
rect 10635 20728 10636 20768
rect 10676 20728 10677 20768
rect 10635 20719 10677 20728
rect 10828 20768 10868 20896
rect 10828 20719 10868 20728
rect 10636 20634 10676 20719
rect 10443 20516 10485 20525
rect 10443 20476 10444 20516
rect 10484 20476 10485 20516
rect 10443 20467 10485 20476
rect 10156 20140 10292 20180
rect 10060 20096 10100 20105
rect 9675 20012 9717 20021
rect 9675 19972 9676 20012
rect 9716 19972 9717 20012
rect 9675 19963 9717 19972
rect 9292 19424 9332 19433
rect 9196 19384 9292 19424
rect 9099 19375 9141 19384
rect 9292 19375 9332 19384
rect 8619 18920 8661 18929
rect 8619 18880 8620 18920
rect 8660 18880 8661 18920
rect 8619 18871 8661 18880
rect 8716 18761 8756 19300
rect 8715 18752 8757 18761
rect 8715 18712 8716 18752
rect 8756 18712 8757 18752
rect 8715 18703 8757 18712
rect 8236 18535 8276 18544
rect 8332 18584 8372 18593
rect 8332 18416 8372 18544
rect 8140 18376 8372 18416
rect 7756 18005 7796 18376
rect 8044 18332 8084 18341
rect 7852 18292 8044 18332
rect 7755 17996 7797 18005
rect 7755 17956 7756 17996
rect 7796 17956 7797 17996
rect 7755 17947 7797 17956
rect 7659 16820 7701 16829
rect 7659 16780 7660 16820
rect 7700 16780 7701 16820
rect 7659 16771 7701 16780
rect 7563 16736 7605 16745
rect 7563 16696 7564 16736
rect 7604 16696 7605 16736
rect 7563 16687 7605 16696
rect 7660 16686 7700 16771
rect 7468 16064 7508 16073
rect 7468 15905 7508 16024
rect 7563 16064 7605 16073
rect 7563 16024 7564 16064
rect 7604 16024 7605 16064
rect 7563 16015 7605 16024
rect 7467 15896 7509 15905
rect 7467 15856 7468 15896
rect 7508 15856 7509 15896
rect 7467 15847 7509 15856
rect 7564 15653 7604 16015
rect 7659 15728 7701 15737
rect 7659 15688 7660 15728
rect 7700 15688 7701 15728
rect 7659 15679 7701 15688
rect 7563 15644 7605 15653
rect 7563 15604 7564 15644
rect 7604 15604 7605 15644
rect 7563 15595 7605 15604
rect 7467 15560 7509 15569
rect 7467 15520 7468 15560
rect 7508 15520 7509 15560
rect 7467 15511 7509 15520
rect 7564 15560 7604 15595
rect 7660 15594 7700 15679
rect 7468 15426 7508 15511
rect 7564 15510 7604 15520
rect 7756 15560 7796 17947
rect 7852 17744 7892 18292
rect 8044 18283 8084 18292
rect 7852 17695 7892 17704
rect 8332 17585 8372 18376
rect 8812 18584 8852 18593
rect 8524 17660 8564 17669
rect 8716 17660 8756 17669
rect 8564 17620 8716 17660
rect 8524 17611 8564 17620
rect 8716 17611 8756 17620
rect 8331 17576 8373 17585
rect 8331 17536 8332 17576
rect 8372 17536 8373 17576
rect 8331 17527 8373 17536
rect 8812 17081 8852 18544
rect 9100 17744 9140 19375
rect 9964 19088 10004 19097
rect 9868 19048 9964 19088
rect 9291 18752 9333 18761
rect 9291 18712 9292 18752
rect 9332 18712 9333 18752
rect 9291 18703 9333 18712
rect 9292 18618 9332 18703
rect 9771 18416 9813 18425
rect 9771 18376 9772 18416
rect 9812 18376 9813 18416
rect 9771 18367 9813 18376
rect 9100 17695 9140 17704
rect 9292 18332 9332 18341
rect 8332 17072 8372 17081
rect 7947 16820 7989 16829
rect 7947 16780 7948 16820
rect 7988 16780 7989 16820
rect 7947 16771 7989 16780
rect 7948 15644 7988 16771
rect 8332 16484 8372 17032
rect 8524 17072 8564 17081
rect 8524 16913 8564 17032
rect 8811 17072 8853 17081
rect 8811 17032 8812 17072
rect 8852 17032 8853 17072
rect 8811 17023 8853 17032
rect 9195 17072 9237 17081
rect 9195 17032 9196 17072
rect 9236 17032 9237 17072
rect 9195 17023 9237 17032
rect 9196 16938 9236 17023
rect 8523 16904 8565 16913
rect 8523 16864 8524 16904
rect 8564 16864 8565 16904
rect 8523 16855 8565 16864
rect 8332 16435 8372 16444
rect 7948 15595 7988 15604
rect 8140 16232 8180 16241
rect 7756 14393 7796 15520
rect 8140 14888 8180 16192
rect 8331 16232 8373 16241
rect 8331 16192 8332 16232
rect 8372 16192 8373 16232
rect 8331 16183 8373 16192
rect 8620 16232 8660 16241
rect 8332 16098 8372 16183
rect 8620 15737 8660 16192
rect 8907 16064 8949 16073
rect 8907 16024 8908 16064
rect 8948 16024 8949 16064
rect 8907 16015 8949 16024
rect 8908 15930 8948 16015
rect 9099 15896 9141 15905
rect 9099 15856 9100 15896
rect 9140 15856 9141 15896
rect 9099 15847 9141 15856
rect 8619 15728 8661 15737
rect 8619 15688 8620 15728
rect 8660 15688 8661 15728
rect 8619 15679 8661 15688
rect 8332 15560 8372 15569
rect 8372 15520 8564 15560
rect 8332 15511 8372 15520
rect 8235 14888 8277 14897
rect 8140 14848 8236 14888
rect 8276 14848 8277 14888
rect 8235 14839 8277 14848
rect 8524 14888 8564 15520
rect 8524 14839 8564 14848
rect 8236 14754 8276 14839
rect 8908 14720 8948 14729
rect 7755 14384 7797 14393
rect 7755 14344 7756 14384
rect 7796 14344 7797 14384
rect 7755 14335 7797 14344
rect 8908 14309 8948 14680
rect 9100 14720 9140 15847
rect 9196 15560 9236 15569
rect 9292 15560 9332 18292
rect 9387 17072 9429 17081
rect 9387 17032 9388 17072
rect 9428 17032 9429 17072
rect 9387 17023 9429 17032
rect 9772 17072 9812 18367
rect 9868 17165 9908 19048
rect 9964 19039 10004 19048
rect 9963 18920 10005 18929
rect 9963 18880 9964 18920
rect 10004 18880 10005 18920
rect 9963 18871 10005 18880
rect 9964 18752 10004 18871
rect 10060 18761 10100 20056
rect 9964 18703 10004 18712
rect 10059 18752 10101 18761
rect 10059 18712 10060 18752
rect 10100 18712 10101 18752
rect 10059 18703 10101 18712
rect 10060 17753 10100 18703
rect 9964 17744 10004 17753
rect 10059 17744 10101 17753
rect 10004 17704 10060 17744
rect 10100 17704 10101 17744
rect 9964 17695 10004 17704
rect 10059 17695 10101 17704
rect 10060 17610 10100 17695
rect 9867 17156 9909 17165
rect 9867 17116 9868 17156
rect 9908 17116 9909 17156
rect 9867 17107 9909 17116
rect 9772 17023 9812 17032
rect 9388 16938 9428 17023
rect 9580 16232 9620 16241
rect 9580 15737 9620 16192
rect 9579 15728 9621 15737
rect 9579 15688 9580 15728
rect 9620 15688 9621 15728
rect 9579 15679 9621 15688
rect 9236 15520 9332 15560
rect 9196 15511 9236 15520
rect 10156 15140 10196 20140
rect 10251 20012 10293 20021
rect 10251 19972 10252 20012
rect 10292 19972 10293 20012
rect 10251 19963 10293 19972
rect 11212 20012 11252 21643
rect 11308 21608 11348 21617
rect 11308 20777 11348 21568
rect 11403 21608 11445 21617
rect 11403 21568 11404 21608
rect 11444 21568 11445 21608
rect 11403 21559 11445 21568
rect 11500 21608 11540 23080
rect 11596 23071 11636 23080
rect 11404 21474 11444 21559
rect 11500 21533 11540 21568
rect 11596 21608 11636 21617
rect 11692 21608 11732 23659
rect 11884 23120 11924 23743
rect 11979 23708 12021 23717
rect 11979 23668 11980 23708
rect 12020 23668 12021 23708
rect 11979 23659 12021 23668
rect 11980 23574 12020 23659
rect 11884 22709 11924 23080
rect 12555 22868 12597 22877
rect 12555 22828 12556 22868
rect 12596 22828 12597 22868
rect 12555 22819 12597 22828
rect 12556 22734 12596 22819
rect 11883 22700 11925 22709
rect 11883 22660 11884 22700
rect 11924 22660 11925 22700
rect 11883 22651 11925 22660
rect 12459 22700 12501 22709
rect 12459 22660 12460 22700
rect 12500 22660 12501 22700
rect 12459 22651 12501 22660
rect 11884 22532 11924 22651
rect 12267 22616 12309 22625
rect 12267 22576 12268 22616
rect 12308 22576 12309 22616
rect 12267 22567 12309 22576
rect 11980 22532 12020 22541
rect 11884 22492 11980 22532
rect 11980 22483 12020 22492
rect 11787 22280 11829 22289
rect 11787 22240 11788 22280
rect 11828 22240 11829 22280
rect 11787 22231 11829 22240
rect 12268 22280 12308 22567
rect 12460 22448 12500 22651
rect 12652 22625 12692 24499
rect 12748 23960 12788 25096
rect 12843 24884 12885 24893
rect 12843 24844 12844 24884
rect 12884 24844 12885 24884
rect 12843 24835 12885 24844
rect 12844 24632 12884 24835
rect 12844 24583 12884 24592
rect 12748 23920 12884 23960
rect 12748 23792 12788 23803
rect 12844 23801 12884 23920
rect 12748 23717 12788 23752
rect 12843 23792 12885 23801
rect 12843 23752 12844 23792
rect 12884 23752 12885 23792
rect 12843 23743 12885 23752
rect 12747 23708 12789 23717
rect 12747 23668 12748 23708
rect 12788 23668 12789 23708
rect 12747 23659 12789 23668
rect 12844 23204 12884 23213
rect 12940 23204 12980 25591
rect 13036 25061 13076 26095
rect 13132 25136 13172 26515
rect 13228 26153 13268 26776
rect 13420 26816 13460 26825
rect 13420 26489 13460 26776
rect 13516 26816 13556 26944
rect 13516 26767 13556 26776
rect 13419 26480 13461 26489
rect 13419 26440 13420 26480
rect 13460 26440 13461 26480
rect 13419 26431 13461 26440
rect 13612 26312 13652 28456
rect 13708 26816 13748 28960
rect 13995 27404 14037 27413
rect 13995 27364 13996 27404
rect 14036 27364 14037 27404
rect 13995 27355 14037 27364
rect 13803 27068 13845 27077
rect 13996 27068 14036 27355
rect 13803 27028 13804 27068
rect 13844 27028 13845 27068
rect 13803 27019 13845 27028
rect 13961 27028 14036 27068
rect 13708 26767 13748 26776
rect 13804 26816 13844 27019
rect 13961 26831 14001 27028
rect 13961 26782 14001 26791
rect 13804 26767 13844 26776
rect 13803 26648 13845 26657
rect 13803 26608 13804 26648
rect 13844 26608 13845 26648
rect 13803 26599 13845 26608
rect 13995 26648 14037 26657
rect 13995 26608 13996 26648
rect 14036 26608 14037 26648
rect 13995 26599 14037 26608
rect 13804 26514 13844 26599
rect 13899 26564 13941 26573
rect 13899 26524 13900 26564
rect 13940 26524 13941 26564
rect 13899 26515 13941 26524
rect 13900 26396 13940 26515
rect 13996 26489 14036 26599
rect 13995 26480 14037 26489
rect 13995 26440 13996 26480
rect 14036 26440 14037 26480
rect 13995 26431 14037 26440
rect 13516 26272 13652 26312
rect 13804 26356 13940 26396
rect 13227 26144 13269 26153
rect 13227 26104 13228 26144
rect 13268 26104 13269 26144
rect 13227 26095 13269 26104
rect 13222 25472 13264 25481
rect 13222 25432 13223 25472
rect 13263 25432 13264 25472
rect 13222 25423 13264 25432
rect 13223 25304 13263 25423
rect 13223 25255 13263 25264
rect 13324 25304 13364 25313
rect 13324 25136 13364 25264
rect 13132 25096 13364 25136
rect 13420 25304 13460 25313
rect 13035 25052 13077 25061
rect 13035 25012 13036 25052
rect 13076 25012 13077 25052
rect 13035 25003 13077 25012
rect 13420 24977 13460 25264
rect 13419 24968 13461 24977
rect 13419 24928 13420 24968
rect 13460 24928 13461 24968
rect 13419 24919 13461 24928
rect 13227 24716 13269 24725
rect 13227 24676 13228 24716
rect 13268 24676 13269 24716
rect 13227 24667 13269 24676
rect 13228 24582 13268 24667
rect 13516 24632 13556 26272
rect 13611 26144 13653 26153
rect 13804 26144 13844 26356
rect 13611 26104 13612 26144
rect 13652 26104 13748 26144
rect 13611 26095 13653 26104
rect 13612 26010 13652 26095
rect 13708 25901 13748 26104
rect 13804 26095 13844 26104
rect 13899 26144 13941 26153
rect 13899 26104 13900 26144
rect 13940 26104 13941 26144
rect 13899 26095 13941 26104
rect 13900 26010 13940 26095
rect 13996 25985 14036 26431
rect 14092 26321 14132 30976
rect 14572 30773 14612 31144
rect 14571 30764 14613 30773
rect 14571 30724 14572 30764
rect 14612 30724 14613 30764
rect 14571 30715 14613 30724
rect 14187 30680 14229 30689
rect 14187 30640 14188 30680
rect 14228 30640 14229 30680
rect 14187 30631 14229 30640
rect 14188 28841 14228 30631
rect 15051 30512 15093 30521
rect 15051 30472 15052 30512
rect 15092 30472 15093 30512
rect 15051 30463 15093 30472
rect 14667 30428 14709 30437
rect 14667 30388 14668 30428
rect 14708 30388 14709 30428
rect 14667 30379 14709 30388
rect 14668 30294 14708 30379
rect 15052 30378 15092 30463
rect 15244 29849 15284 32824
rect 15340 31940 15380 31949
rect 15340 31529 15380 31900
rect 15436 31781 15476 32992
rect 15435 31772 15477 31781
rect 15435 31732 15436 31772
rect 15476 31732 15477 31772
rect 15435 31723 15477 31732
rect 15339 31520 15381 31529
rect 15339 31480 15340 31520
rect 15380 31480 15381 31520
rect 15339 31471 15381 31480
rect 15340 31352 15380 31363
rect 15340 31277 15380 31312
rect 15436 31352 15476 31361
rect 15339 31268 15381 31277
rect 15339 31228 15340 31268
rect 15380 31228 15381 31268
rect 15339 31219 15381 31228
rect 15436 30857 15476 31312
rect 15532 31352 15572 33067
rect 15628 31613 15668 33664
rect 15819 33704 15861 33713
rect 15819 33664 15820 33704
rect 15860 33664 15861 33704
rect 15819 33655 15861 33664
rect 16108 32789 16148 33748
rect 16252 33662 16292 33671
rect 16252 33620 16292 33622
rect 16204 33580 16292 33620
rect 16107 32780 16149 32789
rect 16107 32740 16108 32780
rect 16148 32740 16149 32780
rect 16107 32731 16149 32740
rect 16204 32285 16244 33580
rect 16492 33125 16532 34999
rect 16588 34796 16628 35167
rect 16684 34973 16724 35176
rect 16780 35216 16820 36688
rect 16875 36728 16917 36737
rect 16875 36688 16876 36728
rect 16916 36688 16917 36728
rect 16875 36679 16917 36688
rect 16972 36728 17012 36737
rect 17548 36728 17588 36763
rect 17012 36688 17300 36728
rect 16972 36679 17012 36688
rect 16876 36594 16916 36679
rect 17163 36560 17205 36569
rect 17163 36520 17164 36560
rect 17204 36520 17205 36560
rect 17163 36511 17205 36520
rect 17164 36426 17204 36511
rect 16876 35888 16916 35897
rect 17163 35888 17205 35897
rect 16916 35848 17012 35888
rect 16876 35839 16916 35848
rect 16875 35300 16917 35309
rect 16875 35260 16876 35300
rect 16916 35260 16917 35300
rect 16875 35251 16917 35260
rect 16780 35057 16820 35176
rect 16876 35166 16916 35251
rect 16972 35225 17012 35848
rect 17163 35848 17164 35888
rect 17204 35848 17205 35888
rect 17163 35839 17205 35848
rect 17067 35300 17109 35309
rect 17067 35260 17068 35300
rect 17108 35260 17109 35300
rect 17067 35251 17109 35260
rect 17164 35300 17204 35839
rect 17164 35251 17204 35260
rect 16971 35216 17013 35225
rect 16971 35176 16972 35216
rect 17012 35176 17013 35216
rect 16971 35167 17013 35176
rect 17068 35216 17108 35251
rect 17068 35165 17108 35176
rect 17260 35216 17300 36688
rect 17548 36677 17588 36688
rect 18123 36728 18165 36737
rect 18123 36688 18124 36728
rect 18164 36688 18165 36728
rect 18123 36679 18165 36688
rect 17644 36476 17684 36485
rect 17260 35141 17300 35176
rect 17356 36436 17644 36476
rect 17356 35216 17396 36436
rect 17644 36427 17684 36436
rect 18028 35720 18068 35729
rect 18028 35309 18068 35680
rect 17547 35300 17589 35309
rect 17547 35260 17548 35300
rect 17588 35260 17589 35300
rect 17547 35251 17589 35260
rect 18027 35300 18069 35309
rect 18027 35260 18028 35300
rect 18068 35260 18069 35300
rect 18027 35251 18069 35260
rect 18124 35300 18164 36679
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 18795 36056 18837 36065
rect 18795 36016 18796 36056
rect 18836 36016 18837 36056
rect 18795 36007 18837 36016
rect 19179 36056 19221 36065
rect 19179 36016 19180 36056
rect 19220 36016 19221 36056
rect 19179 36007 19221 36016
rect 18315 35888 18357 35897
rect 18315 35848 18316 35888
rect 18356 35848 18357 35888
rect 18315 35839 18357 35848
rect 18316 35754 18356 35839
rect 18220 35300 18260 35309
rect 18124 35260 18220 35300
rect 17356 35167 17396 35176
rect 17548 35216 17588 35251
rect 17259 35132 17301 35141
rect 17259 35092 17260 35132
rect 17300 35092 17301 35132
rect 17259 35083 17301 35092
rect 16779 35048 16821 35057
rect 16779 35008 16780 35048
rect 16820 35008 16821 35048
rect 16779 34999 16821 35008
rect 16683 34964 16725 34973
rect 16683 34924 16684 34964
rect 16724 34924 16725 34964
rect 16683 34915 16725 34924
rect 16588 34756 16916 34796
rect 16780 33704 16820 33713
rect 16588 33664 16780 33704
rect 16491 33116 16533 33125
rect 16491 33076 16492 33116
rect 16532 33076 16533 33116
rect 16491 33067 16533 33076
rect 16396 32948 16436 32957
rect 16588 32948 16628 33664
rect 16780 33655 16820 33664
rect 16683 33116 16725 33125
rect 16683 33076 16684 33116
rect 16724 33076 16725 33116
rect 16683 33067 16725 33076
rect 16436 32908 16628 32948
rect 16396 32780 16436 32908
rect 16684 32864 16724 33067
rect 16684 32815 16724 32824
rect 16779 32864 16821 32873
rect 16779 32824 16780 32864
rect 16820 32824 16821 32864
rect 16779 32815 16821 32824
rect 16876 32864 16916 34756
rect 16971 34208 17013 34217
rect 17164 34208 17204 34217
rect 16971 34168 16972 34208
rect 17012 34168 17013 34208
rect 16971 34159 17013 34168
rect 17068 34168 17164 34208
rect 16972 34074 17012 34159
rect 16300 32740 16436 32780
rect 16203 32276 16245 32285
rect 16203 32236 16204 32276
rect 16244 32236 16245 32276
rect 16203 32227 16245 32236
rect 16011 32192 16053 32201
rect 16011 32152 16012 32192
rect 16052 32152 16053 32192
rect 16011 32143 16053 32152
rect 16012 32058 16052 32143
rect 16107 31940 16149 31949
rect 16107 31900 16108 31940
rect 16148 31900 16149 31940
rect 16107 31891 16149 31900
rect 15627 31604 15669 31613
rect 15627 31564 15628 31604
rect 15668 31564 15669 31604
rect 15627 31555 15669 31564
rect 16011 31436 16053 31445
rect 16011 31396 16012 31436
rect 16052 31396 16053 31436
rect 16011 31387 16053 31396
rect 15532 30941 15572 31312
rect 15628 31352 15668 31361
rect 15820 31352 15860 31361
rect 15668 31312 15820 31352
rect 15628 31303 15668 31312
rect 15820 31303 15860 31312
rect 16012 31352 16052 31387
rect 16012 31301 16052 31312
rect 16108 31352 16148 31891
rect 16108 31303 16148 31312
rect 15915 31268 15957 31277
rect 15915 31228 15916 31268
rect 15956 31228 15957 31268
rect 15915 31219 15957 31228
rect 15916 31134 15956 31219
rect 16204 31100 16244 32227
rect 16300 32201 16340 32740
rect 16588 32705 16628 32790
rect 16780 32730 16820 32815
rect 16876 32705 16916 32824
rect 16587 32696 16629 32705
rect 16587 32656 16588 32696
rect 16628 32656 16629 32696
rect 16587 32647 16629 32656
rect 16875 32696 16917 32705
rect 16875 32656 16876 32696
rect 16916 32656 16917 32696
rect 16875 32647 16917 32656
rect 17068 32528 17108 34168
rect 17164 34159 17204 34168
rect 17259 34208 17301 34217
rect 17548 34208 17588 35176
rect 17739 34964 17781 34973
rect 17739 34924 17740 34964
rect 17780 34924 17781 34964
rect 17739 34915 17781 34924
rect 17259 34168 17260 34208
rect 17300 34168 17301 34208
rect 17259 34159 17301 34168
rect 17356 34168 17588 34208
rect 17260 33620 17300 34159
rect 17356 33704 17396 34168
rect 17547 34040 17589 34049
rect 17547 34000 17548 34040
rect 17588 34000 17589 34040
rect 17547 33991 17589 34000
rect 17356 33655 17396 33664
rect 17260 32873 17300 33580
rect 17259 32864 17301 32873
rect 17259 32824 17260 32864
rect 17300 32824 17301 32864
rect 17259 32815 17301 32824
rect 17548 32864 17588 33991
rect 17740 33704 17780 34915
rect 17836 34376 17876 34385
rect 17836 34217 17876 34336
rect 17835 34208 17877 34217
rect 17835 34168 17836 34208
rect 17876 34168 17877 34208
rect 17835 34159 17877 34168
rect 17740 33655 17780 33664
rect 17836 33704 17876 33713
rect 17355 32780 17397 32789
rect 17355 32740 17356 32780
rect 17396 32740 17397 32780
rect 17355 32731 17397 32740
rect 16396 32488 17108 32528
rect 16299 32192 16341 32201
rect 16299 32152 16300 32192
rect 16340 32152 16341 32192
rect 16299 32143 16341 32152
rect 16396 32192 16436 32488
rect 16396 32143 16436 32152
rect 16588 32192 16628 32201
rect 16300 31949 16340 32034
rect 16299 31940 16341 31949
rect 16299 31900 16300 31940
rect 16340 31900 16341 31940
rect 16299 31891 16341 31900
rect 16299 31772 16341 31781
rect 16299 31732 16300 31772
rect 16340 31732 16341 31772
rect 16299 31723 16341 31732
rect 16300 31520 16340 31723
rect 16300 31480 16436 31520
rect 16300 31352 16340 31363
rect 16300 31277 16340 31312
rect 16299 31268 16341 31277
rect 16299 31228 16300 31268
rect 16340 31228 16341 31268
rect 16299 31219 16341 31228
rect 16204 31060 16340 31100
rect 15531 30932 15573 30941
rect 15531 30892 15532 30932
rect 15572 30892 15573 30932
rect 15531 30883 15573 30892
rect 15435 30848 15477 30857
rect 15435 30808 15436 30848
rect 15476 30808 15477 30848
rect 15435 30799 15477 30808
rect 15819 30848 15861 30857
rect 15819 30808 15820 30848
rect 15860 30808 15861 30848
rect 15819 30799 15861 30808
rect 15532 30680 15572 30691
rect 15532 30605 15572 30640
rect 15820 30680 15860 30799
rect 15820 30631 15860 30640
rect 15916 30680 15956 30689
rect 15531 30596 15573 30605
rect 15531 30556 15532 30596
rect 15572 30556 15573 30596
rect 15531 30547 15573 30556
rect 15435 30512 15477 30521
rect 15435 30472 15436 30512
rect 15476 30472 15477 30512
rect 15435 30463 15477 30472
rect 14379 29840 14421 29849
rect 14571 29840 14613 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14476 29800 14572 29840
rect 14612 29800 14613 29840
rect 14380 28916 14420 29791
rect 14476 29093 14516 29800
rect 14571 29791 14613 29800
rect 15243 29840 15285 29849
rect 15243 29800 15244 29840
rect 15284 29800 15285 29840
rect 15243 29791 15285 29800
rect 15436 29840 15476 30463
rect 15819 30428 15861 30437
rect 15819 30388 15820 30428
rect 15860 30388 15861 30428
rect 15819 30379 15861 30388
rect 15436 29791 15476 29800
rect 15820 29840 15860 30379
rect 15916 30269 15956 30640
rect 16204 30428 16244 30437
rect 15915 30260 15957 30269
rect 15915 30220 15916 30260
rect 15956 30220 15957 30260
rect 15915 30211 15957 30220
rect 15820 29791 15860 29800
rect 14572 29706 14612 29791
rect 15819 29420 15861 29429
rect 15819 29380 15820 29420
rect 15860 29380 15861 29420
rect 15819 29371 15861 29380
rect 14859 29336 14901 29345
rect 14859 29296 14860 29336
rect 14900 29296 14901 29336
rect 14859 29287 14901 29296
rect 14571 29252 14613 29261
rect 14571 29212 14572 29252
rect 14612 29212 14613 29252
rect 14571 29203 14613 29212
rect 14572 29168 14612 29203
rect 14572 29117 14612 29128
rect 14860 29168 14900 29287
rect 14860 29119 14900 29128
rect 14475 29084 14517 29093
rect 14475 29044 14476 29084
rect 14516 29044 14517 29084
rect 14475 29035 14517 29044
rect 15820 29000 15860 29371
rect 16108 29168 16148 29177
rect 15436 28960 15860 29000
rect 15916 29000 15956 29009
rect 14476 28916 14516 28925
rect 14380 28876 14476 28916
rect 14476 28867 14516 28876
rect 14667 28916 14709 28925
rect 14667 28876 14668 28916
rect 14708 28876 14709 28916
rect 14667 28867 14709 28876
rect 14764 28916 14804 28925
rect 14187 28832 14229 28841
rect 14187 28792 14188 28832
rect 14228 28792 14229 28832
rect 14187 28783 14229 28792
rect 14188 28328 14228 28783
rect 14188 27656 14228 28288
rect 14572 27656 14612 27665
rect 14188 27607 14228 27616
rect 14489 27616 14572 27656
rect 14489 27497 14529 27616
rect 14572 27607 14612 27616
rect 14475 27488 14529 27497
rect 14475 27448 14476 27488
rect 14516 27448 14529 27488
rect 14475 27439 14517 27448
rect 14572 27413 14612 27498
rect 14571 27404 14613 27413
rect 14571 27364 14572 27404
rect 14612 27364 14613 27404
rect 14571 27355 14613 27364
rect 14668 27236 14708 28867
rect 14764 27833 14804 28876
rect 15339 28664 15381 28673
rect 15339 28624 15340 28664
rect 15380 28624 15381 28664
rect 15339 28615 15381 28624
rect 15243 28580 15285 28589
rect 15243 28540 15244 28580
rect 15284 28540 15285 28580
rect 15243 28531 15285 28540
rect 15244 28446 15284 28531
rect 14763 27824 14805 27833
rect 14763 27784 14764 27824
rect 14804 27784 14805 27824
rect 14763 27775 14805 27784
rect 15340 27740 15380 28615
rect 15340 27691 15380 27700
rect 14476 27196 14708 27236
rect 14764 27656 14804 27665
rect 14188 26816 14228 26827
rect 14188 26741 14228 26776
rect 14284 26816 14324 26825
rect 14187 26732 14229 26741
rect 14187 26692 14188 26732
rect 14228 26692 14229 26732
rect 14187 26683 14229 26692
rect 14284 26657 14324 26776
rect 14476 26816 14516 27196
rect 14764 26984 14804 27616
rect 14860 27656 14900 27665
rect 14860 27413 14900 27616
rect 15436 27656 15476 28960
rect 15724 28328 15764 28337
rect 15819 28328 15861 28337
rect 15764 28288 15820 28328
rect 15860 28288 15861 28328
rect 15724 28279 15764 28288
rect 15819 28279 15861 28288
rect 15436 27607 15476 27616
rect 15724 27656 15764 27665
rect 15627 27488 15669 27497
rect 15627 27448 15628 27488
rect 15668 27448 15669 27488
rect 15627 27439 15669 27448
rect 14859 27404 14901 27413
rect 14859 27364 14860 27404
rect 14900 27364 14901 27404
rect 14859 27355 14901 27364
rect 15052 27404 15092 27413
rect 15092 27364 15380 27404
rect 15052 27355 15092 27364
rect 14764 26944 14900 26984
rect 14476 26767 14516 26776
rect 14572 26816 14612 26825
rect 14283 26648 14325 26657
rect 14283 26608 14284 26648
rect 14324 26608 14325 26648
rect 14283 26599 14325 26608
rect 14380 26648 14420 26657
rect 14187 26564 14229 26573
rect 14187 26524 14188 26564
rect 14228 26524 14229 26564
rect 14187 26515 14229 26524
rect 14091 26312 14133 26321
rect 14091 26272 14092 26312
rect 14132 26272 14133 26312
rect 14091 26263 14133 26272
rect 14092 26144 14132 26153
rect 13803 25976 13845 25985
rect 13803 25936 13804 25976
rect 13844 25936 13845 25976
rect 13803 25927 13845 25936
rect 13995 25976 14037 25985
rect 13995 25936 13996 25976
rect 14036 25936 14037 25976
rect 13995 25927 14037 25936
rect 13612 25892 13652 25901
rect 13612 25481 13652 25852
rect 13707 25892 13749 25901
rect 13707 25852 13708 25892
rect 13748 25852 13749 25892
rect 13707 25843 13749 25852
rect 13708 25565 13748 25650
rect 13707 25556 13749 25565
rect 13707 25516 13708 25556
rect 13748 25516 13749 25556
rect 13707 25507 13749 25516
rect 13611 25472 13653 25481
rect 13611 25432 13612 25472
rect 13652 25432 13653 25472
rect 13611 25423 13653 25432
rect 13611 25304 13653 25313
rect 13611 25264 13612 25304
rect 13652 25264 13653 25304
rect 13611 25255 13653 25264
rect 13708 25304 13748 25313
rect 13804 25304 13844 25927
rect 13748 25264 13844 25304
rect 13900 25304 13940 25313
rect 13708 25255 13748 25264
rect 13612 25170 13652 25255
rect 13900 25145 13940 25264
rect 13899 25136 13941 25145
rect 12884 23164 12980 23204
rect 12844 23155 12884 23164
rect 13035 22868 13077 22877
rect 13035 22828 13036 22868
rect 13076 22828 13077 22868
rect 13035 22819 13077 22828
rect 12651 22616 12693 22625
rect 12651 22576 12652 22616
rect 12692 22576 12693 22616
rect 12651 22567 12693 22576
rect 12939 22448 12981 22457
rect 12460 22408 12692 22448
rect 12268 22231 12308 22240
rect 12555 22280 12597 22289
rect 12555 22240 12556 22280
rect 12596 22240 12597 22280
rect 12555 22231 12597 22240
rect 12652 22280 12692 22408
rect 12939 22408 12940 22448
rect 12980 22408 12981 22448
rect 12939 22399 12981 22408
rect 12940 22314 12980 22399
rect 12652 22231 12692 22240
rect 11788 21701 11828 22231
rect 12556 22146 12596 22231
rect 11787 21692 11829 21701
rect 11787 21652 11788 21692
rect 11828 21652 11829 21692
rect 11787 21643 11829 21652
rect 11636 21568 11732 21608
rect 11788 21608 11828 21643
rect 11596 21559 11636 21568
rect 11788 21558 11828 21568
rect 13036 21608 13076 22819
rect 13516 22793 13556 24592
rect 13804 25096 13900 25136
rect 13940 25096 13941 25136
rect 13804 24632 13844 25096
rect 13899 25087 13941 25096
rect 13804 24583 13844 24592
rect 13900 24632 13940 24641
rect 13803 24380 13845 24389
rect 13803 24340 13804 24380
rect 13844 24340 13845 24380
rect 13803 24331 13845 24340
rect 13804 23792 13844 24331
rect 13900 24053 13940 24592
rect 14092 24464 14132 26104
rect 14188 26144 14228 26515
rect 14380 26489 14420 26608
rect 14379 26480 14421 26489
rect 14379 26440 14380 26480
rect 14420 26440 14421 26480
rect 14379 26431 14421 26440
rect 14572 26312 14612 26776
rect 14727 26816 14767 26827
rect 14727 26741 14767 26776
rect 14726 26732 14768 26741
rect 14726 26692 14727 26732
rect 14767 26692 14768 26732
rect 14726 26683 14768 26692
rect 14860 26573 14900 26944
rect 15148 26825 15188 26910
rect 14955 26816 14997 26825
rect 14955 26776 14956 26816
rect 14996 26776 14997 26816
rect 14955 26767 14997 26776
rect 15147 26816 15189 26825
rect 15147 26776 15148 26816
rect 15188 26776 15189 26816
rect 15147 26767 15189 26776
rect 15340 26816 15380 27364
rect 15340 26767 15380 26776
rect 15435 26816 15477 26825
rect 15435 26776 15436 26816
rect 15476 26776 15477 26816
rect 15435 26767 15477 26776
rect 15628 26816 15668 27439
rect 15724 27329 15764 27616
rect 15820 27488 15860 28279
rect 15916 27665 15956 28960
rect 16108 28337 16148 29128
rect 16107 28328 16149 28337
rect 16107 28288 16108 28328
rect 16148 28288 16149 28328
rect 16107 28279 16149 28288
rect 16012 28244 16052 28253
rect 16012 27749 16052 28204
rect 16011 27740 16053 27749
rect 16011 27700 16012 27740
rect 16052 27700 16053 27740
rect 16011 27691 16053 27700
rect 15915 27656 15957 27665
rect 15915 27616 15916 27656
rect 15956 27616 15957 27656
rect 15915 27607 15957 27616
rect 16204 27572 16244 30388
rect 16012 27532 16244 27572
rect 15820 27448 15956 27488
rect 15723 27320 15765 27329
rect 15723 27280 15724 27320
rect 15764 27280 15765 27320
rect 15723 27271 15765 27280
rect 14956 26682 14996 26767
rect 15052 26732 15092 26741
rect 15052 26648 15092 26692
rect 15052 26608 15188 26648
rect 14667 26564 14709 26573
rect 14667 26524 14668 26564
rect 14708 26524 14709 26564
rect 14667 26515 14709 26524
rect 14859 26564 14901 26573
rect 14859 26524 14860 26564
rect 14900 26524 14901 26564
rect 14859 26515 14901 26524
rect 14476 26272 14612 26312
rect 14380 26144 14420 26153
rect 14188 26095 14228 26104
rect 14284 26104 14380 26144
rect 14284 25817 14324 26104
rect 14380 26095 14420 26104
rect 14380 25892 14420 25901
rect 14283 25808 14325 25817
rect 14283 25768 14284 25808
rect 14324 25768 14325 25808
rect 14283 25759 14325 25768
rect 14380 25313 14420 25852
rect 14379 25304 14421 25313
rect 14379 25264 14380 25304
rect 14420 25264 14421 25304
rect 14379 25255 14421 25264
rect 14476 25229 14516 26272
rect 14571 26144 14613 26153
rect 14571 26104 14572 26144
rect 14612 26104 14613 26144
rect 14571 26095 14613 26104
rect 14668 26144 14708 26515
rect 15051 26480 15093 26489
rect 15051 26440 15052 26480
rect 15092 26440 15093 26480
rect 15051 26431 15093 26440
rect 14763 26312 14805 26321
rect 14763 26272 14764 26312
rect 14804 26272 14805 26312
rect 14763 26263 14805 26272
rect 14955 26312 14997 26321
rect 14955 26272 14956 26312
rect 14996 26272 14997 26312
rect 14955 26263 14997 26272
rect 14764 26178 14804 26263
rect 14859 26228 14901 26237
rect 14859 26188 14860 26228
rect 14900 26188 14901 26228
rect 14859 26179 14901 26188
rect 14668 26095 14708 26104
rect 14860 26144 14900 26179
rect 14572 26010 14612 26095
rect 14860 25901 14900 26104
rect 14859 25892 14901 25901
rect 14859 25852 14860 25892
rect 14900 25852 14901 25892
rect 14859 25843 14901 25852
rect 14956 25556 14996 26263
rect 15052 25733 15092 26431
rect 15051 25724 15093 25733
rect 15051 25684 15052 25724
rect 15092 25684 15093 25724
rect 15051 25675 15093 25684
rect 14956 25516 15092 25556
rect 15052 25397 15092 25516
rect 15148 25481 15188 26608
rect 15436 26573 15476 26767
rect 15531 26732 15573 26741
rect 15531 26692 15532 26732
rect 15572 26692 15573 26732
rect 15531 26683 15573 26692
rect 15532 26598 15572 26683
rect 15435 26564 15477 26573
rect 15435 26524 15436 26564
rect 15476 26524 15477 26564
rect 15435 26515 15477 26524
rect 15339 26480 15381 26489
rect 15339 26440 15340 26480
rect 15380 26440 15381 26480
rect 15339 26431 15381 26440
rect 15340 26321 15380 26431
rect 15339 26312 15381 26321
rect 15339 26272 15340 26312
rect 15380 26272 15381 26312
rect 15339 26263 15381 26272
rect 15244 26144 15284 26155
rect 15244 26069 15284 26104
rect 15339 26144 15381 26153
rect 15339 26104 15340 26144
rect 15380 26104 15381 26144
rect 15339 26095 15381 26104
rect 15436 26144 15476 26515
rect 15628 26396 15668 26776
rect 15436 26095 15476 26104
rect 15532 26356 15668 26396
rect 15243 26060 15285 26069
rect 15243 26020 15244 26060
rect 15284 26020 15285 26060
rect 15243 26011 15285 26020
rect 15340 26010 15380 26095
rect 15532 25817 15572 26356
rect 15628 26272 15860 26312
rect 15531 25808 15573 25817
rect 15531 25768 15532 25808
rect 15572 25768 15573 25808
rect 15531 25759 15573 25768
rect 15244 25556 15284 25565
rect 15628 25556 15668 26272
rect 15724 26144 15764 26155
rect 15724 26069 15764 26104
rect 15820 26144 15860 26272
rect 15820 26095 15860 26104
rect 15723 26060 15765 26069
rect 15723 26020 15724 26060
rect 15764 26020 15765 26060
rect 15723 26011 15765 26020
rect 15916 25976 15956 27448
rect 16012 26816 16052 27532
rect 16300 27488 16340 31060
rect 16396 30596 16436 31480
rect 16588 31445 16628 32152
rect 16587 31436 16629 31445
rect 16587 31396 16588 31436
rect 16628 31396 16629 31436
rect 16587 31387 16629 31396
rect 17163 31352 17205 31361
rect 17163 31312 17164 31352
rect 17204 31312 17205 31352
rect 17163 31303 17205 31312
rect 17164 31218 17204 31303
rect 16972 31184 17012 31193
rect 16491 30848 16533 30857
rect 16491 30808 16492 30848
rect 16532 30808 16533 30848
rect 16491 30799 16533 30808
rect 16492 30714 16532 30799
rect 16972 30773 17012 31144
rect 16971 30764 17013 30773
rect 16971 30724 16972 30764
rect 17012 30724 17013 30764
rect 16971 30715 17013 30724
rect 16491 30596 16533 30605
rect 16396 30556 16492 30596
rect 16532 30556 16533 30596
rect 16491 30547 16533 30556
rect 16492 30092 16532 30547
rect 16492 30043 16532 30052
rect 16684 29968 17012 30008
rect 16684 29336 16724 29968
rect 16684 29287 16724 29296
rect 16876 29840 16916 29849
rect 16972 29840 17012 29968
rect 17260 29840 17300 29849
rect 16972 29800 17260 29840
rect 16491 29168 16533 29177
rect 16491 29128 16492 29168
rect 16532 29128 16533 29168
rect 16491 29119 16533 29128
rect 16588 29168 16628 29177
rect 16492 29034 16532 29119
rect 16012 26767 16052 26776
rect 16108 27448 16340 27488
rect 16396 28328 16436 28337
rect 16396 27488 16436 28288
rect 16588 27581 16628 29128
rect 16779 29168 16821 29177
rect 16779 29128 16780 29168
rect 16820 29128 16821 29168
rect 16779 29119 16821 29128
rect 16780 29034 16820 29119
rect 16876 28841 16916 29800
rect 17260 29791 17300 29800
rect 16971 29252 17013 29261
rect 16971 29212 16972 29252
rect 17012 29212 17013 29252
rect 16971 29203 17013 29212
rect 16972 29118 17012 29203
rect 16875 28832 16917 28841
rect 16875 28792 16876 28832
rect 16916 28792 16917 28832
rect 16875 28783 16917 28792
rect 17356 28580 17396 32731
rect 17451 32696 17493 32705
rect 17451 32656 17452 32696
rect 17492 32656 17493 32696
rect 17451 32647 17493 32656
rect 17452 32201 17492 32647
rect 17451 32192 17493 32201
rect 17451 32152 17452 32192
rect 17492 32152 17493 32192
rect 17451 32143 17493 32152
rect 17452 31865 17492 32143
rect 17451 31856 17493 31865
rect 17451 31816 17452 31856
rect 17492 31816 17493 31856
rect 17451 31807 17493 31816
rect 17548 31688 17588 32824
rect 17836 32612 17876 33664
rect 18027 33704 18069 33713
rect 18027 33664 18028 33704
rect 18068 33664 18069 33704
rect 18124 33704 18164 35260
rect 18220 35251 18260 35260
rect 18411 35300 18453 35309
rect 18411 35260 18412 35300
rect 18452 35260 18453 35300
rect 18411 35251 18453 35260
rect 18412 35166 18452 35251
rect 18796 35216 18836 36007
rect 19180 35922 19220 36007
rect 21100 35888 21140 35897
rect 18988 35720 19028 35729
rect 18988 35309 19028 35680
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 21100 35384 21140 35848
rect 21195 35720 21237 35729
rect 21195 35680 21196 35720
rect 21236 35680 21237 35720
rect 21195 35671 21237 35680
rect 22347 35720 22389 35729
rect 22347 35680 22348 35720
rect 22388 35680 22389 35720
rect 22347 35671 22389 35680
rect 21196 35586 21236 35671
rect 21100 35335 21140 35344
rect 18987 35300 19029 35309
rect 18987 35260 18988 35300
rect 19028 35260 19029 35300
rect 18987 35251 19029 35260
rect 18796 35167 18836 35176
rect 19659 35216 19701 35225
rect 19659 35176 19660 35216
rect 19700 35176 19701 35216
rect 19659 35167 19701 35176
rect 20043 35216 20085 35225
rect 20043 35176 20044 35216
rect 20084 35176 20085 35216
rect 20043 35167 20085 35176
rect 21772 35216 21812 35225
rect 19660 35082 19700 35167
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 18316 34553 18356 34638
rect 18796 34553 18836 34638
rect 18315 34544 18357 34553
rect 18315 34504 18316 34544
rect 18356 34504 18357 34544
rect 18315 34495 18357 34504
rect 18795 34544 18837 34553
rect 18795 34504 18796 34544
rect 18836 34504 18837 34544
rect 18795 34495 18837 34504
rect 19659 34544 19701 34553
rect 19659 34504 19660 34544
rect 19700 34504 19701 34544
rect 19659 34495 19701 34504
rect 19947 34544 19989 34553
rect 19947 34504 19948 34544
rect 19988 34504 19989 34544
rect 20044 34544 20084 35167
rect 21772 34973 21812 35176
rect 21964 35048 22004 35057
rect 20811 34964 20853 34973
rect 20811 34924 20812 34964
rect 20852 34924 20853 34964
rect 20811 34915 20853 34924
rect 21771 34964 21813 34973
rect 21771 34924 21772 34964
rect 21812 34924 21813 34964
rect 21771 34915 21813 34924
rect 20812 34830 20852 34915
rect 21675 34544 21717 34553
rect 20044 34504 20276 34544
rect 19947 34495 19989 34504
rect 19371 34460 19413 34469
rect 19371 34420 19372 34460
rect 19412 34420 19413 34460
rect 19371 34411 19413 34420
rect 18508 34376 18548 34385
rect 18316 34336 18508 34376
rect 18316 33872 18356 34336
rect 18508 34327 18548 34336
rect 18603 34376 18645 34385
rect 18603 34336 18604 34376
rect 18644 34336 18645 34376
rect 18603 34327 18645 34336
rect 18795 34376 18837 34385
rect 18795 34336 18796 34376
rect 18836 34336 18837 34376
rect 18795 34327 18837 34336
rect 18604 34242 18644 34327
rect 18796 34242 18836 34327
rect 18316 33823 18356 33832
rect 18988 34208 19028 34217
rect 18988 33788 19028 34168
rect 18988 33739 19028 33748
rect 18220 33704 18260 33713
rect 18508 33704 18548 33713
rect 18124 33664 18220 33704
rect 18027 33655 18069 33664
rect 18220 33655 18260 33664
rect 18316 33664 18508 33704
rect 18028 32705 18068 33655
rect 18316 33452 18356 33664
rect 18508 33655 18548 33664
rect 18699 33704 18741 33713
rect 18699 33664 18700 33704
rect 18740 33664 18741 33704
rect 18699 33655 18741 33664
rect 18796 33704 18836 33713
rect 18700 33570 18740 33655
rect 18124 33412 18356 33452
rect 18508 33452 18548 33461
rect 18548 33412 18740 33452
rect 18027 32696 18069 32705
rect 18027 32656 18028 32696
rect 18068 32656 18069 32696
rect 18027 32647 18069 32656
rect 17452 31648 17588 31688
rect 17740 32572 17876 32612
rect 17452 28589 17492 31648
rect 17740 31520 17780 32572
rect 17931 32444 17973 32453
rect 17931 32404 17932 32444
rect 17972 32404 17973 32444
rect 17931 32395 17973 32404
rect 17835 32192 17877 32201
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 17932 32192 17972 32395
rect 18124 32360 18164 33412
rect 18508 33403 18548 33412
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 18219 33116 18261 33125
rect 18219 33076 18220 33116
rect 18260 33076 18261 33116
rect 18219 33067 18261 33076
rect 18124 32311 18164 32320
rect 17932 32143 17972 32152
rect 18028 32192 18068 32201
rect 18220 32192 18260 33067
rect 18411 32864 18453 32873
rect 18411 32824 18412 32864
rect 18452 32824 18453 32864
rect 18411 32815 18453 32824
rect 18604 32864 18644 32873
rect 18700 32864 18740 33412
rect 18796 33125 18836 33664
rect 19372 33704 19412 34411
rect 19660 34376 19700 34495
rect 19660 34327 19700 34336
rect 19851 34376 19893 34385
rect 19851 34336 19852 34376
rect 19892 34336 19893 34376
rect 19851 34327 19893 34336
rect 19948 34376 19988 34495
rect 19948 34327 19988 34336
rect 20043 34376 20085 34385
rect 20043 34336 20044 34376
rect 20084 34336 20085 34376
rect 20043 34327 20085 34336
rect 20140 34355 20180 34387
rect 19852 34242 19892 34327
rect 20044 34242 20084 34327
rect 20140 34301 20180 34315
rect 20139 34292 20181 34301
rect 20139 34252 20140 34292
rect 20180 34252 20181 34292
rect 20139 34243 20181 34252
rect 19947 34208 19989 34217
rect 19947 34168 19948 34208
rect 19988 34168 19989 34208
rect 19947 34159 19989 34168
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 19372 33655 19412 33664
rect 18795 33116 18837 33125
rect 18795 33076 18796 33116
rect 18836 33076 18837 33116
rect 18795 33067 18837 33076
rect 19851 33116 19893 33125
rect 19851 33076 19852 33116
rect 19892 33076 19893 33116
rect 19851 33067 19893 33076
rect 19659 33032 19701 33041
rect 19659 32992 19660 33032
rect 19700 32992 19701 33032
rect 19659 32983 19701 32992
rect 19275 32948 19317 32957
rect 19275 32908 19276 32948
rect 19316 32908 19317 32948
rect 19275 32899 19317 32908
rect 18644 32824 18740 32864
rect 18604 32815 18644 32824
rect 18412 32730 18452 32815
rect 19276 32814 19316 32899
rect 19660 32898 19700 32983
rect 19852 32982 19892 33067
rect 19371 32864 19413 32873
rect 19371 32824 19372 32864
rect 19412 32824 19413 32864
rect 19371 32815 19413 32824
rect 19948 32864 19988 34159
rect 20236 33713 20276 34504
rect 21675 34504 21676 34544
rect 21716 34504 21717 34544
rect 21675 34495 21717 34504
rect 21195 34376 21237 34385
rect 21195 34336 21196 34376
rect 21236 34336 21332 34376
rect 21195 34327 21237 34336
rect 21196 34242 21236 34327
rect 20523 34208 20565 34217
rect 20523 34168 20524 34208
rect 20564 34168 20565 34208
rect 20523 34159 20565 34168
rect 20524 34074 20564 34159
rect 21292 33872 21332 34336
rect 21387 34292 21429 34301
rect 21387 34252 21388 34292
rect 21428 34252 21429 34292
rect 21387 34243 21429 34252
rect 21388 34158 21428 34243
rect 21579 34208 21621 34217
rect 21579 34168 21580 34208
rect 21620 34168 21621 34208
rect 21579 34159 21621 34168
rect 21388 33872 21428 33881
rect 21292 33832 21388 33872
rect 21388 33823 21428 33832
rect 21580 33797 21620 34159
rect 21676 33872 21716 34495
rect 21772 34376 21812 34385
rect 21964 34376 22004 35008
rect 21812 34336 22004 34376
rect 21772 34327 21812 34336
rect 22155 34292 22197 34301
rect 22155 34252 22156 34292
rect 22196 34252 22197 34292
rect 22155 34243 22197 34252
rect 21771 33872 21813 33881
rect 21676 33832 21772 33872
rect 21812 33832 21813 33872
rect 21771 33823 21813 33832
rect 22156 33872 22196 34243
rect 22156 33823 22196 33832
rect 21579 33788 21621 33797
rect 21579 33748 21580 33788
rect 21620 33748 21621 33788
rect 21579 33739 21621 33748
rect 20235 33704 20277 33713
rect 20235 33664 20236 33704
rect 20276 33664 20277 33704
rect 20235 33655 20277 33664
rect 21580 33704 21620 33739
rect 19948 32815 19988 32824
rect 18411 32444 18453 32453
rect 18411 32404 18412 32444
rect 18452 32404 18453 32444
rect 18411 32395 18453 32404
rect 18068 32152 18260 32192
rect 18412 32192 18452 32395
rect 19372 32192 19412 32815
rect 20236 32789 20276 33655
rect 21580 33654 21620 33664
rect 21676 33704 21716 33713
rect 21388 33452 21428 33461
rect 21428 33412 21620 33452
rect 21388 33403 21428 33412
rect 20523 33032 20565 33041
rect 20523 32992 20524 33032
rect 20564 32992 20565 33032
rect 20523 32983 20565 32992
rect 21291 33032 21333 33041
rect 21291 32992 21292 33032
rect 21332 32992 21333 33032
rect 21291 32983 21333 32992
rect 20235 32780 20277 32789
rect 20235 32740 20236 32780
rect 20276 32740 20277 32780
rect 20235 32731 20277 32740
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 19660 32192 19700 32201
rect 19372 32152 19660 32192
rect 18028 32143 18068 32152
rect 18412 32143 18452 32152
rect 19660 32143 19700 32152
rect 20524 32192 20564 32983
rect 20907 32948 20949 32957
rect 20907 32908 20908 32948
rect 20948 32908 20949 32948
rect 20907 32899 20949 32908
rect 20524 32143 20564 32152
rect 20908 32192 20948 32899
rect 21292 32898 21332 32983
rect 21580 32864 21620 33412
rect 21676 33041 21716 33664
rect 21772 33704 21812 33823
rect 22251 33788 22293 33797
rect 22251 33748 22252 33788
rect 22292 33748 22293 33788
rect 22251 33739 22293 33748
rect 21772 33655 21812 33664
rect 21868 33704 21908 33713
rect 22060 33704 22100 33713
rect 21908 33664 22060 33704
rect 21868 33655 21908 33664
rect 22060 33655 22100 33664
rect 22252 33704 22292 33739
rect 21771 33536 21813 33545
rect 21771 33496 21772 33536
rect 21812 33496 21813 33536
rect 21771 33487 21813 33496
rect 21675 33032 21717 33041
rect 21675 32992 21676 33032
rect 21716 32992 21717 33032
rect 21675 32983 21717 32992
rect 21580 32815 21620 32824
rect 21676 32864 21716 32873
rect 21772 32864 21812 33487
rect 21716 32824 21812 32864
rect 21963 32864 22005 32873
rect 21963 32824 21964 32864
rect 22004 32824 22005 32864
rect 21676 32815 21716 32824
rect 21963 32815 22005 32824
rect 21964 32730 22004 32815
rect 22252 32789 22292 33664
rect 22348 33704 22388 35671
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 23115 35216 23157 35225
rect 23115 35176 23116 35216
rect 23156 35176 23157 35216
rect 23115 35167 23157 35176
rect 24075 35216 24117 35225
rect 24075 35176 24076 35216
rect 24116 35176 24117 35216
rect 24075 35167 24117 35176
rect 26476 35216 26516 35225
rect 22636 34376 22676 34385
rect 22636 33713 22676 34336
rect 23116 33872 23156 35167
rect 24076 35082 24116 35167
rect 26187 35048 26229 35057
rect 26187 35008 26188 35048
rect 26228 35008 26229 35048
rect 26187 34999 26229 35008
rect 23116 33823 23156 33832
rect 23404 34964 23444 34973
rect 25804 34964 25844 34973
rect 23404 33788 23444 34924
rect 25612 34924 25804 34964
rect 24844 34544 24884 34553
rect 24652 34376 24692 34385
rect 23788 34208 23828 34217
rect 23692 34168 23788 34208
rect 23692 33965 23732 34168
rect 23788 34159 23828 34168
rect 23980 34208 24020 34217
rect 23787 34040 23829 34049
rect 23787 34000 23788 34040
rect 23828 34000 23829 34040
rect 23787 33991 23829 34000
rect 23691 33956 23733 33965
rect 23691 33916 23692 33956
rect 23732 33916 23733 33956
rect 23691 33907 23733 33916
rect 23404 33739 23444 33748
rect 22348 33655 22388 33664
rect 22635 33704 22677 33713
rect 22635 33664 22636 33704
rect 22676 33664 22677 33704
rect 22635 33655 22677 33664
rect 22924 33704 22964 33713
rect 22251 32780 22293 32789
rect 22251 32740 22252 32780
rect 22292 32740 22293 32780
rect 22251 32731 22293 32740
rect 22156 32360 22196 32369
rect 22252 32360 22292 32731
rect 22196 32320 22292 32360
rect 22156 32311 22196 32320
rect 20908 32143 20948 32152
rect 22540 32192 22580 32201
rect 17836 32058 17876 32143
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 22540 31529 22580 32152
rect 18220 31520 18260 31529
rect 17548 31480 17780 31520
rect 18124 31480 18220 31520
rect 17548 30605 17588 31480
rect 17836 31352 17876 31361
rect 17836 30857 17876 31312
rect 17835 30848 17877 30857
rect 17835 30808 17836 30848
rect 17876 30808 17877 30848
rect 17835 30799 17877 30808
rect 17644 30680 17684 30689
rect 17684 30640 17780 30680
rect 17644 30631 17684 30640
rect 17547 30596 17589 30605
rect 17547 30556 17548 30596
rect 17588 30556 17589 30596
rect 17547 30547 17589 30556
rect 17643 29672 17685 29681
rect 17643 29632 17644 29672
rect 17684 29632 17685 29672
rect 17643 29623 17685 29632
rect 17644 29429 17684 29623
rect 17643 29420 17685 29429
rect 17643 29380 17644 29420
rect 17684 29380 17685 29420
rect 17643 29371 17685 29380
rect 17644 29168 17684 29371
rect 17644 29119 17684 29128
rect 16684 28540 17396 28580
rect 17451 28580 17493 28589
rect 17451 28540 17452 28580
rect 17492 28540 17493 28580
rect 16587 27572 16629 27581
rect 16587 27532 16588 27572
rect 16628 27532 16629 27572
rect 16587 27523 16629 27532
rect 16492 27488 16532 27497
rect 16396 27448 16492 27488
rect 16108 26816 16148 27448
rect 16492 27439 16532 27448
rect 16108 26489 16148 26776
rect 16300 26816 16340 26825
rect 16204 26648 16244 26657
rect 16107 26480 16149 26489
rect 16107 26440 16108 26480
rect 16148 26440 16149 26480
rect 16107 26431 16149 26440
rect 16107 26312 16149 26321
rect 16107 26272 16108 26312
rect 16148 26272 16149 26312
rect 16107 26263 16149 26272
rect 16011 26144 16053 26153
rect 16011 26104 16012 26144
rect 16052 26104 16053 26144
rect 16011 26095 16053 26104
rect 16108 26144 16148 26263
rect 16204 26153 16244 26608
rect 16300 26312 16340 26776
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16588 26682 16628 26767
rect 16300 26272 16436 26312
rect 16396 26153 16436 26272
rect 16204 26144 16249 26153
rect 16204 26104 16209 26144
rect 16108 26095 16148 26104
rect 16209 26095 16249 26104
rect 16395 26144 16437 26153
rect 16395 26104 16396 26144
rect 16436 26104 16437 26144
rect 16395 26095 16437 26104
rect 16587 26144 16629 26153
rect 16587 26104 16588 26144
rect 16628 26104 16629 26144
rect 16587 26095 16629 26104
rect 16684 26144 16724 28540
rect 17451 28531 17493 28540
rect 17260 28328 17300 28337
rect 17260 27833 17300 28288
rect 17740 27833 17780 30640
rect 18124 30092 18164 31480
rect 18220 31471 18260 31480
rect 18412 31520 18452 31529
rect 20715 31520 20757 31529
rect 18452 31480 18548 31520
rect 18412 31471 18452 31480
rect 18508 30680 18548 31480
rect 20715 31480 20716 31520
rect 20756 31480 20757 31520
rect 20715 31471 20757 31480
rect 21099 31520 21141 31529
rect 21099 31480 21100 31520
rect 21140 31480 21141 31520
rect 21099 31471 21141 31480
rect 21676 31520 21716 31529
rect 22059 31520 22101 31529
rect 21716 31480 21812 31520
rect 21676 31471 21716 31480
rect 20716 31352 20756 31471
rect 20716 31303 20756 31312
rect 20908 31352 20948 31361
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 18891 30764 18933 30773
rect 18891 30724 18892 30764
rect 18932 30724 18933 30764
rect 18891 30715 18933 30724
rect 18508 30631 18548 30640
rect 18892 30630 18932 30715
rect 19084 30680 19124 30689
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 18124 30052 18548 30092
rect 18508 29840 18548 30052
rect 18508 29791 18548 29800
rect 17932 29756 17972 29765
rect 18124 29756 18164 29765
rect 17972 29716 18124 29756
rect 17932 29707 17972 29716
rect 18124 29707 18164 29716
rect 18699 29336 18741 29345
rect 18699 29296 18700 29336
rect 18740 29296 18741 29336
rect 18699 29287 18741 29296
rect 18700 29202 18740 29287
rect 19084 29177 19124 30640
rect 19179 30680 19221 30689
rect 19179 30640 19180 30680
rect 19220 30640 19221 30680
rect 19179 30631 19221 30640
rect 19276 30680 19316 30689
rect 19180 30546 19220 30631
rect 19276 29924 19316 30640
rect 19372 30680 19412 30691
rect 19372 30605 19412 30640
rect 19660 30680 19700 30689
rect 19371 30596 19413 30605
rect 19371 30556 19372 30596
rect 19412 30556 19413 30596
rect 19371 30547 19413 30556
rect 19180 29884 19316 29924
rect 19180 29681 19220 29884
rect 19372 29840 19412 29849
rect 19276 29800 19372 29840
rect 19179 29672 19221 29681
rect 19179 29632 19180 29672
rect 19220 29632 19221 29672
rect 19179 29623 19221 29632
rect 17836 29168 17876 29177
rect 17836 29000 17876 29128
rect 19083 29168 19125 29177
rect 19083 29128 19084 29168
rect 19124 29128 19125 29168
rect 19083 29119 19125 29128
rect 18795 29084 18837 29093
rect 18795 29044 18796 29084
rect 18836 29044 18837 29084
rect 18795 29035 18837 29044
rect 17836 28960 18164 29000
rect 18124 28580 18164 28960
rect 18508 28916 18548 28925
rect 18548 28876 18740 28916
rect 18508 28867 18548 28876
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 18412 28580 18452 28589
rect 18124 28540 18412 28580
rect 17259 27824 17301 27833
rect 17259 27784 17260 27824
rect 17300 27784 17301 27824
rect 17259 27775 17301 27784
rect 17739 27824 17781 27833
rect 17739 27784 17740 27824
rect 17780 27784 17781 27824
rect 17739 27775 17781 27784
rect 17451 27740 17493 27749
rect 17451 27700 17452 27740
rect 17492 27700 17493 27740
rect 17451 27691 17493 27700
rect 17356 27656 17396 27665
rect 17356 27497 17396 27616
rect 17452 27606 17492 27691
rect 17548 27656 17588 27667
rect 17548 27581 17588 27616
rect 17644 27656 17684 27665
rect 17547 27572 17589 27581
rect 17547 27532 17548 27572
rect 17588 27532 17589 27572
rect 17547 27523 17589 27532
rect 17355 27488 17397 27497
rect 17355 27448 17356 27488
rect 17396 27448 17397 27488
rect 17355 27439 17397 27448
rect 17644 27068 17684 27616
rect 18124 27656 18164 27665
rect 17835 27404 17877 27413
rect 17835 27364 17836 27404
rect 17876 27364 17877 27404
rect 17835 27355 17877 27364
rect 17836 27270 17876 27355
rect 18124 27077 18164 27616
rect 18220 27656 18260 28540
rect 18412 28531 18452 28540
rect 18603 28580 18645 28589
rect 18603 28540 18604 28580
rect 18644 28540 18645 28580
rect 18603 28531 18645 28540
rect 18604 28446 18644 28531
rect 18700 28328 18740 28876
rect 18796 28589 18836 29035
rect 18795 28580 18837 28589
rect 18795 28540 18796 28580
rect 18836 28540 18837 28580
rect 18795 28531 18837 28540
rect 19083 28412 19125 28421
rect 19083 28372 19084 28412
rect 19124 28372 19125 28412
rect 19083 28363 19125 28372
rect 18700 28076 18740 28288
rect 18987 28328 19029 28337
rect 18987 28288 18988 28328
rect 19028 28288 19029 28328
rect 18987 28279 19029 28288
rect 18988 28194 19028 28279
rect 18700 28036 19028 28076
rect 18220 27607 18260 27616
rect 18508 27656 18548 27665
rect 18508 27413 18548 27616
rect 18796 27656 18836 27665
rect 18796 27497 18836 27616
rect 18892 27656 18932 27665
rect 18795 27488 18837 27497
rect 18795 27448 18796 27488
rect 18836 27448 18837 27488
rect 18795 27439 18837 27448
rect 18507 27404 18549 27413
rect 18507 27364 18508 27404
rect 18548 27364 18549 27404
rect 18507 27355 18549 27364
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 17740 27068 17780 27077
rect 17644 27028 17740 27068
rect 17740 27019 17780 27028
rect 18123 27068 18165 27077
rect 18123 27028 18124 27068
rect 18164 27028 18165 27068
rect 18123 27019 18165 27028
rect 18699 27068 18741 27077
rect 18699 27028 18700 27068
rect 18740 27028 18741 27068
rect 18699 27019 18741 27028
rect 18603 26984 18645 26993
rect 18603 26944 18604 26984
rect 18644 26944 18645 26984
rect 18603 26935 18645 26944
rect 16972 26825 17012 26910
rect 16779 26816 16821 26825
rect 16779 26776 16780 26816
rect 16820 26776 16821 26816
rect 16779 26767 16821 26776
rect 16971 26816 17013 26825
rect 16971 26776 16972 26816
rect 17012 26776 17013 26816
rect 16971 26767 17013 26776
rect 17163 26816 17205 26825
rect 17163 26776 17164 26816
rect 17204 26776 17205 26816
rect 17163 26767 17205 26776
rect 17835 26816 17877 26825
rect 17835 26776 17836 26816
rect 17876 26776 17877 26816
rect 17835 26767 17877 26776
rect 18124 26816 18164 26825
rect 16780 26682 16820 26767
rect 17068 26732 17108 26741
rect 17068 26321 17108 26692
rect 17164 26682 17204 26767
rect 17836 26682 17876 26767
rect 18124 26657 18164 26776
rect 18220 26816 18260 26825
rect 18028 26648 18068 26657
rect 17932 26608 18028 26648
rect 17163 26396 17205 26405
rect 17163 26356 17164 26396
rect 17204 26356 17205 26396
rect 17163 26347 17205 26356
rect 17067 26312 17109 26321
rect 17067 26272 17068 26312
rect 17108 26272 17109 26312
rect 17067 26263 17109 26272
rect 16684 26095 16724 26104
rect 16780 26144 16820 26155
rect 16012 26010 16052 26095
rect 16588 26010 16628 26095
rect 16780 26069 16820 26104
rect 16876 26144 16916 26153
rect 16779 26060 16821 26069
rect 16779 26020 16780 26060
rect 16820 26020 16821 26060
rect 16779 26011 16821 26020
rect 15820 25936 15956 25976
rect 15284 25516 15668 25556
rect 15724 25892 15764 25901
rect 15244 25507 15284 25516
rect 15147 25472 15189 25481
rect 15147 25432 15148 25472
rect 15188 25432 15189 25472
rect 15147 25423 15189 25432
rect 15724 25397 15764 25852
rect 15051 25388 15093 25397
rect 15051 25348 15052 25388
rect 15092 25348 15093 25388
rect 15051 25339 15093 25348
rect 15531 25388 15573 25397
rect 15531 25348 15532 25388
rect 15572 25348 15573 25388
rect 15531 25339 15573 25348
rect 15723 25388 15765 25397
rect 15723 25348 15724 25388
rect 15764 25348 15765 25388
rect 15723 25339 15765 25348
rect 14956 25304 14996 25313
rect 14475 25220 14517 25229
rect 14475 25180 14476 25220
rect 14516 25180 14517 25220
rect 14475 25171 14517 25180
rect 14572 25136 14612 25145
rect 14476 24632 14516 24641
rect 14572 24632 14612 25096
rect 14516 24592 14612 24632
rect 14476 24583 14516 24592
rect 14188 24464 14228 24473
rect 14764 24464 14804 24473
rect 14092 24424 14188 24464
rect 14188 24415 14228 24424
rect 14668 24424 14764 24464
rect 14379 24380 14421 24389
rect 14379 24340 14380 24380
rect 14420 24340 14421 24380
rect 14379 24331 14421 24340
rect 14380 24246 14420 24331
rect 13899 24044 13941 24053
rect 13899 24004 13900 24044
rect 13940 24004 13941 24044
rect 13899 23995 13941 24004
rect 13995 23960 14037 23969
rect 13995 23920 13996 23960
rect 14036 23920 14037 23960
rect 13995 23911 14037 23920
rect 14092 23960 14132 23969
rect 14132 23920 14324 23960
rect 14092 23911 14132 23920
rect 13804 23743 13844 23752
rect 13899 23792 13941 23801
rect 13899 23752 13900 23792
rect 13940 23752 13941 23792
rect 13996 23792 14036 23911
rect 14092 23792 14132 23801
rect 13996 23752 14092 23792
rect 13899 23743 13941 23752
rect 14092 23743 14132 23752
rect 14284 23792 14324 23920
rect 14284 23743 14324 23752
rect 14668 23792 14708 24424
rect 14764 24415 14804 24424
rect 14956 23876 14996 25264
rect 15052 25304 15092 25339
rect 15052 25253 15092 25264
rect 15244 25304 15284 25315
rect 15244 25229 15284 25264
rect 15243 25220 15285 25229
rect 15243 25180 15244 25220
rect 15284 25180 15285 25220
rect 15243 25171 15285 25180
rect 15243 24632 15285 24641
rect 15436 24632 15476 24641
rect 15243 24592 15244 24632
rect 15284 24592 15285 24632
rect 15243 24583 15285 24592
rect 15340 24592 15436 24632
rect 14668 23743 14708 23752
rect 14764 23836 14996 23876
rect 13900 23658 13940 23743
rect 13708 23120 13748 23129
rect 14476 23120 14516 23129
rect 13708 22793 13748 23080
rect 13996 23080 14476 23120
rect 13515 22784 13557 22793
rect 13515 22744 13516 22784
rect 13556 22744 13557 22784
rect 13515 22735 13557 22744
rect 13707 22784 13749 22793
rect 13707 22744 13708 22784
rect 13748 22744 13749 22784
rect 13707 22735 13749 22744
rect 13515 22616 13557 22625
rect 13515 22576 13516 22616
rect 13556 22576 13557 22616
rect 13515 22567 13557 22576
rect 13516 22280 13556 22567
rect 13516 22231 13556 22240
rect 13804 22280 13844 22289
rect 13036 21559 13076 21568
rect 13707 21608 13749 21617
rect 13707 21568 13708 21608
rect 13748 21568 13749 21608
rect 13707 21559 13749 21568
rect 11499 21524 11541 21533
rect 11499 21484 11500 21524
rect 11540 21484 11541 21524
rect 11499 21475 11541 21484
rect 12075 21440 12117 21449
rect 12075 21400 12076 21440
rect 12116 21400 12117 21440
rect 12075 21391 12117 21400
rect 12651 21440 12693 21449
rect 12651 21400 12652 21440
rect 12692 21400 12693 21440
rect 12651 21391 12693 21400
rect 11307 20768 11349 20777
rect 11307 20728 11308 20768
rect 11348 20728 11349 20768
rect 11307 20719 11349 20728
rect 12076 20768 12116 21391
rect 12076 20719 12116 20728
rect 12460 21356 12500 21365
rect 11500 20684 11540 20693
rect 11692 20684 11732 20693
rect 11540 20644 11692 20684
rect 11500 20635 11540 20644
rect 11692 20635 11732 20644
rect 11595 20516 11637 20525
rect 11595 20476 11596 20516
rect 11636 20476 11637 20516
rect 11595 20467 11637 20476
rect 11404 20096 11444 20105
rect 11596 20096 11636 20467
rect 11444 20056 11540 20096
rect 11404 20047 11444 20056
rect 11212 19963 11252 19972
rect 10252 19181 10292 19963
rect 11211 19844 11253 19853
rect 11211 19804 11212 19844
rect 11252 19804 11253 19844
rect 11211 19795 11253 19804
rect 11404 19844 11444 19855
rect 10636 19256 10676 19265
rect 10251 19172 10293 19181
rect 10251 19132 10252 19172
rect 10292 19132 10293 19172
rect 10251 19123 10293 19132
rect 10252 16400 10292 19123
rect 10636 18929 10676 19216
rect 11019 19256 11061 19265
rect 11019 19216 11020 19256
rect 11060 19216 11061 19256
rect 11019 19207 11061 19216
rect 11116 19256 11156 19267
rect 11020 19122 11060 19207
rect 11116 19181 11156 19216
rect 11212 19256 11252 19795
rect 11404 19769 11444 19804
rect 11403 19760 11445 19769
rect 11403 19720 11404 19760
rect 11444 19720 11445 19760
rect 11403 19711 11445 19720
rect 11500 19265 11540 20056
rect 11212 19207 11252 19216
rect 11308 19256 11348 19265
rect 11115 19172 11157 19181
rect 11115 19132 11116 19172
rect 11156 19132 11157 19172
rect 11115 19123 11157 19132
rect 11308 19088 11348 19216
rect 11499 19256 11541 19265
rect 11499 19216 11500 19256
rect 11540 19216 11541 19256
rect 11499 19207 11541 19216
rect 11596 19088 11636 20056
rect 11692 20096 11732 20107
rect 12460 20105 12500 21316
rect 12652 21306 12692 21391
rect 13131 21356 13173 21365
rect 13131 21316 13132 21356
rect 13172 21316 13173 21356
rect 13131 21307 13173 21316
rect 13132 21222 13172 21307
rect 12940 20768 12980 20777
rect 12940 20180 12980 20728
rect 12940 20140 13076 20180
rect 11692 20021 11732 20056
rect 12459 20096 12501 20105
rect 12459 20056 12460 20096
rect 12500 20056 12501 20096
rect 12459 20047 12501 20056
rect 12556 20096 12596 20105
rect 11691 20012 11733 20021
rect 11691 19972 11692 20012
rect 11732 19972 11733 20012
rect 11691 19963 11733 19972
rect 12267 19928 12309 19937
rect 12267 19888 12268 19928
rect 12308 19888 12309 19928
rect 12267 19879 12309 19888
rect 11884 19844 11924 19853
rect 11884 19256 11924 19804
rect 11884 19207 11924 19216
rect 12268 19256 12308 19879
rect 12556 19769 12596 20056
rect 12747 19928 12789 19937
rect 12747 19888 12748 19928
rect 12788 19888 12789 19928
rect 12747 19879 12789 19888
rect 12748 19794 12788 19879
rect 12555 19760 12597 19769
rect 12555 19720 12556 19760
rect 12596 19720 12597 19760
rect 12555 19711 12597 19720
rect 13036 19256 13076 20140
rect 13708 20105 13748 21559
rect 13131 20096 13173 20105
rect 13131 20056 13132 20096
rect 13172 20056 13173 20096
rect 13131 20047 13173 20056
rect 13420 20096 13460 20105
rect 13132 19962 13172 20047
rect 13227 20012 13269 20021
rect 13227 19972 13228 20012
rect 13268 19972 13269 20012
rect 13227 19963 13269 19972
rect 13228 19878 13268 19963
rect 13420 19853 13460 20056
rect 13707 20096 13749 20105
rect 13707 20056 13708 20096
rect 13748 20056 13749 20096
rect 13707 20047 13749 20056
rect 13419 19844 13461 19853
rect 13419 19804 13420 19844
rect 13460 19804 13461 19844
rect 13419 19795 13461 19804
rect 13132 19256 13172 19265
rect 13036 19216 13132 19256
rect 13172 19216 13364 19256
rect 12268 19207 12308 19216
rect 13132 19207 13172 19216
rect 13324 19097 13364 19216
rect 11308 19048 11636 19088
rect 13323 19088 13365 19097
rect 13323 19048 13324 19088
rect 13364 19048 13365 19088
rect 13323 19039 13365 19048
rect 10635 18920 10677 18929
rect 10635 18880 10636 18920
rect 10676 18880 10677 18920
rect 10635 18871 10677 18880
rect 11403 18920 11445 18929
rect 11403 18880 11404 18920
rect 11444 18880 11445 18920
rect 11403 18871 11445 18880
rect 10636 18584 10676 18593
rect 10676 18544 11156 18584
rect 10636 18535 10676 18544
rect 10827 18416 10869 18425
rect 10827 18376 10828 18416
rect 10868 18376 10869 18416
rect 10827 18367 10869 18376
rect 10828 18282 10868 18367
rect 11116 17996 11156 18544
rect 11116 17947 11156 17956
rect 11404 17837 11444 18871
rect 12556 18416 12596 18425
rect 12075 17912 12117 17921
rect 12075 17872 12076 17912
rect 12116 17872 12117 17912
rect 12075 17863 12117 17872
rect 11403 17828 11445 17837
rect 11403 17788 11404 17828
rect 11444 17788 11445 17828
rect 11403 17779 11445 17788
rect 11787 17828 11829 17837
rect 11787 17788 11788 17828
rect 11828 17788 11829 17828
rect 11787 17779 11829 17788
rect 10635 17744 10677 17753
rect 10635 17704 10636 17744
rect 10676 17704 10677 17744
rect 10635 17695 10677 17704
rect 10636 17072 10676 17695
rect 10636 17023 10676 17032
rect 11788 17072 11828 17779
rect 12076 17744 12116 17863
rect 12076 17695 12116 17704
rect 12460 17744 12500 17753
rect 12556 17744 12596 18376
rect 12500 17704 12596 17744
rect 13324 17744 13364 19039
rect 12460 17695 12500 17704
rect 13324 17695 13364 17704
rect 11788 17023 11828 17032
rect 10252 16351 10292 16360
rect 12076 16904 12116 16913
rect 10924 16232 10964 16241
rect 10347 15728 10389 15737
rect 10347 15688 10348 15728
rect 10388 15688 10389 15728
rect 10347 15679 10389 15688
rect 10348 15594 10388 15679
rect 10924 15485 10964 16192
rect 11596 16232 11636 16241
rect 12076 16232 12116 16864
rect 13611 16400 13653 16409
rect 13611 16360 13612 16400
rect 13652 16360 13653 16400
rect 13611 16351 13653 16360
rect 13612 16266 13652 16351
rect 12460 16232 12500 16241
rect 11636 16192 12116 16232
rect 12172 16192 12460 16232
rect 11596 16183 11636 16192
rect 11212 16148 11252 16157
rect 11020 16108 11212 16148
rect 10923 15476 10965 15485
rect 10923 15436 10924 15476
rect 10964 15436 10965 15476
rect 10923 15427 10965 15436
rect 10060 15100 10196 15140
rect 9867 14888 9909 14897
rect 9867 14848 9868 14888
rect 9908 14848 9909 14888
rect 9867 14839 9909 14848
rect 9868 14754 9908 14839
rect 10060 14804 10100 15100
rect 10060 14729 10100 14764
rect 9100 14671 9140 14680
rect 10059 14720 10101 14729
rect 10059 14680 10060 14720
rect 10100 14680 10101 14720
rect 10059 14671 10101 14680
rect 10444 14720 10484 14729
rect 9004 14552 9044 14561
rect 8907 14300 8949 14309
rect 8907 14260 8908 14300
rect 8948 14260 8949 14300
rect 8907 14251 8949 14260
rect 8619 14216 8661 14225
rect 8619 14176 8620 14216
rect 8660 14176 8661 14216
rect 8619 14167 8661 14176
rect 7851 14048 7893 14057
rect 7851 14008 7852 14048
rect 7892 14008 7893 14048
rect 7851 13999 7893 14008
rect 8043 14048 8085 14057
rect 8043 14008 8044 14048
rect 8084 14008 8085 14048
rect 8043 13999 8085 14008
rect 7372 13831 7412 13840
rect 6891 13292 6933 13301
rect 6796 13252 6892 13292
rect 6932 13252 6933 13292
rect 6699 13208 6741 13217
rect 6699 13168 6700 13208
rect 6740 13168 6741 13208
rect 6699 13159 6741 13168
rect 6700 13074 6740 13159
rect 6068 12496 6164 12536
rect 6028 12487 6068 12496
rect 6411 11948 6453 11957
rect 6411 11908 6412 11948
rect 6452 11908 6453 11948
rect 6411 11899 6453 11908
rect 6412 11814 6452 11899
rect 5835 11780 5877 11789
rect 5835 11740 5836 11780
rect 5876 11740 5877 11780
rect 5835 11731 5877 11740
rect 6219 11780 6261 11789
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 5548 11621 5588 11656
rect 5739 11696 5781 11705
rect 5739 11656 5740 11696
rect 5780 11656 5781 11696
rect 5739 11647 5781 11656
rect 5547 11612 5589 11621
rect 5547 11572 5548 11612
rect 5588 11572 5589 11612
rect 5547 11563 5589 11572
rect 4340 11488 4820 11528
rect 5356 11528 5396 11537
rect 5548 11532 5588 11563
rect 4300 11479 4340 11488
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4683 11192 4725 11201
rect 4683 11152 4684 11192
rect 4724 11152 4725 11192
rect 4683 11143 4725 11152
rect 4300 11024 4340 11033
rect 4108 10984 4300 11024
rect 4300 10975 4340 10984
rect 4107 10856 4149 10865
rect 4107 10816 4108 10856
rect 4148 10816 4149 10856
rect 4107 10807 4149 10816
rect 4108 10722 4148 10807
rect 3723 10436 3765 10445
rect 4203 10436 4245 10445
rect 3723 10396 3724 10436
rect 3764 10396 3860 10436
rect 3723 10387 3765 10396
rect 3532 8884 3668 8924
rect 3532 8681 3572 8884
rect 3724 8849 3764 8934
rect 3723 8840 3765 8849
rect 3723 8800 3724 8840
rect 3764 8800 3765 8840
rect 3723 8791 3765 8800
rect 3627 8756 3669 8765
rect 3627 8716 3628 8756
rect 3668 8716 3669 8756
rect 3627 8707 3669 8716
rect 3436 8672 3476 8681
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 3436 8093 3476 8632
rect 3531 8672 3573 8681
rect 3531 8632 3532 8672
rect 3572 8632 3573 8672
rect 3531 8623 3573 8632
rect 3531 8504 3573 8513
rect 3531 8464 3532 8504
rect 3572 8464 3573 8504
rect 3531 8455 3573 8464
rect 3435 8084 3477 8093
rect 3435 8044 3436 8084
rect 3476 8044 3477 8084
rect 3435 8035 3477 8044
rect 2476 8000 2516 8009
rect 2476 7841 2516 7960
rect 2859 8000 2901 8009
rect 2859 7960 2860 8000
rect 2900 7960 2901 8000
rect 2859 7951 2901 7960
rect 3532 8000 3572 8455
rect 3628 8168 3668 8707
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3820 8672 3860 10396
rect 4203 10396 4204 10436
rect 4244 10396 4245 10436
rect 4203 10387 4245 10396
rect 4204 10302 4244 10387
rect 3915 10268 3957 10277
rect 3915 10228 3916 10268
rect 3956 10228 3957 10268
rect 3915 10219 3957 10228
rect 3916 10134 3956 10219
rect 4684 10109 4724 11143
rect 5259 11024 5301 11033
rect 5259 10984 5260 11024
rect 5300 10984 5301 11024
rect 5259 10975 5301 10984
rect 5260 10890 5300 10975
rect 4972 10772 5012 10781
rect 4779 10688 4821 10697
rect 4779 10648 4780 10688
rect 4820 10648 4821 10688
rect 4779 10639 4821 10648
rect 4683 10100 4725 10109
rect 4683 10060 4684 10100
rect 4724 10060 4725 10100
rect 4683 10051 4725 10060
rect 3915 10016 3957 10025
rect 3915 9976 3916 10016
rect 3956 9976 3957 10016
rect 3915 9967 3957 9976
rect 3916 8924 3956 9967
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4204 9521 4244 9606
rect 4203 9512 4245 9521
rect 4203 9472 4204 9512
rect 4244 9472 4245 9512
rect 4203 9463 4245 9472
rect 4300 9512 4340 9523
rect 4300 9437 4340 9472
rect 4588 9512 4628 9523
rect 4588 9437 4628 9472
rect 4780 9512 4820 10639
rect 4875 10268 4917 10277
rect 4875 10228 4876 10268
rect 4916 10228 4917 10268
rect 4875 10219 4917 10228
rect 4876 10184 4916 10219
rect 4972 10193 5012 10732
rect 5356 10697 5396 11488
rect 5547 11192 5589 11201
rect 5547 11152 5548 11192
rect 5588 11152 5589 11192
rect 5547 11143 5589 11152
rect 5548 11058 5588 11143
rect 5740 11024 5780 11647
rect 5740 10975 5780 10984
rect 5836 11024 5876 11731
rect 6220 11646 6260 11731
rect 6603 11696 6645 11705
rect 6603 11656 6604 11696
rect 6644 11656 6645 11696
rect 6603 11647 6645 11656
rect 6604 11562 6644 11647
rect 6027 11528 6069 11537
rect 6027 11488 6028 11528
rect 6068 11488 6069 11528
rect 6027 11479 6069 11488
rect 6699 11528 6741 11537
rect 6796 11528 6836 13252
rect 6891 13243 6933 13252
rect 7852 13208 7892 13999
rect 8044 13914 8084 13999
rect 7852 13159 7892 13168
rect 8043 13208 8085 13217
rect 8043 13168 8044 13208
rect 8084 13168 8085 13208
rect 8043 13159 8085 13168
rect 7372 13040 7412 13049
rect 6699 11488 6700 11528
rect 6740 11488 6836 11528
rect 6892 12536 6932 12545
rect 6699 11479 6741 11488
rect 5932 11117 5972 11148
rect 5931 11108 5973 11117
rect 5931 11068 5932 11108
rect 5972 11068 5973 11108
rect 5931 11059 5973 11068
rect 5451 10856 5493 10865
rect 5451 10816 5452 10856
rect 5492 10816 5493 10856
rect 5451 10807 5493 10816
rect 5355 10688 5397 10697
rect 5355 10648 5356 10688
rect 5396 10648 5397 10688
rect 5355 10639 5397 10648
rect 4876 10133 4916 10144
rect 4971 10184 5013 10193
rect 4971 10144 4972 10184
rect 5012 10144 5013 10184
rect 4971 10135 5013 10144
rect 5068 10184 5108 10193
rect 4875 10016 4917 10025
rect 4875 9976 4876 10016
rect 4916 9976 4917 10016
rect 4875 9967 4917 9976
rect 4780 9463 4820 9472
rect 4876 9512 4916 9967
rect 5068 9680 5108 10144
rect 5355 10184 5397 10193
rect 5355 10144 5356 10184
rect 5396 10144 5397 10184
rect 5355 10135 5397 10144
rect 5452 10184 5492 10807
rect 5452 10135 5492 10144
rect 5068 9631 5108 9640
rect 4876 9463 4916 9472
rect 5259 9512 5301 9521
rect 5259 9472 5260 9512
rect 5300 9472 5301 9512
rect 5259 9463 5301 9472
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 4299 9379 4341 9388
rect 4587 9428 4629 9437
rect 4587 9388 4588 9428
rect 4628 9388 4629 9428
rect 4587 9379 4629 9388
rect 4012 9344 4052 9353
rect 4875 9344 4917 9353
rect 4052 9304 4244 9344
rect 4012 9295 4052 9304
rect 4011 8924 4053 8933
rect 3916 8884 4012 8924
rect 4052 8884 4053 8924
rect 4011 8875 4053 8884
rect 3916 8672 3956 8681
rect 3820 8632 3916 8672
rect 3723 8623 3765 8632
rect 3916 8623 3956 8632
rect 3724 8538 3764 8623
rect 4012 8504 4052 8875
rect 4107 8840 4149 8849
rect 4107 8800 4108 8840
rect 4148 8800 4149 8840
rect 4107 8791 4149 8800
rect 4108 8672 4148 8791
rect 4204 8672 4244 9304
rect 4875 9304 4876 9344
rect 4916 9304 4917 9344
rect 4875 9295 4917 9304
rect 4876 9210 4916 9295
rect 4971 8756 5013 8765
rect 4971 8716 4972 8756
rect 5012 8716 5013 8756
rect 4971 8707 5013 8716
rect 4492 8672 4532 8681
rect 4204 8632 4492 8672
rect 4108 8623 4148 8632
rect 4492 8623 4532 8632
rect 3820 8464 4052 8504
rect 3724 8168 3764 8177
rect 3628 8128 3724 8168
rect 3724 8119 3764 8128
rect 2475 7832 2517 7841
rect 2475 7792 2476 7832
rect 2516 7792 2517 7832
rect 2475 7783 2517 7792
rect 2860 7757 2900 7951
rect 2859 7748 2901 7757
rect 2859 7708 2860 7748
rect 2900 7708 2901 7748
rect 2859 7699 2901 7708
rect 2860 7614 2900 7699
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 2763 7328 2805 7337
rect 2763 7288 2764 7328
rect 2804 7288 2805 7328
rect 2763 7279 2805 7288
rect 2132 7120 2324 7160
rect 2092 7111 2132 7120
rect 2188 6488 2228 6497
rect 1996 6448 2188 6488
rect 2188 6439 2228 6448
rect 2380 6488 2420 6497
rect 2284 6404 2324 6413
rect 2380 6404 2420 6448
rect 2764 6488 2804 7279
rect 3340 7160 3380 7169
rect 3532 7160 3572 7960
rect 3627 7748 3669 7757
rect 3627 7708 3628 7748
rect 3668 7708 3669 7748
rect 3627 7699 3669 7708
rect 3724 7748 3764 7757
rect 3380 7120 3572 7160
rect 3340 7111 3380 7120
rect 3531 6992 3573 7001
rect 3531 6952 3532 6992
rect 3572 6952 3573 6992
rect 3628 6992 3668 7699
rect 3724 7160 3764 7708
rect 3724 7111 3764 7120
rect 3820 7160 3860 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4876 8168 4916 8177
rect 4395 8084 4437 8093
rect 4395 8044 4396 8084
rect 4436 8044 4437 8084
rect 4395 8035 4437 8044
rect 4396 8000 4436 8035
rect 4876 8009 4916 8128
rect 4972 8093 5012 8707
rect 5067 8420 5109 8429
rect 5067 8380 5068 8420
rect 5108 8380 5109 8420
rect 5067 8371 5109 8380
rect 4971 8084 5013 8093
rect 4971 8044 4972 8084
rect 5012 8044 5013 8084
rect 4971 8035 5013 8044
rect 4684 8000 4724 8009
rect 4396 7949 4436 7960
rect 4588 7960 4684 8000
rect 4011 7328 4053 7337
rect 3820 7111 3860 7120
rect 3916 7288 4012 7328
rect 4052 7288 4053 7328
rect 3724 6992 3764 7001
rect 3628 6952 3724 6992
rect 3531 6943 3573 6952
rect 3724 6943 3764 6952
rect 2764 6439 2804 6448
rect 2859 6488 2901 6497
rect 2859 6448 2860 6488
rect 2900 6448 2901 6488
rect 2859 6439 2901 6448
rect 2572 6404 2612 6413
rect 2380 6364 2572 6404
rect 2284 6320 2324 6364
rect 2572 6355 2612 6364
rect 2860 6354 2900 6439
rect 1324 6271 1364 6280
rect 1708 6280 2324 6320
rect 1035 5648 1077 5657
rect 1035 5608 1036 5648
rect 1076 5608 1077 5648
rect 1035 5599 1077 5608
rect 652 5431 692 5440
rect 1036 5480 1076 5599
rect 1036 5431 1076 5440
rect 652 5144 692 5153
rect 652 4817 692 5104
rect 1708 4976 1748 6280
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 2284 5816 2324 5825
rect 1708 4927 1748 4936
rect 2092 5776 2284 5816
rect 2092 4976 2132 5776
rect 2284 5767 2324 5776
rect 3532 5648 3572 6943
rect 3628 6488 3668 6497
rect 3628 5732 3668 6448
rect 3628 5683 3668 5692
rect 3532 5599 3572 5608
rect 3724 5648 3764 5657
rect 3724 5069 3764 5608
rect 3916 5648 3956 7288
rect 4011 7279 4053 7288
rect 4012 7194 4052 7279
rect 4588 7001 4628 7960
rect 4684 7951 4724 7960
rect 4875 8000 4917 8009
rect 4875 7960 4876 8000
rect 4916 7960 4917 8000
rect 4875 7951 4917 7960
rect 5068 8000 5108 8371
rect 5068 7951 5108 7960
rect 5260 7925 5300 9463
rect 5356 8672 5396 10135
rect 5836 10025 5876 10984
rect 5932 11024 5972 11059
rect 5932 10697 5972 10984
rect 6028 11024 6068 11479
rect 6700 11394 6740 11479
rect 6028 10975 6068 10984
rect 6316 10772 6356 10783
rect 6316 10697 6356 10732
rect 5931 10688 5973 10697
rect 5931 10648 5932 10688
rect 5972 10648 5973 10688
rect 5931 10639 5973 10648
rect 6315 10688 6357 10697
rect 6315 10648 6316 10688
rect 6356 10648 6357 10688
rect 6315 10639 6357 10648
rect 6892 10193 6932 12496
rect 7083 11948 7125 11957
rect 7083 11908 7084 11948
rect 7124 11908 7125 11948
rect 7083 11899 7125 11908
rect 6988 11024 7028 11033
rect 6988 10445 7028 10984
rect 6987 10436 7029 10445
rect 6987 10396 6988 10436
rect 7028 10396 7029 10436
rect 6987 10387 7029 10396
rect 6315 10184 6357 10193
rect 6315 10144 6316 10184
rect 6356 10144 6357 10184
rect 6315 10135 6357 10144
rect 6891 10184 6933 10193
rect 6891 10144 6892 10184
rect 6932 10144 6933 10184
rect 6891 10135 6933 10144
rect 6316 10050 6356 10135
rect 5835 10016 5877 10025
rect 5835 9976 5836 10016
rect 5876 9976 5877 10016
rect 5835 9967 5877 9976
rect 7084 9680 7124 11899
rect 7372 11033 7412 13000
rect 8044 12536 8084 13159
rect 8140 13040 8180 13049
rect 8140 12545 8180 13000
rect 8044 11873 8084 12496
rect 8139 12536 8181 12545
rect 8524 12536 8564 12545
rect 8139 12496 8140 12536
rect 8180 12496 8181 12536
rect 8139 12487 8181 12496
rect 8428 12496 8524 12536
rect 8043 11864 8085 11873
rect 8043 11824 8044 11864
rect 8084 11824 8085 11864
rect 8043 11815 8085 11824
rect 7948 11696 7988 11705
rect 7564 11656 7948 11696
rect 7371 11024 7413 11033
rect 7371 10984 7372 11024
rect 7412 10984 7413 11024
rect 7371 10975 7413 10984
rect 7084 9631 7124 9640
rect 7179 9680 7221 9689
rect 7179 9640 7180 9680
rect 7220 9640 7221 9680
rect 7179 9631 7221 9640
rect 5740 9512 5780 9521
rect 5932 9512 5972 9521
rect 5740 9353 5780 9472
rect 5836 9472 5932 9512
rect 5739 9344 5781 9353
rect 5739 9304 5740 9344
rect 5780 9304 5781 9344
rect 5739 9295 5781 9304
rect 5356 8623 5396 8632
rect 5548 8168 5588 8177
rect 5836 8168 5876 9472
rect 5932 9463 5972 9472
rect 6124 9512 6164 9523
rect 6124 9437 6164 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7180 9512 7220 9631
rect 7180 9463 7220 9472
rect 7276 9512 7316 9521
rect 6123 9428 6165 9437
rect 6123 9388 6124 9428
rect 6164 9388 6165 9428
rect 6123 9379 6165 9388
rect 6988 9378 7028 9463
rect 7276 9353 7316 9472
rect 7275 9344 7317 9353
rect 7275 9304 7276 9344
rect 7316 9304 7317 9344
rect 7275 9295 7317 9304
rect 5932 9260 5972 9269
rect 5932 8849 5972 9220
rect 7372 9185 7412 10975
rect 7467 10436 7509 10445
rect 7467 10396 7468 10436
rect 7508 10396 7509 10436
rect 7467 10387 7509 10396
rect 7468 10302 7508 10387
rect 7564 10361 7604 11656
rect 7948 11647 7988 11656
rect 8236 11696 8276 11705
rect 8428 11696 8468 12496
rect 8524 12487 8564 12496
rect 8620 12536 8660 14167
rect 9004 14141 9044 14512
rect 9771 14216 9813 14225
rect 9771 14176 9772 14216
rect 9812 14176 9813 14216
rect 9771 14167 9813 14176
rect 9003 14132 9045 14141
rect 9003 14092 9004 14132
rect 9044 14092 9045 14132
rect 9003 14083 9045 14092
rect 9772 14082 9812 14167
rect 8811 13880 8853 13889
rect 8811 13840 8812 13880
rect 8852 13840 8853 13880
rect 8811 13831 8853 13840
rect 8812 13746 8852 13831
rect 10060 13217 10100 14671
rect 10444 14225 10484 14680
rect 10923 14720 10965 14729
rect 10923 14680 10924 14720
rect 10964 14680 10965 14720
rect 10923 14671 10965 14680
rect 10443 14216 10485 14225
rect 10443 14176 10444 14216
rect 10484 14176 10485 14216
rect 10443 14167 10485 14176
rect 10924 14048 10964 14671
rect 10924 13999 10964 14008
rect 10155 13880 10197 13889
rect 10155 13840 10156 13880
rect 10196 13840 10197 13880
rect 10155 13831 10197 13840
rect 9291 13208 9333 13217
rect 9291 13168 9292 13208
rect 9332 13168 9333 13208
rect 9291 13159 9333 13168
rect 10059 13208 10101 13217
rect 10059 13168 10060 13208
rect 10100 13168 10101 13208
rect 10059 13159 10101 13168
rect 10156 13208 10196 13831
rect 10156 13159 10196 13168
rect 9292 13074 9332 13159
rect 10540 13124 10580 13133
rect 10732 13124 10772 13133
rect 10580 13084 10732 13124
rect 10540 13075 10580 13084
rect 10732 13075 10772 13084
rect 10251 13040 10293 13049
rect 10251 13000 10252 13040
rect 10292 13000 10293 13040
rect 10251 12991 10293 13000
rect 8907 12956 8949 12965
rect 8907 12916 8908 12956
rect 8948 12916 8949 12956
rect 8907 12907 8949 12916
rect 8812 12704 8852 12713
rect 8660 12496 8756 12536
rect 8620 12487 8660 12496
rect 8276 11656 8372 11696
rect 8236 11647 8276 11656
rect 8043 11612 8085 11621
rect 8043 11572 8044 11612
rect 8084 11572 8085 11612
rect 8043 11563 8085 11572
rect 7947 11528 7989 11537
rect 7947 11488 7948 11528
rect 7988 11488 7989 11528
rect 7947 11479 7989 11488
rect 7851 11192 7893 11201
rect 7851 11152 7852 11192
rect 7892 11152 7893 11192
rect 7851 11143 7893 11152
rect 7755 11108 7797 11117
rect 7755 11068 7756 11108
rect 7796 11068 7797 11108
rect 7755 11059 7797 11068
rect 7660 11024 7700 11033
rect 7563 10352 7605 10361
rect 7563 10312 7564 10352
rect 7604 10312 7605 10352
rect 7563 10303 7605 10312
rect 7660 10277 7700 10984
rect 7756 11024 7796 11059
rect 7756 10973 7796 10984
rect 7852 11024 7892 11143
rect 7852 10975 7892 10984
rect 7948 11024 7988 11479
rect 7948 10975 7988 10984
rect 8044 10856 8084 11563
rect 8140 11528 8180 11537
rect 8140 11444 8180 11488
rect 8235 11444 8277 11453
rect 8140 11404 8236 11444
rect 8276 11404 8277 11444
rect 8235 11395 8277 11404
rect 8332 11285 8372 11656
rect 8428 11621 8468 11656
rect 8619 11696 8661 11705
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 8716 11696 8756 12496
rect 8812 11789 8852 12664
rect 8908 12284 8948 12907
rect 10155 12872 10197 12881
rect 10155 12832 10156 12872
rect 10196 12832 10197 12872
rect 10155 12823 10197 12832
rect 9003 12536 9045 12545
rect 9675 12536 9717 12545
rect 9868 12536 9908 12545
rect 9003 12496 9004 12536
rect 9044 12496 9140 12536
rect 9003 12487 9045 12496
rect 9004 12402 9044 12487
rect 8908 12244 9044 12284
rect 8907 11864 8949 11873
rect 8907 11824 8908 11864
rect 8948 11824 8949 11864
rect 8907 11815 8949 11824
rect 8811 11780 8853 11789
rect 8811 11740 8812 11780
rect 8852 11740 8853 11780
rect 8811 11731 8853 11740
rect 8716 11647 8756 11656
rect 8908 11696 8948 11815
rect 8427 11612 8469 11621
rect 8427 11572 8428 11612
rect 8468 11572 8469 11612
rect 8427 11563 8469 11572
rect 8620 11562 8660 11647
rect 8908 11612 8948 11656
rect 9004 11696 9044 12244
rect 9004 11647 9044 11656
rect 8812 11572 8948 11612
rect 8331 11276 8373 11285
rect 8331 11236 8332 11276
rect 8372 11236 8373 11276
rect 8331 11227 8373 11236
rect 8715 11276 8757 11285
rect 8715 11236 8716 11276
rect 8756 11236 8757 11276
rect 8715 11227 8757 11236
rect 8140 11033 8180 11118
rect 8139 11024 8181 11033
rect 8139 10984 8140 11024
rect 8180 10984 8181 11024
rect 8139 10975 8181 10984
rect 8428 11024 8468 11033
rect 8620 11024 8660 11033
rect 8468 10984 8620 11024
rect 8428 10975 8468 10984
rect 8427 10856 8469 10865
rect 8044 10816 8372 10856
rect 8236 10352 8276 10361
rect 7659 10268 7701 10277
rect 7659 10228 7660 10268
rect 7700 10228 7701 10268
rect 7659 10219 7701 10228
rect 8236 10193 8276 10312
rect 8332 10268 8372 10816
rect 8427 10816 8428 10856
rect 8468 10816 8469 10856
rect 8427 10807 8469 10816
rect 8428 10722 8468 10807
rect 8620 10445 8660 10984
rect 8427 10436 8469 10445
rect 8427 10396 8428 10436
rect 8468 10396 8469 10436
rect 8427 10387 8469 10396
rect 8619 10436 8661 10445
rect 8619 10396 8620 10436
rect 8660 10396 8661 10436
rect 8619 10387 8661 10396
rect 8332 10219 8372 10228
rect 8235 10184 8277 10193
rect 8235 10144 8236 10184
rect 8276 10144 8277 10184
rect 8235 10135 8277 10144
rect 8428 10184 8468 10387
rect 8523 10352 8565 10361
rect 8523 10312 8524 10352
rect 8564 10312 8565 10352
rect 8523 10303 8565 10312
rect 8428 10135 8468 10144
rect 8524 10184 8564 10303
rect 8716 10193 8756 11227
rect 8524 10135 8564 10144
rect 8715 10184 8757 10193
rect 8715 10144 8716 10184
rect 8756 10144 8757 10184
rect 8715 10135 8757 10144
rect 8812 10109 8852 11572
rect 9100 11528 9140 12496
rect 9675 12496 9676 12536
rect 9716 12496 9717 12536
rect 9675 12487 9717 12496
rect 9772 12496 9868 12536
rect 9676 12402 9716 12487
rect 9772 11957 9812 12496
rect 9868 12487 9908 12496
rect 9867 12368 9909 12377
rect 9867 12328 9868 12368
rect 9908 12328 9909 12368
rect 9867 12319 9909 12328
rect 9771 11948 9813 11957
rect 9771 11908 9772 11948
rect 9812 11908 9813 11948
rect 9771 11899 9813 11908
rect 9675 11780 9717 11789
rect 9675 11740 9676 11780
rect 9716 11740 9717 11780
rect 9675 11731 9717 11740
rect 9387 11696 9429 11705
rect 9387 11656 9388 11696
rect 9428 11656 9429 11696
rect 9387 11647 9429 11656
rect 9580 11696 9620 11705
rect 9388 11562 9428 11647
rect 9484 11537 9524 11622
rect 8908 11488 9140 11528
rect 9196 11528 9236 11537
rect 8908 11033 8948 11488
rect 9196 11369 9236 11488
rect 9483 11528 9525 11537
rect 9483 11488 9484 11528
rect 9524 11488 9525 11528
rect 9483 11479 9525 11488
rect 9195 11360 9237 11369
rect 9195 11320 9196 11360
rect 9236 11320 9237 11360
rect 9195 11311 9237 11320
rect 9387 11360 9429 11369
rect 9387 11320 9388 11360
rect 9428 11320 9429 11360
rect 9387 11311 9429 11320
rect 9100 11201 9140 11286
rect 9099 11192 9141 11201
rect 9099 11152 9100 11192
rect 9140 11152 9141 11192
rect 9099 11143 9141 11152
rect 8907 11024 8949 11033
rect 9291 11024 9333 11033
rect 8907 10984 8908 11024
rect 8948 10984 8949 11024
rect 8907 10975 8949 10984
rect 9004 10984 9292 11024
rect 9332 10984 9333 11024
rect 8908 10890 8948 10975
rect 8908 10772 8948 10781
rect 9004 10772 9044 10984
rect 9291 10975 9333 10984
rect 9388 11024 9428 11311
rect 9580 11285 9620 11656
rect 9676 11696 9716 11731
rect 9676 11645 9716 11656
rect 9868 11696 9908 12319
rect 10156 11948 10196 12823
rect 10156 11899 10196 11908
rect 10155 11780 10197 11789
rect 10155 11740 10156 11780
rect 10196 11740 10197 11780
rect 10155 11731 10197 11740
rect 9868 11360 9908 11656
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10156 11696 10196 11731
rect 9964 11562 10004 11647
rect 10156 11645 10196 11656
rect 9963 11444 10005 11453
rect 9963 11404 9964 11444
rect 10004 11404 10005 11444
rect 9963 11395 10005 11404
rect 9772 11320 9908 11360
rect 9579 11276 9621 11285
rect 9579 11236 9580 11276
rect 9620 11236 9621 11276
rect 9579 11227 9621 11236
rect 9676 11024 9716 11033
rect 9388 10975 9428 10984
rect 9484 10982 9524 10991
rect 9292 10890 9332 10975
rect 8948 10732 9044 10772
rect 9387 10772 9429 10781
rect 9387 10732 9388 10772
rect 9428 10732 9429 10772
rect 8908 10723 8948 10732
rect 9387 10723 9429 10732
rect 9291 10688 9333 10697
rect 9291 10648 9292 10688
rect 9332 10648 9333 10688
rect 9291 10639 9333 10648
rect 8907 10436 8949 10445
rect 8907 10396 8908 10436
rect 8948 10396 8949 10436
rect 8907 10387 8949 10396
rect 8811 10100 8853 10109
rect 8811 10060 8812 10100
rect 8852 10060 8853 10100
rect 8811 10051 8853 10060
rect 8428 10016 8468 10025
rect 7948 9976 8428 10016
rect 7659 9596 7701 9605
rect 7659 9556 7660 9596
rect 7700 9556 7701 9596
rect 7659 9547 7701 9556
rect 7468 9512 7508 9521
rect 7371 9176 7413 9185
rect 7371 9136 7372 9176
rect 7412 9136 7413 9176
rect 7371 9127 7413 9136
rect 5931 8840 5973 8849
rect 7468 8840 7508 9472
rect 7564 9512 7604 9521
rect 7564 9344 7604 9472
rect 7660 9438 7700 9547
rect 7660 9389 7700 9398
rect 7756 9344 7796 9353
rect 7564 9304 7700 9344
rect 7563 9176 7605 9185
rect 7563 9136 7564 9176
rect 7604 9136 7605 9176
rect 7563 9127 7605 9136
rect 5931 8800 5932 8840
rect 5972 8800 5973 8840
rect 5931 8791 5973 8800
rect 7372 8800 7508 8840
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6604 8538 6644 8623
rect 6796 8504 6836 8515
rect 6796 8429 6836 8464
rect 6795 8420 6837 8429
rect 6795 8380 6796 8420
rect 6836 8380 6837 8420
rect 6795 8371 6837 8380
rect 6027 8336 6069 8345
rect 6027 8296 6028 8336
rect 6068 8296 6069 8336
rect 6027 8287 6069 8296
rect 5588 8128 5876 8168
rect 5548 8119 5588 8128
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5835 8000 5877 8009
rect 5835 7960 5836 8000
rect 5876 7960 5877 8000
rect 5835 7951 5877 7960
rect 6028 8000 6068 8287
rect 5259 7916 5301 7925
rect 5259 7876 5260 7916
rect 5300 7876 5301 7916
rect 5259 7867 5301 7876
rect 4684 7832 4724 7841
rect 4724 7792 5012 7832
rect 4684 7783 4724 7792
rect 4876 7160 4916 7169
rect 4972 7160 5012 7792
rect 5068 7160 5108 7169
rect 4972 7120 5068 7160
rect 4203 6992 4245 7001
rect 4203 6952 4204 6992
rect 4244 6952 4245 6992
rect 4203 6943 4245 6952
rect 4587 6992 4629 7001
rect 4587 6952 4588 6992
rect 4628 6952 4629 6992
rect 4587 6943 4629 6952
rect 4204 6858 4244 6943
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 4011 6488 4053 6497
rect 4011 6448 4012 6488
rect 4052 6448 4053 6488
rect 4011 6439 4053 6448
rect 4491 6488 4533 6497
rect 4491 6448 4492 6488
rect 4532 6448 4533 6488
rect 4491 6439 4533 6448
rect 3916 5144 3956 5608
rect 4012 5648 4052 6439
rect 4492 6354 4532 6439
rect 4203 6320 4245 6329
rect 4203 6280 4204 6320
rect 4244 6280 4245 6320
rect 4203 6271 4245 6280
rect 4012 5599 4052 5608
rect 4204 5648 4244 6271
rect 4300 6236 4340 6245
rect 4300 5648 4340 6196
rect 4396 5648 4436 5657
rect 4300 5608 4396 5648
rect 4204 5599 4244 5608
rect 4396 5599 4436 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 4780 5514 4820 5599
rect 4203 5480 4245 5489
rect 4203 5440 4204 5480
rect 4244 5440 4245 5480
rect 4203 5431 4245 5440
rect 4204 5346 4244 5431
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4683 5144 4725 5153
rect 4876 5144 4916 7120
rect 4971 6320 5013 6329
rect 4971 6280 4972 6320
rect 5012 6280 5013 6320
rect 4971 6271 5013 6280
rect 3916 5104 4628 5144
rect 3723 5060 3765 5069
rect 3723 5020 3724 5060
rect 3764 5020 3765 5060
rect 3723 5011 3765 5020
rect 2092 4927 2132 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 4204 4976 4244 4987
rect 2956 4842 2996 4927
rect 4204 4901 4244 4936
rect 4588 4976 4628 5104
rect 4683 5104 4684 5144
rect 4724 5104 4725 5144
rect 4683 5095 4725 5104
rect 4780 5104 4916 5144
rect 4588 4927 4628 4936
rect 4684 4976 4724 5095
rect 4780 5060 4820 5104
rect 4780 5011 4820 5020
rect 4684 4901 4724 4936
rect 4876 4976 4916 4985
rect 4972 4976 5012 6271
rect 5068 5489 5108 7120
rect 5164 6488 5204 6499
rect 5164 6413 5204 6448
rect 5163 6404 5205 6413
rect 5163 6364 5164 6404
rect 5204 6364 5205 6404
rect 5163 6355 5205 6364
rect 5067 5480 5109 5489
rect 5067 5440 5068 5480
rect 5108 5440 5109 5480
rect 5067 5431 5109 5440
rect 4916 4936 5012 4976
rect 5068 4976 5108 5431
rect 5164 5237 5204 6355
rect 5163 5228 5205 5237
rect 5163 5188 5164 5228
rect 5204 5188 5205 5228
rect 5163 5179 5205 5188
rect 5163 5060 5205 5069
rect 5163 5020 5164 5060
rect 5204 5020 5205 5060
rect 5163 5011 5205 5020
rect 4876 4927 4916 4936
rect 5068 4927 5108 4936
rect 5164 4926 5204 5011
rect 5260 4976 5300 7867
rect 5356 7866 5396 7951
rect 5836 7866 5876 7951
rect 6028 7925 6068 7960
rect 6027 7916 6069 7925
rect 6027 7876 6028 7916
rect 6068 7876 6069 7916
rect 6027 7867 6069 7876
rect 6412 7832 6452 7841
rect 5932 7748 5972 7757
rect 5836 7708 5932 7748
rect 5740 6992 5780 7001
rect 5452 6952 5740 6992
rect 5452 6488 5492 6952
rect 5740 6943 5780 6952
rect 5547 6824 5589 6833
rect 5547 6784 5548 6824
rect 5588 6784 5589 6824
rect 5547 6775 5589 6784
rect 5452 6439 5492 6448
rect 5548 6488 5588 6775
rect 5548 6439 5588 6448
rect 5740 6488 5780 6497
rect 5836 6488 5876 7708
rect 5932 7699 5972 7708
rect 6316 7160 6356 7169
rect 6412 7160 6452 7792
rect 7084 7748 7124 7757
rect 7084 7160 7124 7708
rect 7180 7160 7220 7169
rect 6356 7120 6452 7160
rect 6988 7120 7180 7160
rect 6316 7111 6356 7120
rect 5780 6448 5876 6488
rect 5932 7076 5972 7085
rect 5740 6439 5780 6448
rect 5932 6404 5972 7036
rect 6027 6992 6069 7001
rect 6027 6952 6028 6992
rect 6068 6952 6069 6992
rect 6027 6943 6069 6952
rect 5836 6364 5972 6404
rect 5740 6320 5780 6329
rect 5836 6320 5876 6364
rect 6028 6329 6068 6943
rect 6604 6488 6644 6497
rect 6796 6488 6836 6497
rect 6988 6488 7028 7120
rect 7180 7111 7220 7120
rect 6604 6329 6644 6448
rect 6700 6448 6796 6488
rect 6836 6448 7028 6488
rect 7083 6488 7125 6497
rect 7083 6448 7084 6488
rect 7124 6448 7125 6488
rect 6027 6320 6069 6329
rect 5780 6280 5876 6320
rect 5932 6280 6028 6320
rect 6068 6280 6069 6320
rect 5740 6271 5780 6280
rect 5932 6236 5972 6280
rect 6027 6271 6069 6280
rect 6603 6320 6645 6329
rect 6603 6280 6604 6320
rect 6644 6280 6645 6320
rect 6603 6271 6645 6280
rect 5932 6187 5972 6196
rect 6028 6186 6068 6271
rect 5451 5648 5493 5657
rect 5644 5648 5684 5657
rect 5451 5608 5452 5648
rect 5492 5608 5493 5648
rect 5451 5599 5493 5608
rect 5548 5608 5644 5648
rect 5260 4927 5300 4936
rect 4203 4892 4245 4901
rect 4203 4852 4204 4892
rect 4244 4852 4245 4892
rect 4203 4843 4245 4852
rect 4683 4892 4725 4901
rect 4683 4852 4684 4892
rect 4724 4852 4725 4892
rect 4683 4843 4725 4852
rect 651 4808 693 4817
rect 4684 4812 4724 4843
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 5452 4808 5492 5599
rect 5548 4985 5588 5608
rect 5644 5599 5684 5608
rect 5547 4976 5589 4985
rect 5547 4936 5548 4976
rect 5588 4936 5589 4976
rect 5547 4927 5589 4936
rect 6603 4976 6645 4985
rect 6603 4936 6604 4976
rect 6644 4936 6645 4976
rect 6603 4927 6645 4936
rect 5452 4759 5492 4768
rect 4299 4724 4341 4733
rect 4299 4684 4300 4724
rect 4340 4684 4341 4724
rect 4299 4675 4341 4684
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4300 4136 4340 4675
rect 5548 4145 5588 4927
rect 6604 4842 6644 4927
rect 5931 4724 5973 4733
rect 5931 4684 5932 4724
rect 5972 4684 5973 4724
rect 5931 4675 5973 4684
rect 5932 4590 5972 4675
rect 4300 4087 4340 4096
rect 4684 4136 4724 4145
rect 5547 4136 5589 4145
rect 4724 4096 4820 4136
rect 4684 4087 4724 4096
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 652 3632 692 3641
rect 652 3137 692 3592
rect 4780 3296 4820 4096
rect 5547 4096 5548 4136
rect 5588 4096 5589 4136
rect 5547 4087 5589 4096
rect 6603 4136 6645 4145
rect 6700 4136 6740 6448
rect 6796 6439 6836 6448
rect 7083 6439 7125 6448
rect 7276 6488 7316 6497
rect 7084 6354 7124 6439
rect 6795 6320 6837 6329
rect 6795 6280 6796 6320
rect 6836 6280 6837 6320
rect 6795 6271 6837 6280
rect 6796 5900 6836 6271
rect 7179 6236 7221 6245
rect 7179 6196 7180 6236
rect 7220 6196 7221 6236
rect 7179 6187 7221 6196
rect 7180 6102 7220 6187
rect 6796 5851 6836 5860
rect 7179 5480 7221 5489
rect 7276 5480 7316 6448
rect 7372 6329 7412 8800
rect 7467 8672 7509 8681
rect 7467 8632 7468 8672
rect 7508 8632 7509 8672
rect 7467 8623 7509 8632
rect 7468 8177 7508 8623
rect 7467 8168 7509 8177
rect 7467 8128 7468 8168
rect 7508 8128 7509 8168
rect 7467 8119 7509 8128
rect 7467 8000 7509 8009
rect 7467 7960 7468 8000
rect 7508 7960 7509 8000
rect 7467 7951 7509 7960
rect 7564 8000 7604 9127
rect 7660 9008 7700 9304
rect 7756 9185 7796 9304
rect 7852 9269 7892 9354
rect 7851 9260 7893 9269
rect 7851 9220 7852 9260
rect 7892 9220 7893 9260
rect 7851 9211 7893 9220
rect 7755 9176 7797 9185
rect 7755 9136 7756 9176
rect 7796 9136 7797 9176
rect 7755 9127 7797 9136
rect 7660 8968 7892 9008
rect 7659 8840 7701 8849
rect 7659 8800 7660 8840
rect 7700 8800 7701 8840
rect 7659 8791 7701 8800
rect 7660 8672 7700 8791
rect 7660 8623 7700 8632
rect 7756 8672 7796 8681
rect 7564 7951 7604 7960
rect 7468 6740 7508 7951
rect 7756 6824 7796 8632
rect 7852 8009 7892 8968
rect 7948 8672 7988 9976
rect 8428 9967 8468 9976
rect 8043 9596 8085 9605
rect 8043 9556 8044 9596
rect 8084 9556 8085 9596
rect 8043 9547 8085 9556
rect 8044 8765 8084 9547
rect 8331 9512 8373 9521
rect 8331 9472 8332 9512
rect 8372 9472 8373 9512
rect 8331 9463 8373 9472
rect 8332 9378 8372 9463
rect 8908 8924 8948 10387
rect 9099 10352 9141 10361
rect 9099 10312 9100 10352
rect 9140 10312 9141 10352
rect 9099 10303 9141 10312
rect 9100 10184 9140 10303
rect 9100 10135 9140 10144
rect 9195 10184 9237 10193
rect 9195 10144 9196 10184
rect 9236 10144 9237 10184
rect 9195 10135 9237 10144
rect 9196 10050 9236 10135
rect 9292 9932 9332 10639
rect 9388 10016 9428 10723
rect 9484 10436 9524 10942
rect 9676 10865 9716 10984
rect 9675 10856 9717 10865
rect 9675 10816 9676 10856
rect 9716 10816 9717 10856
rect 9675 10807 9717 10816
rect 9772 10445 9812 11320
rect 9867 11024 9909 11033
rect 9867 10984 9868 11024
rect 9908 10984 9909 11024
rect 9867 10975 9909 10984
rect 9964 11024 10004 11395
rect 10155 11108 10197 11117
rect 10155 11068 10156 11108
rect 10196 11068 10197 11108
rect 10155 11059 10197 11068
rect 9964 10975 10004 10984
rect 10060 11024 10100 11033
rect 9868 10890 9908 10975
rect 10060 10781 10100 10984
rect 10156 10974 10196 11059
rect 10059 10772 10101 10781
rect 10059 10732 10060 10772
rect 10100 10732 10101 10772
rect 10059 10723 10101 10732
rect 10252 10520 10292 12991
rect 11020 12704 11060 16108
rect 11212 16099 11252 16108
rect 11980 15560 12020 15569
rect 11211 15476 11253 15485
rect 11211 15436 11212 15476
rect 11252 15436 11253 15476
rect 11211 15427 11253 15436
rect 11115 15308 11157 15317
rect 11115 15268 11116 15308
rect 11156 15268 11157 15308
rect 11115 15259 11157 15268
rect 11116 14972 11156 15259
rect 11116 14923 11156 14932
rect 11212 13049 11252 15427
rect 11980 15149 12020 15520
rect 11499 15140 11541 15149
rect 11499 15100 11500 15140
rect 11540 15100 11541 15140
rect 11499 15091 11541 15100
rect 11979 15140 12021 15149
rect 11979 15100 11980 15140
rect 12020 15100 12021 15140
rect 11979 15091 12021 15100
rect 11307 14720 11349 14729
rect 11307 14680 11308 14720
rect 11348 14680 11349 14720
rect 11307 14671 11349 14680
rect 11308 14586 11348 14671
rect 11500 14141 11540 15091
rect 11980 14972 12020 14981
rect 12172 14972 12212 16192
rect 12460 16183 12500 16192
rect 12556 15560 12596 15569
rect 12556 15317 12596 15520
rect 12555 15308 12597 15317
rect 12555 15268 12556 15308
rect 12596 15268 12597 15308
rect 12555 15259 12597 15268
rect 12652 15308 12692 15317
rect 12020 14932 12212 14972
rect 12267 14972 12309 14981
rect 12652 14972 12692 15268
rect 13227 15308 13269 15317
rect 13227 15268 13228 15308
rect 13268 15268 13269 15308
rect 13227 15259 13269 15268
rect 13228 15174 13268 15259
rect 13227 15056 13269 15065
rect 13227 15016 13228 15056
rect 13268 15016 13269 15056
rect 13227 15007 13269 15016
rect 12267 14932 12268 14972
rect 12308 14932 12309 14972
rect 11980 14923 12020 14932
rect 12267 14923 12309 14932
rect 12460 14932 12692 14972
rect 11883 14888 11925 14897
rect 11883 14848 11884 14888
rect 11924 14848 11925 14888
rect 11883 14839 11925 14848
rect 11788 14552 11828 14561
rect 11692 14512 11788 14552
rect 11499 14132 11541 14141
rect 11499 14092 11500 14132
rect 11540 14092 11541 14132
rect 11499 14083 11541 14092
rect 11404 13208 11444 13217
rect 11211 13040 11253 13049
rect 11211 13000 11212 13040
rect 11252 13000 11253 13040
rect 11211 12991 11253 13000
rect 11404 12881 11444 13168
rect 11403 12872 11445 12881
rect 11403 12832 11404 12872
rect 11444 12832 11445 12872
rect 11403 12823 11445 12832
rect 11500 12704 11540 14083
rect 11692 13049 11732 14512
rect 11788 14503 11828 14512
rect 11788 14048 11828 14057
rect 11884 14048 11924 14839
rect 12268 14720 12308 14923
rect 12268 14671 12308 14680
rect 12460 14216 12500 14932
rect 12843 14888 12885 14897
rect 12748 14848 12844 14888
rect 12884 14848 12885 14888
rect 12748 14804 12788 14848
rect 12843 14839 12885 14848
rect 12652 14764 12788 14804
rect 12652 14699 12692 14764
rect 12843 14720 12885 14729
rect 12652 14650 12692 14659
rect 12748 14699 12788 14708
rect 12843 14680 12844 14720
rect 12884 14680 12885 14720
rect 12843 14671 12885 14680
rect 13228 14720 13268 15007
rect 12556 14552 12596 14561
rect 12596 14512 12692 14552
rect 12556 14503 12596 14512
rect 12460 14176 12596 14216
rect 11828 14008 11924 14048
rect 12172 14048 12212 14057
rect 12460 14048 12500 14057
rect 12212 14008 12460 14048
rect 11788 13999 11828 14008
rect 12172 13999 12212 14008
rect 12460 13999 12500 14008
rect 12556 13973 12596 14176
rect 12555 13964 12597 13973
rect 12555 13924 12556 13964
rect 12596 13924 12597 13964
rect 12555 13915 12597 13924
rect 12459 13880 12501 13889
rect 12459 13840 12460 13880
rect 12500 13840 12501 13880
rect 12459 13831 12501 13840
rect 12363 13712 12405 13721
rect 12363 13672 12364 13712
rect 12404 13672 12405 13712
rect 12363 13663 12405 13672
rect 11884 13208 11924 13217
rect 11691 13040 11733 13049
rect 11691 13000 11692 13040
rect 11732 13000 11733 13040
rect 11691 12991 11733 13000
rect 10540 12664 11060 12704
rect 11212 12664 11540 12704
rect 10540 12620 10580 12664
rect 10540 12571 10580 12580
rect 10731 12536 10773 12545
rect 10731 12496 10732 12536
rect 10772 12496 10773 12536
rect 10731 12487 10773 12496
rect 11116 12536 11156 12545
rect 10732 12402 10772 12487
rect 10828 12284 10868 12293
rect 10828 11705 10868 12244
rect 11116 11789 11156 12496
rect 11212 12536 11252 12664
rect 11212 12487 11252 12496
rect 11308 12536 11348 12545
rect 11308 12293 11348 12496
rect 11404 12536 11444 12545
rect 11404 12377 11444 12496
rect 11691 12536 11733 12545
rect 11691 12496 11692 12536
rect 11732 12496 11733 12536
rect 11691 12487 11733 12496
rect 11692 12402 11732 12487
rect 11403 12368 11445 12377
rect 11403 12328 11404 12368
rect 11444 12328 11445 12368
rect 11403 12319 11445 12328
rect 11884 12293 11924 13168
rect 11979 13208 12021 13217
rect 11979 13168 11980 13208
rect 12020 13168 12021 13208
rect 11979 13159 12021 13168
rect 12172 13208 12212 13217
rect 11980 13074 12020 13159
rect 12076 13040 12116 13049
rect 12076 12629 12116 13000
rect 12075 12620 12117 12629
rect 12075 12580 12076 12620
rect 12116 12580 12117 12620
rect 12075 12571 12117 12580
rect 11307 12284 11349 12293
rect 11307 12244 11308 12284
rect 11348 12244 11349 12284
rect 11307 12235 11349 12244
rect 11883 12284 11925 12293
rect 11883 12244 11884 12284
rect 11924 12244 11925 12284
rect 11883 12235 11925 12244
rect 12172 11873 12212 13168
rect 12364 13208 12404 13663
rect 12267 12284 12309 12293
rect 12364 12284 12404 13168
rect 12460 13208 12500 13831
rect 12555 13796 12597 13805
rect 12555 13756 12556 13796
rect 12596 13756 12597 13796
rect 12555 13747 12597 13756
rect 12460 13159 12500 13168
rect 12556 13124 12596 13747
rect 12652 13208 12692 14512
rect 12748 13721 12788 14659
rect 12844 14586 12884 14671
rect 13228 14057 13268 14680
rect 13708 14132 13748 20047
rect 13804 19853 13844 22240
rect 13900 22196 13940 22205
rect 13900 21533 13940 22156
rect 13996 21692 14036 23080
rect 14476 23071 14516 23080
rect 14284 22952 14324 22961
rect 14324 22912 14420 22952
rect 14284 22903 14324 22912
rect 14187 22532 14229 22541
rect 14187 22492 14188 22532
rect 14228 22492 14229 22532
rect 14187 22483 14229 22492
rect 14188 22398 14228 22483
rect 13996 21643 14036 21652
rect 14380 21608 14420 22912
rect 14764 22541 14804 23836
rect 15148 23120 15188 23129
rect 14860 23080 15148 23120
rect 14763 22532 14805 22541
rect 14763 22492 14764 22532
rect 14804 22492 14805 22532
rect 14763 22483 14805 22492
rect 14860 22532 14900 23080
rect 15148 23071 15188 23080
rect 15147 22952 15189 22961
rect 15147 22912 15148 22952
rect 15188 22912 15189 22952
rect 15147 22903 15189 22912
rect 14955 22700 14997 22709
rect 14955 22660 14956 22700
rect 14996 22660 14997 22700
rect 14955 22651 14997 22660
rect 14860 22483 14900 22492
rect 14380 21559 14420 21568
rect 14572 22280 14612 22289
rect 13899 21524 13941 21533
rect 13899 21484 13900 21524
rect 13940 21484 13941 21524
rect 13899 21475 13941 21484
rect 13900 21020 13940 21475
rect 14092 21020 14132 21029
rect 13900 20980 14092 21020
rect 14572 21020 14612 22240
rect 14667 22280 14709 22289
rect 14667 22240 14668 22280
rect 14708 22240 14709 22280
rect 14667 22231 14709 22240
rect 14860 22280 14900 22289
rect 14956 22280 14996 22651
rect 15148 22289 15188 22903
rect 14900 22240 14996 22280
rect 15147 22280 15189 22289
rect 15147 22240 15148 22280
rect 15188 22240 15189 22280
rect 14860 22231 14900 22240
rect 15147 22231 15189 22240
rect 14668 22146 14708 22231
rect 15148 22146 15188 22231
rect 15244 21608 15284 24583
rect 15340 22457 15380 24592
rect 15436 24583 15476 24592
rect 15532 24632 15572 25339
rect 15627 25304 15669 25313
rect 15627 25264 15628 25304
rect 15668 25264 15669 25304
rect 15627 25255 15669 25264
rect 15532 24053 15572 24592
rect 15531 24044 15573 24053
rect 15531 24004 15532 24044
rect 15572 24004 15573 24044
rect 15531 23995 15573 24004
rect 15435 23876 15477 23885
rect 15435 23836 15436 23876
rect 15476 23836 15477 23876
rect 15435 23827 15477 23836
rect 15436 23288 15476 23827
rect 15532 23792 15572 23801
rect 15628 23792 15668 25255
rect 15723 25220 15765 25229
rect 15723 25180 15724 25220
rect 15764 25180 15765 25220
rect 15723 25171 15765 25180
rect 15724 24632 15764 25171
rect 15724 24583 15764 24592
rect 15723 24464 15765 24473
rect 15723 24424 15724 24464
rect 15764 24424 15765 24464
rect 15723 24415 15765 24424
rect 15724 24330 15764 24415
rect 15572 23752 15668 23792
rect 15532 23743 15572 23752
rect 15436 23248 15668 23288
rect 15436 23120 15476 23129
rect 15436 22709 15476 23080
rect 15531 23120 15573 23129
rect 15531 23080 15532 23120
rect 15572 23080 15573 23120
rect 15531 23071 15573 23080
rect 15628 23120 15668 23248
rect 15532 22986 15572 23071
rect 15531 22784 15573 22793
rect 15531 22744 15532 22784
rect 15572 22744 15573 22784
rect 15531 22735 15573 22744
rect 15435 22700 15477 22709
rect 15435 22660 15436 22700
rect 15476 22660 15477 22700
rect 15435 22651 15477 22660
rect 15339 22448 15381 22457
rect 15339 22408 15340 22448
rect 15380 22408 15381 22448
rect 15339 22399 15381 22408
rect 15532 22205 15572 22735
rect 15628 22709 15668 23080
rect 15724 23120 15764 23129
rect 15724 22961 15764 23080
rect 15723 22952 15765 22961
rect 15723 22912 15724 22952
rect 15764 22912 15765 22952
rect 15723 22903 15765 22912
rect 15627 22700 15669 22709
rect 15627 22660 15628 22700
rect 15668 22660 15669 22700
rect 15627 22651 15669 22660
rect 15531 22196 15573 22205
rect 15531 22156 15532 22196
rect 15572 22156 15573 22196
rect 15531 22147 15573 22156
rect 15244 21559 15284 21568
rect 14668 21020 14708 21029
rect 14572 20980 14668 21020
rect 15532 21020 15572 22147
rect 15628 21020 15668 21029
rect 15532 20980 15628 21020
rect 14092 20971 14132 20980
rect 14668 20971 14708 20980
rect 15628 20971 15668 20980
rect 15147 20936 15189 20945
rect 15147 20896 15148 20936
rect 15188 20896 15189 20936
rect 15147 20887 15189 20896
rect 14572 20768 14612 20777
rect 14380 20728 14572 20768
rect 14092 20264 14132 20273
rect 14380 20264 14420 20728
rect 14572 20719 14612 20728
rect 15148 20768 15188 20887
rect 14132 20224 14420 20264
rect 14092 20215 14132 20224
rect 15148 20180 15188 20728
rect 15148 20140 15284 20180
rect 14283 20096 14325 20105
rect 14283 20056 14284 20096
rect 14324 20056 14325 20096
rect 14283 20047 14325 20056
rect 15244 20096 15284 20140
rect 15628 20096 15668 20105
rect 15284 20056 15628 20096
rect 15244 20047 15284 20056
rect 15628 20047 15668 20056
rect 14284 19962 14324 20047
rect 15820 19853 15860 25936
rect 15915 25808 15957 25817
rect 15915 25768 15916 25808
rect 15956 25768 15957 25808
rect 15915 25759 15957 25768
rect 15916 25229 15956 25759
rect 16396 25481 16436 25566
rect 16203 25472 16245 25481
rect 16203 25432 16204 25472
rect 16244 25432 16245 25472
rect 16203 25423 16245 25432
rect 16395 25472 16437 25481
rect 16395 25432 16396 25472
rect 16436 25432 16437 25472
rect 16395 25423 16437 25432
rect 16108 25304 16148 25313
rect 15915 25220 15957 25229
rect 15915 25180 15916 25220
rect 15956 25180 15957 25220
rect 15915 25171 15957 25180
rect 16108 24800 16148 25264
rect 16204 25304 16244 25423
rect 16204 25255 16244 25264
rect 16396 25304 16436 25313
rect 16876 25304 16916 26104
rect 16971 26144 17013 26153
rect 17068 26144 17108 26153
rect 16971 26104 16972 26144
rect 17012 26104 17068 26144
rect 16971 26095 17013 26104
rect 17068 26095 17108 26104
rect 17164 26144 17204 26347
rect 17643 26228 17685 26237
rect 17643 26188 17644 26228
rect 17684 26188 17685 26228
rect 17643 26179 17685 26188
rect 17835 26228 17877 26237
rect 17835 26188 17836 26228
rect 17876 26188 17877 26228
rect 17835 26179 17877 26188
rect 17164 26095 17204 26104
rect 17260 26144 17300 26155
rect 16436 25264 16916 25304
rect 16396 25255 16436 25264
rect 16972 24893 17012 26095
rect 17260 26069 17300 26104
rect 17356 26144 17396 26153
rect 17548 26144 17588 26153
rect 17396 26104 17548 26144
rect 17356 26095 17396 26104
rect 17548 26095 17588 26104
rect 17644 26094 17684 26179
rect 17740 26144 17780 26153
rect 17259 26060 17301 26069
rect 17259 26020 17260 26060
rect 17300 26020 17301 26060
rect 17259 26011 17301 26020
rect 17643 25892 17685 25901
rect 17643 25852 17644 25892
rect 17684 25852 17685 25892
rect 17643 25843 17685 25852
rect 17548 25304 17588 25313
rect 17068 25264 17548 25304
rect 16971 24884 17013 24893
rect 16971 24844 16972 24884
rect 17012 24844 17013 24884
rect 16971 24835 17013 24844
rect 17068 24800 17108 25264
rect 17548 25255 17588 25264
rect 17644 25304 17684 25843
rect 17740 25649 17780 26104
rect 17836 26144 17876 26179
rect 17836 26093 17876 26104
rect 17739 25640 17781 25649
rect 17739 25600 17740 25640
rect 17780 25600 17781 25640
rect 17739 25591 17781 25600
rect 17836 25565 17876 25650
rect 17835 25556 17877 25565
rect 17835 25516 17836 25556
rect 17876 25516 17877 25556
rect 17835 25507 17877 25516
rect 16108 24760 16340 24800
rect 15916 24632 15956 24641
rect 15916 23969 15956 24592
rect 16012 24632 16052 24641
rect 15915 23960 15957 23969
rect 15915 23920 15916 23960
rect 15956 23920 15957 23960
rect 15915 23911 15957 23920
rect 16012 23129 16052 24592
rect 16107 24632 16149 24641
rect 16107 24592 16108 24632
rect 16148 24592 16149 24632
rect 16107 24583 16149 24592
rect 16204 24632 16244 24641
rect 16108 24498 16148 24583
rect 16204 23969 16244 24592
rect 16300 24473 16340 24760
rect 17068 24751 17108 24760
rect 17644 24716 17684 25264
rect 17836 25304 17876 25313
rect 17932 25304 17972 26608
rect 18028 26599 18068 26608
rect 18123 26648 18165 26657
rect 18123 26608 18124 26648
rect 18164 26608 18165 26648
rect 18123 26599 18165 26608
rect 18220 26153 18260 26776
rect 18316 26816 18356 26825
rect 18219 26144 18261 26153
rect 18219 26104 18220 26144
rect 18260 26104 18261 26144
rect 18219 26095 18261 26104
rect 18123 26060 18165 26069
rect 18123 26020 18124 26060
rect 18164 26020 18165 26060
rect 18123 26011 18165 26020
rect 17876 25264 17972 25304
rect 18028 25892 18068 25901
rect 18028 25304 18068 25852
rect 17836 25255 17876 25264
rect 18028 25255 18068 25264
rect 18124 25145 18164 26011
rect 18316 25901 18356 26776
rect 18604 26816 18644 26935
rect 18604 26767 18644 26776
rect 18700 26816 18740 27019
rect 18892 26984 18932 27616
rect 18988 27656 19028 28036
rect 18988 27607 19028 27616
rect 19084 27656 19124 28363
rect 19276 27833 19316 29800
rect 19372 29791 19412 29800
rect 19660 29672 19700 30640
rect 19755 30680 19797 30689
rect 19755 30640 19756 30680
rect 19796 30640 19797 30680
rect 19755 30631 19797 30640
rect 19852 30680 19892 30689
rect 20140 30680 20180 30689
rect 19756 30546 19796 30631
rect 19372 29632 19700 29672
rect 19852 29672 19892 30640
rect 19948 30635 19988 30644
rect 19947 30556 19948 30605
rect 20044 30640 20140 30680
rect 19988 30596 19989 30605
rect 20044 30596 20084 30640
rect 20140 30612 20180 30640
rect 19988 30556 20084 30596
rect 19947 30547 19989 30556
rect 19948 30462 19988 30547
rect 19852 29632 19988 29672
rect 19372 29336 19412 29632
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 19755 29336 19797 29345
rect 19372 29296 19604 29336
rect 19372 29168 19412 29177
rect 19564 29168 19604 29296
rect 19755 29296 19756 29336
rect 19796 29296 19797 29336
rect 19755 29287 19797 29296
rect 19412 29128 19508 29168
rect 19372 29119 19412 29128
rect 19371 29000 19413 29009
rect 19371 28960 19372 29000
rect 19412 28960 19413 29000
rect 19371 28951 19413 28960
rect 19275 27824 19317 27833
rect 19275 27784 19276 27824
rect 19316 27784 19317 27824
rect 19275 27775 19317 27784
rect 19372 27656 19412 28951
rect 19468 28925 19508 29128
rect 19564 29119 19604 29128
rect 19756 29168 19796 29287
rect 19467 28916 19509 28925
rect 19467 28876 19468 28916
rect 19508 28876 19509 28916
rect 19467 28867 19509 28876
rect 19564 28916 19604 28925
rect 19468 28673 19508 28867
rect 19467 28664 19509 28673
rect 19467 28624 19468 28664
rect 19508 28624 19509 28664
rect 19467 28615 19509 28624
rect 19564 28337 19604 28876
rect 19756 28421 19796 29128
rect 19852 29168 19892 29177
rect 19948 29168 19988 29632
rect 20044 29345 20084 30556
rect 20620 30428 20660 30437
rect 20523 29672 20565 29681
rect 20523 29632 20524 29672
rect 20564 29632 20565 29672
rect 20523 29623 20565 29632
rect 20524 29538 20564 29623
rect 20043 29336 20085 29345
rect 20043 29296 20044 29336
rect 20084 29296 20085 29336
rect 20043 29287 20085 29296
rect 20620 29168 20660 30388
rect 19948 29128 20180 29168
rect 19852 29084 19892 29128
rect 19852 29044 19990 29084
rect 19950 29000 19990 29044
rect 19948 28960 19990 29000
rect 19755 28412 19797 28421
rect 19755 28372 19756 28412
rect 19796 28372 19797 28412
rect 19755 28363 19797 28372
rect 19563 28328 19605 28337
rect 19563 28288 19564 28328
rect 19604 28288 19605 28328
rect 19563 28279 19605 28288
rect 19660 28244 19700 28253
rect 19852 28244 19892 28253
rect 19700 28204 19852 28244
rect 19660 28195 19700 28204
rect 19852 28195 19892 28204
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 19467 27824 19509 27833
rect 19467 27784 19468 27824
rect 19508 27784 19509 27824
rect 19467 27775 19509 27784
rect 19084 27581 19124 27616
rect 19276 27616 19412 27656
rect 19083 27572 19125 27581
rect 19083 27532 19084 27572
rect 19124 27532 19125 27572
rect 19083 27523 19125 27532
rect 18987 27404 19029 27413
rect 18987 27364 18988 27404
rect 19028 27364 19029 27404
rect 18987 27355 19029 27364
rect 18700 26767 18740 26776
rect 18796 26944 18932 26984
rect 18796 26816 18836 26944
rect 18796 26657 18836 26776
rect 18795 26648 18837 26657
rect 18795 26608 18796 26648
rect 18836 26608 18837 26648
rect 18795 26599 18837 26608
rect 18892 26648 18932 26659
rect 18700 26144 18740 26153
rect 18315 25892 18357 25901
rect 18315 25852 18316 25892
rect 18356 25852 18357 25892
rect 18315 25843 18357 25852
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 18700 25565 18740 26104
rect 18699 25556 18741 25565
rect 18699 25516 18700 25556
rect 18740 25516 18741 25556
rect 18699 25507 18741 25516
rect 18412 25304 18452 25313
rect 18412 25220 18452 25264
rect 18507 25220 18549 25229
rect 18412 25180 18508 25220
rect 18548 25180 18549 25220
rect 18507 25171 18549 25180
rect 18123 25136 18165 25145
rect 18123 25096 18124 25136
rect 18164 25096 18165 25136
rect 18123 25087 18165 25096
rect 18315 25136 18357 25145
rect 18315 25096 18316 25136
rect 18356 25096 18357 25136
rect 18315 25087 18357 25096
rect 18219 24800 18261 24809
rect 18219 24760 18220 24800
rect 18260 24760 18261 24800
rect 18219 24751 18261 24760
rect 17548 24676 17684 24716
rect 16971 24632 17013 24641
rect 16971 24592 16972 24632
rect 17012 24592 17013 24632
rect 16971 24583 17013 24592
rect 17259 24632 17301 24641
rect 17259 24592 17260 24632
rect 17300 24592 17301 24632
rect 17259 24583 17301 24592
rect 16972 24498 17012 24583
rect 17260 24498 17300 24583
rect 16299 24464 16341 24473
rect 16299 24424 16300 24464
rect 16340 24424 16341 24464
rect 16299 24415 16341 24424
rect 16683 24212 16725 24221
rect 16683 24172 16684 24212
rect 16724 24172 16725 24212
rect 16683 24163 16725 24172
rect 17067 24212 17109 24221
rect 17067 24172 17068 24212
rect 17108 24172 17109 24212
rect 17067 24163 17109 24172
rect 16203 23960 16245 23969
rect 16203 23920 16204 23960
rect 16244 23920 16245 23960
rect 16203 23911 16245 23920
rect 16684 23960 16724 24163
rect 16684 23911 16724 23920
rect 16204 23801 16244 23911
rect 16203 23792 16245 23801
rect 16203 23752 16204 23792
rect 16244 23752 16245 23792
rect 16203 23743 16245 23752
rect 16491 23792 16533 23801
rect 16491 23752 16492 23792
rect 16532 23752 16533 23792
rect 16491 23743 16533 23752
rect 16972 23792 17012 23801
rect 16107 23708 16149 23717
rect 16107 23668 16108 23708
rect 16148 23668 16149 23708
rect 16107 23659 16149 23668
rect 16108 23549 16148 23659
rect 16107 23540 16149 23549
rect 16107 23500 16108 23540
rect 16148 23500 16149 23540
rect 16107 23491 16149 23500
rect 16011 23120 16053 23129
rect 16011 23080 16012 23120
rect 16052 23080 16053 23120
rect 16011 23071 16053 23080
rect 15915 22952 15957 22961
rect 15915 22912 15916 22952
rect 15956 22912 15957 22952
rect 15915 22903 15957 22912
rect 15916 22818 15956 22903
rect 16012 22625 16052 23071
rect 16108 23036 16148 23491
rect 16204 23045 16244 23743
rect 16395 23624 16437 23633
rect 16395 23584 16396 23624
rect 16436 23584 16437 23624
rect 16395 23575 16437 23584
rect 16299 23120 16341 23129
rect 16299 23080 16300 23120
rect 16340 23080 16341 23120
rect 16299 23071 16341 23080
rect 16396 23120 16436 23575
rect 16492 23204 16532 23743
rect 16972 23633 17012 23752
rect 17068 23792 17108 24163
rect 17548 23969 17588 24676
rect 17932 24632 17972 24641
rect 18124 24632 18164 24641
rect 17932 24221 17972 24592
rect 18028 24592 18124 24632
rect 17931 24212 17973 24221
rect 17931 24172 17932 24212
rect 17972 24172 17973 24212
rect 17931 24163 17973 24172
rect 17740 24044 17780 24053
rect 18028 24044 18068 24592
rect 18124 24583 18164 24592
rect 18220 24632 18260 24751
rect 18220 24583 18260 24592
rect 18316 24632 18356 25087
rect 18316 24583 18356 24592
rect 18411 24632 18453 24641
rect 18411 24592 18412 24632
rect 18452 24592 18453 24632
rect 18411 24583 18453 24592
rect 18700 24632 18740 24641
rect 18412 24498 18452 24583
rect 18604 24380 18644 24389
rect 17780 24004 18068 24044
rect 18124 24340 18604 24380
rect 17740 23995 17780 24004
rect 17547 23960 17589 23969
rect 17547 23920 17548 23960
rect 17588 23920 17589 23960
rect 17547 23911 17589 23920
rect 17740 23803 17780 23887
rect 17835 23876 17877 23885
rect 17835 23836 17836 23876
rect 17876 23836 17877 23876
rect 17835 23827 17877 23836
rect 17068 23743 17108 23752
rect 17452 23792 17492 23801
rect 16971 23624 17013 23633
rect 16971 23584 16972 23624
rect 17012 23584 17013 23624
rect 16971 23575 17013 23584
rect 17260 23624 17300 23633
rect 17452 23624 17492 23752
rect 17547 23792 17589 23801
rect 17547 23752 17548 23792
rect 17588 23752 17589 23792
rect 17547 23743 17589 23752
rect 17739 23752 17740 23801
rect 17780 23752 17781 23801
rect 17739 23743 17781 23752
rect 17548 23658 17588 23743
rect 17300 23584 17492 23624
rect 17260 23575 17300 23584
rect 17836 23540 17876 23827
rect 17644 23500 17876 23540
rect 17932 23792 17972 23801
rect 17547 23372 17589 23381
rect 17547 23332 17548 23372
rect 17588 23332 17589 23372
rect 17547 23323 17589 23332
rect 16492 23155 16532 23164
rect 16587 23204 16629 23213
rect 16587 23164 16588 23204
rect 16628 23164 16629 23204
rect 16587 23155 16629 23164
rect 16396 23071 16436 23080
rect 16588 23120 16628 23155
rect 17548 23141 17588 23323
rect 16108 22987 16148 22996
rect 16203 23036 16245 23045
rect 16203 22996 16204 23036
rect 16244 22996 16245 23036
rect 16203 22987 16245 22996
rect 16204 22868 16244 22987
rect 16108 22828 16244 22868
rect 16011 22616 16053 22625
rect 16011 22576 16012 22616
rect 16052 22576 16053 22616
rect 16011 22567 16053 22576
rect 16108 22280 16148 22828
rect 16203 22700 16245 22709
rect 16203 22660 16204 22700
rect 16244 22660 16245 22700
rect 16203 22651 16245 22660
rect 16108 22231 16148 22240
rect 16204 22112 16244 22651
rect 16300 22532 16340 23071
rect 16588 23069 16628 23080
rect 16779 23120 16821 23129
rect 16779 23080 16780 23120
rect 16820 23080 16821 23120
rect 16779 23071 16821 23080
rect 16876 23120 16916 23131
rect 16780 22986 16820 23071
rect 16876 23045 16916 23080
rect 17068 23120 17108 23129
rect 17452 23120 17492 23129
rect 17108 23080 17396 23120
rect 17068 23071 17108 23080
rect 16875 23036 16917 23045
rect 16875 22996 16876 23036
rect 16916 22996 16917 23036
rect 16875 22987 16917 22996
rect 17068 22868 17108 22877
rect 16300 22483 16340 22492
rect 16684 22828 17068 22868
rect 16396 22280 16436 22289
rect 16588 22280 16628 22289
rect 16436 22240 16588 22280
rect 16396 22231 16436 22240
rect 16588 22231 16628 22240
rect 16204 22072 16436 22112
rect 16396 21776 16436 22072
rect 16396 21727 16436 21736
rect 16588 21692 16628 21701
rect 16684 21692 16724 22828
rect 17068 22819 17108 22828
rect 17259 22700 17301 22709
rect 17259 22660 17260 22700
rect 17300 22660 17301 22700
rect 17259 22651 17301 22660
rect 17260 22280 17300 22651
rect 17356 22280 17396 23080
rect 17548 23092 17588 23101
rect 17644 23120 17684 23500
rect 17932 23288 17972 23752
rect 18124 23708 18164 24340
rect 18604 24331 18644 24340
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 18124 23668 18260 23708
rect 18028 23288 18068 23297
rect 17932 23248 18028 23288
rect 18028 23239 18068 23248
rect 17452 22961 17492 23080
rect 17644 23036 17684 23080
rect 17740 23120 17780 23129
rect 17932 23120 17972 23129
rect 17780 23080 17932 23120
rect 17740 23071 17780 23080
rect 17932 23071 17972 23080
rect 18124 23120 18164 23131
rect 18124 23045 18164 23080
rect 18220 23120 18260 23668
rect 18604 23624 18644 23633
rect 18412 23204 18452 23213
rect 18604 23204 18644 23584
rect 18452 23164 18644 23204
rect 18700 23624 18740 24592
rect 18796 23885 18836 26599
rect 18892 26573 18932 26608
rect 18891 26564 18933 26573
rect 18891 26524 18892 26564
rect 18932 26524 18933 26564
rect 18891 26515 18933 26524
rect 18988 26144 19028 27355
rect 19084 26993 19124 27523
rect 19083 26984 19125 26993
rect 19083 26944 19084 26984
rect 19124 26944 19125 26984
rect 19083 26935 19125 26944
rect 19084 26816 19124 26825
rect 19084 26573 19124 26776
rect 19276 26816 19316 27616
rect 19468 27404 19508 27775
rect 19948 27749 19988 28960
rect 20140 28925 20180 29128
rect 20620 29119 20660 29128
rect 20716 30008 20756 30017
rect 20716 29000 20756 29968
rect 20812 29093 20852 29095
rect 20811 29084 20853 29093
rect 20811 29044 20812 29084
rect 20852 29044 20853 29084
rect 20811 29035 20853 29044
rect 20236 28960 20756 29000
rect 20139 28916 20181 28925
rect 20139 28876 20140 28916
rect 20180 28876 20181 28916
rect 20139 28867 20181 28876
rect 20236 28328 20276 28960
rect 20812 28916 20852 29035
rect 20908 29000 20948 31312
rect 21100 30680 21140 31471
rect 21387 30764 21429 30773
rect 21387 30724 21388 30764
rect 21428 30724 21429 30764
rect 21387 30715 21429 30724
rect 21100 30631 21140 30640
rect 21388 30630 21428 30715
rect 21772 30680 21812 31480
rect 22059 31480 22060 31520
rect 22100 31480 22101 31520
rect 22059 31471 22101 31480
rect 22539 31520 22581 31529
rect 22539 31480 22540 31520
rect 22580 31480 22581 31520
rect 22539 31471 22581 31480
rect 21868 31184 21908 31193
rect 21868 30773 21908 31144
rect 21867 30764 21909 30773
rect 21867 30724 21868 30764
rect 21908 30724 21909 30764
rect 21867 30715 21909 30724
rect 21772 30631 21812 30640
rect 21772 29849 21812 29934
rect 21771 29840 21813 29849
rect 21771 29800 21772 29840
rect 21812 29800 21813 29840
rect 21771 29791 21813 29800
rect 21964 29840 22004 29849
rect 21676 29672 21716 29681
rect 21964 29672 22004 29800
rect 22060 29840 22100 31471
rect 22540 31352 22580 31361
rect 22252 31312 22540 31352
rect 22252 30092 22292 31312
rect 22540 31303 22580 31312
rect 22347 31184 22389 31193
rect 22347 31144 22348 31184
rect 22388 31144 22389 31184
rect 22347 31135 22389 31144
rect 22252 30043 22292 30052
rect 22060 29791 22100 29800
rect 22252 29840 22292 29849
rect 22348 29840 22388 31135
rect 22636 30680 22676 33655
rect 22924 33116 22964 33664
rect 23019 33704 23061 33713
rect 23019 33664 23020 33704
rect 23060 33664 23061 33704
rect 23019 33655 23061 33664
rect 23212 33704 23252 33713
rect 23252 33664 23348 33704
rect 23212 33655 23252 33664
rect 23020 33570 23060 33655
rect 23308 33284 23348 33664
rect 23692 33545 23732 33907
rect 23788 33704 23828 33991
rect 23883 33872 23925 33881
rect 23883 33832 23884 33872
rect 23924 33832 23925 33872
rect 23883 33823 23925 33832
rect 23788 33655 23828 33664
rect 23691 33536 23733 33545
rect 23691 33496 23692 33536
rect 23732 33496 23733 33536
rect 23691 33487 23733 33496
rect 23308 33244 23828 33284
rect 23500 33116 23540 33125
rect 22924 33076 23500 33116
rect 23500 33067 23540 33076
rect 23595 33032 23637 33041
rect 23595 32992 23596 33032
rect 23636 32992 23637 33032
rect 23595 32983 23637 32992
rect 23499 32864 23541 32873
rect 23499 32824 23500 32864
rect 23540 32824 23541 32864
rect 23499 32815 23541 32824
rect 23596 32864 23636 32983
rect 23596 32815 23636 32824
rect 23788 32864 23828 33244
rect 23788 32815 23828 32824
rect 23884 32864 23924 33823
rect 23980 33041 24020 34168
rect 24652 33965 24692 34336
rect 24844 34049 24884 34504
rect 25612 34376 25652 34924
rect 25804 34915 25844 34924
rect 25612 34327 25652 34336
rect 26188 34376 26228 34999
rect 26188 34327 26228 34336
rect 25804 34292 25844 34301
rect 25516 34208 25556 34217
rect 24843 34040 24885 34049
rect 24843 34000 24844 34040
rect 24884 34000 24885 34040
rect 24843 33991 24885 34000
rect 24651 33956 24693 33965
rect 24651 33916 24652 33956
rect 24692 33916 24693 33956
rect 24651 33907 24693 33916
rect 25516 33713 25556 34168
rect 25804 33872 25844 34252
rect 26092 33872 26132 33881
rect 25804 33832 26092 33872
rect 26092 33823 26132 33832
rect 24075 33704 24117 33713
rect 24075 33664 24076 33704
rect 24116 33664 24117 33704
rect 24075 33655 24117 33664
rect 24652 33704 24692 33713
rect 24076 33125 24116 33655
rect 24171 33620 24213 33629
rect 24171 33580 24172 33620
rect 24212 33580 24213 33620
rect 24171 33571 24213 33580
rect 24075 33116 24117 33125
rect 24075 33076 24076 33116
rect 24116 33076 24117 33116
rect 24075 33067 24117 33076
rect 23979 33032 24021 33041
rect 23979 32992 23980 33032
rect 24020 32992 24021 33032
rect 23979 32983 24021 32992
rect 23212 32192 23252 32201
rect 23212 31529 23252 32152
rect 22731 31520 22773 31529
rect 22731 31480 22732 31520
rect 22772 31480 22773 31520
rect 22731 31471 22773 31480
rect 23211 31520 23253 31529
rect 23211 31480 23212 31520
rect 23252 31480 23253 31520
rect 23211 31471 23253 31480
rect 22732 31352 22772 31471
rect 22923 31436 22965 31445
rect 22923 31396 22924 31436
rect 22964 31396 22965 31436
rect 22923 31387 22965 31396
rect 22732 31303 22772 31312
rect 22828 31352 22868 31361
rect 22636 30631 22676 30640
rect 22828 30269 22868 31312
rect 22924 31352 22964 31387
rect 22827 30260 22869 30269
rect 22827 30220 22828 30260
rect 22868 30220 22869 30260
rect 22827 30211 22869 30220
rect 22924 30092 22964 31312
rect 23019 31184 23061 31193
rect 23019 31144 23020 31184
rect 23060 31144 23061 31184
rect 23019 31135 23061 31144
rect 23020 31050 23060 31135
rect 23500 30932 23540 32815
rect 23788 31940 23828 31949
rect 23788 31445 23828 31900
rect 23884 31529 23924 32824
rect 23979 32864 24021 32873
rect 23979 32824 23980 32864
rect 24020 32824 24021 32864
rect 23979 32815 24021 32824
rect 24076 32864 24116 33067
rect 24172 32873 24212 33571
rect 24076 32815 24116 32824
rect 24171 32864 24213 32873
rect 24171 32824 24172 32864
rect 24212 32824 24213 32864
rect 24171 32815 24213 32824
rect 24364 32864 24404 32875
rect 24652 32873 24692 33664
rect 25515 33704 25557 33713
rect 25515 33664 25516 33704
rect 25556 33664 25557 33704
rect 25515 33655 25557 33664
rect 25996 33704 26036 33713
rect 26188 33704 26228 33713
rect 26036 33664 26132 33704
rect 25996 33655 26036 33664
rect 25803 33620 25845 33629
rect 25803 33580 25804 33620
rect 25844 33580 25845 33620
rect 25803 33571 25845 33580
rect 25707 33536 25749 33545
rect 25707 33496 25708 33536
rect 25748 33496 25749 33536
rect 25707 33487 25749 33496
rect 24843 33116 24885 33125
rect 24843 33076 24844 33116
rect 24884 33076 24885 33116
rect 24843 33067 24885 33076
rect 24844 32982 24884 33067
rect 23980 32730 24020 32815
rect 24364 32789 24404 32824
rect 24651 32864 24693 32873
rect 24651 32824 24652 32864
rect 24692 32824 24693 32864
rect 24651 32815 24693 32824
rect 25324 32864 25364 32873
rect 24363 32780 24405 32789
rect 24363 32740 24364 32780
rect 24404 32740 24405 32780
rect 24363 32731 24405 32740
rect 25324 32201 25364 32824
rect 25708 32864 25748 33487
rect 25804 33486 25844 33571
rect 25803 33284 25845 33293
rect 25803 33244 25804 33284
rect 25844 33244 25845 33284
rect 25803 33235 25845 33244
rect 25708 32789 25748 32824
rect 25804 32864 25844 33235
rect 25804 32815 25844 32824
rect 25900 32864 25940 32873
rect 25707 32780 25749 32789
rect 25707 32740 25708 32780
rect 25748 32740 25749 32780
rect 25707 32731 25749 32740
rect 25900 32621 25940 32824
rect 25996 32864 26036 32873
rect 26092 32864 26132 33664
rect 26188 33545 26228 33664
rect 26283 33704 26325 33713
rect 26283 33664 26284 33704
rect 26324 33664 26325 33704
rect 26283 33655 26325 33664
rect 26284 33570 26324 33655
rect 26476 33629 26516 35176
rect 30220 35216 30260 35225
rect 29356 35092 29684 35132
rect 26667 35048 26709 35057
rect 26667 35008 26668 35048
rect 26708 35008 26709 35048
rect 26667 34999 26709 35008
rect 29356 35048 29396 35092
rect 29356 34999 29396 35008
rect 26668 34914 26708 34999
rect 29548 34964 29588 34973
rect 29452 34924 29548 34964
rect 27051 34376 27093 34385
rect 26956 34336 27052 34376
rect 27092 34336 27093 34376
rect 26764 33704 26804 33713
rect 26804 33664 26900 33704
rect 26764 33655 26804 33664
rect 26475 33620 26517 33629
rect 26475 33580 26476 33620
rect 26516 33580 26517 33620
rect 26475 33571 26517 33580
rect 26187 33536 26229 33545
rect 26187 33496 26188 33536
rect 26228 33496 26229 33536
rect 26187 33487 26229 33496
rect 26036 32824 26132 32864
rect 25996 32815 26036 32824
rect 26188 32780 26228 32789
rect 26228 32740 26420 32780
rect 26188 32731 26228 32740
rect 25899 32612 25941 32621
rect 25899 32572 25900 32612
rect 25940 32572 25941 32612
rect 25899 32563 25941 32572
rect 26380 32360 26420 32740
rect 26380 32311 26420 32320
rect 26188 32201 26228 32286
rect 25323 32192 25365 32201
rect 25323 32152 25324 32192
rect 25364 32152 25365 32192
rect 25323 32143 25365 32152
rect 25612 32192 25652 32201
rect 25900 32192 25940 32201
rect 25652 32152 25844 32192
rect 25612 32143 25652 32152
rect 24268 32024 24308 32033
rect 23883 31520 23925 31529
rect 23883 31480 23884 31520
rect 23924 31480 24020 31520
rect 23883 31471 23925 31480
rect 23787 31436 23829 31445
rect 23787 31396 23788 31436
rect 23828 31396 23829 31436
rect 23787 31387 23829 31396
rect 23884 31386 23924 31471
rect 23788 31268 23828 31277
rect 23828 31228 23924 31268
rect 23788 31219 23828 31228
rect 23500 30892 23636 30932
rect 22732 30052 22964 30092
rect 22292 29800 22388 29840
rect 22635 29840 22677 29849
rect 22635 29800 22636 29840
rect 22676 29800 22677 29840
rect 22252 29791 22292 29800
rect 22635 29791 22677 29800
rect 21716 29632 22004 29672
rect 22540 29756 22580 29765
rect 21676 29623 21716 29632
rect 22540 29345 22580 29716
rect 22539 29336 22581 29345
rect 22539 29296 22540 29336
rect 22580 29296 22581 29336
rect 22539 29287 22581 29296
rect 22636 29261 22676 29791
rect 22635 29252 22677 29261
rect 22635 29212 22636 29252
rect 22676 29212 22677 29252
rect 22635 29203 22677 29212
rect 21483 29168 21525 29177
rect 21483 29128 21484 29168
rect 21524 29128 21525 29168
rect 21483 29119 21525 29128
rect 22539 29168 22581 29177
rect 22539 29128 22540 29168
rect 22580 29128 22581 29168
rect 22539 29119 22581 29128
rect 22636 29168 22676 29203
rect 21484 29034 21524 29119
rect 22540 29034 22580 29119
rect 22636 29118 22676 29128
rect 22732 29168 22772 30052
rect 22924 29840 22964 29849
rect 22964 29800 23444 29840
rect 22924 29791 22964 29800
rect 23307 29420 23349 29429
rect 23307 29380 23308 29420
rect 23348 29380 23349 29420
rect 23307 29371 23349 29380
rect 23115 29336 23157 29345
rect 23115 29296 23116 29336
rect 23156 29296 23157 29336
rect 23115 29287 23157 29296
rect 23116 29202 23156 29287
rect 22732 29119 22772 29128
rect 22828 29168 22868 29177
rect 23020 29168 23060 29177
rect 22868 29128 23020 29168
rect 22828 29119 22868 29128
rect 23020 29119 23060 29128
rect 23211 29168 23253 29177
rect 23211 29128 23212 29168
rect 23252 29128 23253 29168
rect 23211 29119 23253 29128
rect 23308 29168 23348 29371
rect 23308 29119 23348 29128
rect 23212 29034 23252 29119
rect 23404 29000 23444 29800
rect 23499 29252 23541 29261
rect 23499 29212 23500 29252
rect 23540 29212 23541 29252
rect 23499 29203 23541 29212
rect 23500 29118 23540 29203
rect 20908 28960 21428 29000
rect 23404 28960 23540 29000
rect 20812 28867 20852 28876
rect 20236 28279 20276 28288
rect 20523 28328 20565 28337
rect 20523 28288 20524 28328
rect 20564 28288 20565 28328
rect 20523 28279 20565 28288
rect 21099 28328 21141 28337
rect 21099 28288 21100 28328
rect 21140 28288 21141 28328
rect 21099 28279 21141 28288
rect 19947 27740 19989 27749
rect 19947 27700 19948 27740
rect 19988 27700 19989 27740
rect 19947 27691 19989 27700
rect 19563 27656 19605 27665
rect 19563 27616 19564 27656
rect 19604 27616 19605 27656
rect 19563 27607 19605 27616
rect 20524 27656 20564 28279
rect 21100 28194 21140 28279
rect 20715 27740 20757 27749
rect 20715 27700 20716 27740
rect 20756 27700 20757 27740
rect 20715 27691 20757 27700
rect 20524 27607 20564 27616
rect 19564 27522 19604 27607
rect 20716 27606 20756 27691
rect 20812 27656 20852 27665
rect 21004 27656 21044 27665
rect 20852 27616 21004 27656
rect 20812 27607 20852 27616
rect 21004 27607 21044 27616
rect 19852 27404 19892 27413
rect 19468 27364 19852 27404
rect 19371 26984 19413 26993
rect 19371 26944 19372 26984
rect 19412 26944 19413 26984
rect 19371 26935 19413 26944
rect 19276 26767 19316 26776
rect 19372 26816 19412 26935
rect 19372 26767 19412 26776
rect 19179 26648 19221 26657
rect 19468 26648 19508 27364
rect 19852 27355 19892 27364
rect 20043 27236 20085 27245
rect 20043 27196 20044 27236
rect 20084 27196 20085 27236
rect 20043 27187 20085 27196
rect 19563 26816 19605 26825
rect 19563 26776 19564 26816
rect 19604 26776 19605 26816
rect 19563 26767 19605 26776
rect 19564 26682 19604 26767
rect 20044 26741 20084 27187
rect 20523 27068 20565 27077
rect 20523 27028 20524 27068
rect 20564 27028 20565 27068
rect 20523 27019 20565 27028
rect 20524 26934 20564 27019
rect 20619 26984 20661 26993
rect 20619 26944 20620 26984
rect 20660 26944 20661 26984
rect 20619 26935 20661 26944
rect 20236 26816 20276 26825
rect 20276 26776 20372 26816
rect 20236 26767 20276 26776
rect 20043 26732 20085 26741
rect 20043 26692 20044 26732
rect 20084 26692 20085 26732
rect 20043 26683 20085 26692
rect 19179 26608 19180 26648
rect 19220 26608 19221 26648
rect 19179 26599 19221 26608
rect 19276 26608 19508 26648
rect 19083 26564 19125 26573
rect 19083 26524 19084 26564
rect 19124 26524 19125 26564
rect 19083 26515 19125 26524
rect 19180 26514 19220 26599
rect 19084 26144 19124 26153
rect 18988 26104 19084 26144
rect 18892 24464 18932 24473
rect 18795 23876 18837 23885
rect 18795 23836 18796 23876
rect 18836 23836 18837 23876
rect 18795 23827 18837 23836
rect 18796 23624 18836 23633
rect 18700 23584 18796 23624
rect 18412 23155 18452 23164
rect 18220 23071 18260 23080
rect 17548 22996 17684 23036
rect 18123 23036 18165 23045
rect 18123 22996 18124 23036
rect 18164 22996 18165 23036
rect 17451 22952 17493 22961
rect 17451 22912 17452 22952
rect 17492 22912 17493 22952
rect 17451 22903 17493 22912
rect 17548 22625 17588 22996
rect 18123 22987 18165 22996
rect 17739 22952 17781 22961
rect 17739 22912 17740 22952
rect 17780 22912 17781 22952
rect 17739 22903 17781 22912
rect 17643 22784 17685 22793
rect 17643 22744 17644 22784
rect 17684 22744 17685 22784
rect 17643 22735 17685 22744
rect 17547 22616 17589 22625
rect 17547 22576 17548 22616
rect 17588 22576 17589 22616
rect 17547 22567 17589 22576
rect 17452 22280 17492 22289
rect 17356 22240 17452 22280
rect 17260 22231 17300 22240
rect 17452 22231 17492 22240
rect 17548 22280 17588 22567
rect 17548 22121 17588 22240
rect 17644 22280 17684 22735
rect 17644 22231 17684 22240
rect 17740 22280 17780 22903
rect 18700 22793 18740 23584
rect 18796 23575 18836 23584
rect 18892 23456 18932 24424
rect 18987 23792 19029 23801
rect 18987 23752 18988 23792
rect 19028 23752 19029 23792
rect 18987 23743 19029 23752
rect 18796 23416 18932 23456
rect 18796 23120 18836 23416
rect 18988 23213 19028 23743
rect 19084 23633 19124 26104
rect 19276 25313 19316 26608
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19468 26144 19508 26153
rect 19372 26010 19412 26095
rect 19275 25304 19317 25313
rect 19275 25264 19276 25304
rect 19316 25264 19317 25304
rect 19275 25255 19317 25264
rect 19179 25220 19221 25229
rect 19179 25180 19180 25220
rect 19220 25180 19221 25220
rect 19179 25171 19221 25180
rect 19180 24464 19220 25171
rect 19276 25170 19316 25255
rect 19468 25136 19508 26104
rect 19948 26144 19988 26153
rect 19756 25976 19796 25985
rect 19948 25976 19988 26104
rect 20044 26144 20084 26683
rect 20139 26228 20181 26237
rect 20139 26188 20140 26228
rect 20180 26188 20181 26228
rect 20139 26179 20181 26188
rect 20044 26095 20084 26104
rect 20140 26094 20180 26179
rect 20332 26153 20372 26776
rect 20427 26648 20469 26657
rect 20427 26608 20428 26648
rect 20468 26608 20469 26648
rect 20427 26599 20469 26608
rect 20236 26144 20276 26153
rect 19796 25936 19988 25976
rect 19756 25927 19796 25936
rect 20236 25817 20276 26104
rect 20331 26144 20373 26153
rect 20331 26104 20332 26144
rect 20372 26104 20373 26144
rect 20331 26095 20373 26104
rect 20428 26144 20468 26599
rect 20428 26095 20468 26104
rect 20235 25808 20277 25817
rect 20235 25768 20236 25808
rect 20276 25768 20277 25808
rect 20235 25759 20277 25768
rect 20332 25556 20372 26095
rect 20428 25556 20468 25565
rect 20332 25516 20428 25556
rect 20428 25507 20468 25516
rect 20620 25556 20660 26935
rect 21099 26312 21141 26321
rect 21099 26272 21100 26312
rect 21140 26272 21141 26312
rect 21099 26263 21141 26272
rect 21100 26178 21140 26263
rect 21099 25892 21141 25901
rect 21099 25852 21100 25892
rect 21140 25852 21141 25892
rect 21099 25843 21141 25852
rect 20620 25507 20660 25516
rect 20716 25304 20756 25313
rect 20908 25304 20948 25313
rect 20756 25264 20908 25304
rect 20716 25255 20756 25264
rect 20908 25255 20948 25264
rect 19372 25096 19508 25136
rect 19276 24464 19316 24473
rect 19180 24424 19276 24464
rect 19276 24415 19316 24424
rect 19083 23624 19125 23633
rect 19083 23584 19084 23624
rect 19124 23584 19125 23624
rect 19083 23575 19125 23584
rect 19372 23381 19412 25096
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 20908 24632 20948 24641
rect 20908 24305 20948 24592
rect 21003 24632 21045 24641
rect 21003 24592 21004 24632
rect 21044 24592 21045 24632
rect 21003 24583 21045 24592
rect 21100 24632 21140 25843
rect 21100 24583 21140 24592
rect 21195 24632 21237 24641
rect 21195 24592 21196 24632
rect 21236 24592 21237 24632
rect 21195 24583 21237 24592
rect 21004 24498 21044 24583
rect 21196 24498 21236 24583
rect 20907 24296 20949 24305
rect 20907 24256 20908 24296
rect 20948 24256 20949 24296
rect 20907 24247 20949 24256
rect 20811 23960 20853 23969
rect 20811 23920 20812 23960
rect 20852 23920 20853 23960
rect 20811 23911 20853 23920
rect 21388 23960 21428 28960
rect 22251 28916 22293 28925
rect 22251 28876 22252 28916
rect 22292 28876 22293 28916
rect 22251 28867 22293 28876
rect 21867 28832 21909 28841
rect 21867 28792 21868 28832
rect 21908 28792 21909 28832
rect 21867 28783 21909 28792
rect 21676 27656 21716 27665
rect 21676 27077 21716 27616
rect 21868 27656 21908 28783
rect 22252 28580 22292 28867
rect 22252 28531 22292 28540
rect 23500 28496 23540 28960
rect 23500 28447 23540 28456
rect 23596 27824 23636 30892
rect 23788 30428 23828 30437
rect 23788 30269 23828 30388
rect 23787 30260 23829 30269
rect 23787 30220 23788 30260
rect 23828 30220 23829 30260
rect 23787 30211 23829 30220
rect 23788 29840 23828 29849
rect 23788 28337 23828 29800
rect 23884 29765 23924 31228
rect 23980 30689 24020 31480
rect 24172 31352 24212 31361
rect 24268 31352 24308 31984
rect 24940 31940 24980 31949
rect 24980 31900 25268 31940
rect 24940 31891 24980 31900
rect 25228 31613 25268 31900
rect 25227 31604 25269 31613
rect 25227 31564 25228 31604
rect 25268 31564 25269 31604
rect 25227 31555 25269 31564
rect 25035 31520 25077 31529
rect 25035 31480 25036 31520
rect 25076 31480 25077 31520
rect 25035 31471 25077 31480
rect 24939 31436 24981 31445
rect 24939 31396 24940 31436
rect 24980 31396 24981 31436
rect 24939 31387 24981 31396
rect 24212 31312 24308 31352
rect 24172 31303 24212 31312
rect 23979 30680 24021 30689
rect 23979 30640 23980 30680
rect 24020 30640 24021 30680
rect 23979 30631 24021 30640
rect 23883 29756 23925 29765
rect 23883 29716 23884 29756
rect 23924 29716 23925 29756
rect 23883 29707 23925 29716
rect 23980 29000 24020 30631
rect 24940 30521 24980 31387
rect 25036 31352 25076 31471
rect 25036 31303 25076 31312
rect 25036 30680 25076 30689
rect 24939 30512 24981 30521
rect 24939 30472 24940 30512
rect 24980 30472 24981 30512
rect 24939 30463 24981 30472
rect 24940 30260 24980 30463
rect 25036 30344 25076 30640
rect 25132 30680 25172 30689
rect 25132 30521 25172 30640
rect 25228 30680 25268 31555
rect 25228 30631 25268 30640
rect 25324 30680 25364 32143
rect 25804 31604 25844 32152
rect 25900 31781 25940 32152
rect 25995 32192 26037 32201
rect 25995 32152 25996 32192
rect 26036 32152 26037 32192
rect 25995 32143 26037 32152
rect 26187 32192 26229 32201
rect 26476 32192 26516 33571
rect 26572 32864 26612 32873
rect 26572 32780 26612 32824
rect 26667 32780 26709 32789
rect 26572 32740 26668 32780
rect 26708 32740 26709 32780
rect 26667 32731 26709 32740
rect 26667 32612 26709 32621
rect 26667 32572 26668 32612
rect 26708 32572 26709 32612
rect 26667 32563 26709 32572
rect 26571 32276 26613 32285
rect 26571 32236 26572 32276
rect 26612 32236 26613 32276
rect 26571 32227 26613 32236
rect 26187 32152 26188 32192
rect 26228 32152 26229 32192
rect 26187 32143 26229 32152
rect 26284 32152 26516 32192
rect 25996 32058 26036 32143
rect 26187 32024 26229 32033
rect 26187 31984 26188 32024
rect 26228 31984 26229 32024
rect 26187 31975 26229 31984
rect 26188 31890 26228 31975
rect 25899 31772 25941 31781
rect 25899 31732 25900 31772
rect 25940 31732 25941 31772
rect 25899 31723 25941 31732
rect 26188 31604 26228 31613
rect 25804 31564 26188 31604
rect 25612 30680 25652 30689
rect 25364 30640 25460 30680
rect 25324 30631 25364 30640
rect 25131 30512 25173 30521
rect 25131 30472 25132 30512
rect 25172 30472 25173 30512
rect 25131 30463 25173 30472
rect 25036 30304 25268 30344
rect 24940 30220 25076 30260
rect 24171 29672 24213 29681
rect 24171 29632 24172 29672
rect 24212 29632 24213 29672
rect 24171 29623 24213 29632
rect 24939 29672 24981 29681
rect 24939 29632 24940 29672
rect 24980 29632 24981 29672
rect 24939 29623 24981 29632
rect 24172 29168 24212 29623
rect 24940 29538 24980 29623
rect 24172 29119 24212 29128
rect 24940 29168 24980 29177
rect 24748 29000 24788 29009
rect 23980 28960 24116 29000
rect 23787 28328 23829 28337
rect 23787 28288 23788 28328
rect 23828 28288 23829 28328
rect 23787 28279 23829 28288
rect 23596 27775 23636 27784
rect 23787 27740 23829 27749
rect 23787 27700 23788 27740
rect 23828 27700 23829 27740
rect 23787 27691 23829 27700
rect 21868 27607 21908 27616
rect 22827 27656 22869 27665
rect 22827 27616 22828 27656
rect 22868 27616 22869 27656
rect 22827 27607 22869 27616
rect 22828 27522 22868 27607
rect 23788 27488 23828 27691
rect 23883 27656 23925 27665
rect 23980 27656 24020 27665
rect 23883 27616 23884 27656
rect 23924 27616 23980 27656
rect 23883 27607 23925 27616
rect 23980 27607 24020 27616
rect 23788 27439 23828 27448
rect 21675 27068 21717 27077
rect 21675 27028 21676 27068
rect 21716 27028 21717 27068
rect 21675 27019 21717 27028
rect 23403 26984 23445 26993
rect 23403 26944 23404 26984
rect 23444 26944 23445 26984
rect 23403 26935 23445 26944
rect 23404 26850 23444 26935
rect 21676 26816 21716 26825
rect 21676 26153 21716 26776
rect 22540 26816 22580 26825
rect 22155 26480 22197 26489
rect 22155 26440 22156 26480
rect 22196 26440 22197 26480
rect 22155 26431 22197 26440
rect 21675 26144 21717 26153
rect 21675 26104 21676 26144
rect 21716 26104 21717 26144
rect 21675 26095 21717 26104
rect 21964 26144 22004 26155
rect 21483 25976 21525 25985
rect 21483 25936 21484 25976
rect 21524 25936 21525 25976
rect 21483 25927 21525 25936
rect 21484 25842 21524 25927
rect 21580 25304 21620 25313
rect 21483 24380 21525 24389
rect 21483 24340 21484 24380
rect 21524 24340 21525 24380
rect 21483 24331 21525 24340
rect 21484 24246 21524 24331
rect 21580 23969 21620 25264
rect 21388 23911 21428 23920
rect 21579 23960 21621 23969
rect 21579 23920 21580 23960
rect 21620 23920 21621 23960
rect 21579 23911 21621 23920
rect 19467 23792 19509 23801
rect 19467 23752 19468 23792
rect 19508 23752 19509 23792
rect 19467 23743 19509 23752
rect 20716 23792 20756 23801
rect 19468 23658 19508 23743
rect 20716 23549 20756 23752
rect 20715 23540 20757 23549
rect 20715 23500 20716 23540
rect 20756 23500 20757 23540
rect 20715 23491 20757 23500
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 20812 23381 20852 23911
rect 21580 23792 21620 23801
rect 21580 23465 21620 23752
rect 21579 23456 21621 23465
rect 21484 23416 21580 23456
rect 21620 23416 21621 23456
rect 19371 23372 19413 23381
rect 19371 23332 19372 23372
rect 19412 23332 19413 23372
rect 19371 23323 19413 23332
rect 20811 23372 20853 23381
rect 20811 23332 20812 23372
rect 20852 23332 20853 23372
rect 20811 23323 20853 23332
rect 20812 23288 20852 23323
rect 20812 23238 20852 23248
rect 18987 23204 19029 23213
rect 18987 23164 18988 23204
rect 19028 23164 19029 23204
rect 18987 23155 19029 23164
rect 18796 23071 18836 23080
rect 18699 22784 18741 22793
rect 18699 22744 18700 22784
rect 18740 22744 18741 22784
rect 18699 22735 18741 22744
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 18220 22373 18260 22404
rect 18219 22364 18261 22373
rect 18219 22324 18220 22364
rect 18260 22324 18261 22364
rect 18219 22315 18261 22324
rect 17740 22231 17780 22240
rect 17835 22280 17877 22289
rect 17835 22240 17836 22280
rect 17876 22240 17877 22280
rect 17835 22231 17877 22240
rect 18220 22280 18260 22315
rect 17547 22112 17589 22121
rect 17547 22072 17548 22112
rect 17588 22072 17589 22112
rect 17547 22063 17589 22072
rect 16628 21652 16724 21692
rect 16588 21643 16628 21652
rect 16972 21608 17012 21617
rect 17836 21608 17876 22231
rect 18220 22205 18260 22240
rect 18219 22196 18261 22205
rect 18219 22156 18220 22196
rect 18260 22156 18261 22196
rect 18219 22147 18261 22156
rect 18699 22112 18741 22121
rect 18699 22072 18700 22112
rect 18740 22072 18741 22112
rect 18699 22063 18741 22072
rect 18700 21978 18740 22063
rect 18988 21776 19028 23155
rect 19659 23120 19701 23129
rect 18988 21727 19028 21736
rect 19372 23080 19660 23120
rect 19700 23080 19701 23120
rect 17012 21568 17108 21608
rect 16972 21559 17012 21568
rect 16492 20936 16532 20945
rect 13803 19844 13845 19853
rect 13803 19804 13804 19844
rect 13844 19804 13845 19844
rect 13803 19795 13845 19804
rect 14283 19844 14325 19853
rect 15819 19844 15861 19853
rect 14283 19804 14284 19844
rect 14324 19804 14325 19844
rect 14283 19795 14325 19804
rect 15724 19804 15820 19844
rect 15860 19804 15861 19844
rect 14284 19508 14324 19795
rect 14284 19459 14324 19468
rect 14763 19256 14805 19265
rect 14763 19216 14764 19256
rect 14804 19216 14805 19256
rect 14763 19207 14805 19216
rect 14860 19256 14900 19265
rect 14379 19088 14421 19097
rect 14379 19048 14380 19088
rect 14420 19048 14421 19088
rect 14379 19039 14421 19048
rect 13996 17072 14036 17081
rect 13996 16409 14036 17032
rect 13995 16400 14037 16409
rect 13995 16360 13996 16400
rect 14036 16360 14037 16400
rect 13995 16351 14037 16360
rect 14187 16232 14229 16241
rect 14187 16192 14188 16232
rect 14228 16192 14229 16232
rect 14187 16183 14229 16192
rect 14188 16098 14228 16183
rect 14380 15560 14420 19039
rect 14764 18752 14804 19207
rect 14764 18703 14804 18712
rect 14475 18080 14517 18089
rect 14475 18040 14476 18080
rect 14516 18040 14517 18080
rect 14475 18031 14517 18040
rect 14476 17996 14516 18031
rect 14476 17945 14516 17956
rect 14763 17660 14805 17669
rect 14763 17620 14764 17660
rect 14804 17620 14805 17660
rect 14763 17611 14805 17620
rect 14764 17526 14804 17611
rect 14668 16820 14708 16829
rect 14668 16241 14708 16780
rect 14667 16232 14709 16241
rect 14667 16192 14668 16232
rect 14708 16192 14709 16232
rect 14667 16183 14709 16192
rect 14380 15511 14420 15520
rect 14763 15056 14805 15065
rect 14763 15016 14764 15056
rect 14804 15016 14805 15056
rect 14763 15007 14805 15016
rect 13803 14972 13845 14981
rect 13803 14932 13804 14972
rect 13844 14932 13845 14972
rect 13803 14923 13845 14932
rect 13804 14838 13844 14923
rect 14091 14888 14133 14897
rect 14091 14848 14092 14888
rect 14132 14848 14133 14888
rect 14091 14839 14133 14848
rect 13803 14132 13845 14141
rect 13708 14092 13804 14132
rect 13844 14092 13845 14132
rect 13803 14083 13845 14092
rect 13132 14048 13172 14057
rect 13132 13889 13172 14008
rect 13227 14048 13269 14057
rect 13227 14008 13228 14048
rect 13268 14008 13269 14048
rect 13227 13999 13269 14008
rect 13804 14048 13844 14083
rect 13804 13997 13844 14008
rect 13131 13880 13173 13889
rect 13131 13840 13132 13880
rect 13172 13840 13173 13880
rect 13131 13831 13173 13840
rect 14092 13880 14132 14839
rect 14764 14804 14804 15007
rect 14860 14981 14900 19216
rect 15243 19088 15285 19097
rect 15243 19048 15244 19088
rect 15284 19048 15285 19088
rect 15243 19039 15285 19048
rect 15244 18954 15284 19039
rect 15148 17744 15188 17753
rect 15148 16904 15188 17704
rect 15244 16904 15284 16913
rect 15148 16864 15244 16904
rect 15244 16855 15284 16864
rect 15339 16400 15381 16409
rect 15339 16360 15340 16400
rect 15380 16360 15381 16400
rect 15339 16351 15381 16360
rect 15051 16316 15093 16325
rect 15051 16276 15052 16316
rect 15092 16276 15093 16316
rect 15051 16267 15093 16276
rect 15052 16232 15092 16267
rect 15052 16181 15092 16192
rect 15244 15560 15284 15569
rect 15148 15520 15244 15560
rect 14955 15308 14997 15317
rect 14955 15268 14956 15308
rect 14996 15268 14997 15308
rect 14955 15259 14997 15268
rect 14859 14972 14901 14981
rect 14859 14932 14860 14972
rect 14900 14932 14901 14972
rect 14859 14923 14901 14932
rect 14764 14764 14900 14804
rect 14283 14720 14325 14729
rect 14283 14680 14284 14720
rect 14324 14680 14325 14720
rect 14283 14671 14325 14680
rect 14092 13831 14132 13840
rect 14284 14552 14324 14671
rect 12747 13712 12789 13721
rect 12747 13672 12748 13712
rect 12788 13672 12789 13712
rect 12747 13663 12789 13672
rect 14284 13544 14324 14512
rect 14763 14048 14805 14057
rect 14763 14008 14764 14048
rect 14804 14008 14805 14048
rect 14763 13999 14805 14008
rect 14764 13914 14804 13999
rect 14476 13796 14516 13805
rect 13996 13504 14324 13544
rect 14380 13756 14476 13796
rect 12939 13376 12981 13385
rect 12939 13336 12940 13376
rect 12980 13336 12981 13376
rect 12939 13327 12981 13336
rect 12652 13159 12692 13168
rect 12843 13208 12885 13217
rect 12843 13168 12844 13208
rect 12884 13168 12885 13208
rect 12843 13159 12885 13168
rect 12556 13075 12596 13084
rect 12459 13040 12501 13049
rect 12459 13000 12460 13040
rect 12500 13000 12501 13040
rect 12459 12991 12501 13000
rect 12267 12244 12268 12284
rect 12308 12244 12364 12284
rect 12267 12235 12309 12244
rect 12364 12235 12404 12244
rect 11404 11864 11444 11873
rect 12171 11864 12213 11873
rect 11115 11780 11157 11789
rect 11115 11740 11116 11780
rect 11156 11740 11157 11780
rect 11115 11731 11157 11740
rect 10827 11696 10869 11705
rect 10827 11656 10828 11696
rect 10868 11656 10869 11696
rect 10827 11647 10869 11656
rect 11404 11621 11444 11824
rect 11596 11824 12020 11864
rect 11596 11696 11636 11824
rect 11596 11647 11636 11656
rect 11692 11696 11732 11705
rect 11403 11612 11445 11621
rect 11403 11572 11404 11612
rect 11444 11572 11445 11612
rect 11403 11563 11445 11572
rect 11307 11192 11349 11201
rect 11307 11152 11308 11192
rect 11348 11152 11349 11192
rect 11307 11143 11349 11152
rect 11308 11058 11348 11143
rect 10156 10480 10292 10520
rect 11308 10772 11348 10781
rect 9580 10436 9620 10445
rect 9484 10396 9580 10436
rect 9580 10387 9620 10396
rect 9771 10436 9813 10445
rect 9771 10396 9772 10436
rect 9812 10396 9813 10436
rect 9771 10387 9813 10396
rect 9675 10352 9717 10361
rect 9675 10312 9676 10352
rect 9716 10312 9717 10352
rect 9675 10303 9717 10312
rect 9388 9967 9428 9976
rect 9580 10184 9620 10193
rect 9676 10184 9716 10303
rect 9771 10268 9813 10277
rect 9771 10228 9772 10268
rect 9812 10228 9813 10268
rect 9771 10219 9813 10228
rect 9620 10144 9716 10184
rect 9196 9892 9332 9932
rect 8908 8875 8948 8884
rect 9004 9512 9044 9521
rect 9004 8849 9044 9472
rect 9196 9512 9236 9892
rect 9580 9848 9620 10144
rect 9675 10016 9717 10025
rect 9675 9976 9676 10016
rect 9716 9976 9717 10016
rect 9675 9967 9717 9976
rect 9196 9463 9236 9472
rect 9292 9808 9620 9848
rect 9292 9512 9332 9808
rect 9484 9680 9524 9689
rect 9292 9463 9332 9472
rect 9388 9596 9428 9605
rect 9291 9344 9333 9353
rect 9291 9304 9292 9344
rect 9332 9304 9333 9344
rect 9291 9295 9333 9304
rect 9292 9210 9332 9295
rect 9388 9185 9428 9556
rect 9387 9176 9429 9185
rect 9387 9136 9388 9176
rect 9428 9136 9429 9176
rect 9387 9127 9429 9136
rect 8331 8840 8373 8849
rect 8331 8800 8332 8840
rect 8372 8800 8373 8840
rect 8331 8791 8373 8800
rect 9003 8840 9045 8849
rect 9003 8800 9004 8840
rect 9044 8800 9045 8840
rect 9003 8791 9045 8800
rect 8043 8756 8085 8765
rect 8043 8716 8044 8756
rect 8084 8716 8085 8756
rect 8043 8707 8085 8716
rect 7948 8623 7988 8632
rect 8236 8672 8276 8681
rect 7948 8504 7988 8513
rect 8236 8504 8276 8632
rect 7988 8464 8276 8504
rect 7948 8455 7988 8464
rect 8139 8168 8181 8177
rect 8139 8128 8140 8168
rect 8180 8128 8181 8168
rect 8139 8119 8181 8128
rect 8236 8168 8276 8177
rect 8332 8168 8372 8791
rect 8907 8672 8949 8681
rect 8907 8632 8908 8672
rect 8948 8632 8949 8672
rect 8907 8623 8949 8632
rect 8619 8420 8661 8429
rect 8619 8380 8620 8420
rect 8660 8380 8661 8420
rect 8619 8371 8661 8380
rect 8276 8128 8372 8168
rect 8523 8168 8565 8177
rect 8523 8128 8524 8168
rect 8564 8128 8565 8168
rect 8236 8119 8276 8128
rect 8523 8119 8565 8128
rect 8044 8084 8084 8093
rect 7851 8000 7893 8009
rect 7851 7960 7852 8000
rect 7892 7960 7893 8000
rect 7851 7951 7893 7960
rect 7948 8000 7988 8009
rect 7852 7866 7892 7951
rect 7948 7001 7988 7960
rect 8044 7757 8084 8044
rect 8140 8034 8180 8119
rect 8043 7748 8085 7757
rect 8043 7708 8044 7748
rect 8084 7708 8085 7748
rect 8043 7699 8085 7708
rect 8427 7748 8469 7757
rect 8427 7708 8428 7748
rect 8468 7708 8469 7748
rect 8427 7699 8469 7708
rect 8428 7614 8468 7699
rect 8332 7001 8372 7086
rect 7947 6992 7989 7001
rect 7947 6952 7948 6992
rect 7988 6952 7989 6992
rect 7947 6943 7989 6952
rect 8331 6992 8373 7001
rect 8331 6952 8332 6992
rect 8372 6952 8373 6992
rect 8524 6992 8564 8119
rect 8620 7160 8660 8371
rect 8715 7580 8757 7589
rect 8715 7540 8716 7580
rect 8756 7540 8757 7580
rect 8715 7531 8757 7540
rect 8620 7111 8660 7120
rect 8716 7001 8756 7531
rect 8812 7421 8852 7506
rect 8811 7412 8853 7421
rect 8811 7372 8812 7412
rect 8852 7372 8853 7412
rect 8811 7363 8853 7372
rect 8908 7244 8948 8623
rect 9100 8588 9140 8597
rect 9004 8548 9100 8588
rect 9004 7673 9044 8548
rect 9100 8539 9140 8548
rect 9388 8177 9428 9127
rect 9484 8849 9524 9640
rect 9676 9512 9716 9967
rect 9772 9932 9812 10219
rect 9867 10184 9909 10193
rect 9867 10144 9868 10184
rect 9908 10144 9909 10184
rect 9867 10135 9909 10144
rect 9868 10050 9908 10135
rect 9963 10100 10005 10109
rect 9963 10060 9964 10100
rect 10004 10060 10005 10100
rect 9963 10051 10005 10060
rect 9772 9892 9908 9932
rect 9772 9689 9812 9774
rect 9771 9680 9813 9689
rect 9771 9640 9772 9680
rect 9812 9640 9813 9680
rect 9771 9631 9813 9640
rect 9772 9512 9812 9521
rect 9676 9472 9772 9512
rect 9772 9463 9812 9472
rect 9483 8840 9525 8849
rect 9483 8800 9484 8840
rect 9524 8800 9525 8840
rect 9868 8840 9908 9892
rect 9964 9512 10004 10051
rect 9964 9463 10004 9472
rect 10060 9512 10100 9521
rect 10156 9512 10196 10480
rect 10635 10436 10677 10445
rect 10635 10396 10636 10436
rect 10676 10396 10677 10436
rect 10635 10387 10677 10396
rect 10252 10352 10292 10361
rect 10252 9848 10292 10312
rect 10539 10184 10581 10193
rect 10539 10144 10540 10184
rect 10580 10144 10581 10184
rect 10539 10135 10581 10144
rect 10636 10184 10676 10387
rect 11308 10361 11348 10732
rect 11307 10352 11349 10361
rect 11307 10312 11308 10352
rect 11348 10312 11349 10352
rect 11307 10303 11349 10312
rect 10636 10135 10676 10144
rect 10731 10184 10773 10193
rect 11596 10184 11636 10193
rect 10731 10144 10732 10184
rect 10772 10144 10773 10184
rect 10731 10135 10773 10144
rect 11404 10144 11596 10184
rect 10540 10050 10580 10135
rect 10732 10050 10772 10135
rect 10444 10016 10484 10025
rect 10444 9932 10484 9976
rect 10924 10016 10964 10025
rect 10444 9892 10772 9932
rect 10252 9808 10676 9848
rect 10251 9596 10293 9605
rect 10251 9556 10252 9596
rect 10292 9556 10293 9596
rect 10251 9547 10293 9556
rect 10100 9472 10196 9512
rect 10060 9463 10100 9472
rect 10059 8840 10101 8849
rect 9868 8800 10004 8840
rect 9483 8791 9525 8800
rect 9676 8672 9716 8681
rect 9676 8429 9716 8632
rect 9867 8672 9909 8681
rect 9867 8632 9868 8672
rect 9908 8632 9909 8672
rect 9867 8623 9909 8632
rect 9772 8588 9812 8597
rect 9675 8420 9717 8429
rect 9675 8380 9676 8420
rect 9716 8380 9717 8420
rect 9675 8371 9717 8380
rect 9772 8252 9812 8548
rect 9868 8538 9908 8623
rect 9676 8212 9812 8252
rect 9387 8168 9429 8177
rect 9387 8128 9388 8168
rect 9428 8128 9429 8168
rect 9387 8119 9429 8128
rect 9100 8000 9140 8009
rect 9484 8000 9524 8009
rect 9003 7664 9045 7673
rect 9003 7624 9004 7664
rect 9044 7624 9045 7664
rect 9003 7615 9045 7624
rect 9100 7589 9140 7960
rect 9196 7960 9484 8000
rect 9099 7580 9141 7589
rect 9099 7540 9100 7580
rect 9140 7540 9141 7580
rect 9099 7531 9141 7540
rect 9196 7412 9236 7960
rect 9484 7951 9524 7960
rect 9580 8000 9620 8009
rect 9291 7748 9333 7757
rect 9291 7708 9292 7748
rect 9332 7708 9333 7748
rect 9291 7699 9333 7708
rect 8812 7204 8948 7244
rect 9004 7372 9236 7412
rect 8812 7160 8852 7204
rect 9004 7160 9044 7372
rect 9195 7244 9237 7253
rect 9195 7204 9196 7244
rect 9236 7204 9237 7244
rect 9195 7195 9237 7204
rect 8812 7111 8852 7120
rect 8908 7120 9004 7160
rect 8715 6992 8757 7001
rect 8524 6952 8660 6992
rect 8331 6943 8373 6952
rect 7756 6784 8564 6824
rect 7465 6700 7508 6740
rect 7465 6656 7505 6700
rect 7756 6656 7796 6665
rect 7465 6616 7508 6656
rect 7468 6488 7508 6616
rect 7468 6413 7508 6448
rect 7564 6488 7604 6497
rect 7467 6404 7509 6413
rect 7467 6364 7468 6404
rect 7508 6364 7509 6404
rect 7467 6355 7509 6364
rect 7371 6320 7413 6329
rect 7371 6280 7372 6320
rect 7412 6280 7413 6320
rect 7371 6271 7413 6280
rect 7372 5657 7412 6271
rect 7468 5825 7508 6355
rect 7467 5816 7509 5825
rect 7467 5776 7468 5816
rect 7508 5776 7509 5816
rect 7467 5767 7509 5776
rect 7371 5648 7413 5657
rect 7371 5608 7372 5648
rect 7412 5608 7413 5648
rect 7371 5599 7413 5608
rect 7468 5648 7508 5659
rect 7372 5514 7412 5599
rect 7468 5573 7508 5608
rect 7467 5564 7509 5573
rect 7467 5524 7468 5564
rect 7508 5524 7509 5564
rect 7467 5515 7509 5524
rect 7179 5440 7180 5480
rect 7220 5440 7316 5480
rect 7179 5431 7221 5440
rect 7180 5346 7220 5431
rect 7371 4976 7413 4985
rect 7371 4936 7372 4976
rect 7412 4936 7413 4976
rect 7371 4927 7413 4936
rect 7468 4976 7508 4985
rect 7564 4976 7604 6448
rect 7756 6152 7796 6616
rect 8331 6656 8373 6665
rect 8331 6616 8332 6656
rect 8372 6616 8373 6656
rect 8331 6607 8373 6616
rect 8332 6522 8372 6607
rect 8428 6497 8468 6582
rect 8236 6488 8276 6497
rect 8236 6329 8276 6448
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8331 6404 8373 6413
rect 8331 6364 8332 6404
rect 8372 6364 8373 6404
rect 8331 6355 8373 6364
rect 8235 6320 8277 6329
rect 8235 6280 8236 6320
rect 8276 6280 8277 6320
rect 8235 6271 8277 6280
rect 7756 6112 8276 6152
rect 7659 5648 7701 5657
rect 7659 5608 7660 5648
rect 7700 5608 7701 5648
rect 7659 5599 7701 5608
rect 7756 5648 7796 5657
rect 7660 5514 7700 5599
rect 7756 5573 7796 5608
rect 7947 5648 7989 5657
rect 7947 5608 7948 5648
rect 7988 5608 7989 5648
rect 7947 5599 7989 5608
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8236 5648 8276 6112
rect 8236 5599 8276 5608
rect 7755 5564 7797 5573
rect 7755 5524 7756 5564
rect 7796 5524 7797 5564
rect 7755 5515 7797 5524
rect 7756 5228 7796 5515
rect 7948 5480 7988 5599
rect 8140 5514 8180 5599
rect 8332 5564 8372 6355
rect 8427 6320 8469 6329
rect 8427 6280 8428 6320
rect 8468 6280 8469 6320
rect 8524 6320 8564 6784
rect 8620 6488 8660 6952
rect 8715 6952 8716 6992
rect 8756 6952 8757 6992
rect 8715 6943 8757 6952
rect 8716 6572 8756 6943
rect 8812 6581 8852 6612
rect 8811 6572 8853 6581
rect 8716 6532 8812 6572
rect 8852 6532 8853 6572
rect 8800 6523 8853 6532
rect 8800 6488 8852 6523
rect 8800 6448 8812 6488
rect 8620 6439 8660 6448
rect 8812 6439 8852 6448
rect 8812 6320 8852 6329
rect 8524 6280 8812 6320
rect 8908 6320 8948 7120
rect 9004 7111 9044 7120
rect 9196 7160 9236 7195
rect 9196 7109 9236 7120
rect 9100 7076 9140 7085
rect 9003 6572 9045 6581
rect 9003 6532 9004 6572
rect 9044 6532 9045 6572
rect 9003 6523 9045 6532
rect 9004 6488 9044 6523
rect 9100 6497 9140 7036
rect 9004 6437 9044 6448
rect 9099 6488 9141 6497
rect 9099 6448 9100 6488
rect 9140 6448 9141 6488
rect 9099 6439 9141 6448
rect 9196 6488 9236 6497
rect 9292 6488 9332 7699
rect 9388 7337 9428 7422
rect 9580 7421 9620 7960
rect 9676 8000 9716 8212
rect 9964 8168 10004 8800
rect 10059 8800 10060 8840
rect 10100 8800 10101 8840
rect 10059 8791 10101 8800
rect 9868 8128 10004 8168
rect 9676 7951 9716 7960
rect 9771 8000 9813 8009
rect 9771 7960 9772 8000
rect 9812 7960 9813 8000
rect 9771 7951 9813 7960
rect 9772 7866 9812 7951
rect 9579 7412 9621 7421
rect 9579 7372 9580 7412
rect 9620 7372 9621 7412
rect 9579 7363 9621 7372
rect 9387 7328 9429 7337
rect 9387 7288 9388 7328
rect 9428 7288 9429 7328
rect 9387 7279 9429 7288
rect 9387 7160 9429 7169
rect 9387 7120 9388 7160
rect 9428 7120 9429 7160
rect 9387 7111 9429 7120
rect 9580 7160 9620 7169
rect 9388 7026 9428 7111
rect 9483 6908 9525 6917
rect 9580 6908 9620 7120
rect 9675 7160 9717 7169
rect 9675 7120 9676 7160
rect 9716 7120 9717 7160
rect 9675 7111 9717 7120
rect 9676 7026 9716 7111
rect 9771 6992 9813 7001
rect 9771 6952 9772 6992
rect 9812 6952 9813 6992
rect 9771 6943 9813 6952
rect 9483 6868 9484 6908
rect 9524 6868 9620 6908
rect 9483 6859 9525 6868
rect 9484 6656 9524 6859
rect 9579 6740 9621 6749
rect 9579 6700 9580 6740
rect 9620 6700 9621 6740
rect 9579 6691 9621 6700
rect 9484 6607 9524 6616
rect 9388 6488 9428 6497
rect 9292 6448 9388 6488
rect 9196 6329 9236 6448
rect 9388 6439 9428 6448
rect 9483 6488 9525 6497
rect 9483 6448 9484 6488
rect 9524 6448 9525 6488
rect 9483 6439 9525 6448
rect 9100 6320 9140 6329
rect 8908 6280 9100 6320
rect 8427 6271 8469 6280
rect 8812 6271 8852 6280
rect 9100 6271 9140 6280
rect 9195 6320 9237 6329
rect 9195 6280 9196 6320
rect 9236 6280 9237 6320
rect 9195 6271 9237 6280
rect 8428 6152 8468 6271
rect 9291 6236 9333 6245
rect 9291 6196 9292 6236
rect 9332 6196 9333 6236
rect 9291 6187 9333 6196
rect 8428 6112 8948 6152
rect 8908 5900 8948 6112
rect 8908 5851 8948 5860
rect 9003 5816 9045 5825
rect 9003 5776 9004 5816
rect 9044 5776 9045 5816
rect 9003 5767 9045 5776
rect 8908 5648 8948 5659
rect 8908 5573 8948 5608
rect 9004 5648 9044 5767
rect 9004 5599 9044 5608
rect 9196 5648 9236 5657
rect 7948 5431 7988 5440
rect 7756 5188 7892 5228
rect 7756 4985 7796 5070
rect 7660 4976 7700 4985
rect 7564 4936 7660 4976
rect 6603 4096 6604 4136
rect 6644 4096 6740 4136
rect 6796 4724 6836 4733
rect 6603 4087 6645 4096
rect 5548 4002 5588 4087
rect 5355 3800 5397 3809
rect 5355 3760 5356 3800
rect 5396 3760 5397 3800
rect 5355 3751 5397 3760
rect 5356 3548 5396 3751
rect 5356 3499 5396 3508
rect 6604 3473 6644 4087
rect 6699 3968 6741 3977
rect 6699 3928 6700 3968
rect 6740 3928 6741 3968
rect 6699 3919 6741 3928
rect 6700 3834 6740 3919
rect 6796 3809 6836 4684
rect 6988 3968 7028 3977
rect 6795 3800 6837 3809
rect 6795 3760 6796 3800
rect 6836 3760 6837 3800
rect 6795 3751 6837 3760
rect 5740 3464 5780 3473
rect 6603 3464 6645 3473
rect 5780 3424 5876 3464
rect 5740 3415 5780 3424
rect 4780 3247 4820 3256
rect 651 3128 693 3137
rect 651 3088 652 3128
rect 692 3088 693 3128
rect 651 3079 693 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 5836 2792 5876 3424
rect 6603 3424 6604 3464
rect 6644 3424 6645 3464
rect 6603 3415 6645 3424
rect 6604 3330 6644 3415
rect 5836 2743 5876 2752
rect 843 2708 885 2717
rect 843 2668 844 2708
rect 884 2668 885 2708
rect 843 2659 885 2668
rect 844 2574 884 2659
rect 6988 2624 7028 3928
rect 7372 2876 7412 4927
rect 7468 3977 7508 4936
rect 7660 4136 7700 4936
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 7852 4808 7892 5188
rect 7948 5144 7988 5153
rect 8332 5144 8372 5524
rect 8907 5564 8949 5573
rect 8907 5524 8908 5564
rect 8948 5524 8949 5564
rect 8907 5515 8949 5524
rect 8427 5480 8469 5489
rect 8427 5440 8428 5480
rect 8468 5440 8469 5480
rect 8427 5431 8469 5440
rect 8524 5480 8564 5489
rect 8428 5346 8468 5431
rect 7988 5104 8372 5144
rect 7948 5095 7988 5104
rect 8524 4976 8564 5440
rect 9099 5480 9141 5489
rect 9099 5440 9100 5480
rect 9140 5440 9141 5480
rect 9099 5431 9141 5440
rect 8716 5144 8756 5153
rect 8811 5144 8853 5153
rect 8756 5104 8812 5144
rect 8852 5104 8853 5144
rect 8716 5095 8756 5104
rect 8811 5095 8853 5104
rect 8620 4976 8660 4985
rect 8524 4936 8620 4976
rect 7660 4061 7700 4096
rect 7756 4768 7892 4808
rect 7659 4052 7701 4061
rect 7659 4012 7660 4052
rect 7700 4012 7701 4052
rect 7659 4003 7701 4012
rect 7467 3968 7509 3977
rect 7660 3972 7700 4003
rect 7467 3928 7468 3968
rect 7508 3928 7509 3968
rect 7467 3919 7509 3928
rect 7756 3641 7796 4768
rect 7948 4136 7988 4145
rect 8140 4136 8180 4145
rect 7988 4096 8140 4136
rect 7948 4087 7988 4096
rect 8140 4087 8180 4096
rect 7852 3968 7892 3977
rect 8139 3968 8181 3977
rect 7892 3928 8084 3968
rect 7852 3919 7892 3928
rect 7947 3800 7989 3809
rect 7947 3760 7948 3800
rect 7988 3760 7989 3800
rect 7947 3751 7989 3760
rect 7755 3632 7797 3641
rect 7755 3592 7756 3632
rect 7796 3592 7797 3632
rect 7755 3583 7797 3592
rect 7756 3498 7796 3583
rect 7372 2827 7412 2836
rect 7948 3464 7988 3751
rect 7180 2633 7220 2718
rect 7467 2708 7509 2717
rect 7372 2668 7468 2708
rect 7508 2668 7509 2708
rect 7084 2624 7124 2633
rect 6988 2584 7084 2624
rect 7084 2575 7124 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7372 2624 7412 2668
rect 7467 2659 7509 2668
rect 7564 2633 7604 2718
rect 7372 2575 7412 2584
rect 7563 2624 7605 2633
rect 7563 2584 7564 2624
rect 7604 2584 7605 2624
rect 7563 2575 7605 2584
rect 7660 2624 7700 2633
rect 7948 2624 7988 3424
rect 8044 3464 8084 3928
rect 8139 3928 8140 3968
rect 8180 3928 8181 3968
rect 8139 3919 8181 3928
rect 8140 3632 8180 3919
rect 8140 3583 8180 3592
rect 8235 3548 8277 3557
rect 8235 3508 8236 3548
rect 8276 3508 8277 3548
rect 8235 3499 8277 3508
rect 8044 3415 8084 3424
rect 8236 3464 8276 3499
rect 8620 3464 8660 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 8716 4842 8756 4927
rect 8811 4892 8853 4901
rect 9100 4892 9140 5431
rect 9196 5153 9236 5608
rect 9292 5648 9332 6187
rect 9292 5599 9332 5608
rect 9392 5648 9434 5657
rect 9392 5608 9393 5648
rect 9433 5608 9434 5648
rect 9392 5599 9434 5608
rect 9393 5514 9433 5599
rect 9484 5564 9524 6439
rect 9580 5648 9620 6691
rect 9772 6488 9812 6943
rect 9772 6439 9812 6448
rect 9675 6320 9717 6329
rect 9675 6280 9676 6320
rect 9716 6280 9717 6320
rect 9675 6271 9717 6280
rect 9676 6186 9716 6271
rect 9868 5825 9908 8128
rect 9963 8000 10005 8009
rect 9963 7960 9964 8000
rect 10004 7960 10005 8000
rect 9963 7951 10005 7960
rect 9964 7866 10004 7951
rect 10060 6749 10100 8791
rect 10156 8345 10196 9472
rect 10252 9462 10292 9547
rect 10636 9512 10676 9808
rect 10636 9463 10676 9472
rect 10251 8756 10293 8765
rect 10251 8716 10252 8756
rect 10292 8716 10293 8756
rect 10251 8707 10293 8716
rect 10635 8756 10677 8765
rect 10635 8716 10636 8756
rect 10676 8716 10677 8756
rect 10635 8707 10677 8716
rect 10155 8336 10197 8345
rect 10155 8296 10156 8336
rect 10196 8296 10197 8336
rect 10155 8287 10197 8296
rect 10156 8000 10196 8009
rect 10156 7832 10196 7960
rect 10252 8000 10292 8707
rect 10444 8672 10484 8681
rect 10252 7951 10292 7960
rect 10348 8632 10444 8672
rect 10348 7832 10388 8632
rect 10444 8623 10484 8632
rect 10540 8672 10580 8681
rect 10540 8009 10580 8632
rect 10636 8672 10676 8707
rect 10732 8681 10772 9892
rect 10924 9605 10964 9976
rect 10923 9596 10965 9605
rect 10923 9556 10924 9596
rect 10964 9556 10965 9596
rect 10923 9547 10965 9556
rect 11404 8840 11444 10144
rect 11596 10135 11636 10144
rect 11692 10109 11732 11656
rect 11788 11696 11828 11705
rect 11788 11453 11828 11656
rect 11883 11696 11925 11705
rect 11883 11656 11884 11696
rect 11924 11656 11925 11696
rect 11883 11647 11925 11656
rect 11884 11562 11924 11647
rect 11787 11444 11829 11453
rect 11787 11404 11788 11444
rect 11828 11404 11829 11444
rect 11787 11395 11829 11404
rect 11980 10184 12020 11824
rect 12171 11824 12172 11864
rect 12212 11824 12213 11864
rect 12171 11815 12213 11824
rect 12076 11696 12116 11705
rect 12116 11656 12212 11696
rect 12076 11647 12116 11656
rect 12075 11528 12117 11537
rect 12075 11488 12076 11528
rect 12116 11488 12117 11528
rect 12075 11479 12117 11488
rect 11980 10135 12020 10144
rect 11691 10100 11733 10109
rect 11691 10060 11692 10100
rect 11732 10060 11733 10100
rect 11691 10051 11733 10060
rect 12076 10100 12116 11479
rect 12172 11201 12212 11656
rect 12268 11453 12308 12235
rect 12267 11444 12309 11453
rect 12267 11404 12268 11444
rect 12308 11404 12309 11444
rect 12267 11395 12309 11404
rect 12171 11192 12213 11201
rect 12171 11152 12172 11192
rect 12212 11152 12213 11192
rect 12171 11143 12213 11152
rect 12172 10193 12212 10278
rect 12171 10184 12213 10193
rect 12171 10144 12172 10184
rect 12212 10144 12213 10184
rect 12171 10135 12213 10144
rect 12268 10184 12308 11395
rect 12460 11024 12500 12991
rect 12844 11948 12884 13159
rect 12940 12965 12980 13327
rect 12939 12956 12981 12965
rect 12939 12916 12940 12956
rect 12980 12916 12981 12956
rect 12939 12907 12981 12916
rect 12939 12620 12981 12629
rect 12939 12580 12940 12620
rect 12980 12580 12981 12620
rect 12939 12571 12981 12580
rect 13611 12620 13653 12629
rect 13611 12580 13612 12620
rect 13652 12580 13653 12620
rect 13611 12571 13653 12580
rect 12940 12536 12980 12571
rect 12940 12485 12980 12496
rect 13612 12486 13652 12571
rect 12940 11948 12980 11957
rect 12844 11908 12940 11948
rect 12940 11899 12980 11908
rect 13035 11696 13077 11705
rect 13035 11656 13036 11696
rect 13076 11656 13077 11696
rect 13035 11647 13077 11656
rect 13228 11696 13268 11705
rect 13036 11562 13076 11647
rect 13228 11537 13268 11656
rect 13323 11612 13365 11621
rect 13323 11572 13324 11612
rect 13364 11572 13365 11612
rect 13323 11563 13365 11572
rect 12748 11528 12788 11537
rect 12748 11360 12788 11488
rect 13227 11528 13269 11537
rect 13227 11488 13228 11528
rect 13268 11488 13269 11528
rect 13227 11479 13269 11488
rect 12748 11320 12884 11360
rect 12460 10975 12500 10984
rect 12844 10856 12884 11320
rect 13324 11024 13364 11563
rect 13900 11528 13940 11537
rect 13900 11360 13940 11488
rect 13708 11320 13940 11360
rect 13708 11108 13748 11320
rect 13708 11059 13748 11068
rect 13324 10975 13364 10984
rect 13899 11024 13941 11033
rect 13899 10984 13900 11024
rect 13940 10984 13941 11024
rect 13899 10975 13941 10984
rect 13900 10890 13940 10975
rect 12844 10816 13364 10856
rect 13132 10184 13172 10193
rect 12076 10051 12116 10060
rect 11979 10016 12021 10025
rect 11979 9976 11980 10016
rect 12020 9976 12021 10016
rect 11979 9967 12021 9976
rect 11404 8791 11444 8800
rect 11500 9512 11540 9521
rect 10636 8621 10676 8632
rect 10731 8672 10773 8681
rect 10731 8632 10732 8672
rect 10772 8632 10773 8672
rect 10731 8623 10773 8632
rect 11403 8672 11445 8681
rect 11403 8632 11404 8672
rect 11444 8632 11445 8672
rect 11403 8623 11445 8632
rect 11404 8538 11444 8623
rect 10732 8504 10772 8513
rect 10539 8000 10581 8009
rect 10539 7960 10540 8000
rect 10580 7960 10581 8000
rect 10732 8000 10772 8464
rect 10827 8336 10869 8345
rect 10827 8296 10828 8336
rect 10868 8296 10869 8336
rect 10827 8287 10869 8296
rect 10828 8168 10868 8287
rect 10828 8119 10868 8128
rect 11115 8084 11157 8093
rect 11115 8044 11116 8084
rect 11156 8044 11157 8084
rect 11115 8035 11157 8044
rect 10828 8000 10868 8009
rect 10732 7960 10828 8000
rect 10539 7951 10581 7960
rect 10828 7951 10868 7960
rect 10924 8000 10964 8009
rect 10156 7792 10388 7832
rect 10444 7832 10484 7841
rect 10924 7832 10964 7960
rect 11116 7950 11156 8035
rect 10484 7792 10964 7832
rect 10156 6833 10196 7792
rect 10444 7783 10484 7792
rect 11500 7589 11540 9472
rect 11596 8672 11636 8683
rect 11596 8597 11636 8632
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 11980 8672 12020 9967
rect 11980 8623 12020 8632
rect 12172 8840 12212 8849
rect 11595 8588 11637 8597
rect 11595 8548 11596 8588
rect 11636 8548 11637 8588
rect 11595 8539 11637 8548
rect 11692 8538 11732 8623
rect 11883 8588 11925 8597
rect 11883 8548 11884 8588
rect 11924 8548 11925 8588
rect 11883 8539 11925 8548
rect 11884 8454 11924 8539
rect 11691 8084 11733 8093
rect 11691 8044 11692 8084
rect 11732 8044 11733 8084
rect 11691 8035 11733 8044
rect 11692 7950 11732 8035
rect 12076 8000 12116 8009
rect 12172 8000 12212 8800
rect 12268 8681 12308 10144
rect 12652 10144 13132 10184
rect 12459 10016 12501 10025
rect 12459 9976 12460 10016
rect 12500 9976 12501 10016
rect 12459 9967 12501 9976
rect 12460 9882 12500 9967
rect 12652 9680 12692 10144
rect 13132 10135 13172 10144
rect 13324 10184 13364 10816
rect 13996 10436 14036 13504
rect 14092 13208 14132 13217
rect 14092 13049 14132 13168
rect 14380 13124 14420 13756
rect 14476 13747 14516 13756
rect 14188 13084 14420 13124
rect 14091 13040 14133 13049
rect 14091 13000 14092 13040
rect 14132 13000 14133 13040
rect 14091 12991 14133 13000
rect 14091 11864 14133 11873
rect 14091 11824 14092 11864
rect 14132 11824 14133 11864
rect 14091 11815 14133 11824
rect 14092 11696 14132 11815
rect 14092 11647 14132 11656
rect 14188 11696 14228 13084
rect 14860 12536 14900 14764
rect 14956 14720 14996 15259
rect 14956 14671 14996 14680
rect 15148 13880 15188 15520
rect 15244 15511 15284 15520
rect 15340 15224 15380 16351
rect 15627 15560 15669 15569
rect 15627 15520 15628 15560
rect 15668 15520 15669 15560
rect 15627 15511 15669 15520
rect 15628 15426 15668 15511
rect 15244 15184 15380 15224
rect 15244 14720 15284 15184
rect 15435 15140 15477 15149
rect 15435 15100 15436 15140
rect 15476 15100 15477 15140
rect 15435 15091 15477 15100
rect 15244 14141 15284 14680
rect 15340 14720 15380 14731
rect 15340 14645 15380 14680
rect 15339 14636 15381 14645
rect 15339 14596 15340 14636
rect 15380 14596 15381 14636
rect 15339 14587 15381 14596
rect 15436 14636 15476 15091
rect 15724 15065 15764 19804
rect 15819 19795 15861 19804
rect 16300 19844 16340 19853
rect 16300 19760 16340 19804
rect 16395 19760 16437 19769
rect 16300 19720 16396 19760
rect 16436 19720 16437 19760
rect 16395 19711 16437 19720
rect 16107 19256 16149 19265
rect 16107 19216 16108 19256
rect 16148 19216 16149 19256
rect 16107 19207 16149 19216
rect 16108 19122 16148 19207
rect 15915 19088 15957 19097
rect 15915 19048 15916 19088
rect 15956 19048 15957 19088
rect 15915 19039 15957 19048
rect 15916 18584 15956 19039
rect 16492 18584 16532 20896
rect 17068 20936 17108 21568
rect 17836 21559 17876 21568
rect 18891 21608 18933 21617
rect 18891 21568 18892 21608
rect 18932 21568 18933 21608
rect 18891 21559 18933 21568
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 17068 20887 17108 20896
rect 17068 20224 17300 20264
rect 16971 19928 17013 19937
rect 16971 19888 16972 19928
rect 17012 19888 17013 19928
rect 16971 19879 17013 19888
rect 16972 19794 17012 19879
rect 16972 19172 17012 19181
rect 16780 19088 16820 19097
rect 16820 19048 16916 19088
rect 16780 19039 16820 19048
rect 16780 18584 16820 18593
rect 15956 18544 16052 18584
rect 16492 18544 16780 18584
rect 15916 18535 15956 18544
rect 16012 17744 16052 18544
rect 16780 18535 16820 18544
rect 16012 17695 16052 17704
rect 16299 17660 16341 17669
rect 16299 17620 16300 17660
rect 16340 17620 16341 17660
rect 16299 17611 16341 17620
rect 16107 17492 16149 17501
rect 16107 17452 16108 17492
rect 16148 17452 16149 17492
rect 16107 17443 16149 17452
rect 16011 17240 16053 17249
rect 16011 17200 16012 17240
rect 16052 17200 16053 17240
rect 16011 17191 16053 17200
rect 16012 17156 16052 17191
rect 16012 17105 16052 17116
rect 15915 17072 15957 17081
rect 15915 17032 15916 17072
rect 15956 17032 15957 17072
rect 15915 17023 15957 17032
rect 16108 17072 16148 17443
rect 16300 17240 16340 17611
rect 16300 17191 16340 17200
rect 16108 17023 16148 17032
rect 16779 17072 16821 17081
rect 16779 17032 16780 17072
rect 16820 17032 16821 17072
rect 16779 17023 16821 17032
rect 15916 16938 15956 17023
rect 16204 16400 16244 16409
rect 16588 16400 16628 16409
rect 16244 16360 16436 16400
rect 16204 16351 16244 16360
rect 16396 16316 16436 16360
rect 16396 16267 16436 16276
rect 16012 16232 16052 16243
rect 16588 16241 16628 16360
rect 16012 16157 16052 16192
rect 16204 16232 16244 16241
rect 16011 16148 16053 16157
rect 16011 16108 16012 16148
rect 16052 16108 16053 16148
rect 16011 16099 16053 16108
rect 16204 15569 16244 16192
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16780 16232 16820 17023
rect 16780 16183 16820 16192
rect 16876 16232 16916 19048
rect 16972 18761 17012 19132
rect 16971 18752 17013 18761
rect 16971 18712 16972 18752
rect 17012 18712 17013 18752
rect 16971 18703 17013 18712
rect 16971 17576 17013 17585
rect 16971 17536 16972 17576
rect 17012 17536 17013 17576
rect 16971 17527 17013 17536
rect 16972 17072 17012 17527
rect 16972 17023 17012 17032
rect 16971 16316 17013 16325
rect 16971 16276 16972 16316
rect 17012 16276 17013 16316
rect 16971 16267 17013 16276
rect 16395 16148 16437 16157
rect 16395 16108 16396 16148
rect 16436 16108 16437 16148
rect 16395 16099 16437 16108
rect 15819 15560 15861 15569
rect 15819 15520 15820 15560
rect 15860 15520 15861 15560
rect 15819 15511 15861 15520
rect 16203 15560 16245 15569
rect 16203 15520 16204 15560
rect 16244 15520 16245 15560
rect 16203 15511 16245 15520
rect 15820 15426 15860 15511
rect 15723 15056 15765 15065
rect 15723 15016 15724 15056
rect 15764 15016 15765 15056
rect 15723 15007 15765 15016
rect 15724 14729 15764 14814
rect 15436 14587 15476 14596
rect 15532 14720 15572 14729
rect 15532 14216 15572 14680
rect 15723 14720 15765 14729
rect 15723 14680 15724 14720
rect 15764 14680 15765 14720
rect 15723 14671 15765 14680
rect 16204 14720 16244 14729
rect 15819 14636 15861 14645
rect 15819 14596 15820 14636
rect 15860 14596 15861 14636
rect 15819 14587 15861 14596
rect 15820 14502 15860 14587
rect 15628 14216 15668 14225
rect 15532 14176 15628 14216
rect 15628 14167 15668 14176
rect 15243 14132 15285 14141
rect 15243 14092 15244 14132
rect 15284 14092 15285 14132
rect 15243 14083 15285 14092
rect 15819 14132 15861 14141
rect 15819 14092 15820 14132
rect 15860 14092 15861 14132
rect 15819 14083 15861 14092
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 15820 14048 15860 14083
rect 16204 14057 16244 14680
rect 16299 14720 16341 14729
rect 16299 14680 16300 14720
rect 16340 14680 16341 14720
rect 16396 14720 16436 16099
rect 16876 16064 16916 16192
rect 16972 16232 17012 16267
rect 16972 16181 17012 16192
rect 17068 16232 17108 20224
rect 17164 20096 17204 20105
rect 17164 19256 17204 20056
rect 17260 20096 17300 20224
rect 17260 20047 17300 20056
rect 17452 20096 17492 20107
rect 17452 20021 17492 20056
rect 17547 20096 17589 20105
rect 17547 20056 17548 20096
rect 17588 20056 17589 20096
rect 17547 20047 17589 20056
rect 18315 20096 18357 20105
rect 18315 20056 18316 20096
rect 18356 20056 18357 20096
rect 18315 20047 18357 20056
rect 17451 20012 17493 20021
rect 17451 19972 17452 20012
rect 17492 19972 17493 20012
rect 17451 19963 17493 19972
rect 17355 19928 17397 19937
rect 17355 19888 17356 19928
rect 17396 19888 17397 19928
rect 17355 19879 17397 19888
rect 17356 19256 17396 19879
rect 17164 19216 17300 19256
rect 17163 19004 17205 19013
rect 17163 18964 17164 19004
rect 17204 18964 17205 19004
rect 17163 18955 17205 18964
rect 17164 18668 17204 18955
rect 17260 18845 17300 19216
rect 17356 19207 17396 19216
rect 17452 19844 17492 19853
rect 17452 18929 17492 19804
rect 17451 18920 17493 18929
rect 17451 18880 17452 18920
rect 17492 18880 17493 18920
rect 17451 18871 17493 18880
rect 17259 18836 17301 18845
rect 17259 18796 17260 18836
rect 17300 18796 17301 18836
rect 17259 18787 17301 18796
rect 17355 18752 17397 18761
rect 17355 18712 17356 18752
rect 17396 18712 17397 18752
rect 17355 18703 17397 18712
rect 17164 18619 17204 18628
rect 17356 18618 17396 18703
rect 17548 18500 17588 20047
rect 18316 19962 18356 20047
rect 18795 20012 18837 20021
rect 18795 19972 18796 20012
rect 18836 19972 18837 20012
rect 18795 19963 18837 19972
rect 18796 19878 18836 19963
rect 18892 19937 18932 21559
rect 18987 20600 19029 20609
rect 18987 20560 18988 20600
rect 19028 20560 19029 20600
rect 18987 20551 19029 20560
rect 18988 20264 19028 20551
rect 18988 20215 19028 20224
rect 19180 20096 19220 20105
rect 19180 19937 19220 20056
rect 19276 20096 19316 20105
rect 18891 19928 18933 19937
rect 19179 19928 19221 19937
rect 18891 19888 18892 19928
rect 18932 19888 19028 19928
rect 18891 19879 18933 19888
rect 17644 19844 17684 19853
rect 17644 19013 17684 19804
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 18219 19256 18261 19265
rect 18219 19216 18220 19256
rect 18260 19216 18261 19256
rect 18219 19207 18261 19216
rect 18220 19122 18260 19207
rect 17643 19004 17685 19013
rect 17643 18964 17644 19004
rect 17684 18964 17685 19004
rect 17643 18955 17685 18964
rect 18027 18920 18069 18929
rect 18027 18880 18028 18920
rect 18068 18880 18069 18920
rect 18027 18871 18069 18880
rect 17643 18584 17685 18593
rect 17643 18544 17644 18584
rect 17684 18544 17685 18584
rect 17643 18535 17685 18544
rect 18028 18584 18068 18871
rect 18892 18584 18932 18593
rect 18028 18535 18068 18544
rect 18700 18544 18892 18584
rect 17356 18460 17588 18500
rect 17163 17828 17205 17837
rect 17163 17788 17164 17828
rect 17204 17788 17205 17828
rect 17163 17779 17205 17788
rect 17164 17694 17204 17779
rect 17356 17744 17396 18460
rect 17451 18332 17493 18341
rect 17451 18292 17452 18332
rect 17492 18292 17493 18332
rect 17451 18283 17493 18292
rect 17356 17695 17396 17704
rect 17452 17744 17492 18283
rect 17547 17912 17589 17921
rect 17547 17872 17548 17912
rect 17588 17872 17589 17912
rect 17547 17863 17589 17872
rect 17452 17695 17492 17704
rect 17548 17744 17588 17863
rect 17548 17695 17588 17704
rect 17644 17744 17684 18535
rect 18220 18341 18260 18426
rect 18219 18332 18261 18341
rect 18219 18292 18220 18332
rect 18260 18292 18261 18332
rect 18219 18283 18261 18292
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 18700 17912 18740 18544
rect 18892 18535 18932 18544
rect 18988 18341 19028 19888
rect 19179 19888 19180 19928
rect 19220 19888 19221 19928
rect 19179 19879 19221 19888
rect 19276 19013 19316 20056
rect 19372 19265 19412 23080
rect 19659 23071 19701 23080
rect 19660 22986 19700 23071
rect 19755 22448 19797 22457
rect 19755 22408 19756 22448
rect 19796 22408 19797 22448
rect 19755 22399 19797 22408
rect 20331 22448 20373 22457
rect 20331 22408 20332 22448
rect 20372 22408 20373 22448
rect 20331 22399 20373 22408
rect 19756 22314 19796 22399
rect 20332 22280 20372 22399
rect 20332 22231 20372 22240
rect 21195 22280 21237 22289
rect 21195 22240 21196 22280
rect 21236 22240 21237 22280
rect 21195 22231 21237 22240
rect 19948 22196 19988 22205
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 19468 21776 19508 21785
rect 19948 21776 19988 22156
rect 21196 22146 21236 22231
rect 21291 22112 21333 22121
rect 21291 22072 21292 22112
rect 21332 22072 21333 22112
rect 21291 22063 21333 22072
rect 19508 21736 19988 21776
rect 19468 21727 19508 21736
rect 21004 21608 21044 21617
rect 21196 21608 21236 21617
rect 21044 21568 21196 21608
rect 21004 21559 21044 21568
rect 21196 21559 21236 21568
rect 21292 21608 21332 22063
rect 21484 21785 21524 23416
rect 21579 23407 21621 23416
rect 21676 23129 21716 26095
rect 21964 26069 22004 26104
rect 22156 26144 22196 26431
rect 22156 26095 22196 26104
rect 21963 26060 22005 26069
rect 21963 26020 21964 26060
rect 22004 26020 22005 26060
rect 21963 26011 22005 26020
rect 22251 26060 22293 26069
rect 22251 26020 22252 26060
rect 22292 26020 22293 26060
rect 22251 26011 22293 26020
rect 22059 25892 22101 25901
rect 22059 25852 22060 25892
rect 22100 25852 22101 25892
rect 22059 25843 22101 25852
rect 22060 25758 22100 25843
rect 22155 25640 22197 25649
rect 22155 25600 22156 25640
rect 22196 25600 22197 25640
rect 22155 25591 22197 25600
rect 21771 25472 21813 25481
rect 21771 25432 21772 25472
rect 21812 25432 21813 25472
rect 21771 25423 21813 25432
rect 21772 24632 21812 25423
rect 22156 25304 22196 25591
rect 22156 25255 22196 25264
rect 22252 25339 22292 26011
rect 22540 25985 22580 26776
rect 22924 26732 22964 26741
rect 22924 26321 22964 26692
rect 22923 26312 22965 26321
rect 22923 26272 22924 26312
rect 22964 26272 22965 26312
rect 22923 26263 22965 26272
rect 23596 26144 23636 26153
rect 22635 26060 22677 26069
rect 22635 26020 22636 26060
rect 22676 26020 22677 26060
rect 22635 26011 22677 26020
rect 22539 25976 22581 25985
rect 22539 25936 22540 25976
rect 22580 25936 22581 25976
rect 22539 25927 22581 25936
rect 22347 25472 22389 25481
rect 22347 25432 22348 25472
rect 22388 25432 22389 25472
rect 22347 25423 22389 25432
rect 22636 25472 22676 26011
rect 23596 25565 23636 26104
rect 23595 25556 23637 25565
rect 23595 25516 23596 25556
rect 23636 25516 23637 25556
rect 23595 25507 23637 25516
rect 22636 25423 22676 25432
rect 21868 25136 21908 25145
rect 22155 25136 22197 25145
rect 21908 25096 22100 25136
rect 21868 25087 21908 25096
rect 21867 24884 21909 24893
rect 21867 24844 21868 24884
rect 21908 24844 21909 24884
rect 21867 24835 21909 24844
rect 21772 24583 21812 24592
rect 21868 24627 21908 24835
rect 21868 24578 21908 24587
rect 21964 24632 22004 24641
rect 21964 24473 22004 24592
rect 21963 24464 22005 24473
rect 21963 24424 21964 24464
rect 22004 24424 22005 24464
rect 21963 24415 22005 24424
rect 21771 24380 21813 24389
rect 21771 24340 21772 24380
rect 21812 24340 21813 24380
rect 21771 24331 21813 24340
rect 21675 23120 21717 23129
rect 21675 23080 21676 23120
rect 21716 23080 21717 23120
rect 21675 23071 21717 23080
rect 21483 21776 21525 21785
rect 21483 21736 21484 21776
rect 21524 21736 21525 21776
rect 21483 21727 21525 21736
rect 21292 21559 21332 21568
rect 21388 21608 21428 21617
rect 20140 21549 20180 21558
rect 19948 21509 20140 21524
rect 19948 21484 20180 21509
rect 19948 20852 19988 21484
rect 20332 21440 20372 21449
rect 19948 20803 19988 20812
rect 20044 21400 20332 21440
rect 19852 20768 19892 20777
rect 19852 20600 19892 20728
rect 20044 20768 20084 21400
rect 20332 21391 20372 21400
rect 21291 21020 21333 21029
rect 21388 21020 21428 21568
rect 21484 21608 21524 21617
rect 21484 21449 21524 21568
rect 21483 21440 21525 21449
rect 21483 21400 21484 21440
rect 21524 21400 21525 21440
rect 21483 21391 21525 21400
rect 21675 21440 21717 21449
rect 21675 21400 21676 21440
rect 21716 21400 21717 21440
rect 21675 21391 21717 21400
rect 21291 20980 21292 21020
rect 21332 20980 21428 21020
rect 21291 20971 21333 20980
rect 20044 20719 20084 20728
rect 20523 20768 20565 20777
rect 20523 20728 20524 20768
rect 20564 20728 20565 20768
rect 20523 20719 20565 20728
rect 20620 20768 20660 20777
rect 20524 20634 20564 20719
rect 19852 20560 19911 20600
rect 19871 20516 19911 20560
rect 20620 20525 20660 20728
rect 21292 20609 21332 20971
rect 21387 20768 21429 20777
rect 21484 20768 21524 21391
rect 21676 21306 21716 21391
rect 21580 20782 21620 20863
rect 21675 20852 21717 20861
rect 21675 20812 21676 20852
rect 21716 20812 21720 20852
rect 21675 20803 21720 20812
rect 21387 20728 21388 20768
rect 21428 20728 21524 20768
rect 21579 20728 21580 20777
rect 21680 20787 21720 20803
rect 21620 20728 21621 20777
rect 21387 20719 21429 20728
rect 21579 20719 21621 20728
rect 20812 20600 20852 20609
rect 21291 20600 21333 20609
rect 20852 20560 21236 20600
rect 20812 20551 20852 20560
rect 20619 20516 20661 20525
rect 19871 20476 19988 20516
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 19948 20180 19988 20476
rect 20619 20476 20620 20516
rect 20660 20476 20661 20516
rect 20619 20467 20661 20476
rect 20907 20432 20949 20441
rect 20907 20392 20908 20432
rect 20948 20392 20949 20432
rect 20907 20383 20949 20392
rect 19564 20140 19988 20180
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19468 19962 19508 20047
rect 19468 19844 19508 19853
rect 19564 19844 19604 20140
rect 20332 20096 20372 20105
rect 19659 20012 19701 20021
rect 19659 19972 19660 20012
rect 19700 19972 19701 20012
rect 19659 19963 19701 19972
rect 19508 19804 19604 19844
rect 19468 19795 19508 19804
rect 19371 19256 19413 19265
rect 19371 19216 19372 19256
rect 19412 19216 19413 19256
rect 19371 19207 19413 19216
rect 19660 19256 19700 19963
rect 19660 19207 19700 19216
rect 20332 19097 20372 20056
rect 20908 19508 20948 20383
rect 21196 20096 21236 20560
rect 21291 20560 21292 20600
rect 21332 20560 21333 20600
rect 21291 20551 21333 20560
rect 21388 20357 21428 20719
rect 21680 20684 21720 20747
rect 21675 20644 21720 20684
rect 21483 20600 21525 20609
rect 21483 20560 21484 20600
rect 21524 20560 21525 20600
rect 21675 20600 21715 20644
rect 21675 20560 21716 20600
rect 21483 20551 21525 20560
rect 21484 20466 21524 20551
rect 21387 20348 21429 20357
rect 21387 20308 21388 20348
rect 21428 20308 21429 20348
rect 21387 20299 21429 20308
rect 21676 20273 21716 20560
rect 21772 20516 21812 24331
rect 22060 22616 22100 25096
rect 22155 25096 22156 25136
rect 22196 25096 22197 25136
rect 22155 25087 22197 25096
rect 22156 24557 22196 25087
rect 22252 24893 22292 25299
rect 22348 25304 22388 25423
rect 23499 25388 23541 25397
rect 23499 25348 23500 25388
rect 23540 25348 23541 25388
rect 23499 25339 23541 25348
rect 22348 25255 22388 25264
rect 22732 25304 22772 25313
rect 22732 25145 22772 25264
rect 23500 25304 23540 25339
rect 23596 25313 23636 25399
rect 23500 25253 23540 25264
rect 23595 25309 23637 25313
rect 23595 25264 23596 25309
rect 23636 25264 23637 25309
rect 23595 25255 23637 25264
rect 23692 25304 23732 25313
rect 22731 25136 22773 25145
rect 22731 25096 22732 25136
rect 22772 25096 22773 25136
rect 22731 25087 22773 25096
rect 23212 25136 23252 25145
rect 22251 24884 22293 24893
rect 22251 24844 22252 24884
rect 22292 24844 22293 24884
rect 22251 24835 22293 24844
rect 22251 24632 22293 24641
rect 22251 24592 22252 24632
rect 22292 24592 22293 24632
rect 22251 24583 22293 24592
rect 22155 24548 22197 24557
rect 22155 24508 22156 24548
rect 22196 24508 22197 24548
rect 22155 24499 22197 24508
rect 22156 23288 22196 24499
rect 22252 24498 22292 24583
rect 23116 24548 23156 24557
rect 23019 23876 23061 23885
rect 23019 23836 23020 23876
rect 23060 23836 23061 23876
rect 23019 23827 23061 23836
rect 23020 23792 23060 23827
rect 23020 23741 23060 23752
rect 22156 23239 22196 23248
rect 22540 23120 22580 23129
rect 22924 23120 22964 23129
rect 22348 23080 22540 23120
rect 22060 22576 22292 22616
rect 21867 22112 21909 22121
rect 21867 22072 21868 22112
rect 21908 22072 21909 22112
rect 21867 22063 21909 22072
rect 21868 21524 21908 22063
rect 21868 21475 21908 21484
rect 22059 21020 22101 21029
rect 22059 20980 22060 21020
rect 22100 20980 22101 21020
rect 22059 20971 22101 20980
rect 21868 20768 21908 20779
rect 21868 20693 21908 20728
rect 21964 20768 22004 20777
rect 21867 20684 21909 20693
rect 21867 20644 21868 20684
rect 21908 20644 21909 20684
rect 21867 20635 21909 20644
rect 21772 20476 21908 20516
rect 21771 20348 21813 20357
rect 21771 20308 21772 20348
rect 21812 20308 21813 20348
rect 21771 20299 21813 20308
rect 21483 20264 21525 20273
rect 21483 20224 21484 20264
rect 21524 20224 21525 20264
rect 21483 20215 21525 20224
rect 21675 20264 21717 20273
rect 21675 20224 21676 20264
rect 21716 20224 21717 20264
rect 21675 20215 21717 20224
rect 21196 20047 21236 20056
rect 21292 20096 21332 20105
rect 21003 20012 21045 20021
rect 21003 19972 21004 20012
rect 21044 19972 21045 20012
rect 21003 19963 21045 19972
rect 21004 19878 21044 19963
rect 20908 19459 20948 19468
rect 21292 19349 21332 20056
rect 21484 19844 21524 20215
rect 21772 20096 21812 20299
rect 21772 20047 21812 20056
rect 21772 19844 21812 19853
rect 21484 19804 21620 19844
rect 21484 19424 21524 19433
rect 21291 19340 21333 19349
rect 21291 19300 21292 19340
rect 21332 19300 21333 19340
rect 21291 19291 21333 19300
rect 20812 19256 20852 19265
rect 20524 19172 20564 19181
rect 19371 19088 19413 19097
rect 19371 19048 19372 19088
rect 19412 19048 19413 19088
rect 19371 19039 19413 19048
rect 20331 19088 20373 19097
rect 20331 19048 20332 19088
rect 20372 19048 20373 19088
rect 20331 19039 20373 19048
rect 19275 19004 19317 19013
rect 19275 18964 19276 19004
rect 19316 18964 19317 19004
rect 19275 18955 19317 18964
rect 19372 18954 19412 19039
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 19084 18761 19124 18846
rect 19083 18752 19125 18761
rect 19083 18712 19084 18752
rect 19124 18712 19125 18752
rect 19083 18703 19125 18712
rect 19084 18584 19124 18595
rect 19084 18509 19124 18544
rect 19275 18584 19317 18593
rect 19275 18544 19276 18584
rect 19316 18544 19317 18584
rect 19275 18535 19317 18544
rect 19372 18584 19412 18593
rect 19564 18584 19604 18593
rect 19412 18544 19564 18584
rect 19083 18500 19125 18509
rect 19083 18460 19084 18500
rect 19124 18460 19125 18500
rect 19083 18451 19125 18460
rect 18987 18332 19029 18341
rect 18987 18292 18988 18332
rect 19028 18292 19029 18332
rect 18987 18283 19029 18292
rect 18988 18005 19028 18090
rect 18987 17996 19029 18005
rect 18987 17956 18988 17996
rect 19028 17956 19029 17996
rect 18987 17947 19029 17956
rect 18604 17872 18740 17912
rect 17739 17828 17781 17837
rect 17739 17788 17740 17828
rect 17780 17788 17781 17828
rect 17739 17779 17781 17788
rect 17644 17695 17684 17704
rect 17355 17492 17397 17501
rect 17355 17452 17356 17492
rect 17396 17452 17397 17492
rect 17355 17443 17397 17452
rect 17163 17072 17205 17081
rect 17163 17032 17164 17072
rect 17204 17032 17205 17072
rect 17163 17023 17205 17032
rect 17164 16938 17204 17023
rect 17068 16183 17108 16192
rect 17260 16232 17300 16241
rect 17260 16064 17300 16192
rect 17356 16232 17396 17443
rect 17451 17324 17493 17333
rect 17451 17284 17452 17324
rect 17492 17284 17493 17324
rect 17451 17275 17493 17284
rect 17452 16232 17492 17275
rect 17740 17072 17780 17779
rect 17836 17744 17876 17753
rect 17836 17249 17876 17704
rect 18507 17744 18549 17753
rect 18507 17704 18508 17744
rect 18548 17704 18549 17744
rect 18507 17695 18549 17704
rect 18123 17660 18165 17669
rect 18123 17620 18124 17660
rect 18164 17620 18165 17660
rect 18123 17611 18165 17620
rect 18411 17660 18453 17669
rect 18411 17620 18412 17660
rect 18452 17620 18453 17660
rect 18411 17611 18453 17620
rect 18027 17408 18069 17417
rect 18027 17368 18028 17408
rect 18068 17368 18069 17408
rect 18027 17359 18069 17368
rect 17835 17240 17877 17249
rect 17835 17200 17836 17240
rect 17876 17200 17877 17240
rect 17835 17191 17877 17200
rect 17836 17072 17876 17081
rect 17740 17032 17836 17072
rect 17836 17023 17876 17032
rect 18028 17072 18068 17359
rect 17547 16820 17589 16829
rect 17547 16780 17548 16820
rect 17588 16780 17589 16820
rect 17547 16771 17589 16780
rect 17548 16400 17588 16771
rect 17548 16351 17588 16360
rect 18028 16241 18068 17032
rect 18124 17072 18164 17611
rect 18315 17240 18357 17249
rect 18315 17200 18316 17240
rect 18356 17200 18357 17240
rect 18315 17191 18357 17200
rect 18412 17240 18452 17611
rect 18508 17610 18548 17695
rect 18412 17191 18452 17200
rect 18220 17156 18260 17167
rect 18220 17081 18260 17116
rect 18316 17106 18356 17191
rect 18124 16997 18164 17032
rect 18219 17072 18261 17081
rect 18219 17032 18220 17072
rect 18260 17032 18261 17072
rect 18219 17023 18261 17032
rect 18123 16988 18165 16997
rect 18123 16948 18124 16988
rect 18164 16948 18165 16988
rect 18123 16939 18165 16948
rect 18604 16829 18644 17872
rect 18795 17828 18837 17837
rect 18795 17788 18796 17828
rect 18836 17788 18837 17828
rect 18795 17779 18837 17788
rect 18987 17828 19029 17837
rect 18987 17788 18988 17828
rect 19028 17788 19029 17828
rect 18987 17779 19029 17788
rect 18700 17744 18740 17753
rect 18700 17417 18740 17704
rect 18796 17744 18836 17779
rect 18796 17693 18836 17704
rect 18988 17744 19028 17779
rect 18699 17408 18741 17417
rect 18699 17368 18700 17408
rect 18740 17368 18741 17408
rect 18699 17359 18741 17368
rect 18699 17240 18741 17249
rect 18988 17240 19028 17704
rect 19084 17249 19124 18451
rect 19276 18257 19316 18535
rect 19275 18248 19317 18257
rect 19275 18208 19276 18248
rect 19316 18208 19317 18248
rect 19275 18199 19317 18208
rect 19372 18005 19412 18544
rect 19564 18535 19604 18544
rect 19756 18584 19796 18595
rect 19756 18509 19796 18544
rect 20524 18509 20564 19132
rect 20812 18929 20852 19216
rect 21004 19256 21044 19265
rect 21004 19097 21044 19216
rect 21003 19088 21045 19097
rect 21003 19048 21004 19088
rect 21044 19048 21045 19088
rect 21003 19039 21045 19048
rect 21099 19004 21141 19013
rect 21099 18964 21100 19004
rect 21140 18964 21141 19004
rect 21099 18955 21141 18964
rect 20811 18920 20853 18929
rect 20811 18880 20812 18920
rect 20852 18880 20853 18920
rect 20811 18871 20853 18880
rect 20715 18668 20757 18677
rect 20715 18628 20716 18668
rect 20756 18628 20757 18668
rect 20715 18619 20757 18628
rect 20619 18584 20661 18593
rect 20619 18544 20620 18584
rect 20660 18544 20661 18584
rect 20619 18535 20661 18544
rect 20716 18584 20756 18619
rect 19755 18500 19797 18509
rect 19755 18460 19756 18500
rect 19796 18460 19797 18500
rect 19755 18451 19797 18460
rect 20523 18500 20565 18509
rect 20523 18460 20524 18500
rect 20564 18460 20565 18500
rect 20523 18451 20565 18460
rect 19467 18332 19509 18341
rect 19467 18292 19468 18332
rect 19508 18292 19509 18332
rect 19467 18283 19509 18292
rect 19660 18332 19700 18341
rect 19371 17996 19413 18005
rect 19371 17956 19372 17996
rect 19412 17956 19413 17996
rect 19371 17947 19413 17956
rect 19180 17744 19220 17753
rect 19180 17669 19220 17704
rect 19275 17744 19317 17753
rect 19275 17704 19276 17744
rect 19316 17704 19317 17744
rect 19275 17695 19317 17704
rect 19468 17744 19508 18283
rect 19660 17921 19700 18292
rect 20524 18005 20564 18451
rect 20620 18450 20660 18535
rect 20716 18332 20756 18544
rect 20620 18292 20756 18332
rect 20523 17996 20565 18005
rect 20523 17956 20524 17996
rect 20564 17956 20565 17996
rect 20523 17947 20565 17956
rect 19659 17912 19701 17921
rect 19659 17872 19660 17912
rect 19700 17872 19701 17912
rect 19659 17863 19701 17872
rect 19468 17695 19508 17704
rect 19756 17744 19796 17753
rect 20620 17744 20660 18292
rect 20812 18257 20852 18871
rect 20908 18752 20948 18761
rect 20908 18593 20948 18712
rect 21100 18668 21140 18955
rect 21388 18752 21428 18761
rect 21484 18752 21524 19384
rect 21428 18712 21524 18752
rect 21388 18703 21428 18712
rect 21100 18619 21140 18628
rect 21195 18668 21237 18677
rect 21195 18628 21196 18668
rect 21236 18628 21237 18668
rect 21195 18619 21237 18628
rect 20907 18584 20949 18593
rect 20907 18544 20908 18584
rect 20948 18544 20949 18584
rect 20907 18535 20949 18544
rect 20811 18248 20853 18257
rect 20811 18208 20812 18248
rect 20852 18208 20853 18248
rect 20811 18199 20853 18208
rect 20715 18080 20757 18089
rect 20715 18040 20716 18080
rect 20756 18040 20757 18080
rect 20715 18031 20757 18040
rect 19796 17704 19988 17744
rect 19756 17695 19796 17704
rect 19180 17660 19222 17669
rect 19180 17620 19181 17660
rect 19221 17620 19222 17660
rect 19180 17611 19222 17620
rect 19276 17610 19316 17695
rect 19660 17585 19700 17670
rect 19371 17576 19413 17585
rect 19371 17536 19372 17576
rect 19412 17536 19413 17576
rect 19371 17527 19413 17536
rect 19659 17576 19701 17585
rect 19659 17536 19660 17576
rect 19700 17536 19701 17576
rect 19659 17527 19701 17536
rect 19372 17442 19412 17527
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 18699 17200 18700 17240
rect 18740 17200 18741 17240
rect 18699 17191 18741 17200
rect 18892 17200 19028 17240
rect 19083 17240 19125 17249
rect 19083 17200 19084 17240
rect 19124 17200 19125 17240
rect 18700 17106 18740 17191
rect 18795 17156 18837 17165
rect 18795 17116 18796 17156
rect 18836 17116 18837 17156
rect 18795 17107 18837 17116
rect 18796 17022 18836 17107
rect 18892 17081 18932 17200
rect 19083 17191 19125 17200
rect 18891 17072 18933 17081
rect 18891 17032 18892 17072
rect 18932 17032 18933 17072
rect 18891 17023 18933 17032
rect 18988 17072 19028 17081
rect 18892 16938 18932 17023
rect 18603 16820 18645 16829
rect 18603 16780 18604 16820
rect 18644 16780 18645 16820
rect 18603 16771 18645 16780
rect 18700 16820 18740 16829
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 18700 16409 18740 16780
rect 18699 16400 18741 16409
rect 18699 16360 18700 16400
rect 18740 16360 18741 16400
rect 18699 16351 18741 16360
rect 17548 16232 17588 16241
rect 17452 16192 17548 16232
rect 17356 16183 17396 16192
rect 17548 16183 17588 16192
rect 18027 16232 18069 16241
rect 18027 16192 18028 16232
rect 18068 16192 18069 16232
rect 18027 16183 18069 16192
rect 18699 16232 18741 16241
rect 18988 16232 19028 17032
rect 19180 17072 19220 17081
rect 19180 16325 19220 17032
rect 19179 16316 19221 16325
rect 19179 16276 19180 16316
rect 19220 16276 19221 16316
rect 19179 16267 19221 16276
rect 18699 16192 18700 16232
rect 18740 16192 19028 16232
rect 18699 16183 18741 16192
rect 18220 16064 18260 16073
rect 16876 16024 17300 16064
rect 18124 16024 18220 16064
rect 16492 15560 16532 15569
rect 16492 15149 16532 15520
rect 16875 15560 16917 15569
rect 16875 15520 16876 15560
rect 16916 15520 16917 15560
rect 16875 15511 16917 15520
rect 17643 15560 17685 15569
rect 17643 15520 17644 15560
rect 17684 15520 17685 15560
rect 17643 15511 17685 15520
rect 16491 15140 16533 15149
rect 16491 15100 16492 15140
rect 16532 15100 16533 15140
rect 16491 15091 16533 15100
rect 16684 14897 16724 14982
rect 16683 14888 16725 14897
rect 16683 14848 16684 14888
rect 16724 14848 16725 14888
rect 16683 14839 16725 14848
rect 16492 14720 16532 14729
rect 16396 14680 16492 14720
rect 16299 14671 16341 14680
rect 16300 14586 16340 14671
rect 16492 14225 16532 14680
rect 16683 14720 16725 14729
rect 16683 14680 16684 14720
rect 16724 14680 16725 14720
rect 16683 14671 16725 14680
rect 16684 14586 16724 14671
rect 16876 14468 16916 15511
rect 17644 15426 17684 15511
rect 17068 15308 17108 15317
rect 16971 14720 17013 14729
rect 16971 14680 16972 14720
rect 17012 14680 17013 14720
rect 16971 14671 17013 14680
rect 16972 14586 17012 14671
rect 16876 14428 17012 14468
rect 16491 14216 16533 14225
rect 16491 14176 16492 14216
rect 16532 14176 16533 14216
rect 16491 14167 16533 14176
rect 15724 13914 15764 13999
rect 15820 13997 15860 14008
rect 15916 14048 15956 14057
rect 15148 13831 15188 13840
rect 14860 12487 14900 12496
rect 14956 13208 14996 13217
rect 14668 12284 14708 12293
rect 14572 11864 14612 11873
rect 14475 11780 14517 11789
rect 14380 11740 14476 11780
rect 14516 11740 14517 11780
rect 13900 10396 14036 10436
rect 13324 10135 13364 10144
rect 13419 10184 13461 10193
rect 13419 10144 13420 10184
rect 13460 10144 13461 10184
rect 13419 10135 13461 10144
rect 13227 10100 13269 10109
rect 13227 10060 13228 10100
rect 13268 10060 13269 10100
rect 13227 10051 13269 10060
rect 12652 9631 12692 9640
rect 12267 8672 12309 8681
rect 12267 8632 12268 8672
rect 12308 8632 12309 8672
rect 13228 8672 13268 10051
rect 13420 10050 13460 10135
rect 13612 9512 13652 9521
rect 13612 9353 13652 9472
rect 13611 9344 13653 9353
rect 13611 9304 13612 9344
rect 13652 9304 13653 9344
rect 13611 9295 13653 9304
rect 13900 8765 13940 10396
rect 14092 10352 14132 10361
rect 13996 10312 14092 10352
rect 13996 9512 14036 10312
rect 14092 10303 14132 10312
rect 13996 9463 14036 9472
rect 13899 8756 13941 8765
rect 13899 8716 13900 8756
rect 13940 8716 13941 8756
rect 13899 8707 13941 8716
rect 13420 8672 13460 8681
rect 13228 8632 13420 8672
rect 12267 8623 12309 8632
rect 12116 7960 12212 8000
rect 12940 8000 12980 8009
rect 12076 7951 12116 7960
rect 12940 7589 12980 7960
rect 11499 7580 11541 7589
rect 11499 7540 11500 7580
rect 11540 7540 11541 7580
rect 11499 7531 11541 7540
rect 11691 7580 11733 7589
rect 11691 7540 11692 7580
rect 11732 7540 11733 7580
rect 11691 7531 11733 7540
rect 12939 7580 12981 7589
rect 12939 7540 12940 7580
rect 12980 7540 12981 7580
rect 12939 7531 12981 7540
rect 13131 7580 13173 7589
rect 13131 7540 13132 7580
rect 13172 7540 13173 7580
rect 13131 7531 13173 7540
rect 10252 7328 10292 7337
rect 10252 7160 10292 7288
rect 11116 7160 11156 7169
rect 10252 7120 10580 7160
rect 10444 6992 10484 7001
rect 10155 6824 10197 6833
rect 10155 6784 10156 6824
rect 10196 6784 10197 6824
rect 10155 6775 10197 6784
rect 10059 6740 10101 6749
rect 10059 6700 10060 6740
rect 10100 6700 10101 6740
rect 10059 6691 10101 6700
rect 10155 6656 10197 6665
rect 10155 6616 10156 6656
rect 10196 6616 10197 6656
rect 10155 6607 10197 6616
rect 10156 6522 10196 6607
rect 10252 6497 10292 6582
rect 10444 6572 10484 6952
rect 10444 6523 10484 6532
rect 9964 6488 10004 6497
rect 9867 5816 9909 5825
rect 9867 5776 9868 5816
rect 9908 5776 9909 5816
rect 9867 5767 9909 5776
rect 9964 5732 10004 6448
rect 10060 6488 10100 6497
rect 10060 6329 10100 6448
rect 10251 6488 10293 6497
rect 10251 6448 10252 6488
rect 10292 6448 10293 6488
rect 10540 6488 10580 7120
rect 11116 6665 11156 7120
rect 11403 6992 11445 7001
rect 11403 6952 11404 6992
rect 11444 6952 11445 6992
rect 11403 6943 11445 6952
rect 11404 6858 11444 6943
rect 11115 6656 11157 6665
rect 11115 6616 11116 6656
rect 11156 6616 11157 6656
rect 11115 6607 11157 6616
rect 10828 6488 10868 6497
rect 10540 6448 10828 6488
rect 10251 6439 10293 6448
rect 10828 6439 10868 6448
rect 11692 6488 11732 7531
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12843 7160 12885 7169
rect 12843 7120 12844 7160
rect 12884 7120 12885 7160
rect 12843 7111 12885 7120
rect 12076 7026 12116 7111
rect 12844 6656 12884 7111
rect 12844 6607 12884 6616
rect 12940 6497 12980 7531
rect 13132 7160 13172 7531
rect 13132 7111 13172 7120
rect 13420 6992 13460 8632
rect 13995 8672 14037 8681
rect 13995 8632 13996 8672
rect 14036 8632 14037 8672
rect 14188 8672 14228 11656
rect 14284 11696 14324 11705
rect 14284 11453 14324 11656
rect 14380 11696 14420 11740
rect 14475 11731 14517 11740
rect 14380 11647 14420 11656
rect 14283 11444 14325 11453
rect 14283 11404 14284 11444
rect 14324 11404 14325 11444
rect 14283 11395 14325 11404
rect 14284 11024 14324 11033
rect 14572 11024 14612 11824
rect 14324 10984 14612 11024
rect 14284 10975 14324 10984
rect 14668 8681 14708 12244
rect 14956 11864 14996 13168
rect 15340 13124 15380 13133
rect 15340 12629 15380 13084
rect 15532 13040 15572 13049
rect 15339 12620 15381 12629
rect 15339 12580 15340 12620
rect 15380 12580 15381 12620
rect 15339 12571 15381 12580
rect 14956 11815 14996 11824
rect 15532 11705 15572 13000
rect 15531 11696 15573 11705
rect 15531 11656 15532 11696
rect 15572 11656 15573 11696
rect 15531 11647 15573 11656
rect 15148 11024 15188 11033
rect 14860 9512 14900 9521
rect 14860 9101 14900 9472
rect 15148 9101 15188 10984
rect 15435 10268 15477 10277
rect 15435 10228 15436 10268
rect 15476 10228 15477 10268
rect 15435 10219 15477 10228
rect 15436 10134 15476 10219
rect 15916 9857 15956 14008
rect 16203 14048 16245 14057
rect 16203 14008 16204 14048
rect 16244 14008 16245 14048
rect 16203 13999 16245 14008
rect 16876 13796 16916 13805
rect 16780 13756 16876 13796
rect 16203 13376 16245 13385
rect 16203 13336 16204 13376
rect 16244 13336 16245 13376
rect 16203 13327 16245 13336
rect 16204 13208 16244 13327
rect 16683 13292 16725 13301
rect 16683 13252 16684 13292
rect 16724 13252 16725 13292
rect 16683 13243 16725 13252
rect 16204 13159 16244 13168
rect 16395 12620 16437 12629
rect 16395 12580 16396 12620
rect 16436 12580 16437 12620
rect 16395 12571 16437 12580
rect 16684 12620 16724 13243
rect 16684 12571 16724 12580
rect 16107 11696 16149 11705
rect 16107 11656 16108 11696
rect 16148 11656 16149 11696
rect 16107 11647 16149 11656
rect 16396 11696 16436 12571
rect 16780 12545 16820 13756
rect 16876 13747 16916 13756
rect 16875 13208 16917 13217
rect 16875 13168 16876 13208
rect 16916 13168 16917 13208
rect 16875 13159 16917 13168
rect 16588 12536 16628 12545
rect 16588 12377 16628 12496
rect 16779 12536 16821 12545
rect 16779 12496 16780 12536
rect 16820 12496 16821 12536
rect 16779 12487 16821 12496
rect 16780 12402 16820 12487
rect 16587 12368 16629 12377
rect 16587 12328 16588 12368
rect 16628 12328 16629 12368
rect 16587 12319 16629 12328
rect 16779 11864 16821 11873
rect 16779 11824 16780 11864
rect 16820 11824 16821 11864
rect 16779 11815 16821 11824
rect 16780 11730 16820 11815
rect 16108 11562 16148 11647
rect 16299 11192 16341 11201
rect 16299 11152 16300 11192
rect 16340 11152 16341 11192
rect 16299 11143 16341 11152
rect 16300 11058 16340 11143
rect 16012 10352 16052 10361
rect 16396 10352 16436 11656
rect 16492 11612 16532 11621
rect 16492 11024 16532 11572
rect 16876 11360 16916 13159
rect 16684 11320 16916 11360
rect 16684 11192 16724 11320
rect 16780 11192 16820 11201
rect 16684 11152 16780 11192
rect 16780 11143 16820 11152
rect 16972 11033 17012 14428
rect 17068 14057 17108 15268
rect 17643 15056 17685 15065
rect 17643 15016 17644 15056
rect 17684 15016 17685 15056
rect 17643 15007 17685 15016
rect 17547 14720 17589 14729
rect 17547 14680 17548 14720
rect 17588 14680 17589 14720
rect 17547 14671 17589 14680
rect 17452 14552 17492 14561
rect 17356 14512 17452 14552
rect 17163 14216 17205 14225
rect 17163 14176 17164 14216
rect 17204 14176 17205 14216
rect 17163 14167 17205 14176
rect 17164 14082 17204 14167
rect 17067 14048 17109 14057
rect 17067 14008 17068 14048
rect 17108 14008 17109 14048
rect 17067 13999 17109 14008
rect 17068 12536 17108 13999
rect 17163 13964 17205 13973
rect 17163 13924 17164 13964
rect 17204 13924 17205 13964
rect 17163 13915 17205 13924
rect 17068 11705 17108 12496
rect 17067 11696 17109 11705
rect 17067 11656 17068 11696
rect 17108 11656 17109 11696
rect 17067 11647 17109 11656
rect 17067 11528 17109 11537
rect 17067 11488 17068 11528
rect 17108 11488 17109 11528
rect 17067 11479 17109 11488
rect 17068 11192 17108 11479
rect 17164 11192 17204 13915
rect 17356 13217 17396 14512
rect 17452 14503 17492 14512
rect 17451 14048 17493 14057
rect 17451 14008 17452 14048
rect 17492 14008 17493 14048
rect 17451 13999 17493 14008
rect 17452 13914 17492 13999
rect 17548 13880 17588 14671
rect 17644 14225 17684 15007
rect 18124 14720 18164 16024
rect 18220 16015 18260 16024
rect 18603 16064 18645 16073
rect 18603 16024 18604 16064
rect 18644 16024 18645 16064
rect 18603 16015 18645 16024
rect 18412 15560 18452 15569
rect 18412 15308 18452 15520
rect 18507 15560 18549 15569
rect 18507 15520 18508 15560
rect 18548 15520 18549 15560
rect 18507 15511 18549 15520
rect 18604 15560 18644 16015
rect 18700 15653 18740 16183
rect 19180 16073 19220 16267
rect 19948 16241 19988 17704
rect 20620 17695 20660 17704
rect 20716 17744 20756 18031
rect 21099 17912 21141 17921
rect 21099 17872 21100 17912
rect 21140 17872 21141 17912
rect 21099 17863 21141 17872
rect 20811 17828 20853 17837
rect 20811 17788 20812 17828
rect 20852 17788 20853 17828
rect 20811 17779 20853 17788
rect 20716 17695 20756 17704
rect 20812 17694 20852 17779
rect 21100 17778 21140 17863
rect 20907 17744 20949 17753
rect 20907 17704 20908 17744
rect 20948 17704 20949 17744
rect 21196 17744 21236 18619
rect 21291 18584 21333 18593
rect 21291 18544 21292 18584
rect 21332 18544 21333 18584
rect 21291 18535 21333 18544
rect 21388 18584 21428 18593
rect 21292 18450 21332 18535
rect 21388 18425 21428 18544
rect 21387 18416 21429 18425
rect 21387 18376 21388 18416
rect 21428 18376 21429 18416
rect 21387 18367 21429 18376
rect 21388 18089 21428 18367
rect 21387 18080 21429 18089
rect 21387 18040 21388 18080
rect 21428 18040 21429 18080
rect 21387 18031 21429 18040
rect 21484 17837 21524 18712
rect 21580 18173 21620 19804
rect 21772 18929 21812 19804
rect 21771 18920 21813 18929
rect 21771 18880 21772 18920
rect 21812 18880 21813 18920
rect 21771 18871 21813 18880
rect 21868 18677 21908 20476
rect 21964 20441 22004 20728
rect 22060 20768 22100 20971
rect 22060 20719 22100 20728
rect 22156 20600 22196 20609
rect 21963 20432 22005 20441
rect 21963 20392 21964 20432
rect 22004 20392 22005 20432
rect 21963 20383 22005 20392
rect 22059 20264 22101 20273
rect 22059 20224 22060 20264
rect 22100 20224 22101 20264
rect 22059 20215 22101 20224
rect 21964 20096 22004 20107
rect 21964 20021 22004 20056
rect 22060 20096 22100 20215
rect 22156 20105 22196 20560
rect 22060 20045 22100 20056
rect 22155 20096 22197 20105
rect 22155 20056 22156 20096
rect 22196 20056 22197 20096
rect 22155 20047 22197 20056
rect 21963 20012 22005 20021
rect 21963 19972 21964 20012
rect 22004 19972 22005 20012
rect 21963 19963 22005 19972
rect 22156 19256 22196 19265
rect 22252 19256 22292 22576
rect 22348 22541 22388 23080
rect 22540 23071 22580 23080
rect 22636 23080 22924 23120
rect 22443 22700 22485 22709
rect 22443 22660 22444 22700
rect 22484 22660 22485 22700
rect 22443 22651 22485 22660
rect 22347 22532 22389 22541
rect 22347 22492 22348 22532
rect 22388 22492 22389 22532
rect 22347 22483 22389 22492
rect 22348 22398 22388 22483
rect 22444 22196 22484 22651
rect 22348 22156 22484 22196
rect 22348 20180 22388 22156
rect 22539 22112 22581 22121
rect 22539 22072 22540 22112
rect 22580 22072 22581 22112
rect 22539 22063 22581 22072
rect 22540 21978 22580 22063
rect 22636 21776 22676 23080
rect 22924 23071 22964 23080
rect 23116 21785 23156 24508
rect 23212 22709 23252 25096
rect 23692 24893 23732 25264
rect 23691 24884 23733 24893
rect 23691 24844 23692 24884
rect 23732 24844 23733 24884
rect 23691 24835 23733 24844
rect 23787 23960 23829 23969
rect 23787 23920 23788 23960
rect 23828 23920 23829 23960
rect 23787 23911 23829 23920
rect 23788 23876 23828 23911
rect 23884 23885 23924 27607
rect 24076 27068 24116 28960
rect 24940 29000 24980 29128
rect 25036 29168 25076 30220
rect 25228 29840 25268 30304
rect 25228 29791 25268 29800
rect 25420 29840 25460 30640
rect 25420 29791 25460 29800
rect 25516 29840 25556 29849
rect 25323 29756 25365 29765
rect 25323 29716 25324 29756
rect 25364 29716 25365 29756
rect 25323 29707 25365 29716
rect 25324 29622 25364 29707
rect 25516 29345 25556 29800
rect 25515 29336 25557 29345
rect 25515 29296 25516 29336
rect 25556 29296 25557 29336
rect 25515 29287 25557 29296
rect 25036 29119 25076 29128
rect 25131 29168 25173 29177
rect 25131 29128 25132 29168
rect 25172 29128 25173 29168
rect 25131 29119 25173 29128
rect 25228 29168 25268 29208
rect 25132 29034 25172 29119
rect 25228 29093 25268 29128
rect 25516 29168 25556 29177
rect 25612 29168 25652 30640
rect 25900 30680 25940 31564
rect 26188 31555 26228 31564
rect 25996 30764 26036 30773
rect 26284 30764 26324 32152
rect 26475 31772 26517 31781
rect 26475 31732 26476 31772
rect 26516 31732 26517 31772
rect 26475 31723 26517 31732
rect 26379 31604 26421 31613
rect 26379 31564 26380 31604
rect 26420 31564 26421 31604
rect 26379 31555 26421 31564
rect 26380 31352 26420 31555
rect 26476 31520 26516 31723
rect 26476 31471 26516 31480
rect 26380 31303 26420 31312
rect 26572 30848 26612 32227
rect 26036 30724 26324 30764
rect 26476 30808 26612 30848
rect 25996 30715 26036 30724
rect 26476 30689 26516 30808
rect 25900 30631 25940 30640
rect 26475 30680 26517 30689
rect 26475 30640 26476 30680
rect 26516 30640 26517 30680
rect 26475 30631 26517 30640
rect 26572 30680 26612 30689
rect 26476 30546 26516 30631
rect 26284 30428 26324 30437
rect 26092 30388 26284 30428
rect 25707 30260 25749 30269
rect 25707 30220 25708 30260
rect 25748 30220 25749 30260
rect 25707 30211 25749 30220
rect 25708 29849 25748 30211
rect 25707 29840 25749 29849
rect 25707 29800 25708 29840
rect 25748 29800 25749 29840
rect 25707 29791 25749 29800
rect 25708 29706 25748 29791
rect 25899 29672 25941 29681
rect 25899 29632 25900 29672
rect 25940 29632 25941 29672
rect 25899 29623 25941 29632
rect 25900 29252 25940 29623
rect 25995 29420 26037 29429
rect 25995 29380 25996 29420
rect 26036 29380 26037 29420
rect 25995 29371 26037 29380
rect 25900 29203 25940 29212
rect 25556 29128 25652 29168
rect 25803 29168 25845 29177
rect 25803 29128 25804 29168
rect 25844 29128 25845 29168
rect 25227 29084 25269 29093
rect 25227 29044 25228 29084
rect 25268 29044 25269 29084
rect 25227 29035 25269 29044
rect 24940 28960 25076 29000
rect 24748 28328 24788 28960
rect 24844 28328 24884 28337
rect 24748 28288 24844 28328
rect 24844 28279 24884 28288
rect 24460 28244 24500 28253
rect 24500 28204 24788 28244
rect 24460 28195 24500 28204
rect 24748 27824 24788 28204
rect 24748 27784 24980 27824
rect 24747 27656 24789 27665
rect 24747 27616 24748 27656
rect 24788 27616 24789 27656
rect 24747 27607 24789 27616
rect 24844 27656 24884 27665
rect 24748 27522 24788 27607
rect 24844 27068 24884 27616
rect 24940 27488 24980 27784
rect 25036 27656 25076 28960
rect 25036 27607 25076 27616
rect 25228 27656 25268 29035
rect 25516 29000 25556 29128
rect 25803 29119 25845 29128
rect 25804 29034 25844 29119
rect 25420 28960 25556 29000
rect 25228 27581 25268 27616
rect 25323 27656 25365 27665
rect 25323 27616 25324 27656
rect 25364 27616 25365 27656
rect 25323 27607 25365 27616
rect 25227 27572 25269 27581
rect 25227 27532 25228 27572
rect 25268 27532 25269 27572
rect 25227 27523 25269 27532
rect 25036 27488 25076 27497
rect 24940 27448 25036 27488
rect 25036 27439 25076 27448
rect 25228 27404 25268 27523
rect 25324 27522 25364 27607
rect 25132 27364 25268 27404
rect 24844 27028 25076 27068
rect 24076 27019 24116 27028
rect 23979 26984 24021 26993
rect 23979 26944 23980 26984
rect 24020 26944 24021 26984
rect 23979 26935 24021 26944
rect 23980 26144 24020 26935
rect 24460 26816 24500 26825
rect 24940 26816 24980 26825
rect 23980 26095 24020 26104
rect 24268 26776 24460 26816
rect 24500 26776 24940 26816
rect 24171 25304 24213 25313
rect 24171 25264 24172 25304
rect 24212 25264 24213 25304
rect 24171 25255 24213 25264
rect 24075 24800 24117 24809
rect 24075 24760 24076 24800
rect 24116 24760 24117 24800
rect 24075 24751 24117 24760
rect 24076 24666 24116 24751
rect 23403 23624 23445 23633
rect 23403 23584 23404 23624
rect 23444 23584 23445 23624
rect 23403 23575 23445 23584
rect 23404 23490 23444 23575
rect 23308 23120 23348 23129
rect 23348 23080 23444 23120
rect 23308 23071 23348 23080
rect 23211 22700 23253 22709
rect 23211 22660 23212 22700
rect 23252 22660 23253 22700
rect 23211 22651 23253 22660
rect 23211 22532 23253 22541
rect 23211 22492 23212 22532
rect 23252 22492 23253 22532
rect 23211 22483 23253 22492
rect 23212 22280 23252 22483
rect 23404 22448 23444 23080
rect 23788 22709 23828 23836
rect 23883 23876 23925 23885
rect 23883 23836 23884 23876
rect 23924 23836 23925 23876
rect 23883 23827 23925 23836
rect 24172 23624 24212 25255
rect 24172 23575 24212 23584
rect 24171 23120 24213 23129
rect 24171 23080 24172 23120
rect 24212 23080 24213 23120
rect 24171 23071 24213 23080
rect 23787 22700 23829 22709
rect 23787 22660 23788 22700
rect 23828 22660 23829 22700
rect 23787 22651 23829 22660
rect 23404 22399 23444 22408
rect 24172 22289 24212 23071
rect 24268 22373 24308 26776
rect 24460 26767 24500 26776
rect 24940 26767 24980 26776
rect 25036 26816 25076 27028
rect 24844 26648 24884 26657
rect 24652 26608 24844 26648
rect 24652 25304 24692 26608
rect 24844 26599 24884 26608
rect 25036 26573 25076 26776
rect 25132 26816 25172 27364
rect 25420 26984 25460 28960
rect 25707 28328 25749 28337
rect 25707 28288 25708 28328
rect 25748 28288 25749 28328
rect 25707 28279 25749 28288
rect 25708 28194 25748 28279
rect 25611 27740 25653 27749
rect 25611 27700 25612 27740
rect 25652 27700 25653 27740
rect 25611 27691 25653 27700
rect 25612 27656 25652 27691
rect 25900 27665 25940 27750
rect 25996 27740 26036 29371
rect 25996 27691 26036 27700
rect 25612 27605 25652 27616
rect 25899 27656 25941 27665
rect 25899 27616 25900 27656
rect 25940 27616 25941 27656
rect 25899 27607 25941 27616
rect 26092 27488 26132 30388
rect 26284 30379 26324 30388
rect 26572 30269 26612 30640
rect 26668 30680 26708 32563
rect 26860 30932 26900 33664
rect 26956 31529 26996 34336
rect 27051 34327 27093 34336
rect 29068 34376 29108 34385
rect 27052 34242 27092 34327
rect 28204 34208 28244 34217
rect 28204 34049 28244 34168
rect 28396 34208 28436 34217
rect 27147 34040 27189 34049
rect 27147 34000 27148 34040
rect 27188 34000 27189 34040
rect 27147 33991 27189 34000
rect 28203 34040 28245 34049
rect 28203 34000 28204 34040
rect 28244 34000 28245 34040
rect 28203 33991 28245 34000
rect 27148 33788 27188 33991
rect 28396 33872 28436 34168
rect 29068 34049 29108 34336
rect 29260 34376 29300 34385
rect 29452 34376 29492 34924
rect 29548 34915 29588 34924
rect 29300 34336 29492 34376
rect 29644 34376 29684 35092
rect 29260 34327 29300 34336
rect 29644 34327 29684 34336
rect 30027 34376 30069 34385
rect 30027 34336 30028 34376
rect 30068 34336 30069 34376
rect 30027 34327 30069 34336
rect 29067 34040 29109 34049
rect 29067 34000 29068 34040
rect 29108 34000 29109 34040
rect 29067 33991 29109 34000
rect 27148 33739 27188 33748
rect 28108 33832 28436 33872
rect 28971 33872 29013 33881
rect 28971 33832 28972 33872
rect 29012 33832 29013 33872
rect 27052 33704 27092 33713
rect 27052 32957 27092 33664
rect 28108 33704 28148 33832
rect 28971 33823 29013 33832
rect 28972 33738 29012 33823
rect 27436 33452 27476 33461
rect 27476 33412 27668 33452
rect 27436 33403 27476 33412
rect 27051 32948 27093 32957
rect 27051 32908 27052 32948
rect 27092 32908 27093 32948
rect 27051 32899 27093 32908
rect 27052 32528 27092 32899
rect 27435 32864 27477 32873
rect 27435 32824 27436 32864
rect 27476 32824 27477 32864
rect 27435 32815 27477 32824
rect 27436 32730 27476 32815
rect 27052 32488 27380 32528
rect 27243 32276 27285 32285
rect 27243 32236 27244 32276
rect 27284 32236 27285 32276
rect 27243 32227 27285 32236
rect 27052 32192 27092 32201
rect 27052 32033 27092 32152
rect 27244 32192 27284 32227
rect 27244 32141 27284 32152
rect 27340 32192 27380 32488
rect 27340 32143 27380 32152
rect 27436 32192 27476 32201
rect 27051 32024 27093 32033
rect 27051 31984 27052 32024
rect 27092 31984 27093 32024
rect 27051 31975 27093 31984
rect 26955 31520 26997 31529
rect 26955 31480 26956 31520
rect 26996 31480 26997 31520
rect 26955 31471 26997 31480
rect 27339 31352 27381 31361
rect 27339 31312 27340 31352
rect 27380 31312 27381 31352
rect 27436 31352 27476 32152
rect 27531 32192 27573 32201
rect 27531 32152 27532 32192
rect 27572 32152 27573 32192
rect 27531 32143 27573 32152
rect 27532 32058 27572 32143
rect 27436 31312 27572 31352
rect 27339 31303 27381 31312
rect 26860 30892 27188 30932
rect 26763 30764 26805 30773
rect 26763 30724 26764 30764
rect 26804 30724 26805 30764
rect 26763 30715 26805 30724
rect 26668 30521 26708 30640
rect 26764 30630 26804 30715
rect 26956 30680 26996 30689
rect 26860 30640 26956 30680
rect 26667 30512 26709 30521
rect 26667 30472 26668 30512
rect 26708 30472 26709 30512
rect 26667 30463 26709 30472
rect 26571 30260 26613 30269
rect 26571 30220 26572 30260
rect 26612 30220 26613 30260
rect 26571 30211 26613 30220
rect 26764 30092 26804 30101
rect 26860 30092 26900 30640
rect 26956 30631 26996 30640
rect 27051 30680 27093 30689
rect 27051 30640 27052 30680
rect 27092 30640 27093 30680
rect 27051 30631 27093 30640
rect 27052 30546 27092 30631
rect 26804 30052 26900 30092
rect 26764 30043 26804 30052
rect 26668 29840 26708 29849
rect 27052 29840 27092 29849
rect 27148 29840 27188 30892
rect 27243 30764 27285 30773
rect 27243 30724 27244 30764
rect 27284 30724 27285 30764
rect 27243 30715 27285 30724
rect 27244 30680 27284 30715
rect 27244 30629 27284 30640
rect 27244 30512 27284 30521
rect 27340 30512 27380 31303
rect 27436 31184 27476 31193
rect 27436 30764 27476 31144
rect 27436 30715 27476 30724
rect 27532 30521 27572 31312
rect 27284 30472 27380 30512
rect 27531 30512 27573 30521
rect 27531 30472 27532 30512
rect 27572 30472 27573 30512
rect 27244 30463 27284 30472
rect 27531 30463 27573 30472
rect 27628 30344 27668 33412
rect 28108 33293 28148 33664
rect 28204 33704 28244 33713
rect 28780 33704 28820 33713
rect 28244 33664 28780 33704
rect 28204 33655 28244 33664
rect 28780 33655 28820 33664
rect 28876 33704 28916 33713
rect 28587 33536 28629 33545
rect 28587 33496 28588 33536
rect 28628 33496 28629 33536
rect 28587 33487 28629 33496
rect 28588 33402 28628 33487
rect 28876 33377 28916 33664
rect 29067 33704 29109 33713
rect 29932 33704 29972 33713
rect 29067 33664 29068 33704
rect 29108 33664 29109 33704
rect 29067 33655 29109 33664
rect 29836 33664 29932 33704
rect 29068 33570 29108 33655
rect 29163 33536 29205 33545
rect 29163 33496 29164 33536
rect 29204 33496 29205 33536
rect 29163 33487 29205 33496
rect 28875 33368 28917 33377
rect 28875 33328 28876 33368
rect 28916 33328 28917 33368
rect 28875 33319 28917 33328
rect 28107 33284 28149 33293
rect 28107 33244 28108 33284
rect 28148 33244 28149 33284
rect 28107 33235 28149 33244
rect 28587 32948 28629 32957
rect 28587 32908 28588 32948
rect 28628 32908 28629 32948
rect 28587 32899 28629 32908
rect 28491 32864 28533 32873
rect 28491 32824 28492 32864
rect 28532 32824 28533 32864
rect 28491 32815 28533 32824
rect 27723 32780 27765 32789
rect 27723 32740 27724 32780
rect 27764 32740 27765 32780
rect 27723 32731 27765 32740
rect 27724 32024 27764 32731
rect 27724 31975 27764 31984
rect 28300 31520 28340 31529
rect 28107 31352 28149 31361
rect 28107 31312 28108 31352
rect 28148 31312 28149 31352
rect 28107 31303 28149 31312
rect 28108 31218 28148 31303
rect 27820 30680 27860 30689
rect 28300 30680 28340 31480
rect 27860 30640 28340 30680
rect 28492 30680 28532 32815
rect 28588 32814 28628 32899
rect 28779 32864 28821 32873
rect 28779 32824 28780 32864
rect 28820 32824 28821 32864
rect 28779 32815 28821 32824
rect 29164 32864 29204 33487
rect 29260 33452 29300 33461
rect 29260 32873 29300 33412
rect 29451 33368 29493 33377
rect 29451 33328 29452 33368
rect 29492 33328 29493 33368
rect 29451 33319 29493 33328
rect 29164 32815 29204 32824
rect 29259 32864 29301 32873
rect 29259 32824 29260 32864
rect 29300 32824 29301 32864
rect 29259 32815 29301 32824
rect 28780 32730 28820 32815
rect 28780 32192 28820 32201
rect 28972 32192 29012 32201
rect 28820 32152 28972 32192
rect 28780 32143 28820 32152
rect 28972 32143 29012 32152
rect 28683 31940 28725 31949
rect 28683 31900 28684 31940
rect 28724 31900 28725 31940
rect 28683 31891 28725 31900
rect 29355 31940 29397 31949
rect 29355 31900 29356 31940
rect 29396 31900 29397 31940
rect 29355 31891 29397 31900
rect 28684 31806 28724 31891
rect 29356 31352 29396 31891
rect 29356 31303 29396 31312
rect 29452 31352 29492 33319
rect 29643 32948 29685 32957
rect 29643 32908 29644 32948
rect 29684 32908 29685 32948
rect 29643 32899 29685 32908
rect 29644 32192 29684 32899
rect 29644 32143 29684 32152
rect 29644 31604 29684 31613
rect 29836 31604 29876 33664
rect 29932 33655 29972 33664
rect 30028 32864 30068 34327
rect 30220 33881 30260 35176
rect 32140 35216 32180 35225
rect 31468 34964 31508 34973
rect 30892 34924 31468 34964
rect 30507 34376 30549 34385
rect 30507 34336 30508 34376
rect 30548 34336 30549 34376
rect 30507 34327 30549 34336
rect 30508 34242 30548 34327
rect 30219 33872 30261 33881
rect 30219 33832 30220 33872
rect 30260 33832 30261 33872
rect 30219 33823 30261 33832
rect 30795 33872 30837 33881
rect 30795 33832 30796 33872
rect 30836 33832 30837 33872
rect 30795 33823 30837 33832
rect 30796 33738 30836 33823
rect 30892 33704 30932 34924
rect 31468 34915 31508 34924
rect 32140 34637 32180 35176
rect 32716 35048 32756 35057
rect 31275 34628 31317 34637
rect 31275 34588 31276 34628
rect 31316 34588 31317 34628
rect 31275 34579 31317 34588
rect 31659 34628 31701 34637
rect 31659 34588 31660 34628
rect 31700 34588 31701 34628
rect 31659 34579 31701 34588
rect 32139 34628 32181 34637
rect 32139 34588 32140 34628
rect 32180 34588 32181 34628
rect 32139 34579 32181 34588
rect 30987 33872 31029 33881
rect 30987 33832 30988 33872
rect 31028 33832 31029 33872
rect 30987 33823 31029 33832
rect 30892 33655 30932 33664
rect 30219 32948 30261 32957
rect 30219 32908 30220 32948
rect 30260 32908 30261 32948
rect 30219 32899 30261 32908
rect 30028 32780 30068 32824
rect 29684 31564 29876 31604
rect 29932 32740 30068 32780
rect 29644 31555 29684 31564
rect 29643 31436 29685 31445
rect 29643 31396 29644 31436
rect 29684 31396 29685 31436
rect 29643 31387 29685 31396
rect 29452 31303 29492 31312
rect 29644 31352 29684 31387
rect 29932 31361 29972 32740
rect 30028 32192 30068 32201
rect 30028 31445 30068 32152
rect 30124 32192 30164 32201
rect 30124 31529 30164 32152
rect 30220 32192 30260 32899
rect 30315 32360 30357 32369
rect 30315 32320 30316 32360
rect 30356 32320 30357 32360
rect 30315 32311 30357 32320
rect 30699 32360 30741 32369
rect 30699 32320 30700 32360
rect 30740 32320 30741 32360
rect 30699 32311 30741 32320
rect 30123 31520 30165 31529
rect 30123 31480 30124 31520
rect 30164 31480 30165 31520
rect 30123 31471 30165 31480
rect 30027 31436 30069 31445
rect 30027 31396 30028 31436
rect 30068 31396 30069 31436
rect 30027 31387 30069 31396
rect 29644 31301 29684 31312
rect 29931 31352 29973 31361
rect 29931 31312 29932 31352
rect 29972 31312 29973 31352
rect 29931 31303 29973 31312
rect 29836 31184 29876 31193
rect 29876 31144 29972 31184
rect 29836 31135 29876 31144
rect 28684 30680 28724 30689
rect 28492 30640 28684 30680
rect 27820 30631 27860 30640
rect 28203 30512 28245 30521
rect 28203 30472 28204 30512
rect 28244 30472 28245 30512
rect 28203 30463 28245 30472
rect 26708 29800 26900 29840
rect 26668 29791 26708 29800
rect 26379 29672 26421 29681
rect 26379 29632 26380 29672
rect 26420 29632 26421 29672
rect 26379 29623 26421 29632
rect 26380 29538 26420 29623
rect 26667 29588 26709 29597
rect 26667 29548 26668 29588
rect 26708 29548 26709 29588
rect 26667 29539 26709 29548
rect 26571 29336 26613 29345
rect 26571 29296 26572 29336
rect 26612 29296 26613 29336
rect 26571 29287 26613 29296
rect 26572 29202 26612 29287
rect 26668 29168 26708 29539
rect 26860 29261 26900 29800
rect 27092 29800 27188 29840
rect 27244 30304 27668 30344
rect 26859 29252 26901 29261
rect 26859 29212 26860 29252
rect 26900 29212 26901 29252
rect 26859 29203 26901 29212
rect 26668 29119 26708 29128
rect 26763 29168 26805 29177
rect 26763 29128 26764 29168
rect 26804 29128 26805 29168
rect 26763 29119 26805 29128
rect 25900 27448 26132 27488
rect 26188 28916 26228 28925
rect 25611 27068 25653 27077
rect 25611 27028 25612 27068
rect 25652 27028 25653 27068
rect 25611 27019 25653 27028
rect 25035 26564 25077 26573
rect 25035 26524 25036 26564
rect 25076 26524 25077 26564
rect 25035 26515 25077 26524
rect 24843 26144 24885 26153
rect 24843 26104 24844 26144
rect 24884 26104 24885 26144
rect 24843 26095 24885 26104
rect 24844 26010 24884 26095
rect 25132 25892 25172 26776
rect 24844 25852 25172 25892
rect 25228 26944 25460 26984
rect 24747 25556 24789 25565
rect 24747 25516 24748 25556
rect 24788 25516 24789 25556
rect 24747 25507 24789 25516
rect 24652 25255 24692 25264
rect 24748 25220 24788 25507
rect 24844 25304 24884 25852
rect 25131 25640 25173 25649
rect 25131 25600 25132 25640
rect 25172 25600 25173 25640
rect 25131 25591 25173 25600
rect 24844 25255 24884 25264
rect 24939 25304 24981 25313
rect 24939 25264 24940 25304
rect 24980 25264 24981 25304
rect 24939 25255 24981 25264
rect 24748 25171 24788 25180
rect 24940 25170 24980 25255
rect 24555 24800 24597 24809
rect 24555 24760 24556 24800
rect 24596 24760 24597 24800
rect 24555 24751 24597 24760
rect 24363 24632 24405 24641
rect 24363 24592 24364 24632
rect 24404 24592 24405 24632
rect 24363 24583 24405 24592
rect 24556 24632 24596 24751
rect 24556 24583 24596 24592
rect 24364 23792 24404 24583
rect 25132 23960 25172 25591
rect 25228 23969 25268 26944
rect 25420 26816 25460 26825
rect 25324 26776 25420 26816
rect 25324 25817 25364 26776
rect 25420 26767 25460 26776
rect 25612 26816 25652 27019
rect 25612 26767 25652 26776
rect 25708 26816 25748 26825
rect 25900 26816 25940 27448
rect 26188 26909 26228 28876
rect 26764 28580 26804 29119
rect 26860 29118 26900 29203
rect 26860 28580 26900 28589
rect 26764 28540 26860 28580
rect 26860 28531 26900 28540
rect 27052 27749 27092 29800
rect 27051 27740 27093 27749
rect 27051 27700 27052 27740
rect 27092 27700 27093 27740
rect 27051 27691 27093 27700
rect 26284 27404 26324 27413
rect 26324 27364 26516 27404
rect 26284 27355 26324 27364
rect 26379 27068 26421 27077
rect 26379 27028 26380 27068
rect 26420 27028 26421 27068
rect 26379 27019 26421 27028
rect 26187 26900 26229 26909
rect 26187 26860 26188 26900
rect 26228 26860 26229 26900
rect 26187 26851 26229 26860
rect 25748 26776 25940 26816
rect 25995 26816 26037 26825
rect 25995 26776 25996 26816
rect 26036 26776 26037 26816
rect 25708 26767 25748 26776
rect 25995 26767 26037 26776
rect 25515 26648 25557 26657
rect 25515 26608 25516 26648
rect 25556 26608 25557 26648
rect 25515 26599 25557 26608
rect 25900 26648 25940 26659
rect 25516 26514 25556 26599
rect 25900 26573 25940 26608
rect 25899 26564 25941 26573
rect 25899 26524 25900 26564
rect 25940 26524 25941 26564
rect 25899 26515 25941 26524
rect 25996 26312 26036 26767
rect 25996 26263 26036 26272
rect 26380 26144 26420 27019
rect 26380 26095 26420 26104
rect 26476 26144 26516 27364
rect 26955 27068 26997 27077
rect 26955 27028 26956 27068
rect 26996 27028 26997 27068
rect 26955 27019 26997 27028
rect 26572 26825 26612 26910
rect 26571 26816 26613 26825
rect 26571 26776 26572 26816
rect 26612 26776 26613 26816
rect 26571 26767 26613 26776
rect 26956 26816 26996 27019
rect 27051 26900 27093 26909
rect 27051 26860 27052 26900
rect 27092 26860 27093 26900
rect 27244 26900 27284 30304
rect 27339 30176 27381 30185
rect 27339 30136 27340 30176
rect 27380 30136 27381 30176
rect 27339 30127 27381 30136
rect 27340 29840 27380 30127
rect 27724 30008 27764 30017
rect 27764 29968 27956 30008
rect 27724 29959 27764 29968
rect 27340 29791 27380 29800
rect 27435 29840 27477 29849
rect 27435 29800 27436 29840
rect 27476 29800 27477 29840
rect 27435 29791 27477 29800
rect 27436 29706 27476 29791
rect 27723 29672 27765 29681
rect 27723 29632 27724 29672
rect 27764 29632 27765 29672
rect 27723 29623 27765 29632
rect 27435 29168 27477 29177
rect 27532 29168 27572 29177
rect 27435 29128 27436 29168
rect 27476 29128 27532 29168
rect 27435 29119 27477 29128
rect 27532 29119 27572 29128
rect 27627 29168 27669 29177
rect 27627 29128 27628 29168
rect 27668 29128 27669 29168
rect 27627 29119 27669 29128
rect 27724 29168 27764 29623
rect 27724 29119 27764 29128
rect 27339 29084 27381 29093
rect 27339 29044 27340 29084
rect 27380 29044 27381 29084
rect 27339 29035 27381 29044
rect 27340 28328 27380 29035
rect 27340 28279 27380 28288
rect 27436 28328 27476 28337
rect 27436 27581 27476 28288
rect 27628 28328 27668 29119
rect 27820 29093 27860 29178
rect 27819 29084 27861 29093
rect 27819 29044 27820 29084
rect 27860 29044 27861 29084
rect 27819 29035 27861 29044
rect 27628 28279 27668 28288
rect 27820 28244 27860 28253
rect 27532 28160 27572 28169
rect 27820 28160 27860 28204
rect 27572 28120 27860 28160
rect 27532 28111 27572 28120
rect 27916 28076 27956 29968
rect 28107 29168 28149 29177
rect 28107 29128 28108 29168
rect 28148 29128 28149 29168
rect 28107 29119 28149 29128
rect 28204 29168 28244 30463
rect 28204 29119 28244 29128
rect 28300 29168 28340 29177
rect 28108 29034 28148 29119
rect 28300 28589 28340 29128
rect 28396 29168 28436 29177
rect 28299 28580 28341 28589
rect 28299 28540 28300 28580
rect 28340 28540 28341 28580
rect 28299 28531 28341 28540
rect 28396 28505 28436 29128
rect 28395 28496 28437 28505
rect 28395 28456 28396 28496
rect 28436 28456 28437 28496
rect 28395 28447 28437 28456
rect 28684 28337 28724 30640
rect 29836 30428 29876 30437
rect 29836 30269 29876 30388
rect 29835 30260 29877 30269
rect 29835 30220 29836 30260
rect 29876 30220 29877 30260
rect 29835 30211 29877 30220
rect 29260 30008 29300 30017
rect 29300 29968 29876 30008
rect 29260 29959 29300 29968
rect 29836 29840 29876 29968
rect 29836 29791 29876 29800
rect 29452 29756 29492 29765
rect 29259 29672 29301 29681
rect 29259 29632 29260 29672
rect 29300 29632 29301 29672
rect 29452 29672 29492 29716
rect 29932 29672 29972 31144
rect 30220 30848 30260 32152
rect 30316 32192 30356 32311
rect 30316 32143 30356 32152
rect 30508 32192 30548 32201
rect 30700 32192 30740 32311
rect 30548 32152 30644 32192
rect 30508 32143 30548 32152
rect 30508 31940 30548 31949
rect 30508 31352 30548 31900
rect 30604 31529 30644 32152
rect 30700 32143 30740 32152
rect 30795 32192 30837 32201
rect 30795 32152 30796 32192
rect 30836 32152 30837 32192
rect 30795 32143 30837 32152
rect 30796 32058 30836 32143
rect 30603 31520 30645 31529
rect 30603 31480 30604 31520
rect 30644 31480 30645 31520
rect 30603 31471 30645 31480
rect 30508 31303 30548 31312
rect 30699 31352 30741 31361
rect 30699 31312 30700 31352
rect 30740 31312 30741 31352
rect 30699 31303 30741 31312
rect 30700 31218 30740 31303
rect 30220 30808 30356 30848
rect 30028 30680 30068 30689
rect 30028 30269 30068 30640
rect 30027 30260 30069 30269
rect 30027 30220 30028 30260
rect 30068 30220 30069 30260
rect 30027 30211 30069 30220
rect 29452 29632 29972 29672
rect 29259 29623 29301 29632
rect 29260 29168 29300 29623
rect 29260 29119 29300 29128
rect 29452 29168 29492 29177
rect 29163 29084 29205 29093
rect 29163 29044 29164 29084
rect 29204 29044 29205 29084
rect 29163 29035 29205 29044
rect 29164 28950 29204 29035
rect 29452 28337 29492 29128
rect 29931 28916 29973 28925
rect 29931 28876 29932 28916
rect 29972 28876 29973 28916
rect 29931 28867 29973 28876
rect 29739 28580 29781 28589
rect 29739 28540 29740 28580
rect 29780 28540 29781 28580
rect 29739 28531 29781 28540
rect 28204 28328 28244 28337
rect 28683 28328 28725 28337
rect 28244 28288 28628 28328
rect 28204 28279 28244 28288
rect 27820 28036 27956 28076
rect 27820 27656 27860 28036
rect 28588 27908 28628 28288
rect 28683 28288 28684 28328
rect 28724 28288 28725 28328
rect 28683 28279 28725 28288
rect 29067 28328 29109 28337
rect 29067 28288 29068 28328
rect 29108 28288 29109 28328
rect 29067 28279 29109 28288
rect 29451 28328 29493 28337
rect 29451 28288 29452 28328
rect 29492 28288 29493 28328
rect 29451 28279 29493 28288
rect 29068 28194 29108 28279
rect 28588 27868 28916 27908
rect 27820 27607 27860 27616
rect 27916 27656 27956 27665
rect 28108 27656 28148 27665
rect 27435 27572 27477 27581
rect 27435 27532 27436 27572
rect 27476 27532 27477 27572
rect 27435 27523 27477 27532
rect 27916 27245 27956 27616
rect 28012 27616 28108 27656
rect 27915 27236 27957 27245
rect 27915 27196 27916 27236
rect 27956 27196 27957 27236
rect 27915 27187 27957 27196
rect 28012 27068 28052 27616
rect 28108 27607 28148 27616
rect 28683 27572 28725 27581
rect 28683 27532 28684 27572
rect 28724 27532 28725 27572
rect 28683 27523 28725 27532
rect 28684 27438 28724 27523
rect 28876 27488 28916 27868
rect 29740 27656 29780 28531
rect 29835 27740 29877 27749
rect 29835 27700 29836 27740
rect 29876 27700 29877 27740
rect 29835 27691 29877 27700
rect 29740 27607 29780 27616
rect 29836 27606 29876 27691
rect 29259 27572 29301 27581
rect 29259 27532 29260 27572
rect 29300 27532 29301 27572
rect 29259 27523 29301 27532
rect 28876 27439 28916 27448
rect 27916 27028 28052 27068
rect 28108 27404 28148 27413
rect 27436 26900 27476 26909
rect 27244 26860 27436 26900
rect 27051 26851 27093 26860
rect 27436 26851 27476 26860
rect 26956 26767 26996 26776
rect 27052 26816 27092 26851
rect 27052 26765 27092 26776
rect 27532 26816 27572 26825
rect 26571 26648 26613 26657
rect 26571 26608 26572 26648
rect 26612 26608 26613 26648
rect 26571 26599 26613 26608
rect 26476 26095 26516 26104
rect 26572 26144 26612 26599
rect 27532 26405 27572 26776
rect 27531 26396 27573 26405
rect 27531 26356 27532 26396
rect 27572 26356 27573 26396
rect 27531 26347 27573 26356
rect 27916 26237 27956 27028
rect 28108 26909 28148 27364
rect 28492 27404 28532 27413
rect 28492 27245 28532 27364
rect 28491 27236 28533 27245
rect 28491 27196 28492 27236
rect 28532 27196 28533 27236
rect 28491 27187 28533 27196
rect 28875 26984 28917 26993
rect 28875 26944 28876 26984
rect 28916 26944 28917 26984
rect 28875 26935 28917 26944
rect 28107 26900 28149 26909
rect 28107 26860 28108 26900
rect 28148 26860 28149 26900
rect 28107 26851 28149 26860
rect 28779 26900 28821 26909
rect 28779 26860 28780 26900
rect 28820 26860 28821 26900
rect 28779 26851 28821 26860
rect 28011 26816 28053 26825
rect 28011 26776 28012 26816
rect 28052 26776 28053 26816
rect 28011 26767 28053 26776
rect 28492 26821 28532 26830
rect 28012 26682 28052 26767
rect 28107 26564 28149 26573
rect 28107 26524 28108 26564
rect 28148 26524 28149 26564
rect 28107 26515 28149 26524
rect 27915 26228 27957 26237
rect 27915 26188 27916 26228
rect 27956 26188 27957 26228
rect 27915 26179 27957 26188
rect 26572 26095 26612 26104
rect 26668 26144 26708 26153
rect 25323 25808 25365 25817
rect 25323 25768 25324 25808
rect 25364 25768 25365 25808
rect 25323 25759 25365 25768
rect 25324 24800 25364 25759
rect 26668 25640 26708 26104
rect 26859 26144 26901 26153
rect 26859 26104 26860 26144
rect 26900 26104 26901 26144
rect 26859 26095 26901 26104
rect 26956 26144 26996 26153
rect 26572 25600 26708 25640
rect 26475 25472 26517 25481
rect 26475 25432 26476 25472
rect 26516 25432 26517 25472
rect 26475 25423 26517 25432
rect 26379 25304 26421 25313
rect 26379 25264 26380 25304
rect 26420 25264 26421 25304
rect 26379 25255 26421 25264
rect 26476 25304 26516 25423
rect 26572 25339 26612 25600
rect 26860 25388 26900 26095
rect 26956 25817 26996 26104
rect 27916 26144 27956 26179
rect 27916 26093 27956 26104
rect 27244 25892 27284 25901
rect 27148 25852 27244 25892
rect 26955 25808 26997 25817
rect 26955 25768 26956 25808
rect 26996 25768 26997 25808
rect 26955 25759 26997 25768
rect 26860 25313 26900 25348
rect 26572 25290 26612 25299
rect 26668 25304 26708 25313
rect 26859 25304 26901 25313
rect 26476 25255 26516 25264
rect 26708 25264 26804 25304
rect 26668 25255 26708 25264
rect 26187 25220 26229 25229
rect 26187 25180 26188 25220
rect 26228 25180 26229 25220
rect 26187 25171 26229 25180
rect 26188 25086 26228 25171
rect 25324 24751 25364 24760
rect 26091 24800 26133 24809
rect 26091 24760 26092 24800
rect 26132 24760 26133 24800
rect 26091 24751 26133 24760
rect 26380 24800 26420 25255
rect 26571 25220 26613 25229
rect 26571 25180 26572 25220
rect 26612 25180 26613 25220
rect 26571 25171 26613 25180
rect 26380 24751 26420 24760
rect 25707 24632 25749 24641
rect 25707 24592 25708 24632
rect 25748 24592 25749 24632
rect 25707 24583 25749 24592
rect 26092 24632 26132 24751
rect 26475 24716 26517 24725
rect 26475 24676 26476 24716
rect 26516 24676 26517 24716
rect 26475 24667 26517 24676
rect 25708 24498 25748 24583
rect 25515 24128 25557 24137
rect 25515 24088 25516 24128
rect 25556 24088 25557 24128
rect 25515 24079 25557 24088
rect 25132 23911 25172 23920
rect 25227 23960 25269 23969
rect 25227 23920 25228 23960
rect 25268 23920 25269 23960
rect 25227 23911 25269 23920
rect 24364 23743 24404 23752
rect 24460 23792 24500 23801
rect 24652 23792 24692 23801
rect 24500 23752 24596 23792
rect 24460 23743 24500 23752
rect 24363 22700 24405 22709
rect 24363 22660 24364 22700
rect 24404 22660 24405 22700
rect 24363 22651 24405 22660
rect 24267 22364 24309 22373
rect 24267 22324 24268 22364
rect 24308 22324 24309 22364
rect 24267 22315 24309 22324
rect 23212 22231 23252 22240
rect 24171 22280 24213 22289
rect 24171 22240 24172 22280
rect 24212 22240 24213 22280
rect 24171 22231 24213 22240
rect 24364 22280 24404 22651
rect 24364 22231 24404 22240
rect 24172 22112 24212 22121
rect 24460 22112 24500 22121
rect 24212 22072 24308 22112
rect 24172 22063 24212 22072
rect 22636 21727 22676 21736
rect 23115 21776 23157 21785
rect 23115 21736 23116 21776
rect 23156 21736 23157 21776
rect 23115 21727 23157 21736
rect 22540 21617 22580 21702
rect 23980 21617 24020 21702
rect 22539 21608 22581 21617
rect 22539 21568 22540 21608
rect 22580 21568 22581 21608
rect 22539 21559 22581 21568
rect 22732 21608 22772 21617
rect 22924 21608 22964 21617
rect 23596 21608 23636 21617
rect 22772 21568 22924 21608
rect 22732 21559 22772 21568
rect 22924 21559 22964 21568
rect 23020 21568 23596 21608
rect 22635 21440 22677 21449
rect 22635 21400 22636 21440
rect 22676 21400 22677 21440
rect 22635 21391 22677 21400
rect 22539 21020 22581 21029
rect 22539 20980 22540 21020
rect 22580 20980 22581 21020
rect 22539 20971 22581 20980
rect 22540 20861 22580 20971
rect 22539 20852 22581 20861
rect 22539 20812 22540 20852
rect 22580 20812 22581 20852
rect 22539 20803 22581 20812
rect 22540 20768 22580 20803
rect 22636 20777 22676 21391
rect 23020 21104 23060 21568
rect 23596 21559 23636 21568
rect 23788 21608 23828 21617
rect 23403 21440 23445 21449
rect 23403 21400 23404 21440
rect 23444 21400 23445 21440
rect 23403 21391 23445 21400
rect 22828 21064 23060 21104
rect 23115 21104 23157 21113
rect 23115 21064 23116 21104
rect 23156 21064 23157 21104
rect 22540 20718 22580 20728
rect 22635 20768 22677 20777
rect 22635 20728 22636 20768
rect 22676 20728 22677 20768
rect 22635 20719 22677 20728
rect 22732 20768 22772 20777
rect 22348 20140 22484 20180
rect 22444 19424 22484 20140
rect 22539 20096 22581 20105
rect 22539 20056 22540 20096
rect 22580 20056 22581 20096
rect 22539 20047 22581 20056
rect 22636 20096 22676 20719
rect 22732 20441 22772 20728
rect 22828 20768 22868 21064
rect 23115 21055 23157 21064
rect 23019 20936 23061 20945
rect 23019 20896 23020 20936
rect 23060 20896 23061 20936
rect 23019 20887 23061 20896
rect 22828 20719 22868 20728
rect 23020 20768 23060 20887
rect 23020 20719 23060 20728
rect 23116 20768 23156 21055
rect 23211 20852 23253 20861
rect 23211 20812 23212 20852
rect 23252 20812 23253 20852
rect 23211 20803 23253 20812
rect 22731 20432 22773 20441
rect 22731 20392 22732 20432
rect 22772 20392 22773 20432
rect 22731 20383 22773 20392
rect 23116 20180 23156 20728
rect 23212 20768 23252 20803
rect 23212 20717 23252 20728
rect 23307 20768 23349 20777
rect 23307 20728 23308 20768
rect 23348 20728 23349 20768
rect 23404 20768 23444 21391
rect 23595 21356 23637 21365
rect 23595 21316 23596 21356
rect 23636 21316 23637 21356
rect 23595 21307 23637 21316
rect 23500 20945 23540 20964
rect 23499 20936 23541 20945
rect 23596 20936 23636 21307
rect 23788 21113 23828 21568
rect 23979 21608 24021 21617
rect 23979 21568 23980 21608
rect 24020 21568 24021 21608
rect 23979 21559 24021 21568
rect 23884 21524 23924 21533
rect 23884 21440 23924 21484
rect 23884 21400 24212 21440
rect 23787 21104 23829 21113
rect 23787 21064 23788 21104
rect 23828 21064 23829 21104
rect 23787 21055 23829 21064
rect 23499 20896 23500 20936
rect 23540 20910 23636 20936
rect 23540 20896 23596 20910
rect 23499 20887 23541 20896
rect 23788 20936 23828 20945
rect 23828 20896 24116 20936
rect 23788 20887 23828 20896
rect 23596 20861 23636 20870
rect 23596 20768 23636 20777
rect 23404 20728 23596 20768
rect 23307 20719 23349 20728
rect 23308 20634 23348 20719
rect 22540 19962 22580 20047
rect 22636 20021 22676 20056
rect 22828 20140 23156 20180
rect 23596 20180 23636 20728
rect 24076 20768 24116 20896
rect 24076 20719 24116 20728
rect 24172 20768 24212 21400
rect 24268 21365 24308 22072
rect 24460 21533 24500 22072
rect 24459 21524 24501 21533
rect 24459 21484 24460 21524
rect 24500 21484 24501 21524
rect 24459 21475 24501 21484
rect 24267 21356 24309 21365
rect 24267 21316 24268 21356
rect 24308 21316 24309 21356
rect 24267 21307 24309 21316
rect 24267 21188 24309 21197
rect 24267 21148 24268 21188
rect 24308 21148 24309 21188
rect 24267 21139 24309 21148
rect 24268 20777 24308 21139
rect 24172 20719 24212 20728
rect 24267 20768 24309 20777
rect 24460 20768 24500 21475
rect 24267 20728 24268 20768
rect 24308 20728 24309 20768
rect 24267 20719 24309 20728
rect 24364 20728 24500 20768
rect 24268 20634 24308 20719
rect 23980 20600 24020 20609
rect 23596 20140 23924 20180
rect 22635 20012 22677 20021
rect 22635 19972 22636 20012
rect 22676 19972 22677 20012
rect 22635 19963 22677 19972
rect 22636 19932 22676 19963
rect 22444 19384 22676 19424
rect 22444 19256 22484 19265
rect 22196 19216 22444 19256
rect 22156 19207 22196 19216
rect 22444 19207 22484 19216
rect 22443 19088 22485 19097
rect 22443 19048 22444 19088
rect 22484 19048 22485 19088
rect 22443 19039 22485 19048
rect 22444 18954 22484 19039
rect 21867 18668 21909 18677
rect 21867 18628 21868 18668
rect 21908 18628 21909 18668
rect 21867 18619 21909 18628
rect 22443 18668 22485 18677
rect 22443 18628 22444 18668
rect 22484 18628 22485 18668
rect 22540 18668 22580 19384
rect 22636 19256 22676 19384
rect 22636 19207 22676 19216
rect 22732 19256 22772 19265
rect 22636 18845 22676 18889
rect 22635 18836 22677 18845
rect 22635 18796 22636 18836
rect 22676 18796 22677 18836
rect 22635 18794 22677 18796
rect 22635 18787 22636 18794
rect 22676 18787 22677 18794
rect 22636 18745 22676 18754
rect 22540 18628 22628 18668
rect 22443 18619 22485 18628
rect 22444 18584 22484 18619
rect 22588 18593 22628 18628
rect 22732 18593 22772 19216
rect 22828 19013 22868 20140
rect 23884 20117 23924 20140
rect 23308 20096 23348 20105
rect 22924 20012 22964 20021
rect 23308 20012 23348 20056
rect 23403 20096 23445 20105
rect 23403 20056 23404 20096
rect 23444 20056 23540 20096
rect 23884 20068 23924 20077
rect 23403 20047 23445 20056
rect 22964 19972 23348 20012
rect 22924 19963 22964 19972
rect 23308 19760 23348 19972
rect 23404 19962 23444 20047
rect 23308 19720 23444 19760
rect 23307 19592 23349 19601
rect 23307 19552 23308 19592
rect 23348 19552 23349 19592
rect 23307 19543 23349 19552
rect 23211 19340 23253 19349
rect 23211 19300 23212 19340
rect 23252 19300 23253 19340
rect 23211 19291 23253 19300
rect 23212 19256 23252 19291
rect 23212 19205 23252 19216
rect 23308 19256 23348 19543
rect 23308 19207 23348 19216
rect 23404 19256 23444 19720
rect 23404 19207 23444 19216
rect 23500 19256 23540 20056
rect 23692 20012 23732 20021
rect 23980 20012 24020 20560
rect 24171 20432 24213 20441
rect 24171 20392 24172 20432
rect 24212 20392 24213 20432
rect 24171 20383 24213 20392
rect 24076 20096 24116 20107
rect 24076 20021 24116 20056
rect 23732 19972 23828 20012
rect 23692 19963 23732 19972
rect 23692 19349 23732 19380
rect 23691 19340 23733 19349
rect 23691 19300 23692 19340
rect 23732 19300 23733 19340
rect 23691 19291 23733 19300
rect 23500 19207 23540 19216
rect 23692 19256 23732 19291
rect 23692 19097 23732 19216
rect 23788 19256 23828 19972
rect 23788 19207 23828 19216
rect 23884 19972 24020 20012
rect 24075 20012 24117 20021
rect 24075 19972 24076 20012
rect 24116 19972 24117 20012
rect 23884 19256 23924 19972
rect 24075 19963 24117 19972
rect 23980 19844 24020 19853
rect 23980 19601 24020 19804
rect 23979 19592 24021 19601
rect 23979 19552 23980 19592
rect 24020 19552 24021 19592
rect 23979 19543 24021 19552
rect 23884 19207 23924 19216
rect 23980 19256 24020 19265
rect 24172 19256 24212 20383
rect 24268 20189 24308 20220
rect 24267 20180 24309 20189
rect 24267 20140 24268 20180
rect 24308 20140 24309 20180
rect 24267 20131 24309 20140
rect 24020 19216 24212 19256
rect 24268 20096 24308 20131
rect 23980 19207 24020 19216
rect 24268 19181 24308 20056
rect 24364 20096 24404 20728
rect 24556 20609 24596 23752
rect 24652 21617 24692 23752
rect 25419 23792 25461 23801
rect 25419 23752 25420 23792
rect 25460 23752 25461 23792
rect 25419 23743 25461 23752
rect 25420 23120 25460 23743
rect 25420 23071 25460 23080
rect 25035 21776 25077 21785
rect 25516 21776 25556 24079
rect 26092 23801 26132 24592
rect 26187 24632 26229 24641
rect 26187 24592 26188 24632
rect 26228 24592 26229 24632
rect 26187 24583 26229 24592
rect 26476 24632 26516 24667
rect 26188 24498 26228 24583
rect 26476 24581 26516 24592
rect 26572 24128 26612 25171
rect 26764 24800 26804 25264
rect 26859 25264 26860 25304
rect 26900 25264 26901 25304
rect 26859 25255 26901 25264
rect 26860 25224 26900 25255
rect 27052 24800 27092 24809
rect 26764 24760 27052 24800
rect 27052 24751 27092 24760
rect 26956 24632 26996 24643
rect 26956 24557 26996 24592
rect 27148 24632 27188 25852
rect 27244 25843 27284 25852
rect 27915 25556 27957 25565
rect 27915 25516 27916 25556
rect 27956 25516 28052 25556
rect 27915 25507 27957 25516
rect 27916 25422 27956 25507
rect 27243 25304 27285 25313
rect 27243 25264 27244 25304
rect 27284 25264 27285 25304
rect 27243 25255 27285 25264
rect 27244 25170 27284 25255
rect 27339 24884 27381 24893
rect 27339 24844 27340 24884
rect 27380 24844 27381 24884
rect 27339 24835 27381 24844
rect 27148 24583 27188 24592
rect 27243 24632 27285 24641
rect 27243 24592 27244 24632
rect 27284 24592 27285 24632
rect 27243 24583 27285 24592
rect 26955 24548 26997 24557
rect 26955 24508 26956 24548
rect 26996 24508 26997 24548
rect 26955 24499 26997 24508
rect 27244 24498 27284 24583
rect 27340 24557 27380 24835
rect 27435 24716 27477 24725
rect 27435 24676 27436 24716
rect 27476 24676 27477 24716
rect 27435 24667 27477 24676
rect 27436 24582 27476 24667
rect 27339 24548 27381 24557
rect 27339 24508 27340 24548
rect 27380 24508 27381 24548
rect 27339 24499 27381 24508
rect 26572 24088 26996 24128
rect 26187 23960 26229 23969
rect 26187 23920 26188 23960
rect 26228 23920 26229 23960
rect 26187 23911 26229 23920
rect 26763 23960 26805 23969
rect 26763 23920 26764 23960
rect 26804 23920 26805 23960
rect 26763 23911 26805 23920
rect 25612 23792 25652 23801
rect 25900 23792 25940 23801
rect 25652 23752 25900 23792
rect 25612 23743 25652 23752
rect 25900 23743 25940 23752
rect 26091 23792 26133 23801
rect 26091 23752 26092 23792
rect 26132 23752 26133 23792
rect 26091 23743 26133 23752
rect 25804 23120 25844 23129
rect 26188 23120 26228 23911
rect 26764 23826 26804 23911
rect 26571 23792 26613 23801
rect 26571 23752 26572 23792
rect 26612 23752 26613 23792
rect 26571 23743 26613 23752
rect 26572 23658 26612 23743
rect 25844 23080 25940 23120
rect 25804 23071 25844 23080
rect 25035 21736 25036 21776
rect 25076 21736 25077 21776
rect 25035 21727 25077 21736
rect 25420 21736 25556 21776
rect 25900 21776 25940 23080
rect 26188 23071 26228 23080
rect 24651 21608 24693 21617
rect 24651 21568 24652 21608
rect 24692 21568 24693 21608
rect 24651 21559 24693 21568
rect 24844 21608 24884 21617
rect 24844 20945 24884 21568
rect 24940 21608 24980 21619
rect 24940 21533 24980 21568
rect 25036 21608 25076 21727
rect 25036 21559 25076 21568
rect 25131 21608 25173 21617
rect 25131 21568 25132 21608
rect 25172 21568 25173 21608
rect 25131 21559 25173 21568
rect 25324 21608 25364 21619
rect 24939 21524 24981 21533
rect 24939 21484 24940 21524
rect 24980 21484 24981 21524
rect 24939 21475 24981 21484
rect 25132 21474 25172 21559
rect 25324 21533 25364 21568
rect 25420 21608 25460 21736
rect 25900 21727 25940 21736
rect 26476 21776 26516 21785
rect 26516 21736 26708 21776
rect 26476 21727 26516 21736
rect 25804 21617 25844 21702
rect 26668 21692 26708 21736
rect 26764 21692 26804 21701
rect 26668 21652 26764 21692
rect 26764 21643 26804 21652
rect 25323 21524 25365 21533
rect 25323 21484 25324 21524
rect 25364 21484 25365 21524
rect 25323 21475 25365 21484
rect 24843 20936 24885 20945
rect 24843 20896 24844 20936
rect 24884 20896 24885 20936
rect 24843 20887 24885 20896
rect 25036 20768 25076 20777
rect 24748 20728 25036 20768
rect 24555 20600 24597 20609
rect 24555 20560 24556 20600
rect 24596 20560 24597 20600
rect 24555 20551 24597 20560
rect 24460 20189 24500 20274
rect 24459 20180 24501 20189
rect 24748 20180 24788 20728
rect 25036 20719 25076 20728
rect 25228 20768 25268 20777
rect 25035 20348 25077 20357
rect 25035 20308 25036 20348
rect 25076 20308 25077 20348
rect 25035 20299 25077 20308
rect 25036 20264 25076 20299
rect 25036 20213 25076 20224
rect 24459 20140 24460 20180
rect 24500 20140 24501 20180
rect 24459 20131 24501 20140
rect 24556 20140 24748 20180
rect 24364 19937 24404 20056
rect 24556 20096 24596 20140
rect 24748 20131 24788 20140
rect 24556 20047 24596 20056
rect 24939 20096 24981 20105
rect 24939 20056 24940 20096
rect 24980 20056 24981 20096
rect 24939 20047 24981 20056
rect 25036 20096 25076 20105
rect 24940 19962 24980 20047
rect 24363 19928 24405 19937
rect 24363 19888 24364 19928
rect 24404 19888 24405 19928
rect 24363 19879 24405 19888
rect 25036 19265 25076 20056
rect 25228 19517 25268 20728
rect 25324 20768 25364 20777
rect 25420 20768 25460 21568
rect 25516 21608 25556 21617
rect 25516 21197 25556 21568
rect 25612 21608 25652 21617
rect 25612 21440 25652 21568
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 25803 21559 25845 21568
rect 25996 21608 26036 21617
rect 25996 21440 26036 21568
rect 25612 21400 26036 21440
rect 26092 21608 26132 21617
rect 26380 21608 26420 21617
rect 25515 21188 25557 21197
rect 25515 21148 25516 21188
rect 25556 21148 25557 21188
rect 25515 21139 25557 21148
rect 25516 21020 25556 21029
rect 26092 21020 26132 21568
rect 25556 20980 26132 21020
rect 26188 21568 26380 21608
rect 25516 20971 25556 20980
rect 25708 20768 25748 20777
rect 25420 20728 25708 20768
rect 25227 19508 25269 19517
rect 25227 19468 25228 19508
rect 25268 19468 25269 19508
rect 25227 19459 25269 19468
rect 25324 19349 25364 20728
rect 25708 20357 25748 20728
rect 26092 20768 26132 20777
rect 25707 20348 25749 20357
rect 25707 20308 25708 20348
rect 25748 20308 25749 20348
rect 25707 20299 25749 20308
rect 25612 20189 25652 20220
rect 25516 20180 25556 20189
rect 25516 20105 25556 20140
rect 25611 20180 25653 20189
rect 25611 20140 25612 20180
rect 25652 20140 25653 20180
rect 25708 20180 25748 20299
rect 25708 20140 25940 20180
rect 25611 20131 25653 20140
rect 25515 20096 25557 20105
rect 25515 20056 25516 20096
rect 25556 20056 25557 20096
rect 25515 20047 25557 20056
rect 25612 20096 25652 20131
rect 25323 19340 25365 19349
rect 25323 19300 25324 19340
rect 25364 19300 25365 19340
rect 25323 19291 25365 19300
rect 24363 19256 24405 19265
rect 24363 19216 24364 19256
rect 24404 19216 24405 19256
rect 24363 19207 24405 19216
rect 25035 19256 25077 19265
rect 25035 19216 25036 19256
rect 25076 19216 25077 19256
rect 25035 19207 25077 19216
rect 25227 19256 25269 19265
rect 25227 19216 25228 19256
rect 25268 19216 25269 19256
rect 25227 19207 25269 19216
rect 25324 19256 25364 19291
rect 24267 19172 24309 19181
rect 24267 19132 24268 19172
rect 24308 19132 24309 19172
rect 24267 19123 24309 19132
rect 23691 19088 23733 19097
rect 23691 19048 23692 19088
rect 23732 19048 23733 19088
rect 23691 19039 23733 19048
rect 23883 19088 23925 19097
rect 23883 19048 23884 19088
rect 23924 19048 23925 19088
rect 23883 19039 23925 19048
rect 22827 19004 22869 19013
rect 22827 18964 22828 19004
rect 22868 18964 22869 19004
rect 22827 18955 22869 18964
rect 22588 18584 22663 18593
rect 22731 18584 22773 18593
rect 22588 18544 22623 18584
rect 22663 18544 22676 18584
rect 22059 18416 22101 18425
rect 22059 18376 22060 18416
rect 22100 18376 22101 18416
rect 22059 18367 22101 18376
rect 21579 18164 21621 18173
rect 21579 18124 21580 18164
rect 21620 18124 21621 18164
rect 21579 18115 21621 18124
rect 21579 17996 21621 18005
rect 21579 17956 21580 17996
rect 21620 17956 21621 17996
rect 21579 17947 21621 17956
rect 21483 17828 21525 17837
rect 21483 17788 21484 17828
rect 21524 17788 21525 17828
rect 21483 17779 21525 17788
rect 21292 17744 21332 17753
rect 21196 17704 21292 17744
rect 20907 17695 20949 17704
rect 21292 17695 21332 17704
rect 21387 17744 21429 17753
rect 21387 17704 21388 17744
rect 21428 17704 21429 17744
rect 21387 17695 21429 17704
rect 21484 17744 21524 17779
rect 20908 17610 20948 17695
rect 21388 17610 21428 17695
rect 21484 17693 21524 17704
rect 21580 17744 21620 17947
rect 21963 17828 22005 17837
rect 21963 17788 21964 17828
rect 22004 17788 22005 17828
rect 21963 17779 22005 17788
rect 21580 17695 21620 17704
rect 21867 17744 21909 17753
rect 21867 17704 21868 17744
rect 21908 17704 21909 17744
rect 21867 17695 21909 17704
rect 21964 17744 22004 17779
rect 21868 17240 21908 17695
rect 21964 17693 22004 17704
rect 21868 17191 21908 17200
rect 20043 17156 20085 17165
rect 20043 17116 20044 17156
rect 20084 17116 20085 17156
rect 20043 17107 20085 17116
rect 20044 17072 20084 17107
rect 20044 17021 20084 17032
rect 21004 17072 21044 17081
rect 20427 16400 20469 16409
rect 20427 16360 20428 16400
rect 20468 16360 20469 16400
rect 20427 16351 20469 16360
rect 20235 16316 20277 16325
rect 20235 16276 20236 16316
rect 20276 16276 20277 16316
rect 20235 16267 20277 16276
rect 19947 16232 19989 16241
rect 19947 16192 19948 16232
rect 19988 16192 19989 16232
rect 19947 16183 19989 16192
rect 20139 16232 20181 16241
rect 20139 16192 20140 16232
rect 20180 16192 20181 16232
rect 20139 16183 20181 16192
rect 20236 16232 20276 16267
rect 20140 16098 20180 16183
rect 20236 16181 20276 16192
rect 20428 16232 20468 16351
rect 20907 16316 20949 16325
rect 20907 16276 20908 16316
rect 20948 16276 20949 16316
rect 20907 16267 20949 16276
rect 20620 16232 20660 16241
rect 20428 16183 20468 16192
rect 20524 16192 20620 16232
rect 19179 16064 19221 16073
rect 20428 16064 20468 16073
rect 19179 16024 19180 16064
rect 19220 16024 19221 16064
rect 19179 16015 19221 16024
rect 20236 16024 20428 16064
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 20140 15737 20180 15822
rect 20139 15728 20181 15737
rect 19660 15688 19892 15728
rect 18699 15644 18741 15653
rect 18699 15604 18700 15644
rect 18740 15604 18741 15644
rect 18699 15595 18741 15604
rect 18604 15511 18644 15520
rect 18796 15560 18836 15569
rect 18508 15426 18548 15511
rect 18699 15308 18741 15317
rect 18412 15268 18700 15308
rect 18740 15268 18741 15308
rect 18699 15259 18741 15268
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 18603 14972 18645 14981
rect 18603 14932 18604 14972
rect 18644 14932 18645 14972
rect 18603 14923 18645 14932
rect 18028 14680 18124 14720
rect 17643 14216 17685 14225
rect 17643 14176 17644 14216
rect 17684 14176 17685 14216
rect 17643 14167 17685 14176
rect 17644 13964 17684 14167
rect 17931 14048 17973 14057
rect 18028 14048 18068 14680
rect 18124 14671 18164 14680
rect 18507 14720 18549 14729
rect 18507 14680 18508 14720
rect 18548 14680 18549 14720
rect 18507 14671 18549 14680
rect 18508 14586 18548 14671
rect 18604 14636 18644 14923
rect 18700 14729 18740 15259
rect 18699 14720 18741 14729
rect 18699 14680 18700 14720
rect 18740 14680 18741 14720
rect 18699 14671 18741 14680
rect 18411 14216 18453 14225
rect 18604 14216 18644 14596
rect 18796 14477 18836 15520
rect 18892 15560 18932 15571
rect 18892 15485 18932 15520
rect 18988 15560 19028 15569
rect 18891 15476 18933 15485
rect 18891 15436 18892 15476
rect 18932 15436 18933 15476
rect 18891 15427 18933 15436
rect 18988 15317 19028 15520
rect 19084 15560 19124 15569
rect 19275 15560 19317 15569
rect 19124 15520 19220 15560
rect 19084 15511 19124 15520
rect 18987 15308 19029 15317
rect 18987 15268 18988 15308
rect 19028 15268 19029 15308
rect 18987 15259 19029 15268
rect 19180 14897 19220 15520
rect 19275 15520 19276 15560
rect 19316 15520 19317 15560
rect 19275 15511 19317 15520
rect 19468 15560 19508 15569
rect 19660 15560 19700 15688
rect 19508 15520 19604 15560
rect 19468 15511 19508 15520
rect 19276 15149 19316 15511
rect 19467 15392 19509 15401
rect 19467 15352 19468 15392
rect 19508 15352 19509 15392
rect 19564 15392 19604 15520
rect 19660 15511 19700 15520
rect 19756 15560 19796 15569
rect 19660 15392 19700 15401
rect 19564 15352 19660 15392
rect 19467 15343 19509 15352
rect 19660 15343 19700 15352
rect 19468 15258 19508 15343
rect 19756 15317 19796 15520
rect 19755 15308 19797 15317
rect 19755 15268 19756 15308
rect 19796 15268 19797 15308
rect 19755 15259 19797 15268
rect 19275 15140 19317 15149
rect 19275 15100 19276 15140
rect 19316 15100 19317 15140
rect 19275 15091 19317 15100
rect 19755 15140 19797 15149
rect 19755 15100 19756 15140
rect 19796 15100 19797 15140
rect 19755 15091 19797 15100
rect 18987 14888 19029 14897
rect 18987 14848 18988 14888
rect 19028 14848 19029 14888
rect 18987 14839 19029 14848
rect 19084 14888 19124 14897
rect 18892 14729 18932 14814
rect 18988 14804 19028 14839
rect 18988 14753 19028 14764
rect 18891 14720 18933 14729
rect 18891 14680 18892 14720
rect 18932 14680 18933 14720
rect 18891 14671 18933 14680
rect 19084 14645 19124 14848
rect 19179 14888 19221 14897
rect 19179 14848 19180 14888
rect 19220 14848 19221 14888
rect 19179 14846 19221 14848
rect 19179 14839 19180 14846
rect 19220 14839 19221 14846
rect 19180 14753 19220 14806
rect 19276 14720 19316 14729
rect 19083 14636 19125 14645
rect 19276 14636 19316 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19756 14720 19796 15091
rect 19852 15056 19892 15688
rect 20139 15688 20140 15728
rect 20180 15688 20181 15728
rect 20139 15679 20181 15688
rect 19948 15560 19988 15569
rect 19948 15233 19988 15520
rect 20139 15560 20181 15569
rect 20139 15520 20140 15560
rect 20180 15520 20181 15560
rect 20139 15511 20181 15520
rect 20140 15426 20180 15511
rect 19947 15224 19989 15233
rect 19947 15184 19948 15224
rect 19988 15184 19989 15224
rect 19947 15175 19989 15184
rect 19852 15016 19988 15056
rect 19851 14804 19893 14813
rect 19851 14764 19852 14804
rect 19892 14764 19893 14804
rect 19851 14755 19893 14764
rect 19756 14671 19796 14680
rect 19852 14720 19892 14755
rect 19948 14729 19988 15016
rect 20139 14804 20181 14813
rect 20139 14764 20140 14804
rect 20180 14764 20181 14804
rect 20139 14755 20181 14764
rect 19083 14596 19084 14636
rect 19124 14596 19125 14636
rect 19083 14587 19125 14596
rect 19180 14596 19316 14636
rect 18795 14468 18837 14477
rect 19180 14468 19220 14596
rect 18795 14428 18796 14468
rect 18836 14428 18837 14468
rect 18795 14419 18837 14428
rect 19084 14428 19220 14468
rect 19275 14468 19317 14477
rect 19275 14428 19276 14468
rect 19316 14428 19317 14468
rect 18411 14176 18412 14216
rect 18452 14176 18453 14216
rect 18411 14167 18453 14176
rect 18508 14176 18644 14216
rect 18987 14216 19029 14225
rect 18987 14176 18988 14216
rect 19028 14176 19029 14216
rect 18412 14082 18452 14167
rect 17931 14008 17932 14048
rect 17972 14008 18068 14048
rect 18124 14048 18164 14059
rect 17931 13999 17973 14008
rect 17644 13915 17684 13924
rect 17355 13208 17397 13217
rect 17355 13168 17356 13208
rect 17396 13168 17397 13208
rect 17355 13159 17397 13168
rect 17548 13040 17588 13840
rect 17836 13376 17876 13385
rect 17643 13292 17685 13301
rect 17643 13252 17644 13292
rect 17684 13252 17685 13292
rect 17643 13243 17685 13252
rect 17740 13292 17780 13301
rect 17644 13208 17684 13243
rect 17644 13157 17684 13168
rect 17548 13000 17684 13040
rect 17547 12620 17589 12629
rect 17547 12580 17548 12620
rect 17588 12580 17589 12620
rect 17356 12563 17396 12572
rect 17547 12571 17589 12580
rect 17260 12523 17356 12536
rect 17260 12496 17396 12523
rect 17452 12536 17492 12545
rect 17260 11369 17300 12496
rect 17452 12293 17492 12496
rect 17451 12284 17493 12293
rect 17451 12244 17452 12284
rect 17492 12244 17493 12284
rect 17451 12235 17493 12244
rect 17452 11948 17492 12235
rect 17356 11908 17492 11948
rect 17356 11696 17396 11908
rect 17356 11453 17396 11656
rect 17452 11696 17492 11705
rect 17548 11696 17588 12571
rect 17644 11705 17684 13000
rect 17740 12629 17780 13252
rect 17739 12620 17781 12629
rect 17739 12580 17740 12620
rect 17780 12580 17781 12620
rect 17739 12571 17781 12580
rect 17740 12284 17780 12295
rect 17740 12209 17780 12244
rect 17739 12200 17781 12209
rect 17739 12160 17740 12200
rect 17780 12160 17781 12200
rect 17739 12151 17781 12160
rect 17739 11948 17781 11957
rect 17739 11908 17740 11948
rect 17780 11908 17781 11948
rect 17739 11899 17781 11908
rect 17740 11814 17780 11899
rect 17492 11656 17588 11696
rect 17643 11696 17685 11705
rect 17643 11656 17644 11696
rect 17684 11656 17685 11696
rect 17836 11696 17876 13336
rect 17932 13292 17972 13999
rect 18124 13973 18164 14008
rect 18123 13964 18165 13973
rect 18123 13924 18124 13964
rect 18164 13924 18165 13964
rect 18123 13915 18165 13924
rect 18508 13889 18548 14176
rect 18987 14167 19029 14176
rect 18699 14132 18741 14141
rect 18699 14092 18700 14132
rect 18740 14092 18836 14132
rect 18699 14083 18745 14092
rect 18705 14057 18745 14083
rect 18603 14048 18645 14057
rect 18603 14008 18604 14048
rect 18644 14008 18645 14048
rect 18603 13999 18645 14008
rect 18705 14002 18745 14017
rect 18604 13914 18644 13999
rect 18507 13880 18549 13889
rect 18507 13840 18508 13880
rect 18548 13840 18549 13880
rect 18507 13831 18549 13840
rect 18699 13880 18741 13889
rect 18699 13840 18700 13880
rect 18740 13840 18741 13880
rect 18699 13831 18741 13840
rect 18220 13796 18260 13805
rect 17932 12881 17972 13252
rect 18124 13756 18220 13796
rect 18028 13208 18068 13217
rect 17931 12872 17973 12881
rect 17931 12832 17932 12872
rect 17972 12832 17973 12872
rect 17931 12823 17973 12832
rect 18028 12629 18068 13168
rect 18124 12797 18164 13756
rect 18220 13747 18260 13756
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18700 13460 18740 13831
rect 18508 13420 18740 13460
rect 18412 13217 18452 13302
rect 18411 13208 18453 13217
rect 18411 13168 18412 13208
rect 18452 13168 18453 13208
rect 18411 13159 18453 13168
rect 18219 12872 18261 12881
rect 18219 12832 18220 12872
rect 18260 12832 18261 12872
rect 18219 12823 18261 12832
rect 18123 12788 18165 12797
rect 18123 12748 18124 12788
rect 18164 12748 18165 12788
rect 18123 12739 18165 12748
rect 18027 12620 18069 12629
rect 18027 12580 18028 12620
rect 18068 12580 18069 12620
rect 18027 12571 18069 12580
rect 17931 12536 17973 12545
rect 17931 12496 17932 12536
rect 17972 12496 17973 12536
rect 17931 12487 17973 12496
rect 17932 12402 17972 12487
rect 18220 12461 18260 12823
rect 18315 12704 18357 12713
rect 18315 12664 18316 12704
rect 18356 12664 18357 12704
rect 18315 12655 18357 12664
rect 18316 12536 18356 12655
rect 18316 12487 18356 12496
rect 18508 12536 18548 13420
rect 18699 13208 18741 13217
rect 18699 13168 18700 13208
rect 18740 13168 18741 13208
rect 18699 13159 18741 13168
rect 18796 13208 18836 14092
rect 18892 14048 18932 14057
rect 18892 13469 18932 14008
rect 18988 14048 19028 14167
rect 18988 13999 19028 14008
rect 19084 14048 19124 14428
rect 19275 14419 19317 14428
rect 19084 13889 19124 14008
rect 19179 14048 19221 14057
rect 19179 14008 19180 14048
rect 19220 14008 19221 14048
rect 19179 13999 19221 14008
rect 19180 13914 19220 13999
rect 19083 13880 19125 13889
rect 19083 13840 19084 13880
rect 19124 13840 19125 13880
rect 19083 13831 19125 13840
rect 18891 13460 18933 13469
rect 18891 13420 18892 13460
rect 18932 13420 18933 13460
rect 18891 13411 18933 13420
rect 19083 13376 19125 13385
rect 19083 13336 19084 13376
rect 19124 13336 19125 13376
rect 19083 13327 19125 13336
rect 19084 13242 19124 13327
rect 19276 13208 19316 14419
rect 19372 14057 19412 14671
rect 19852 14669 19892 14680
rect 19947 14720 19989 14729
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 19947 14671 19989 14680
rect 20044 14720 20084 14729
rect 19947 14552 19989 14561
rect 19947 14512 19948 14552
rect 19988 14512 19989 14552
rect 19947 14503 19989 14512
rect 19948 14418 19988 14503
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 20044 14309 20084 14680
rect 20043 14300 20085 14309
rect 20043 14260 20044 14300
rect 20084 14260 20085 14300
rect 20043 14251 20085 14260
rect 19659 14216 19701 14225
rect 19659 14176 19660 14216
rect 19700 14176 19701 14216
rect 19659 14167 19701 14176
rect 19947 14216 19989 14225
rect 19947 14176 19948 14216
rect 19988 14176 19989 14216
rect 19947 14167 19989 14176
rect 19371 14048 19413 14057
rect 19371 14008 19372 14048
rect 19412 14008 19413 14048
rect 19371 13999 19413 14008
rect 19660 14048 19700 14167
rect 19948 14048 19988 14167
rect 20043 14132 20085 14141
rect 20043 14092 20044 14132
rect 20084 14092 20085 14132
rect 20043 14083 20085 14092
rect 19660 13999 19700 14008
rect 19756 14008 19948 14048
rect 19756 13880 19796 14008
rect 19948 13999 19988 14008
rect 20044 13998 20084 14083
rect 19660 13840 19796 13880
rect 19947 13880 19989 13889
rect 19947 13840 19948 13880
rect 19988 13840 19989 13880
rect 19467 13460 19509 13469
rect 19467 13420 19468 13460
rect 19508 13420 19509 13460
rect 19467 13411 19509 13420
rect 18836 13168 19028 13208
rect 18796 13159 18836 13168
rect 18700 13074 18740 13159
rect 18603 12788 18645 12797
rect 18603 12748 18604 12788
rect 18644 12748 18645 12788
rect 18603 12739 18645 12748
rect 18508 12461 18548 12496
rect 18604 12536 18644 12739
rect 18604 12487 18644 12496
rect 18700 12536 18740 12545
rect 18028 12452 18068 12461
rect 18028 12293 18068 12412
rect 18219 12452 18261 12461
rect 18219 12412 18220 12452
rect 18260 12412 18261 12452
rect 18219 12403 18261 12412
rect 18507 12452 18549 12461
rect 18507 12412 18508 12452
rect 18548 12412 18549 12452
rect 18507 12403 18549 12412
rect 18124 12368 18164 12377
rect 18027 12284 18069 12293
rect 18027 12244 18028 12284
rect 18068 12244 18069 12284
rect 18124 12284 18164 12328
rect 18700 12284 18740 12496
rect 18796 12536 18836 12545
rect 18988 12536 19028 13168
rect 19276 13159 19316 13168
rect 19468 13208 19508 13411
rect 19468 13159 19508 13168
rect 19660 13208 19700 13840
rect 19947 13831 19989 13840
rect 19948 13385 19988 13831
rect 20140 13385 20180 14755
rect 19852 13376 19892 13385
rect 19755 13292 19797 13301
rect 19755 13252 19756 13292
rect 19796 13252 19797 13292
rect 19755 13243 19797 13252
rect 19660 13159 19700 13168
rect 19756 13158 19796 13243
rect 19372 13040 19412 13049
rect 19852 13040 19892 13336
rect 19947 13376 19989 13385
rect 19947 13336 19948 13376
rect 19988 13336 19989 13376
rect 19947 13327 19989 13336
rect 20139 13376 20181 13385
rect 20139 13336 20140 13376
rect 20180 13336 20181 13376
rect 20139 13327 20181 13336
rect 19948 13292 19988 13327
rect 19948 13241 19988 13252
rect 20044 13208 20084 13217
rect 19852 13000 19988 13040
rect 19372 12629 19412 13000
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 19563 12704 19605 12713
rect 19563 12664 19564 12704
rect 19604 12664 19605 12704
rect 19563 12655 19605 12664
rect 19371 12620 19413 12629
rect 19371 12580 19372 12620
rect 19412 12580 19413 12620
rect 19371 12571 19413 12580
rect 19180 12536 19220 12545
rect 18836 12496 18932 12536
rect 18988 12496 19180 12536
rect 18796 12487 18836 12496
rect 18124 12244 18740 12284
rect 18027 12235 18069 12244
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 18892 11780 18932 12496
rect 19180 12487 19220 12496
rect 19564 12536 19604 12655
rect 19564 12487 19604 12496
rect 19948 12536 19988 13000
rect 20044 12881 20084 13168
rect 20139 13040 20181 13049
rect 20139 13000 20140 13040
rect 20180 13000 20181 13040
rect 20139 12991 20181 13000
rect 20043 12872 20085 12881
rect 20043 12832 20044 12872
rect 20084 12832 20085 12872
rect 20043 12823 20085 12832
rect 20043 12704 20085 12713
rect 20043 12664 20044 12704
rect 20084 12664 20085 12704
rect 20043 12655 20085 12664
rect 19948 12487 19988 12496
rect 20044 12536 20084 12655
rect 20044 12487 20084 12496
rect 19276 12452 19316 12461
rect 19083 12368 19125 12377
rect 19083 12328 19084 12368
rect 19124 12328 19125 12368
rect 19083 12319 19125 12328
rect 18892 11731 18932 11740
rect 18988 11864 19028 11873
rect 18220 11696 18260 11705
rect 17836 11656 18220 11696
rect 17452 11647 17492 11656
rect 17643 11647 17685 11656
rect 18220 11647 18260 11656
rect 18315 11696 18357 11705
rect 18315 11656 18316 11696
rect 18356 11656 18357 11696
rect 18315 11647 18357 11656
rect 18412 11696 18452 11705
rect 18316 11562 18356 11647
rect 18124 11528 18164 11537
rect 18028 11488 18124 11528
rect 17355 11444 17397 11453
rect 17355 11404 17356 11444
rect 17396 11404 17397 11444
rect 17355 11395 17397 11404
rect 17259 11360 17301 11369
rect 17259 11320 17260 11360
rect 17300 11320 17301 11360
rect 17259 11311 17301 11320
rect 17643 11276 17685 11285
rect 17643 11236 17644 11276
rect 17684 11236 17685 11276
rect 17643 11227 17685 11236
rect 17260 11192 17300 11201
rect 17164 11152 17260 11192
rect 17068 11143 17108 11152
rect 17260 11143 17300 11152
rect 16876 11024 16916 11033
rect 16492 10984 16876 11024
rect 16779 10436 16821 10445
rect 16779 10396 16780 10436
rect 16820 10396 16821 10436
rect 16779 10387 16821 10396
rect 16052 10312 16244 10352
rect 16396 10312 16724 10352
rect 16012 10303 16052 10312
rect 15531 9848 15573 9857
rect 15531 9808 15532 9848
rect 15572 9808 15573 9848
rect 15531 9799 15573 9808
rect 15915 9848 15957 9857
rect 15915 9808 15916 9848
rect 15956 9808 15957 9848
rect 15915 9799 15957 9808
rect 14859 9092 14901 9101
rect 14859 9052 14860 9092
rect 14900 9052 14901 9092
rect 14859 9043 14901 9052
rect 15147 9092 15189 9101
rect 15147 9052 15148 9092
rect 15188 9052 15189 9092
rect 15147 9043 15189 9052
rect 14380 8672 14420 8681
rect 14188 8632 14380 8672
rect 13995 8623 14037 8632
rect 13996 7160 14036 8623
rect 14380 8009 14420 8632
rect 14667 8672 14709 8681
rect 14667 8632 14668 8672
rect 14708 8632 14709 8672
rect 14667 8623 14709 8632
rect 15532 8672 15572 9799
rect 15723 9680 15765 9689
rect 15723 9640 15724 9680
rect 15764 9640 15765 9680
rect 15723 9631 15765 9640
rect 16011 9680 16053 9689
rect 16011 9640 16012 9680
rect 16052 9640 16053 9680
rect 16011 9631 16053 9640
rect 15627 9512 15669 9521
rect 15627 9472 15628 9512
rect 15668 9472 15669 9512
rect 15627 9463 15669 9472
rect 15628 8756 15668 9463
rect 15628 8707 15668 8716
rect 15532 8623 15572 8632
rect 15724 8672 15764 9631
rect 16012 9546 16052 9631
rect 16204 9344 16244 10312
rect 16300 10184 16340 10193
rect 16588 10184 16628 10193
rect 16340 10144 16588 10184
rect 16300 10135 16340 10144
rect 16588 10135 16628 10144
rect 16587 10016 16629 10025
rect 16587 9976 16588 10016
rect 16628 9976 16629 10016
rect 16587 9967 16629 9976
rect 16395 9764 16437 9773
rect 16395 9724 16396 9764
rect 16436 9724 16437 9764
rect 16395 9715 16437 9724
rect 16396 9512 16436 9715
rect 16491 9596 16533 9605
rect 16491 9556 16492 9596
rect 16532 9556 16533 9596
rect 16491 9547 16533 9556
rect 16396 9463 16436 9472
rect 16492 9462 16532 9547
rect 16588 9512 16628 9967
rect 16588 9463 16628 9472
rect 16204 9304 16628 9344
rect 16491 9092 16533 9101
rect 16491 9052 16492 9092
rect 16532 9052 16533 9092
rect 16491 9043 16533 9052
rect 16492 8840 16532 9043
rect 15724 8623 15764 8632
rect 16011 8672 16053 8681
rect 16011 8632 16012 8672
rect 16052 8632 16053 8672
rect 16011 8623 16053 8632
rect 16395 8672 16437 8681
rect 16395 8632 16396 8672
rect 16436 8632 16437 8672
rect 16395 8623 16437 8632
rect 16012 8538 16052 8623
rect 15915 8420 15957 8429
rect 15915 8380 15916 8420
rect 15956 8380 15957 8420
rect 15915 8371 15957 8380
rect 15819 8168 15861 8177
rect 15819 8128 15820 8168
rect 15860 8128 15861 8168
rect 15819 8119 15861 8128
rect 15916 8168 15956 8371
rect 15916 8119 15956 8128
rect 14379 8000 14421 8009
rect 14379 7960 14380 8000
rect 14420 7960 14421 8000
rect 14379 7951 14421 7960
rect 15820 8000 15860 8119
rect 14860 7832 14900 7841
rect 14092 7748 14132 7757
rect 14379 7748 14421 7757
rect 14132 7708 14324 7748
rect 14092 7699 14132 7708
rect 13996 7111 14036 7120
rect 13132 6952 13460 6992
rect 11692 6439 11732 6448
rect 11883 6488 11925 6497
rect 12939 6488 12981 6497
rect 11883 6448 11884 6488
rect 11924 6448 11925 6488
rect 11883 6439 11925 6448
rect 12844 6448 12940 6488
rect 12980 6448 12981 6488
rect 10059 6320 10101 6329
rect 10059 6280 10060 6320
rect 10100 6280 10101 6320
rect 10059 6271 10101 6280
rect 9964 5692 10100 5732
rect 9676 5648 9716 5657
rect 9580 5608 9676 5648
rect 9484 5524 9620 5564
rect 9387 5396 9429 5405
rect 9387 5356 9388 5396
rect 9428 5356 9429 5396
rect 9387 5347 9429 5356
rect 9195 5144 9237 5153
rect 9195 5104 9196 5144
rect 9236 5104 9237 5144
rect 9195 5095 9237 5104
rect 9195 4976 9237 4985
rect 9195 4936 9196 4976
rect 9236 4936 9237 4976
rect 9195 4927 9237 4936
rect 8811 4852 8812 4892
rect 8852 4852 8853 4892
rect 8811 4843 8853 4852
rect 8908 4852 9140 4892
rect 8908 4850 8948 4852
rect 8812 4758 8852 4843
rect 8908 4801 8948 4810
rect 9003 4640 9045 4649
rect 9003 4600 9004 4640
rect 9044 4600 9045 4640
rect 9003 4591 9045 4600
rect 8812 4136 8852 4145
rect 8716 4096 8812 4136
rect 8716 3641 8756 4096
rect 8812 4087 8852 4096
rect 8811 3968 8853 3977
rect 8811 3928 8812 3968
rect 8852 3928 8853 3968
rect 8811 3919 8853 3928
rect 8715 3632 8757 3641
rect 8715 3592 8716 3632
rect 8756 3592 8757 3632
rect 8715 3583 8757 3592
rect 8812 3632 8852 3919
rect 9004 3809 9044 4591
rect 9003 3800 9045 3809
rect 9003 3760 9004 3800
rect 9044 3760 9045 3800
rect 9003 3751 9045 3760
rect 8812 3583 8852 3592
rect 8716 3464 8756 3473
rect 8620 3424 8716 3464
rect 8236 3413 8276 3424
rect 8716 3415 8756 3424
rect 8908 3464 8948 3475
rect 8908 3389 8948 3424
rect 9004 3464 9044 3473
rect 9100 3464 9140 4852
rect 9196 4808 9236 4927
rect 9196 4759 9236 4768
rect 9196 4304 9236 4313
rect 9196 3977 9236 4264
rect 9388 4136 9428 5347
rect 9580 5069 9620 5524
rect 9676 5405 9716 5608
rect 9868 5648 9908 5657
rect 9908 5608 10004 5648
rect 9868 5599 9908 5608
rect 9771 5480 9813 5489
rect 9771 5440 9772 5480
rect 9812 5440 9813 5480
rect 9771 5431 9813 5440
rect 9675 5396 9717 5405
rect 9675 5356 9676 5396
rect 9716 5356 9717 5396
rect 9675 5347 9717 5356
rect 9772 5346 9812 5431
rect 9676 5148 9716 5157
rect 9579 5060 9621 5069
rect 9579 5020 9580 5060
rect 9620 5020 9621 5060
rect 9579 5011 9621 5020
rect 9484 4976 9524 4985
rect 9484 4808 9524 4936
rect 9580 4976 9620 5011
rect 9676 4985 9716 5108
rect 9580 4926 9620 4936
rect 9675 4976 9717 4985
rect 9868 4976 9908 4985
rect 9675 4936 9676 4976
rect 9716 4936 9717 4976
rect 9675 4927 9717 4936
rect 9772 4936 9868 4976
rect 9772 4808 9812 4936
rect 9868 4927 9908 4936
rect 9484 4768 9812 4808
rect 9484 4220 9524 4768
rect 9868 4724 9908 4733
rect 9772 4684 9868 4724
rect 9580 4220 9620 4229
rect 9484 4180 9580 4220
rect 9580 4171 9620 4180
rect 9388 4087 9428 4096
rect 9676 4136 9716 4145
rect 9195 3968 9237 3977
rect 9195 3928 9196 3968
rect 9236 3928 9237 3968
rect 9195 3919 9237 3928
rect 9676 3809 9716 4096
rect 9195 3800 9237 3809
rect 9195 3760 9196 3800
rect 9236 3760 9237 3800
rect 9195 3751 9237 3760
rect 9675 3800 9717 3809
rect 9675 3760 9676 3800
rect 9716 3760 9717 3800
rect 9675 3751 9717 3760
rect 9044 3424 9140 3464
rect 9196 3464 9236 3751
rect 9004 3415 9044 3424
rect 8907 3380 8949 3389
rect 8907 3340 8908 3380
rect 8948 3340 8949 3380
rect 8907 3331 8949 3340
rect 9196 2885 9236 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 8235 2876 8277 2885
rect 8235 2836 8236 2876
rect 8276 2836 8277 2876
rect 8235 2827 8277 2836
rect 9195 2876 9237 2885
rect 9195 2836 9196 2876
rect 9236 2836 9237 2876
rect 9195 2827 9237 2836
rect 8236 2742 8276 2827
rect 7700 2584 7988 2624
rect 9388 2624 9428 3415
rect 9772 3389 9812 4684
rect 9868 4675 9908 4684
rect 9867 4304 9909 4313
rect 9867 4264 9868 4304
rect 9908 4264 9909 4304
rect 9867 4255 9909 4264
rect 9868 4136 9908 4255
rect 9868 4087 9908 4096
rect 9964 4136 10004 5608
rect 10060 5144 10100 5692
rect 11884 5648 11924 6439
rect 11884 5599 11924 5608
rect 11979 5648 12021 5657
rect 11979 5608 11980 5648
rect 12020 5608 12021 5648
rect 11979 5599 12021 5608
rect 12076 5648 12116 5657
rect 10060 5104 10292 5144
rect 10060 4976 10100 4985
rect 10060 4817 10100 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10156 4842 10196 4927
rect 10059 4808 10101 4817
rect 10059 4768 10060 4808
rect 10100 4768 10101 4808
rect 10059 4759 10101 4768
rect 10252 4313 10292 5104
rect 10347 5060 10389 5069
rect 10347 5020 10348 5060
rect 10388 5020 10389 5060
rect 10347 5011 10389 5020
rect 10348 4976 10388 5011
rect 10348 4817 10388 4936
rect 10539 4976 10581 4985
rect 10539 4936 10540 4976
rect 10580 4936 10581 4976
rect 10539 4927 10581 4936
rect 11596 4976 11636 4985
rect 10443 4892 10485 4901
rect 10443 4852 10444 4892
rect 10484 4852 10485 4892
rect 10443 4843 10485 4852
rect 10347 4808 10389 4817
rect 10347 4768 10348 4808
rect 10388 4768 10389 4808
rect 10347 4759 10389 4768
rect 10444 4758 10484 4843
rect 10540 4842 10580 4927
rect 11596 4817 11636 4936
rect 11595 4808 11637 4817
rect 11595 4768 11596 4808
rect 11636 4768 11637 4808
rect 11595 4759 11637 4768
rect 11884 4724 11924 4733
rect 11788 4684 11884 4724
rect 11595 4388 11637 4397
rect 11595 4348 11596 4388
rect 11636 4348 11637 4388
rect 11595 4339 11637 4348
rect 10251 4304 10293 4313
rect 10251 4264 10252 4304
rect 10292 4264 10293 4304
rect 10251 4255 10293 4264
rect 10539 4304 10581 4313
rect 10539 4264 10540 4304
rect 10580 4264 10581 4304
rect 10539 4255 10581 4264
rect 11019 4304 11061 4313
rect 11019 4264 11020 4304
rect 11060 4264 11061 4304
rect 11019 4255 11061 4264
rect 11499 4304 11541 4313
rect 11499 4264 11500 4304
rect 11540 4264 11541 4304
rect 11499 4255 11541 4264
rect 10443 4220 10485 4229
rect 10443 4180 10444 4220
rect 10484 4180 10485 4220
rect 10443 4171 10485 4180
rect 9964 3809 10004 4096
rect 10156 4136 10196 4145
rect 10348 4136 10388 4145
rect 10196 4096 10348 4136
rect 10156 4087 10196 4096
rect 10348 4087 10388 4096
rect 10444 4136 10484 4171
rect 10444 4085 10484 4096
rect 10540 4136 10580 4255
rect 10923 4220 10965 4229
rect 10923 4180 10924 4220
rect 10964 4180 10965 4220
rect 10923 4171 10965 4180
rect 10540 4087 10580 4096
rect 10636 4136 10676 4145
rect 10060 3968 10100 3977
rect 9963 3800 10005 3809
rect 9963 3760 9964 3800
rect 10004 3760 10005 3800
rect 9963 3751 10005 3760
rect 10060 3641 10100 3928
rect 10251 3968 10293 3977
rect 10251 3928 10252 3968
rect 10292 3928 10293 3968
rect 10251 3919 10293 3928
rect 10155 3800 10197 3809
rect 10155 3760 10156 3800
rect 10196 3760 10197 3800
rect 10155 3751 10197 3760
rect 10059 3632 10101 3641
rect 10059 3592 10060 3632
rect 10100 3592 10101 3632
rect 10059 3583 10101 3592
rect 10156 3632 10196 3751
rect 10156 3583 10196 3592
rect 9868 3464 9908 3473
rect 10060 3464 10100 3473
rect 9908 3424 10060 3464
rect 9868 3415 9908 3424
rect 10060 3415 10100 3424
rect 9771 3380 9813 3389
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 7660 2575 7700 2584
rect 9388 2575 9428 2584
rect 10252 2624 10292 3919
rect 10636 3893 10676 4096
rect 10924 4136 10964 4171
rect 10924 4085 10964 4096
rect 11020 4136 11060 4255
rect 11403 4220 11445 4229
rect 11403 4180 11404 4220
rect 11444 4180 11445 4220
rect 11403 4171 11445 4180
rect 11020 4087 11060 4096
rect 11116 4136 11156 4145
rect 11116 3977 11156 4096
rect 11404 4136 11444 4171
rect 11404 4085 11444 4096
rect 11500 4136 11540 4255
rect 11500 4087 11540 4096
rect 11596 4136 11636 4339
rect 11788 4313 11828 4684
rect 11884 4675 11924 4684
rect 11980 4556 12020 5599
rect 12076 5144 12116 5608
rect 12172 5648 12212 5659
rect 12172 5573 12212 5608
rect 12171 5564 12213 5573
rect 12171 5524 12172 5564
rect 12212 5524 12213 5564
rect 12171 5515 12213 5524
rect 12076 5095 12116 5104
rect 11884 4516 12020 4556
rect 12748 4808 12788 4817
rect 11787 4304 11829 4313
rect 11787 4264 11788 4304
rect 11828 4264 11829 4304
rect 11787 4255 11829 4264
rect 11884 4229 11924 4516
rect 11979 4304 12021 4313
rect 11979 4264 11980 4304
rect 12020 4264 12021 4304
rect 11979 4255 12021 4264
rect 11883 4220 11925 4229
rect 11883 4180 11884 4220
rect 11924 4180 11925 4220
rect 11883 4171 11925 4180
rect 11596 4087 11636 4096
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 11884 4136 11924 4171
rect 11788 4002 11828 4087
rect 11884 4086 11924 4096
rect 11980 4136 12020 4255
rect 12171 4220 12213 4229
rect 11980 4087 12020 4096
rect 12076 4180 12172 4220
rect 12212 4180 12213 4220
rect 12076 4136 12116 4180
rect 12171 4171 12213 4180
rect 12076 4087 12116 4096
rect 11320 3977 11360 3996
rect 10828 3968 10868 3977
rect 10635 3884 10677 3893
rect 10635 3844 10636 3884
rect 10676 3844 10677 3884
rect 10635 3835 10677 3844
rect 10828 3557 10868 3928
rect 11115 3968 11157 3977
rect 11115 3928 11116 3968
rect 11156 3928 11157 3968
rect 11115 3919 11157 3928
rect 11308 3968 11360 3977
rect 12268 3968 12308 3977
rect 11348 3928 11444 3968
rect 11308 3919 11348 3928
rect 11307 3632 11349 3641
rect 11307 3592 11308 3632
rect 11348 3592 11349 3632
rect 11307 3583 11349 3592
rect 10827 3548 10869 3557
rect 10827 3508 10828 3548
rect 10868 3508 10869 3548
rect 10827 3499 10869 3508
rect 11308 3464 11348 3583
rect 11308 3415 11348 3424
rect 10252 2575 10292 2584
rect 10636 3212 10676 3221
rect 10636 2624 10676 3172
rect 11404 2717 11444 3928
rect 11884 3928 12268 3968
rect 11884 3716 11924 3928
rect 12268 3919 12308 3928
rect 12748 3809 12788 4768
rect 12075 3800 12117 3809
rect 12075 3760 12076 3800
rect 12116 3760 12117 3800
rect 12075 3751 12117 3760
rect 12747 3800 12789 3809
rect 12747 3760 12748 3800
rect 12788 3760 12789 3800
rect 12747 3751 12789 3760
rect 11692 3676 11924 3716
rect 11692 3548 11732 3676
rect 11692 3499 11732 3508
rect 12076 3464 12116 3751
rect 12844 3464 12884 6448
rect 12939 6439 12981 6448
rect 12940 6354 12980 6439
rect 12940 5648 12980 5659
rect 13132 5657 13172 6952
rect 13612 6488 13652 6497
rect 13228 6448 13612 6488
rect 12940 5573 12980 5608
rect 13036 5648 13076 5657
rect 12939 5564 12981 5573
rect 12939 5524 12940 5564
rect 12980 5524 12981 5564
rect 12939 5515 12981 5524
rect 13036 5153 13076 5608
rect 13131 5648 13173 5657
rect 13131 5608 13132 5648
rect 13172 5608 13173 5648
rect 13131 5599 13173 5608
rect 13228 5648 13268 6448
rect 13612 6439 13652 6448
rect 13900 6488 13940 6497
rect 13940 6448 14228 6488
rect 13900 6439 13940 6448
rect 14092 6320 14132 6329
rect 13804 6280 14092 6320
rect 13612 6236 13652 6245
rect 13228 5599 13268 5608
rect 13420 6196 13612 6236
rect 13420 5648 13460 6196
rect 13612 6187 13652 6196
rect 13420 5599 13460 5608
rect 13804 5648 13844 6280
rect 14092 6271 14132 6280
rect 13804 5599 13844 5608
rect 13132 5514 13172 5599
rect 14188 5489 14228 6448
rect 14187 5480 14229 5489
rect 14187 5440 14188 5480
rect 14228 5440 14229 5480
rect 14187 5431 14229 5440
rect 13035 5144 13077 5153
rect 13035 5104 13036 5144
rect 13076 5104 13077 5144
rect 13035 5095 13077 5104
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 13132 4304 13172 4313
rect 12940 4264 13132 4304
rect 12940 4136 12980 4264
rect 13132 4255 13172 4264
rect 13324 4145 13364 4927
rect 14187 4808 14229 4817
rect 14187 4768 14188 4808
rect 14228 4768 14229 4808
rect 14187 4759 14229 4768
rect 13996 4724 14036 4733
rect 13804 4684 13996 4724
rect 13419 4304 13461 4313
rect 13419 4264 13420 4304
rect 13460 4264 13461 4304
rect 13419 4255 13461 4264
rect 12940 4087 12980 4096
rect 13131 4136 13173 4145
rect 13131 4096 13132 4136
rect 13172 4096 13173 4136
rect 13131 4087 13173 4096
rect 13323 4136 13365 4145
rect 13323 4096 13324 4136
rect 13364 4096 13365 4136
rect 13323 4087 13365 4096
rect 13420 4136 13460 4255
rect 13420 4087 13460 4096
rect 13611 4136 13653 4145
rect 13611 4096 13612 4136
rect 13652 4096 13653 4136
rect 13611 4087 13653 4096
rect 13804 4136 13844 4684
rect 13996 4675 14036 4684
rect 14188 4388 14228 4759
rect 14188 4339 14228 4348
rect 13804 4087 13844 4096
rect 13132 4002 13172 4087
rect 13324 4002 13364 4087
rect 13612 4002 13652 4087
rect 14091 3632 14133 3641
rect 14091 3592 14092 3632
rect 14132 3592 14133 3632
rect 14091 3583 14133 3592
rect 14092 3498 14132 3583
rect 12940 3464 12980 3473
rect 12844 3424 12940 3464
rect 12076 3415 12116 3424
rect 12940 3415 12980 3424
rect 14284 2801 14324 7708
rect 14379 7708 14380 7748
rect 14420 7708 14421 7748
rect 14379 7699 14421 7708
rect 14380 7160 14420 7699
rect 14380 7111 14420 7120
rect 14764 7160 14804 7169
rect 14860 7160 14900 7792
rect 14804 7120 14900 7160
rect 15628 7160 15668 7169
rect 14764 7111 14804 7120
rect 15628 7001 15668 7120
rect 14667 6992 14709 7001
rect 14667 6952 14668 6992
rect 14708 6952 14709 6992
rect 14667 6943 14709 6952
rect 15627 6992 15669 7001
rect 15627 6952 15628 6992
rect 15668 6952 15669 6992
rect 15627 6943 15669 6952
rect 14668 6497 14708 6943
rect 14667 6488 14709 6497
rect 14667 6448 14668 6488
rect 14708 6448 14709 6488
rect 14667 6439 14709 6448
rect 15532 6488 15572 6497
rect 14668 5648 14708 6439
rect 14668 5599 14708 5608
rect 15532 5573 15572 6448
rect 15820 6320 15860 7960
rect 16203 7748 16245 7757
rect 16203 7708 16204 7748
rect 16244 7708 16245 7748
rect 16203 7699 16245 7708
rect 16204 7614 16244 7699
rect 16107 6908 16149 6917
rect 16396 6908 16436 8623
rect 16107 6868 16108 6908
rect 16148 6868 16149 6908
rect 16107 6859 16149 6868
rect 16204 6868 16436 6908
rect 15820 6280 16052 6320
rect 15819 5900 15861 5909
rect 15819 5860 15820 5900
rect 15860 5860 15861 5900
rect 15819 5851 15861 5860
rect 15820 5766 15860 5851
rect 15531 5564 15573 5573
rect 15531 5524 15532 5564
rect 15572 5524 15573 5564
rect 15531 5515 15573 5524
rect 16012 5396 16052 6280
rect 16108 5648 16148 6859
rect 16204 6320 16244 6868
rect 16299 6656 16341 6665
rect 16299 6616 16300 6656
rect 16340 6616 16341 6656
rect 16299 6607 16341 6616
rect 16204 5825 16244 6280
rect 16203 5816 16245 5825
rect 16203 5776 16204 5816
rect 16244 5776 16245 5816
rect 16203 5767 16245 5776
rect 16108 5599 16148 5608
rect 16204 5648 16244 5657
rect 16204 5405 16244 5608
rect 16300 5564 16340 6607
rect 16395 6488 16437 6497
rect 16395 6448 16396 6488
rect 16436 6448 16437 6488
rect 16395 6439 16437 6448
rect 16396 6354 16436 6439
rect 16300 5515 16340 5524
rect 16396 5648 16436 5657
rect 16203 5396 16245 5405
rect 16012 5356 16148 5396
rect 16011 5060 16053 5069
rect 16011 5020 16012 5060
rect 16052 5020 16053 5060
rect 16011 5011 16053 5020
rect 14668 4976 14708 4985
rect 14668 3641 14708 4936
rect 15916 4976 15956 4985
rect 15052 4808 15092 4817
rect 15052 4061 15092 4768
rect 15339 4136 15381 4145
rect 15339 4096 15340 4136
rect 15380 4096 15381 4136
rect 15339 4087 15381 4096
rect 15051 4052 15093 4061
rect 15051 4012 15052 4052
rect 15092 4012 15093 4052
rect 15051 4003 15093 4012
rect 15340 4002 15380 4087
rect 15723 3968 15765 3977
rect 15723 3928 15724 3968
rect 15764 3928 15765 3968
rect 15723 3919 15765 3928
rect 14667 3632 14709 3641
rect 14667 3592 14668 3632
rect 14708 3592 14709 3632
rect 14667 3583 14709 3592
rect 15724 3137 15764 3919
rect 15916 3641 15956 4936
rect 16012 4926 16052 5011
rect 16108 4985 16148 5356
rect 16203 5356 16204 5396
rect 16244 5356 16245 5396
rect 16203 5347 16245 5356
rect 16396 5312 16436 5608
rect 16300 5272 16436 5312
rect 16107 4976 16149 4985
rect 16107 4936 16108 4976
rect 16148 4936 16149 4976
rect 16107 4927 16149 4936
rect 16108 4842 16148 4927
rect 16300 4892 16340 5272
rect 16395 5144 16437 5153
rect 16395 5104 16396 5144
rect 16436 5104 16437 5144
rect 16395 5095 16437 5104
rect 16396 5060 16436 5095
rect 16396 5009 16436 5020
rect 16395 4892 16437 4901
rect 16300 4852 16396 4892
rect 16436 4852 16437 4892
rect 16395 4843 16437 4852
rect 16395 4472 16437 4481
rect 16395 4432 16396 4472
rect 16436 4432 16437 4472
rect 16395 4423 16437 4432
rect 16396 4229 16436 4423
rect 16395 4220 16437 4229
rect 16395 4180 16396 4220
rect 16436 4180 16437 4220
rect 16395 4171 16437 4180
rect 16204 4136 16244 4145
rect 16107 4052 16149 4061
rect 16204 4052 16244 4096
rect 16107 4012 16108 4052
rect 16148 4012 16244 4052
rect 16107 4003 16149 4012
rect 16299 3884 16341 3893
rect 16299 3844 16300 3884
rect 16340 3844 16341 3884
rect 16299 3835 16341 3844
rect 15820 3632 15860 3641
rect 15820 3305 15860 3592
rect 15915 3632 15957 3641
rect 15915 3592 15916 3632
rect 15956 3592 16052 3632
rect 15915 3583 15957 3592
rect 15916 3464 15956 3473
rect 15916 3380 15956 3424
rect 16012 3380 16052 3592
rect 16300 3473 16340 3835
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 16299 3415 16341 3424
rect 16396 3464 16436 4171
rect 16492 4145 16532 8800
rect 16588 8261 16628 9304
rect 16684 9269 16724 10312
rect 16780 10025 16820 10387
rect 16779 10016 16821 10025
rect 16779 9976 16780 10016
rect 16820 9976 16821 10016
rect 16779 9967 16821 9976
rect 16876 9680 16916 10984
rect 16971 11024 17013 11033
rect 16971 10984 16972 11024
rect 17012 10984 17013 11024
rect 16971 10975 17013 10984
rect 17356 11024 17396 11033
rect 16972 9773 17012 10975
rect 17260 10184 17300 10193
rect 17067 9848 17109 9857
rect 17067 9808 17068 9848
rect 17108 9808 17109 9848
rect 17067 9799 17109 9808
rect 16971 9764 17013 9773
rect 16971 9724 16972 9764
rect 17012 9724 17013 9764
rect 16971 9715 17013 9724
rect 16876 9631 16916 9640
rect 17068 9521 17108 9799
rect 17260 9689 17300 10144
rect 17259 9680 17301 9689
rect 17259 9640 17260 9680
rect 17300 9640 17301 9680
rect 17259 9631 17301 9640
rect 17356 9605 17396 10984
rect 17452 11024 17492 11033
rect 17452 10865 17492 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 17548 10890 17588 10975
rect 17451 10856 17493 10865
rect 17451 10816 17452 10856
rect 17492 10816 17493 10856
rect 17451 10807 17493 10816
rect 17644 10445 17684 11227
rect 17931 11108 17973 11117
rect 17931 11068 17932 11108
rect 17972 11068 17973 11108
rect 17931 11059 17973 11068
rect 17739 10940 17781 10949
rect 17739 10900 17740 10940
rect 17780 10900 17781 10940
rect 17739 10891 17781 10900
rect 17740 10806 17780 10891
rect 17643 10436 17685 10445
rect 17643 10396 17644 10436
rect 17684 10396 17685 10436
rect 17643 10387 17685 10396
rect 17739 10184 17781 10193
rect 17739 10144 17740 10184
rect 17780 10144 17781 10184
rect 17739 10135 17781 10144
rect 17932 10184 17972 11059
rect 18028 11033 18068 11488
rect 18124 11479 18164 11488
rect 18123 11360 18165 11369
rect 18123 11320 18124 11360
rect 18164 11320 18165 11360
rect 18412 11360 18452 11656
rect 18795 11696 18837 11705
rect 18795 11656 18796 11696
rect 18836 11656 18837 11696
rect 18795 11647 18837 11656
rect 18796 11562 18836 11647
rect 18412 11320 18836 11360
rect 18123 11311 18165 11320
rect 18027 11024 18069 11033
rect 18027 10984 18028 11024
rect 18068 10984 18069 11024
rect 18027 10975 18069 10984
rect 17932 10135 17972 10144
rect 18028 10184 18068 10975
rect 18124 10184 18164 11311
rect 18603 11192 18645 11201
rect 18603 11152 18604 11192
rect 18644 11152 18645 11192
rect 18603 11143 18645 11152
rect 18412 11024 18452 11033
rect 18412 10781 18452 10984
rect 18604 11024 18644 11143
rect 18604 10975 18644 10984
rect 18796 10865 18836 11320
rect 18795 10856 18837 10865
rect 18795 10816 18796 10856
rect 18836 10816 18837 10856
rect 18795 10807 18837 10816
rect 18411 10772 18453 10781
rect 18411 10732 18412 10772
rect 18452 10732 18453 10772
rect 18411 10723 18453 10732
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 18219 10436 18261 10445
rect 18219 10396 18220 10436
rect 18260 10396 18261 10436
rect 18219 10387 18261 10396
rect 18699 10436 18741 10445
rect 18699 10396 18700 10436
rect 18740 10396 18741 10436
rect 18699 10387 18741 10396
rect 18220 10302 18260 10387
rect 18603 10352 18645 10361
rect 18603 10312 18604 10352
rect 18644 10312 18645 10352
rect 18603 10303 18645 10312
rect 18604 10184 18644 10303
rect 18124 10144 18260 10184
rect 18028 10135 18068 10144
rect 17740 10050 17780 10135
rect 17836 10016 17876 10025
rect 17876 9976 17972 10016
rect 17836 9967 17876 9976
rect 17355 9596 17397 9605
rect 17355 9556 17356 9596
rect 17396 9556 17397 9596
rect 17355 9547 17397 9556
rect 16779 9512 16821 9521
rect 16779 9472 16780 9512
rect 16820 9472 16821 9512
rect 16779 9463 16821 9472
rect 16972 9512 17012 9521
rect 16780 9378 16820 9463
rect 16683 9260 16725 9269
rect 16683 9220 16684 9260
rect 16724 9220 16725 9260
rect 16683 9211 16725 9220
rect 16972 8513 17012 9472
rect 17067 9512 17109 9521
rect 17260 9512 17300 9521
rect 17067 9472 17068 9512
rect 17108 9472 17109 9512
rect 17067 9463 17109 9472
rect 17164 9472 17260 9512
rect 17068 8672 17108 9463
rect 17164 8924 17204 9472
rect 17260 9463 17300 9472
rect 17452 9512 17492 9521
rect 17259 9260 17301 9269
rect 17259 9220 17260 9260
rect 17300 9220 17301 9260
rect 17259 9211 17301 9220
rect 17260 9126 17300 9211
rect 17164 8875 17204 8884
rect 17452 8840 17492 9472
rect 17547 9512 17589 9521
rect 17547 9472 17548 9512
rect 17588 9472 17589 9512
rect 17547 9463 17589 9472
rect 17739 9512 17781 9521
rect 17739 9472 17740 9512
rect 17780 9472 17781 9512
rect 17739 9463 17781 9472
rect 17836 9512 17876 9521
rect 17548 9378 17588 9463
rect 17740 9378 17780 9463
rect 17643 9344 17685 9353
rect 17643 9304 17644 9344
rect 17684 9304 17685 9344
rect 17643 9295 17685 9304
rect 17260 8800 17492 8840
rect 17164 8672 17204 8681
rect 17068 8632 17164 8672
rect 17164 8623 17204 8632
rect 16971 8504 17013 8513
rect 16971 8464 16972 8504
rect 17012 8464 17013 8504
rect 16971 8455 17013 8464
rect 17260 8429 17300 8800
rect 17355 8672 17397 8681
rect 17548 8672 17588 8681
rect 17355 8632 17356 8672
rect 17396 8632 17397 8672
rect 17355 8623 17397 8632
rect 17452 8632 17548 8672
rect 17356 8538 17396 8623
rect 17259 8420 17301 8429
rect 17259 8380 17260 8420
rect 17300 8380 17301 8420
rect 17259 8371 17301 8380
rect 16587 8252 16629 8261
rect 16587 8212 16588 8252
rect 16628 8212 16629 8252
rect 16587 8203 16629 8212
rect 17067 8252 17109 8261
rect 17067 8212 17068 8252
rect 17108 8212 17109 8252
rect 17067 8203 17109 8212
rect 16876 8000 16916 8009
rect 17068 8000 17108 8203
rect 17356 8168 17396 8177
rect 17452 8168 17492 8632
rect 17548 8623 17588 8632
rect 17644 8588 17684 9295
rect 17836 8849 17876 9472
rect 17835 8840 17877 8849
rect 17835 8800 17836 8840
rect 17876 8800 17877 8840
rect 17835 8791 17877 8800
rect 17644 8539 17684 8548
rect 17740 8672 17780 8681
rect 17740 8168 17780 8632
rect 17836 8672 17876 8681
rect 17932 8672 17972 9976
rect 18028 9512 18068 9521
rect 18068 9472 18164 9512
rect 18028 9463 18068 9472
rect 18027 9344 18069 9353
rect 18027 9304 18028 9344
rect 18068 9304 18069 9344
rect 18027 9295 18069 9304
rect 18028 9210 18068 9295
rect 18124 8924 18164 9472
rect 18220 9353 18260 10144
rect 18604 10135 18644 10144
rect 18507 10100 18549 10109
rect 18507 10060 18508 10100
rect 18548 10060 18549 10100
rect 18507 10051 18549 10060
rect 18508 9966 18548 10051
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18316 9378 18356 9463
rect 18219 9344 18261 9353
rect 18219 9304 18220 9344
rect 18260 9304 18261 9344
rect 18219 9295 18261 9304
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 18316 8924 18356 8933
rect 18124 8884 18316 8924
rect 18316 8875 18356 8884
rect 18700 8840 18740 10387
rect 18796 9773 18836 10807
rect 18988 10445 19028 11824
rect 19084 11780 19124 12319
rect 19179 12116 19221 12125
rect 19179 12076 19180 12116
rect 19220 12076 19221 12116
rect 19179 12067 19221 12076
rect 19084 11117 19124 11740
rect 19180 11696 19220 12067
rect 19180 11537 19220 11656
rect 19179 11528 19221 11537
rect 19179 11488 19180 11528
rect 19220 11488 19221 11528
rect 19179 11479 19221 11488
rect 19276 11285 19316 12412
rect 19468 12452 19508 12461
rect 19372 12368 19412 12377
rect 19372 11711 19412 12328
rect 19468 12293 19508 12412
rect 19947 12368 19989 12377
rect 20140 12368 20180 12991
rect 20236 12881 20276 16024
rect 20428 16015 20468 16024
rect 20428 15569 20468 15654
rect 20332 15560 20372 15569
rect 20332 15392 20372 15520
rect 20427 15560 20469 15569
rect 20524 15560 20564 16192
rect 20620 16183 20660 16192
rect 20811 16232 20853 16241
rect 20811 16192 20812 16232
rect 20852 16192 20853 16232
rect 20811 16183 20853 16192
rect 20908 16232 20948 16267
rect 20812 16098 20852 16183
rect 20908 16181 20948 16192
rect 20907 16064 20949 16073
rect 20907 16024 20908 16064
rect 20948 16024 20949 16064
rect 20907 16015 20949 16024
rect 20908 15930 20948 16015
rect 20427 15520 20428 15560
rect 20468 15520 20564 15560
rect 20620 15560 20660 15569
rect 20427 15511 20469 15520
rect 20620 15392 20660 15520
rect 20332 15352 20660 15392
rect 20716 15560 20756 15569
rect 20332 14720 20372 15352
rect 20619 15140 20661 15149
rect 20619 15100 20620 15140
rect 20660 15100 20661 15140
rect 20619 15091 20661 15100
rect 20620 14813 20660 15091
rect 20716 14981 20756 15520
rect 20812 15560 20852 15569
rect 20812 15401 20852 15520
rect 20907 15560 20949 15569
rect 20907 15520 20908 15560
rect 20948 15520 20949 15560
rect 20907 15511 20949 15520
rect 20908 15426 20948 15511
rect 20811 15392 20853 15401
rect 20811 15352 20812 15392
rect 20852 15352 20853 15392
rect 20811 15343 20853 15352
rect 20715 14972 20757 14981
rect 20715 14932 20716 14972
rect 20756 14932 20757 14972
rect 20715 14923 20757 14932
rect 21004 14888 21044 17032
rect 21196 17072 21236 17081
rect 21099 16820 21141 16829
rect 21099 16780 21100 16820
rect 21140 16780 21141 16820
rect 21099 16771 21141 16780
rect 21100 16686 21140 16771
rect 21196 15737 21236 17032
rect 21675 17072 21717 17081
rect 21675 17032 21676 17072
rect 21716 17032 21717 17072
rect 21675 17023 21717 17032
rect 21964 17072 22004 17081
rect 22060 17072 22100 18367
rect 22251 17744 22293 17753
rect 22251 17704 22252 17744
rect 22292 17704 22293 17744
rect 22251 17695 22293 17704
rect 22156 17576 22196 17585
rect 22156 17081 22196 17536
rect 22252 17156 22292 17695
rect 22348 17576 22388 17585
rect 22444 17576 22484 18544
rect 22623 18535 22676 18544
rect 22731 18544 22732 18584
rect 22772 18544 22773 18584
rect 22731 18535 22773 18544
rect 22636 18425 22676 18535
rect 22635 18416 22677 18425
rect 22635 18376 22636 18416
rect 22676 18376 22677 18416
rect 22635 18367 22677 18376
rect 22827 17744 22869 17753
rect 22827 17704 22828 17744
rect 22868 17704 22869 17744
rect 22827 17695 22869 17704
rect 23787 17744 23829 17753
rect 23787 17704 23788 17744
rect 23828 17704 23829 17744
rect 23787 17695 23829 17704
rect 22539 17660 22581 17669
rect 22539 17620 22540 17660
rect 22580 17620 22581 17660
rect 22539 17611 22581 17620
rect 22388 17536 22484 17576
rect 22348 17527 22388 17536
rect 22540 17240 22580 17611
rect 22828 17610 22868 17695
rect 23788 17610 23828 17695
rect 22252 17107 22292 17116
rect 22348 17200 22540 17240
rect 22004 17032 22100 17072
rect 21964 17023 22004 17032
rect 21579 16400 21621 16409
rect 21579 16360 21580 16400
rect 21620 16360 21621 16400
rect 21579 16351 21621 16360
rect 21580 16316 21620 16351
rect 21580 16073 21620 16276
rect 21676 16241 21716 17023
rect 22060 16409 22100 17032
rect 22155 17072 22197 17081
rect 22155 17032 22156 17072
rect 22196 17032 22197 17072
rect 22155 17023 22197 17032
rect 22348 17072 22388 17200
rect 22540 17191 22580 17200
rect 23884 17165 23924 19039
rect 24364 19004 24404 19207
rect 24076 18964 24404 19004
rect 23883 17156 23925 17165
rect 23883 17116 23884 17156
rect 23924 17116 23925 17156
rect 23883 17107 23925 17116
rect 22348 17023 22388 17032
rect 22636 17072 22676 17083
rect 22636 16997 22676 17032
rect 22635 16988 22677 16997
rect 22635 16948 22636 16988
rect 22676 16948 22677 16988
rect 22635 16939 22677 16948
rect 22828 16820 22868 16829
rect 22828 16736 22868 16780
rect 22923 16736 22965 16745
rect 22828 16696 22924 16736
rect 22964 16696 22965 16736
rect 21772 16400 21812 16409
rect 22059 16400 22101 16409
rect 21812 16360 22004 16400
rect 21772 16351 21812 16360
rect 21675 16232 21717 16241
rect 21772 16232 21812 16241
rect 21675 16192 21676 16232
rect 21716 16192 21772 16232
rect 21675 16183 21717 16192
rect 21772 16183 21812 16192
rect 21676 16098 21716 16183
rect 21579 16064 21621 16073
rect 21579 16024 21580 16064
rect 21620 16024 21621 16064
rect 21579 16015 21621 16024
rect 21195 15728 21237 15737
rect 21195 15688 21196 15728
rect 21236 15688 21237 15728
rect 21195 15679 21237 15688
rect 21772 15732 21812 15741
rect 21772 15485 21812 15692
rect 21867 15560 21909 15569
rect 21867 15520 21868 15560
rect 21908 15520 21909 15560
rect 21867 15511 21909 15520
rect 21964 15560 22004 16360
rect 22059 16360 22060 16400
rect 22100 16360 22101 16400
rect 22059 16351 22101 16360
rect 21771 15476 21813 15485
rect 21771 15436 21772 15476
rect 21812 15436 21813 15476
rect 21771 15427 21813 15436
rect 21868 15426 21908 15511
rect 21387 15224 21429 15233
rect 21387 15184 21388 15224
rect 21428 15184 21429 15224
rect 21387 15175 21429 15184
rect 21291 14972 21333 14981
rect 21291 14932 21292 14972
rect 21332 14932 21333 14972
rect 21291 14923 21333 14932
rect 21004 14839 21044 14848
rect 20619 14804 20661 14813
rect 20619 14764 20620 14804
rect 20660 14764 20661 14804
rect 20619 14755 20661 14764
rect 20908 14804 20948 14813
rect 20332 14671 20372 14680
rect 20427 14720 20469 14729
rect 20427 14680 20428 14720
rect 20468 14680 20469 14720
rect 20427 14671 20469 14680
rect 20524 14720 20564 14729
rect 20428 14586 20468 14671
rect 20427 13964 20469 13973
rect 20427 13924 20428 13964
rect 20468 13924 20469 13964
rect 20427 13915 20469 13924
rect 20332 13796 20372 13807
rect 20332 13721 20372 13756
rect 20331 13712 20373 13721
rect 20331 13672 20332 13712
rect 20372 13672 20373 13712
rect 20331 13663 20373 13672
rect 20428 13208 20468 13915
rect 20524 13469 20564 14680
rect 20620 14720 20660 14755
rect 20812 14720 20852 14729
rect 20620 14669 20660 14680
rect 20716 14680 20812 14720
rect 20619 14552 20661 14561
rect 20619 14512 20620 14552
rect 20660 14512 20661 14552
rect 20619 14503 20661 14512
rect 20620 14048 20660 14503
rect 20716 14141 20756 14680
rect 20812 14671 20852 14680
rect 20908 14216 20948 14764
rect 21100 14804 21140 14813
rect 21003 14468 21045 14477
rect 21100 14468 21140 14764
rect 21196 14720 21236 14731
rect 21196 14645 21236 14680
rect 21195 14636 21237 14645
rect 21195 14596 21196 14636
rect 21236 14596 21237 14636
rect 21195 14587 21237 14596
rect 21003 14428 21004 14468
rect 21044 14428 21140 14468
rect 21003 14419 21045 14428
rect 20812 14176 20948 14216
rect 20715 14132 20757 14141
rect 20715 14092 20716 14132
rect 20756 14092 20757 14132
rect 20715 14083 20757 14092
rect 20620 13999 20660 14008
rect 20716 14048 20756 14083
rect 20523 13460 20565 13469
rect 20716 13460 20756 14008
rect 20812 13721 20852 14176
rect 20908 14048 20948 14057
rect 20908 13805 20948 14008
rect 21004 14048 21044 14419
rect 21100 14225 21140 14310
rect 21099 14216 21141 14225
rect 21099 14176 21100 14216
rect 21140 14176 21141 14216
rect 21099 14167 21141 14176
rect 21004 13999 21044 14008
rect 21105 14048 21145 14057
rect 21105 13889 21145 14008
rect 21104 13880 21146 13889
rect 21104 13840 21105 13880
rect 21145 13840 21146 13880
rect 21104 13831 21146 13840
rect 20907 13796 20949 13805
rect 20907 13756 20908 13796
rect 20948 13756 21044 13796
rect 20907 13747 20949 13756
rect 20811 13712 20853 13721
rect 20811 13672 20812 13712
rect 20852 13672 20853 13712
rect 20811 13663 20853 13672
rect 20523 13420 20524 13460
rect 20564 13420 20565 13460
rect 20523 13411 20565 13420
rect 20620 13420 20756 13460
rect 20620 13292 20660 13420
rect 20908 13385 20948 13470
rect 20907 13376 20949 13385
rect 20907 13336 20908 13376
rect 20948 13336 20949 13376
rect 20907 13327 20949 13336
rect 20531 13252 20660 13292
rect 20715 13292 20757 13301
rect 20715 13252 20716 13292
rect 20756 13252 20757 13292
rect 20531 13208 20571 13252
rect 20715 13243 20757 13252
rect 20428 13159 20468 13168
rect 20524 13168 20571 13208
rect 20716 13208 20756 13243
rect 20620 13193 20660 13202
rect 20332 13049 20372 13134
rect 20331 13040 20373 13049
rect 20331 13000 20332 13040
rect 20372 13000 20373 13040
rect 20331 12991 20373 13000
rect 20235 12872 20277 12881
rect 20235 12832 20236 12872
rect 20276 12832 20277 12872
rect 20235 12823 20277 12832
rect 20236 12536 20276 12823
rect 20428 12536 20468 12545
rect 20236 12487 20276 12496
rect 20332 12496 20428 12536
rect 19947 12328 19948 12368
rect 19988 12328 19989 12368
rect 19947 12319 19989 12328
rect 20044 12328 20180 12368
rect 20236 12368 20276 12377
rect 20332 12368 20372 12496
rect 20428 12487 20468 12496
rect 20524 12536 20564 13168
rect 20716 13157 20756 13168
rect 20908 13208 20948 13217
rect 20620 12797 20660 13153
rect 20908 12881 20948 13168
rect 20907 12872 20949 12881
rect 20907 12832 20908 12872
rect 20948 12832 20949 12872
rect 20907 12823 20949 12832
rect 20619 12788 20661 12797
rect 20619 12748 20620 12788
rect 20660 12748 20661 12788
rect 20619 12739 20661 12748
rect 20812 12629 20852 12660
rect 20811 12620 20853 12629
rect 20811 12580 20812 12620
rect 20852 12580 20853 12620
rect 20811 12571 20853 12580
rect 20276 12328 20372 12368
rect 19467 12284 19509 12293
rect 19467 12244 19468 12284
rect 19508 12244 19509 12284
rect 19467 12235 19509 12244
rect 19372 11696 19892 11711
rect 19372 11671 19852 11696
rect 19852 11647 19892 11656
rect 19948 11696 19988 12319
rect 19948 11647 19988 11656
rect 20044 11696 20084 12328
rect 20236 12319 20276 12328
rect 20428 12293 20468 12378
rect 20427 12284 20469 12293
rect 20427 12244 20428 12284
rect 20468 12244 20469 12284
rect 20427 12235 20469 12244
rect 20524 12116 20564 12496
rect 20716 12536 20756 12545
rect 20716 12125 20756 12496
rect 20812 12536 20852 12571
rect 20913 12536 20953 12545
rect 20332 12076 20564 12116
rect 20715 12116 20757 12125
rect 20715 12076 20716 12116
rect 20756 12076 20757 12116
rect 20235 12032 20277 12041
rect 20235 11992 20236 12032
rect 20276 11992 20277 12032
rect 20235 11983 20277 11992
rect 20044 11647 20084 11656
rect 20236 11696 20276 11983
rect 20332 11705 20372 12076
rect 20715 12067 20757 12076
rect 20523 11948 20565 11957
rect 20812 11948 20852 12496
rect 20908 12496 20913 12536
rect 20908 12487 20953 12496
rect 20908 12041 20948 12487
rect 20907 12032 20949 12041
rect 20907 11992 20908 12032
rect 20948 11992 20949 12032
rect 20907 11983 20949 11992
rect 20523 11908 20524 11948
rect 20564 11908 20565 11948
rect 20523 11899 20565 11908
rect 20620 11908 20852 11948
rect 20524 11711 20564 11899
rect 20620 11789 20660 11908
rect 20907 11864 20949 11873
rect 20907 11824 20908 11864
rect 20948 11824 20949 11864
rect 20907 11815 20949 11824
rect 20619 11780 20661 11789
rect 20619 11740 20620 11780
rect 20660 11740 20661 11780
rect 20619 11731 20661 11740
rect 20776 11780 20818 11789
rect 20776 11740 20777 11780
rect 20817 11740 20818 11780
rect 20776 11731 20818 11740
rect 20236 11647 20276 11656
rect 20331 11696 20373 11705
rect 20331 11656 20332 11696
rect 20372 11656 20373 11696
rect 20524 11662 20564 11671
rect 20620 11696 20660 11731
rect 20331 11647 20373 11656
rect 19756 11537 19796 11622
rect 20332 11562 20372 11647
rect 20620 11612 20660 11656
rect 20777 11711 20817 11731
rect 20777 11645 20817 11671
rect 20524 11572 20660 11612
rect 19755 11528 19797 11537
rect 19755 11488 19756 11528
rect 19796 11488 19797 11528
rect 19755 11479 19797 11488
rect 20428 11528 20468 11537
rect 20428 11369 20468 11488
rect 20524 11453 20564 11572
rect 20715 11528 20757 11537
rect 20620 11488 20716 11528
rect 20756 11488 20757 11528
rect 20523 11444 20565 11453
rect 20523 11404 20524 11444
rect 20564 11404 20565 11444
rect 20523 11395 20565 11404
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 20427 11360 20469 11369
rect 20427 11320 20428 11360
rect 20468 11320 20469 11360
rect 20427 11311 20469 11320
rect 19275 11276 19317 11285
rect 19275 11236 19276 11276
rect 19316 11236 19317 11276
rect 19275 11227 19317 11236
rect 19083 11108 19125 11117
rect 19083 11068 19084 11108
rect 19124 11068 19125 11108
rect 19083 11059 19125 11068
rect 19563 11108 19605 11117
rect 19563 11068 19564 11108
rect 19604 11068 19605 11108
rect 19563 11059 19605 11068
rect 19467 11024 19509 11033
rect 19467 10984 19468 11024
rect 19508 10984 19509 11024
rect 19467 10975 19509 10984
rect 19564 11024 19604 11059
rect 19468 10890 19508 10975
rect 19564 10973 19604 10984
rect 19755 11024 19797 11033
rect 19755 10984 19756 11024
rect 19796 10984 19797 11024
rect 19755 10975 19797 10984
rect 20524 11024 20564 11395
rect 20524 10975 20564 10984
rect 19756 10890 19796 10975
rect 20620 10940 20660 11488
rect 20715 11479 20757 11488
rect 20811 11108 20853 11117
rect 20811 11068 20812 11108
rect 20852 11068 20853 11108
rect 20811 11059 20853 11068
rect 20620 10891 20660 10900
rect 20812 10940 20852 11059
rect 20908 11024 20948 11815
rect 21004 11789 21044 13756
rect 21099 13712 21141 13721
rect 21292 13712 21332 14923
rect 21388 14720 21428 15175
rect 21579 14888 21621 14897
rect 21579 14848 21580 14888
rect 21620 14848 21621 14888
rect 21579 14839 21621 14848
rect 21388 14671 21428 14680
rect 21483 14720 21525 14729
rect 21483 14680 21484 14720
rect 21524 14680 21525 14720
rect 21483 14671 21525 14680
rect 21580 14720 21620 14839
rect 21580 14671 21620 14680
rect 21484 14586 21524 14671
rect 21867 14636 21909 14645
rect 21867 14596 21868 14636
rect 21908 14596 21909 14636
rect 21867 14587 21909 14596
rect 21771 14468 21813 14477
rect 21771 14428 21772 14468
rect 21812 14428 21813 14468
rect 21771 14419 21813 14428
rect 21388 14057 21428 14142
rect 21675 14132 21717 14141
rect 21675 14092 21676 14132
rect 21716 14092 21717 14132
rect 21675 14083 21717 14092
rect 21387 14048 21429 14057
rect 21387 14008 21388 14048
rect 21428 14008 21429 14048
rect 21387 13999 21429 14008
rect 21484 13964 21524 13973
rect 21387 13880 21429 13889
rect 21484 13880 21524 13924
rect 21676 13964 21716 14083
rect 21676 13915 21716 13924
rect 21772 14048 21812 14419
rect 21387 13840 21388 13880
rect 21428 13840 21524 13880
rect 21579 13880 21621 13889
rect 21579 13840 21580 13880
rect 21620 13840 21621 13880
rect 21387 13831 21429 13840
rect 21579 13831 21621 13840
rect 21580 13746 21620 13831
rect 21099 13672 21100 13712
rect 21140 13672 21141 13712
rect 21099 13663 21141 13672
rect 21196 13672 21332 13712
rect 21100 13208 21140 13663
rect 21100 13159 21140 13168
rect 21196 13208 21236 13672
rect 21772 13628 21812 14008
rect 21868 13973 21908 14587
rect 21964 14309 22004 15520
rect 22155 15476 22197 15485
rect 22155 15436 22156 15476
rect 22196 15436 22197 15476
rect 22155 15427 22197 15436
rect 22156 15056 22196 15427
rect 22251 15308 22293 15317
rect 22251 15268 22252 15308
rect 22292 15268 22293 15308
rect 22251 15259 22293 15268
rect 22252 15174 22292 15259
rect 22156 15016 22292 15056
rect 22252 14888 22292 15016
rect 22252 14839 22292 14848
rect 22156 14804 22196 14813
rect 22060 14720 22100 14729
rect 22060 14561 22100 14680
rect 22059 14552 22101 14561
rect 22059 14512 22060 14552
rect 22100 14512 22101 14552
rect 22059 14503 22101 14512
rect 21963 14300 22005 14309
rect 21963 14260 21964 14300
rect 22004 14260 22005 14300
rect 21963 14251 22005 14260
rect 21964 14048 22004 14251
rect 21964 13999 22004 14008
rect 21867 13964 21909 13973
rect 21867 13924 21868 13964
rect 21908 13924 21909 13964
rect 21867 13915 21909 13924
rect 21868 13712 21908 13915
rect 21868 13672 22004 13712
rect 21484 13588 21812 13628
rect 21387 13376 21429 13385
rect 21387 13336 21388 13376
rect 21428 13336 21429 13376
rect 21387 13327 21429 13336
rect 21196 13159 21236 13168
rect 21292 13208 21332 13217
rect 21388 13208 21428 13327
rect 21332 13168 21428 13208
rect 21292 13159 21332 13168
rect 21388 13040 21428 13049
rect 21196 13000 21388 13040
rect 21099 12956 21141 12965
rect 21099 12916 21100 12956
rect 21140 12916 21141 12956
rect 21099 12907 21141 12916
rect 21100 12461 21140 12907
rect 21196 12536 21236 13000
rect 21388 12991 21428 13000
rect 21484 12788 21524 13588
rect 21292 12748 21524 12788
rect 21580 13208 21620 13217
rect 21292 12629 21332 12748
rect 21580 12704 21620 13168
rect 21772 13208 21812 13217
rect 21812 13168 21908 13208
rect 21772 13159 21812 13168
rect 21676 13124 21716 13133
rect 21676 12713 21716 13084
rect 21388 12664 21620 12704
rect 21675 12704 21717 12713
rect 21675 12664 21676 12704
rect 21716 12664 21717 12704
rect 21291 12620 21333 12629
rect 21291 12580 21292 12620
rect 21332 12580 21333 12620
rect 21291 12571 21333 12580
rect 21196 12487 21236 12496
rect 21388 12536 21428 12664
rect 21675 12655 21717 12664
rect 21099 12452 21141 12461
rect 21099 12412 21100 12452
rect 21140 12412 21141 12452
rect 21099 12403 21141 12412
rect 21291 12452 21333 12461
rect 21291 12412 21292 12452
rect 21332 12412 21333 12452
rect 21291 12403 21333 12412
rect 21196 12284 21236 12293
rect 21100 12244 21196 12284
rect 21003 11780 21045 11789
rect 21003 11740 21004 11780
rect 21044 11740 21045 11780
rect 21003 11731 21045 11740
rect 21100 11696 21140 12244
rect 21196 12235 21236 12244
rect 21100 11647 21140 11656
rect 21195 11696 21237 11705
rect 21195 11656 21196 11696
rect 21236 11656 21237 11696
rect 21195 11647 21237 11656
rect 21196 11562 21236 11647
rect 21292 11285 21332 12403
rect 21388 12377 21428 12496
rect 21484 12536 21524 12545
rect 21676 12536 21716 12545
rect 21524 12496 21676 12536
rect 21484 12487 21524 12496
rect 21676 12487 21716 12496
rect 21771 12536 21813 12545
rect 21771 12496 21772 12536
rect 21812 12496 21813 12536
rect 21771 12487 21813 12496
rect 21772 12402 21812 12487
rect 21868 12377 21908 13168
rect 21387 12368 21429 12377
rect 21387 12328 21388 12368
rect 21428 12328 21429 12368
rect 21387 12319 21429 12328
rect 21867 12368 21909 12377
rect 21867 12328 21868 12368
rect 21908 12328 21909 12368
rect 21867 12319 21909 12328
rect 21964 12368 22004 13672
rect 21964 12319 22004 12328
rect 22156 12209 22196 14764
rect 22347 14804 22389 14813
rect 22347 14764 22348 14804
rect 22388 14764 22389 14804
rect 22347 14755 22389 14764
rect 22348 14670 22388 14755
rect 22443 14720 22485 14729
rect 22443 14680 22444 14720
rect 22484 14680 22485 14720
rect 22443 14671 22485 14680
rect 22444 14586 22484 14671
rect 22347 14552 22389 14561
rect 22347 14512 22348 14552
rect 22388 14512 22389 14552
rect 22347 14503 22389 14512
rect 22251 14468 22293 14477
rect 22251 14428 22252 14468
rect 22292 14428 22293 14468
rect 22251 14419 22293 14428
rect 22252 14216 22292 14419
rect 22252 14167 22292 14176
rect 22348 14216 22388 14503
rect 22635 14300 22677 14309
rect 22635 14260 22636 14300
rect 22676 14260 22677 14300
rect 22635 14251 22677 14260
rect 22444 14216 22484 14225
rect 22348 14176 22444 14216
rect 22251 13964 22293 13973
rect 22251 13924 22252 13964
rect 22292 13924 22293 13964
rect 22251 13915 22293 13924
rect 22252 13208 22292 13915
rect 22348 13292 22388 14176
rect 22444 14167 22484 14176
rect 22636 14048 22676 14251
rect 22636 13999 22676 14008
rect 22348 13243 22388 13252
rect 22252 13159 22292 13168
rect 22443 13208 22485 13217
rect 22443 13168 22444 13208
rect 22484 13168 22485 13208
rect 22443 13159 22485 13168
rect 22732 13208 22772 13217
rect 22444 13074 22484 13159
rect 22636 13040 22676 13049
rect 22252 12536 22292 12545
rect 22252 12377 22292 12496
rect 22347 12536 22389 12545
rect 22347 12496 22348 12536
rect 22388 12496 22389 12536
rect 22347 12487 22389 12496
rect 22636 12536 22676 13000
rect 22251 12368 22293 12377
rect 22251 12328 22252 12368
rect 22292 12328 22293 12368
rect 22251 12319 22293 12328
rect 22348 12209 22388 12487
rect 22155 12200 22197 12209
rect 22155 12160 22156 12200
rect 22196 12160 22197 12200
rect 22155 12151 22197 12160
rect 22347 12200 22389 12209
rect 22347 12160 22348 12200
rect 22388 12160 22389 12200
rect 22347 12151 22389 12160
rect 21387 11864 21429 11873
rect 21387 11824 21388 11864
rect 21428 11824 21429 11864
rect 21387 11815 21429 11824
rect 21388 11696 21428 11815
rect 22156 11789 22196 12151
rect 21640 11780 21682 11789
rect 21640 11740 21641 11780
rect 21681 11740 21682 11780
rect 21640 11731 21682 11740
rect 22155 11780 22197 11789
rect 22155 11740 22156 11780
rect 22196 11740 22197 11780
rect 22155 11731 22197 11740
rect 21641 11711 21681 11731
rect 21388 11647 21428 11656
rect 21484 11696 21524 11705
rect 21388 11528 21428 11537
rect 21291 11276 21333 11285
rect 21291 11236 21292 11276
rect 21332 11236 21333 11276
rect 21291 11227 21333 11236
rect 20908 10975 20948 10984
rect 20812 10891 20852 10900
rect 19659 10856 19701 10865
rect 19659 10816 19660 10856
rect 19700 10816 19701 10856
rect 19659 10807 19701 10816
rect 20716 10856 20756 10865
rect 19276 10772 19316 10781
rect 18987 10436 19029 10445
rect 18987 10396 18988 10436
rect 19028 10396 19029 10436
rect 18987 10387 19029 10396
rect 19276 10193 19316 10732
rect 19371 10520 19413 10529
rect 19371 10480 19372 10520
rect 19412 10480 19413 10520
rect 19371 10471 19413 10480
rect 18892 10184 18932 10193
rect 18892 10100 18932 10144
rect 19275 10184 19317 10193
rect 19275 10144 19276 10184
rect 19316 10144 19317 10184
rect 19275 10135 19317 10144
rect 19372 10100 19412 10471
rect 19660 10184 19700 10807
rect 19755 10772 19797 10781
rect 19755 10732 19756 10772
rect 19796 10732 19797 10772
rect 19755 10723 19797 10732
rect 19756 10638 19796 10723
rect 20619 10688 20661 10697
rect 20619 10648 20620 10688
rect 20660 10648 20661 10688
rect 20619 10639 20661 10648
rect 20331 10352 20373 10361
rect 20331 10312 20332 10352
rect 20372 10312 20373 10352
rect 20331 10303 20373 10312
rect 19660 10135 19700 10144
rect 20235 10184 20277 10193
rect 20235 10144 20236 10184
rect 20276 10144 20277 10184
rect 20235 10135 20277 10144
rect 20332 10184 20372 10303
rect 20332 10135 20372 10144
rect 20428 10184 20468 10193
rect 18892 10060 19220 10100
rect 18795 9764 18837 9773
rect 18795 9724 18796 9764
rect 18836 9724 18837 9764
rect 18795 9715 18837 9724
rect 18892 9344 18932 10060
rect 19180 10016 19220 10060
rect 19372 10051 19412 10060
rect 20236 10050 20276 10135
rect 19180 9967 19220 9976
rect 19083 9932 19125 9941
rect 19083 9892 19084 9932
rect 19124 9892 19125 9932
rect 19083 9883 19125 9892
rect 18892 9295 18932 9304
rect 19084 9512 19124 9883
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 20331 9848 20373 9857
rect 20331 9808 20332 9848
rect 20372 9808 20373 9848
rect 20331 9799 20373 9808
rect 20332 9512 20372 9799
rect 18412 8800 18740 8840
rect 18891 8840 18933 8849
rect 18891 8800 18892 8840
rect 18932 8800 18933 8840
rect 17876 8632 17972 8672
rect 18315 8672 18357 8681
rect 18315 8632 18316 8672
rect 18356 8632 18357 8672
rect 17836 8623 17876 8632
rect 18315 8623 18357 8632
rect 18316 8538 18356 8623
rect 17835 8252 17877 8261
rect 17835 8212 17836 8252
rect 17876 8212 17877 8252
rect 17835 8203 17877 8212
rect 17396 8128 17492 8168
rect 17644 8128 17780 8168
rect 17356 8119 17396 8128
rect 16916 7960 17012 8000
rect 16876 7951 16916 7960
rect 16587 7496 16629 7505
rect 16587 7456 16588 7496
rect 16628 7456 16629 7496
rect 16587 7447 16629 7456
rect 16588 5648 16628 7447
rect 16875 7244 16917 7253
rect 16875 7204 16876 7244
rect 16916 7204 16917 7244
rect 16875 7195 16917 7204
rect 16876 7160 16916 7195
rect 16876 7109 16916 7120
rect 16875 6992 16917 7001
rect 16875 6952 16876 6992
rect 16916 6952 16917 6992
rect 16875 6943 16917 6952
rect 16779 6488 16821 6497
rect 16779 6448 16780 6488
rect 16820 6448 16821 6488
rect 16779 6439 16821 6448
rect 16780 6354 16820 6439
rect 16683 5816 16725 5825
rect 16683 5776 16684 5816
rect 16724 5776 16725 5816
rect 16683 5767 16725 5776
rect 16588 5599 16628 5608
rect 16684 5648 16724 5767
rect 16684 5599 16724 5608
rect 16779 5648 16821 5657
rect 16779 5608 16780 5648
rect 16820 5608 16821 5648
rect 16779 5599 16821 5608
rect 16876 5648 16916 6943
rect 16972 5900 17012 7960
rect 17068 7951 17108 7960
rect 17164 8000 17204 8009
rect 17164 7160 17204 7960
rect 17259 8000 17301 8009
rect 17259 7960 17260 8000
rect 17300 7960 17301 8000
rect 17259 7951 17301 7960
rect 17260 7866 17300 7951
rect 17548 7916 17588 7925
rect 17068 7120 17204 7160
rect 17356 7160 17396 7171
rect 17548 7169 17588 7876
rect 17644 7505 17684 8128
rect 17836 8000 17876 8203
rect 17836 7951 17876 7960
rect 17932 8000 17972 8009
rect 17643 7496 17685 7505
rect 17643 7456 17644 7496
rect 17684 7456 17685 7496
rect 17643 7447 17685 7456
rect 17068 6320 17108 7120
rect 17356 7085 17396 7120
rect 17547 7160 17589 7169
rect 17547 7120 17548 7160
rect 17588 7120 17589 7160
rect 17547 7111 17589 7120
rect 17644 7160 17684 7169
rect 17355 7076 17397 7085
rect 17355 7036 17356 7076
rect 17396 7036 17397 7076
rect 17355 7027 17397 7036
rect 17164 6992 17204 7003
rect 17164 6917 17204 6952
rect 17163 6908 17205 6917
rect 17163 6868 17164 6908
rect 17204 6868 17205 6908
rect 17163 6859 17205 6868
rect 17451 6824 17493 6833
rect 17451 6784 17452 6824
rect 17492 6784 17493 6824
rect 17451 6775 17493 6784
rect 17452 6488 17492 6775
rect 17068 6280 17204 6320
rect 17068 5900 17108 5909
rect 16972 5860 17068 5900
rect 17068 5851 17108 5860
rect 16981 5732 17023 5741
rect 16981 5692 16982 5732
rect 17022 5692 17108 5732
rect 16981 5683 17023 5692
rect 16876 5599 16916 5608
rect 17068 5648 17108 5692
rect 17068 5599 17108 5608
rect 16780 5514 16820 5599
rect 16971 5396 17013 5405
rect 16971 5356 16972 5396
rect 17012 5356 17013 5396
rect 17164 5396 17204 6280
rect 17259 6152 17301 6161
rect 17259 6112 17260 6152
rect 17300 6112 17301 6152
rect 17259 6103 17301 6112
rect 17260 5648 17300 6103
rect 17355 5984 17397 5993
rect 17355 5944 17356 5984
rect 17396 5944 17397 5984
rect 17355 5935 17397 5944
rect 17260 5599 17300 5608
rect 17356 5648 17396 5935
rect 17452 5909 17492 6448
rect 17451 5900 17493 5909
rect 17451 5860 17452 5900
rect 17492 5860 17493 5900
rect 17451 5851 17493 5860
rect 17548 5657 17588 7111
rect 17644 6992 17684 7120
rect 17932 7085 17972 7960
rect 18412 7748 18452 8800
rect 18891 8791 18933 8800
rect 18508 8672 18548 8681
rect 18508 8093 18548 8632
rect 18700 8672 18740 8681
rect 18507 8084 18549 8093
rect 18507 8044 18508 8084
rect 18548 8044 18549 8084
rect 18507 8035 18549 8044
rect 18124 7708 18452 7748
rect 17931 7076 17973 7085
rect 17931 7036 17932 7076
rect 17972 7036 17973 7076
rect 17931 7027 17973 7036
rect 17836 6992 17876 7001
rect 17644 6952 17836 6992
rect 17836 6749 17876 6952
rect 17835 6740 17877 6749
rect 17835 6700 17836 6740
rect 17876 6700 17877 6740
rect 18124 6740 18164 7708
rect 18700 7589 18740 8632
rect 18795 8504 18837 8513
rect 18795 8464 18796 8504
rect 18836 8464 18837 8504
rect 18795 8455 18837 8464
rect 18796 8370 18836 8455
rect 18892 8009 18932 8791
rect 19084 8681 19124 9472
rect 20236 9472 20332 9512
rect 20139 9176 20181 9185
rect 20139 9136 20140 9176
rect 20180 9136 20181 9176
rect 20139 9127 20181 9136
rect 20140 8840 20180 9127
rect 19948 8800 20180 8840
rect 19083 8672 19125 8681
rect 19083 8632 19084 8672
rect 19124 8632 19125 8672
rect 19083 8623 19125 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19852 8672 19892 8681
rect 19756 8538 19796 8623
rect 19852 8513 19892 8632
rect 19948 8672 19988 8800
rect 19948 8623 19988 8632
rect 20044 8672 20084 8681
rect 19851 8504 19893 8513
rect 19851 8464 19852 8504
rect 19892 8464 19893 8504
rect 19851 8455 19893 8464
rect 20044 8429 20084 8632
rect 20043 8420 20085 8429
rect 20043 8380 20044 8420
rect 20084 8380 20085 8420
rect 20043 8371 20085 8380
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 20140 8168 20180 8800
rect 20236 8672 20276 9472
rect 20332 9463 20372 9472
rect 20332 9260 20372 9271
rect 20332 9185 20372 9220
rect 20331 9176 20373 9185
rect 20331 9136 20332 9176
rect 20372 9136 20373 9176
rect 20331 9127 20373 9136
rect 20428 9017 20468 10144
rect 20523 10184 20565 10193
rect 20523 10144 20524 10184
rect 20564 10144 20565 10184
rect 20523 10135 20565 10144
rect 20524 10050 20564 10135
rect 20620 10109 20660 10639
rect 20716 10529 20756 10816
rect 20715 10520 20757 10529
rect 20715 10480 20716 10520
rect 20756 10480 20757 10520
rect 20715 10471 20757 10480
rect 21196 10352 21236 10361
rect 20716 10312 21196 10352
rect 20716 10184 20756 10312
rect 21196 10303 21236 10312
rect 20716 10135 20756 10144
rect 20908 10184 20948 10193
rect 20908 10109 20948 10144
rect 21004 10184 21044 10193
rect 20619 10100 20661 10109
rect 20619 10060 20620 10100
rect 20660 10060 20661 10100
rect 20619 10051 20661 10060
rect 20811 10100 20853 10109
rect 20811 10060 20812 10100
rect 20852 10060 20853 10100
rect 20908 10100 20960 10109
rect 20908 10060 20919 10100
rect 20959 10060 20960 10100
rect 20811 10051 20853 10060
rect 20918 10051 20960 10060
rect 20812 9966 20852 10051
rect 21004 9689 21044 10144
rect 21003 9680 21045 9689
rect 21003 9640 21004 9680
rect 21044 9640 21045 9680
rect 21003 9631 21045 9640
rect 20812 9521 20852 9606
rect 20524 9512 20564 9521
rect 20716 9512 20756 9521
rect 20564 9472 20660 9512
rect 20524 9463 20564 9472
rect 20427 9008 20469 9017
rect 20427 8968 20428 9008
rect 20468 8968 20469 9008
rect 20427 8959 20469 8968
rect 20428 8840 20468 8849
rect 20236 8345 20276 8632
rect 20332 8756 20372 8765
rect 20332 8513 20372 8716
rect 20331 8504 20373 8513
rect 20331 8464 20332 8504
rect 20372 8464 20373 8504
rect 20331 8455 20373 8464
rect 20235 8336 20277 8345
rect 20235 8296 20236 8336
rect 20276 8296 20277 8336
rect 20235 8287 20277 8296
rect 20332 8261 20372 8455
rect 20428 8429 20468 8800
rect 20524 8756 20564 8765
rect 20427 8420 20469 8429
rect 20427 8380 20428 8420
rect 20468 8380 20469 8420
rect 20427 8371 20469 8380
rect 20331 8252 20373 8261
rect 20331 8212 20332 8252
rect 20372 8212 20373 8252
rect 20331 8203 20373 8212
rect 20140 8128 20276 8168
rect 18891 8000 18933 8009
rect 18891 7960 18892 8000
rect 18932 7960 18933 8000
rect 18891 7951 18933 7960
rect 18892 7916 18932 7951
rect 20236 7925 20276 8128
rect 20331 8084 20373 8093
rect 20331 8044 20332 8084
rect 20372 8044 20373 8084
rect 20331 8035 20373 8044
rect 20332 8000 20372 8035
rect 20428 8009 20468 8371
rect 18892 7866 18932 7876
rect 20235 7916 20277 7925
rect 20235 7876 20236 7916
rect 20276 7876 20277 7916
rect 20235 7867 20277 7876
rect 19084 7748 19124 7757
rect 19124 7708 19988 7748
rect 19084 7699 19124 7708
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 18699 7580 18741 7589
rect 18699 7540 18700 7580
rect 18740 7540 18741 7580
rect 18699 7531 18741 7540
rect 18507 7412 18549 7421
rect 18507 7372 18508 7412
rect 18548 7372 18549 7412
rect 18507 7363 18549 7372
rect 18508 7253 18548 7363
rect 18507 7244 18549 7253
rect 18507 7204 18508 7244
rect 18548 7204 18549 7244
rect 18507 7195 18549 7204
rect 18508 7160 18548 7195
rect 18988 7169 19028 7254
rect 18508 7110 18548 7120
rect 18699 7160 18741 7169
rect 18699 7120 18700 7160
rect 18740 7120 18741 7160
rect 18699 7111 18741 7120
rect 18796 7160 18836 7169
rect 18700 7026 18740 7111
rect 18796 7001 18836 7120
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 18795 6992 18837 7001
rect 18795 6952 18796 6992
rect 18836 6952 18837 6992
rect 18795 6943 18837 6952
rect 18892 6992 18932 7001
rect 19179 6992 19221 7001
rect 18932 6952 19028 6992
rect 18892 6943 18932 6952
rect 18124 6700 18260 6740
rect 17835 6691 17877 6700
rect 18220 6656 18260 6700
rect 18260 6616 18644 6656
rect 18220 6607 18260 6616
rect 18124 6572 18164 6581
rect 17932 6488 17972 6497
rect 17932 6245 17972 6448
rect 18028 6488 18068 6497
rect 17931 6236 17973 6245
rect 17931 6196 17932 6236
rect 17972 6196 17973 6236
rect 17931 6187 17973 6196
rect 17356 5599 17396 5608
rect 17547 5648 17589 5657
rect 17547 5608 17548 5648
rect 17588 5608 17589 5648
rect 17547 5599 17589 5608
rect 17836 5648 17876 5657
rect 17548 5480 17588 5489
rect 17164 5356 17300 5396
rect 16971 5347 17013 5356
rect 16587 4220 16629 4229
rect 16587 4180 16588 4220
rect 16628 4180 16629 4220
rect 16587 4171 16629 4180
rect 16491 4136 16533 4145
rect 16491 4096 16492 4136
rect 16532 4096 16533 4136
rect 16491 4087 16533 4096
rect 16588 4136 16628 4171
rect 16588 4085 16628 4096
rect 16972 4136 17012 5347
rect 17260 5069 17300 5356
rect 17548 5144 17588 5440
rect 17836 5396 17876 5608
rect 17740 5356 17876 5396
rect 17932 5648 17972 5657
rect 17740 5153 17780 5356
rect 17932 5321 17972 5608
rect 17931 5312 17973 5321
rect 17931 5272 17932 5312
rect 17972 5272 17973 5312
rect 17931 5263 17973 5272
rect 17739 5144 17781 5153
rect 18028 5144 18068 6448
rect 18124 6413 18164 6532
rect 18123 6404 18165 6413
rect 18123 6364 18124 6404
rect 18164 6364 18165 6404
rect 18123 6355 18165 6364
rect 18604 6320 18644 6616
rect 18892 6581 18932 6625
rect 18891 6572 18933 6581
rect 18891 6532 18892 6572
rect 18932 6532 18933 6572
rect 18891 6530 18933 6532
rect 18891 6523 18892 6530
rect 18796 6488 18836 6497
rect 18932 6523 18933 6530
rect 18892 6481 18932 6490
rect 18796 6404 18836 6448
rect 18796 6364 18932 6404
rect 18604 6280 18836 6320
rect 18220 6236 18260 6245
rect 17548 5104 17684 5144
rect 17067 5060 17109 5069
rect 17067 5020 17068 5060
rect 17108 5020 17109 5060
rect 17067 5011 17109 5020
rect 17259 5060 17301 5069
rect 17259 5020 17260 5060
rect 17300 5020 17301 5060
rect 17259 5011 17301 5020
rect 16972 4087 17012 4096
rect 17068 4136 17108 5011
rect 17260 4976 17300 5011
rect 17260 4925 17300 4936
rect 17548 4976 17588 4987
rect 17548 4901 17588 4936
rect 17547 4892 17589 4901
rect 17547 4852 17548 4892
rect 17588 4852 17589 4892
rect 17547 4843 17589 4852
rect 17548 4724 17588 4733
rect 17259 4388 17301 4397
rect 17259 4348 17260 4388
rect 17300 4348 17301 4388
rect 17259 4339 17301 4348
rect 17163 4304 17205 4313
rect 17163 4264 17164 4304
rect 17204 4264 17205 4304
rect 17163 4255 17205 4264
rect 17068 4087 17108 4096
rect 17164 4136 17204 4255
rect 17164 4087 17204 4096
rect 17260 4136 17300 4339
rect 17355 4304 17397 4313
rect 17355 4264 17356 4304
rect 17396 4264 17397 4304
rect 17355 4255 17397 4264
rect 16491 3632 16533 3641
rect 16780 3632 16820 3641
rect 16491 3592 16492 3632
rect 16532 3592 16533 3632
rect 16491 3583 16533 3592
rect 16684 3592 16780 3632
rect 16396 3415 16436 3424
rect 16492 3464 16532 3583
rect 16492 3415 16532 3424
rect 16588 3464 16628 3492
rect 16684 3464 16724 3592
rect 16780 3583 16820 3592
rect 17067 3548 17109 3557
rect 17067 3508 17068 3548
rect 17108 3508 17109 3548
rect 17067 3499 17109 3508
rect 16628 3424 16724 3464
rect 16588 3415 16628 3424
rect 15916 3340 16052 3380
rect 15819 3296 15861 3305
rect 15819 3256 15820 3296
rect 15860 3256 15956 3296
rect 15819 3247 15861 3256
rect 15723 3128 15765 3137
rect 15723 3088 15724 3128
rect 15764 3088 15765 3128
rect 15723 3079 15765 3088
rect 14283 2792 14325 2801
rect 14283 2752 14284 2792
rect 14324 2752 14325 2792
rect 14283 2743 14325 2752
rect 11403 2708 11445 2717
rect 11403 2668 11404 2708
rect 11444 2668 11445 2708
rect 11403 2659 11445 2668
rect 15724 2624 15764 3079
rect 15820 2624 15860 2633
rect 15724 2584 15820 2624
rect 10636 2575 10676 2584
rect 15820 2575 15860 2584
rect 15916 2624 15956 3256
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 15916 1952 15956 2584
rect 16012 2624 16052 3340
rect 16300 3330 16340 3415
rect 16108 3212 16148 3221
rect 16148 3172 16244 3212
rect 16108 3163 16148 3172
rect 16204 2708 16244 3172
rect 16300 2885 16340 2970
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 16587 2792 16629 2801
rect 16587 2752 16588 2792
rect 16628 2752 16629 2792
rect 16587 2743 16629 2752
rect 16204 2668 16436 2708
rect 16012 2129 16052 2584
rect 16107 2624 16149 2633
rect 16107 2584 16108 2624
rect 16148 2584 16149 2624
rect 16107 2575 16149 2584
rect 16300 2624 16340 2668
rect 16300 2575 16340 2584
rect 16108 2490 16148 2575
rect 16396 2549 16436 2668
rect 16492 2624 16532 2635
rect 16395 2540 16437 2549
rect 16395 2500 16396 2540
rect 16436 2500 16437 2540
rect 16395 2491 16437 2500
rect 16492 2213 16532 2584
rect 16588 2624 16628 2743
rect 16588 2575 16628 2584
rect 16684 2297 16724 3424
rect 16876 3464 16916 3473
rect 16779 2876 16821 2885
rect 16779 2836 16780 2876
rect 16820 2836 16821 2876
rect 16779 2827 16821 2836
rect 16780 2742 16820 2827
rect 16876 2633 16916 3424
rect 17068 3414 17108 3499
rect 17260 3464 17300 4096
rect 17260 3415 17300 3424
rect 17356 3464 17396 4255
rect 17548 4061 17588 4684
rect 17644 4313 17684 5104
rect 17739 5104 17740 5144
rect 17780 5104 17781 5144
rect 17739 5095 17781 5104
rect 17932 5104 18068 5144
rect 18124 6196 18220 6236
rect 17835 5060 17877 5069
rect 17835 5020 17836 5060
rect 17876 5020 17877 5060
rect 17835 5011 17877 5020
rect 17740 4976 17780 4987
rect 17740 4901 17780 4936
rect 17836 4976 17876 5011
rect 17836 4925 17876 4936
rect 17739 4892 17781 4901
rect 17739 4852 17740 4892
rect 17780 4852 17781 4892
rect 17739 4843 17781 4852
rect 17835 4808 17877 4817
rect 17835 4768 17836 4808
rect 17876 4768 17877 4808
rect 17835 4759 17877 4768
rect 17739 4388 17781 4397
rect 17739 4348 17740 4388
rect 17780 4348 17781 4388
rect 17739 4339 17781 4348
rect 17643 4304 17685 4313
rect 17643 4264 17644 4304
rect 17684 4264 17685 4304
rect 17643 4255 17685 4264
rect 17644 4136 17684 4255
rect 17644 4087 17684 4096
rect 17740 4136 17780 4339
rect 17836 4313 17876 4759
rect 17835 4304 17877 4313
rect 17835 4264 17836 4304
rect 17876 4264 17877 4304
rect 17932 4304 17972 5104
rect 18027 4976 18069 4985
rect 18027 4936 18028 4976
rect 18068 4936 18069 4976
rect 18027 4927 18069 4936
rect 18028 4842 18068 4927
rect 17932 4264 18068 4304
rect 17835 4255 17877 4264
rect 17836 4136 17876 4255
rect 17932 4136 17972 4145
rect 17836 4096 17932 4136
rect 17740 4087 17780 4096
rect 17547 4052 17589 4061
rect 17547 4012 17548 4052
rect 17588 4012 17589 4052
rect 17547 4003 17589 4012
rect 17451 3968 17493 3977
rect 17451 3928 17452 3968
rect 17492 3928 17493 3968
rect 17451 3919 17493 3928
rect 17835 3968 17877 3977
rect 17835 3928 17836 3968
rect 17876 3928 17877 3968
rect 17835 3919 17877 3928
rect 17356 3415 17396 3424
rect 17452 3464 17492 3919
rect 17739 3884 17781 3893
rect 17739 3844 17740 3884
rect 17780 3844 17781 3884
rect 17739 3835 17781 3844
rect 17547 3800 17589 3809
rect 17547 3760 17548 3800
rect 17588 3760 17589 3800
rect 17547 3751 17589 3760
rect 17548 3632 17588 3751
rect 17548 3583 17588 3592
rect 17740 3632 17780 3835
rect 17836 3834 17876 3919
rect 17932 3725 17972 4096
rect 18028 3809 18068 4264
rect 18124 4136 18164 6196
rect 18220 6187 18260 6196
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18796 5648 18836 6280
rect 18892 5909 18932 6364
rect 18891 5900 18933 5909
rect 18891 5860 18892 5900
rect 18932 5860 18933 5900
rect 18891 5851 18933 5860
rect 18988 5825 19028 6952
rect 19179 6952 19180 6992
rect 19220 6952 19221 6992
rect 19179 6943 19221 6952
rect 19084 6497 19124 6582
rect 19083 6488 19125 6497
rect 19083 6448 19084 6488
rect 19124 6448 19125 6488
rect 19083 6439 19125 6448
rect 19084 6320 19124 6329
rect 19180 6320 19220 6943
rect 19275 6908 19317 6917
rect 19275 6868 19276 6908
rect 19316 6868 19412 6908
rect 19275 6859 19317 6868
rect 19124 6280 19220 6320
rect 19276 6488 19316 6497
rect 19084 6271 19124 6280
rect 19276 6068 19316 6448
rect 19372 6488 19412 6868
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 19467 6656 19509 6665
rect 19467 6616 19468 6656
rect 19508 6616 19509 6656
rect 19467 6607 19509 6616
rect 19755 6656 19797 6665
rect 19755 6616 19756 6656
rect 19796 6616 19797 6656
rect 19755 6607 19797 6616
rect 19372 6439 19412 6448
rect 19468 6488 19508 6607
rect 19468 6439 19508 6448
rect 19564 6488 19604 6497
rect 19564 6161 19604 6448
rect 19756 6488 19796 6607
rect 19756 6439 19796 6448
rect 19852 6488 19892 6499
rect 19852 6413 19892 6448
rect 19948 6488 19988 7708
rect 19851 6404 19893 6413
rect 19851 6364 19852 6404
rect 19892 6364 19893 6404
rect 19851 6355 19893 6364
rect 19563 6152 19605 6161
rect 19563 6112 19564 6152
rect 19604 6112 19605 6152
rect 19563 6103 19605 6112
rect 19755 6152 19797 6161
rect 19948 6152 19988 6448
rect 19755 6112 19756 6152
rect 19796 6112 19797 6152
rect 19755 6103 19797 6112
rect 19852 6112 19988 6152
rect 20044 6488 20084 6497
rect 19084 6028 19316 6068
rect 18987 5816 19029 5825
rect 18987 5776 18988 5816
rect 19028 5776 19029 5816
rect 18987 5767 19029 5776
rect 18796 5599 18836 5608
rect 18892 5648 18932 5657
rect 18700 5564 18740 5573
rect 18507 5480 18549 5489
rect 18507 5440 18508 5480
rect 18548 5440 18549 5480
rect 18507 5431 18549 5440
rect 18604 5480 18644 5489
rect 18508 5346 18548 5431
rect 18604 5237 18644 5440
rect 18603 5228 18645 5237
rect 18603 5188 18604 5228
rect 18644 5188 18645 5228
rect 18603 5179 18645 5188
rect 18700 4892 18740 5524
rect 18892 5489 18932 5608
rect 18891 5480 18933 5489
rect 18891 5440 18892 5480
rect 18932 5440 18933 5480
rect 18891 5431 18933 5440
rect 19084 5405 19124 6028
rect 19179 5900 19221 5909
rect 19179 5860 19180 5900
rect 19220 5860 19221 5900
rect 19179 5851 19221 5860
rect 19180 5564 19220 5851
rect 19275 5816 19317 5825
rect 19275 5776 19276 5816
rect 19316 5776 19317 5816
rect 19275 5767 19317 5776
rect 19083 5396 19125 5405
rect 19083 5356 19084 5396
rect 19124 5356 19125 5396
rect 19083 5347 19125 5356
rect 19180 5228 19220 5524
rect 18892 5188 19220 5228
rect 18892 5069 18932 5188
rect 19276 5144 19316 5767
rect 19660 5657 19700 5742
rect 19372 5648 19412 5657
rect 19372 5480 19412 5608
rect 19659 5648 19701 5657
rect 19756 5648 19796 6103
rect 19852 5825 19892 6112
rect 19947 5984 19989 5993
rect 19947 5944 19948 5984
rect 19988 5944 19989 5984
rect 19947 5935 19989 5944
rect 19851 5816 19893 5825
rect 19851 5776 19852 5816
rect 19892 5776 19893 5816
rect 19851 5767 19893 5776
rect 19659 5608 19660 5648
rect 19700 5608 19796 5648
rect 19948 5648 19988 5935
rect 20044 5825 20084 6448
rect 20043 5816 20085 5825
rect 20043 5776 20044 5816
rect 20084 5776 20085 5816
rect 20043 5767 20085 5776
rect 20140 5648 20180 5657
rect 19659 5599 19701 5608
rect 19948 5599 19988 5608
rect 20044 5608 20140 5648
rect 20044 5480 20084 5608
rect 20140 5580 20180 5608
rect 19372 5440 20084 5480
rect 19371 5312 19413 5321
rect 19371 5272 19372 5312
rect 19412 5272 19413 5312
rect 19371 5263 19413 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 19180 5104 19316 5144
rect 19372 5144 19412 5263
rect 19372 5104 19508 5144
rect 18891 5060 18933 5069
rect 18891 5020 18892 5060
rect 18932 5020 18933 5060
rect 18891 5011 18933 5020
rect 18700 4852 18836 4892
rect 18699 4724 18741 4733
rect 18699 4684 18700 4724
rect 18740 4684 18741 4724
rect 18699 4675 18741 4684
rect 18700 4590 18740 4675
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 18507 4388 18549 4397
rect 18796 4388 18836 4852
rect 18507 4348 18508 4388
rect 18548 4348 18549 4388
rect 18507 4339 18549 4348
rect 18604 4348 18836 4388
rect 18219 4220 18261 4229
rect 18316 4220 18356 4229
rect 18219 4180 18220 4220
rect 18260 4180 18316 4220
rect 18219 4171 18261 4180
rect 18316 4171 18356 4180
rect 18411 4220 18453 4229
rect 18411 4180 18412 4220
rect 18452 4180 18453 4220
rect 18411 4171 18453 4180
rect 18124 4087 18164 4096
rect 18412 4136 18452 4171
rect 18412 4085 18452 4096
rect 18508 3977 18548 4339
rect 18604 4136 18644 4348
rect 18892 4304 18932 5011
rect 19084 4976 19124 4985
rect 18987 4892 19029 4901
rect 18987 4852 18988 4892
rect 19028 4852 19029 4892
rect 18987 4843 19029 4852
rect 18796 4264 18932 4304
rect 18604 4087 18644 4096
rect 18700 4136 18740 4147
rect 18700 4061 18740 4096
rect 18796 4136 18836 4264
rect 18796 4087 18836 4096
rect 18892 4136 18932 4145
rect 18988 4136 19028 4843
rect 19084 4229 19124 4936
rect 19180 4976 19220 5104
rect 19083 4220 19125 4229
rect 19083 4180 19084 4220
rect 19124 4180 19125 4220
rect 19083 4171 19125 4180
rect 18932 4096 19028 4136
rect 18699 4052 18741 4061
rect 18699 4012 18700 4052
rect 18740 4012 18741 4052
rect 18699 4003 18741 4012
rect 18507 3968 18549 3977
rect 18507 3928 18508 3968
rect 18548 3928 18549 3968
rect 18507 3919 18549 3928
rect 18892 3893 18932 4096
rect 18891 3884 18933 3893
rect 18891 3844 18892 3884
rect 18932 3844 18933 3884
rect 18891 3835 18933 3844
rect 18027 3800 18069 3809
rect 18027 3760 18028 3800
rect 18068 3760 18069 3800
rect 18027 3751 18069 3760
rect 17931 3716 17973 3725
rect 17931 3676 17932 3716
rect 17972 3676 17973 3716
rect 17931 3667 17973 3676
rect 18123 3716 18165 3725
rect 18123 3676 18124 3716
rect 18164 3676 18165 3716
rect 18123 3667 18165 3676
rect 17740 3583 17780 3592
rect 17835 3548 17877 3557
rect 17835 3508 17836 3548
rect 17876 3508 17877 3548
rect 17835 3499 17877 3508
rect 18027 3548 18069 3557
rect 18027 3508 18028 3548
rect 18068 3508 18069 3548
rect 18027 3499 18069 3508
rect 17452 3415 17492 3424
rect 17836 3464 17876 3499
rect 17836 3413 17876 3424
rect 17932 3464 17972 3473
rect 17739 3044 17781 3053
rect 17739 3004 17740 3044
rect 17780 3004 17781 3044
rect 17739 2995 17781 3004
rect 17451 2792 17493 2801
rect 17451 2752 17452 2792
rect 17492 2752 17493 2792
rect 17451 2743 17493 2752
rect 16875 2624 16917 2633
rect 16875 2584 16876 2624
rect 16916 2584 16917 2624
rect 16875 2575 16917 2584
rect 16972 2624 17012 2633
rect 16683 2288 16725 2297
rect 16683 2248 16684 2288
rect 16724 2248 16725 2288
rect 16683 2239 16725 2248
rect 16491 2204 16533 2213
rect 16972 2204 17012 2584
rect 17068 2624 17108 2635
rect 17164 2633 17204 2719
rect 17259 2708 17301 2717
rect 17259 2668 17260 2708
rect 17300 2668 17301 2708
rect 17259 2659 17301 2668
rect 17068 2549 17108 2584
rect 17163 2626 17205 2633
rect 17163 2584 17164 2626
rect 17204 2584 17205 2626
rect 17163 2575 17205 2584
rect 17067 2540 17109 2549
rect 17067 2500 17068 2540
rect 17108 2500 17109 2540
rect 17067 2491 17109 2500
rect 17163 2456 17205 2465
rect 17163 2416 17164 2456
rect 17204 2416 17205 2456
rect 17163 2407 17205 2416
rect 16491 2164 16492 2204
rect 16532 2164 16533 2204
rect 16491 2155 16533 2164
rect 16780 2164 17012 2204
rect 16011 2120 16053 2129
rect 16011 2080 16012 2120
rect 16052 2080 16053 2120
rect 16011 2071 16053 2080
rect 16491 2036 16533 2045
rect 16491 1996 16492 2036
rect 16532 1996 16533 2036
rect 16491 1987 16533 1996
rect 16300 1952 16340 1961
rect 15916 1912 16300 1952
rect 16300 1903 16340 1912
rect 16492 1952 16532 1987
rect 16492 1901 16532 1912
rect 16780 1709 16820 2164
rect 16875 2036 16917 2045
rect 17067 2036 17109 2045
rect 16875 1996 16876 2036
rect 16916 1996 16917 2036
rect 16875 1987 16917 1996
rect 16972 1996 17068 2036
rect 17108 1996 17109 2036
rect 16876 1952 16916 1987
rect 16972 1962 17012 1996
rect 17067 1987 17109 1996
rect 16972 1913 17012 1922
rect 16876 1901 16916 1912
rect 17164 1784 17204 2407
rect 17260 2045 17300 2659
rect 17356 2624 17396 2633
rect 17356 2549 17396 2584
rect 17355 2540 17397 2549
rect 17452 2540 17492 2743
rect 17355 2500 17356 2540
rect 17396 2500 17397 2540
rect 17355 2491 17397 2500
rect 17449 2500 17492 2540
rect 17548 2624 17588 2633
rect 17356 2460 17396 2491
rect 17449 2372 17489 2500
rect 17548 2465 17588 2584
rect 17643 2624 17685 2633
rect 17643 2584 17644 2624
rect 17684 2584 17685 2624
rect 17643 2575 17685 2584
rect 17547 2456 17589 2465
rect 17547 2416 17548 2456
rect 17588 2416 17589 2456
rect 17547 2407 17589 2416
rect 17449 2332 17492 2372
rect 17355 2204 17397 2213
rect 17355 2164 17356 2204
rect 17396 2164 17397 2204
rect 17355 2155 17397 2164
rect 17259 2036 17301 2045
rect 17259 1996 17260 2036
rect 17300 1996 17301 2036
rect 17259 1987 17301 1996
rect 17164 1735 17204 1744
rect 16491 1700 16533 1709
rect 16491 1660 16492 1700
rect 16532 1660 16533 1700
rect 16491 1651 16533 1660
rect 16779 1700 16821 1709
rect 16779 1660 16780 1700
rect 16820 1660 16821 1700
rect 16779 1651 16821 1660
rect 16492 1566 16532 1651
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 17356 1196 17396 2155
rect 17452 2120 17492 2332
rect 17547 2288 17589 2297
rect 17547 2248 17548 2288
rect 17588 2248 17589 2288
rect 17547 2239 17589 2248
rect 17452 2071 17492 2080
rect 17548 1952 17588 2239
rect 17548 1903 17588 1912
rect 17644 1952 17684 2575
rect 17644 1903 17684 1912
rect 17740 1952 17780 2995
rect 17932 2885 17972 3424
rect 18028 3464 18068 3499
rect 18028 3053 18068 3424
rect 18027 3044 18069 3053
rect 18027 3004 18028 3044
rect 18068 3004 18069 3044
rect 18027 2995 18069 3004
rect 17931 2876 17973 2885
rect 17931 2836 17932 2876
rect 17972 2836 17973 2876
rect 18124 2876 18164 3667
rect 19180 3389 19220 4936
rect 19275 4976 19317 4985
rect 19275 4936 19276 4976
rect 19316 4936 19317 4976
rect 19275 4927 19317 4936
rect 19372 4976 19412 4985
rect 19276 4842 19316 4927
rect 19372 4817 19412 4936
rect 19371 4808 19413 4817
rect 19371 4768 19372 4808
rect 19412 4768 19413 4808
rect 19371 4759 19413 4768
rect 19372 4136 19412 4145
rect 19468 4136 19508 5104
rect 20044 4976 20084 5440
rect 20044 4229 20084 4936
rect 20236 4976 20276 4985
rect 20139 4892 20181 4901
rect 20139 4852 20140 4892
rect 20180 4852 20181 4892
rect 20139 4843 20181 4852
rect 20140 4758 20180 4843
rect 20236 4481 20276 4936
rect 20235 4472 20277 4481
rect 20235 4432 20236 4472
rect 20276 4432 20277 4472
rect 20235 4423 20277 4432
rect 20332 4313 20372 7960
rect 20427 8000 20469 8009
rect 20427 7960 20428 8000
rect 20468 7960 20469 8000
rect 20427 7951 20469 7960
rect 20427 7832 20469 7841
rect 20427 7792 20428 7832
rect 20468 7792 20469 7832
rect 20427 7783 20469 7792
rect 20428 7698 20468 7783
rect 20524 7673 20564 8716
rect 20620 8672 20660 9472
rect 20716 8933 20756 9472
rect 20811 9512 20853 9521
rect 21004 9512 21044 9521
rect 20811 9472 20812 9512
rect 20852 9472 20853 9512
rect 20811 9463 20853 9472
rect 20908 9472 21004 9512
rect 20811 9344 20853 9353
rect 20811 9304 20812 9344
rect 20852 9304 20853 9344
rect 20811 9295 20853 9304
rect 20715 8924 20757 8933
rect 20715 8884 20716 8924
rect 20756 8884 20757 8924
rect 20715 8875 20757 8884
rect 20620 8597 20660 8632
rect 20619 8588 20661 8597
rect 20619 8548 20620 8588
rect 20660 8548 20661 8588
rect 20619 8539 20661 8548
rect 20620 8429 20660 8539
rect 20619 8420 20661 8429
rect 20619 8380 20620 8420
rect 20660 8380 20661 8420
rect 20619 8371 20661 8380
rect 20812 8168 20852 9295
rect 20908 8849 20948 9472
rect 21004 9463 21044 9472
rect 21004 9260 21044 9269
rect 21044 9220 21236 9260
rect 21004 9211 21044 9220
rect 21003 9092 21045 9101
rect 21003 9052 21004 9092
rect 21044 9052 21045 9092
rect 21003 9043 21045 9052
rect 20907 8840 20949 8849
rect 20907 8800 20908 8840
rect 20948 8800 20949 8840
rect 20907 8791 20949 8800
rect 20908 8672 20948 8681
rect 20908 8513 20948 8632
rect 21004 8672 21044 9043
rect 21004 8623 21044 8632
rect 21100 8672 21140 8681
rect 21196 8672 21236 9220
rect 21292 9101 21332 11227
rect 21388 9437 21428 11488
rect 21484 11453 21524 11656
rect 21641 11645 21681 11671
rect 22636 11621 22676 12496
rect 22635 11612 22677 11621
rect 22635 11572 22636 11612
rect 22676 11572 22677 11612
rect 22635 11563 22677 11572
rect 21483 11444 21525 11453
rect 21483 11404 21484 11444
rect 21524 11404 21525 11444
rect 21483 11395 21525 11404
rect 22732 11360 22772 13168
rect 22636 11320 22772 11360
rect 22347 10940 22389 10949
rect 22347 10900 22348 10940
rect 22388 10900 22389 10940
rect 22347 10891 22389 10900
rect 21579 10352 21621 10361
rect 21579 10312 21580 10352
rect 21620 10312 21621 10352
rect 21579 10303 21621 10312
rect 22155 10352 22197 10361
rect 22155 10312 22156 10352
rect 22196 10312 22197 10352
rect 22155 10303 22197 10312
rect 21387 9428 21429 9437
rect 21387 9388 21388 9428
rect 21428 9388 21429 9428
rect 21387 9379 21429 9388
rect 21291 9092 21333 9101
rect 21291 9052 21292 9092
rect 21332 9052 21333 9092
rect 21291 9043 21333 9052
rect 21388 8672 21428 8681
rect 21196 8632 21388 8672
rect 21100 8513 21140 8632
rect 21388 8623 21428 8632
rect 21483 8672 21525 8681
rect 21483 8632 21484 8672
rect 21524 8632 21525 8672
rect 21483 8623 21525 8632
rect 21580 8672 21620 10303
rect 22059 10268 22101 10277
rect 22059 10228 22060 10268
rect 22100 10228 22101 10268
rect 22059 10219 22101 10228
rect 21867 10184 21909 10193
rect 21867 10144 21868 10184
rect 21908 10144 21909 10184
rect 21867 10135 21909 10144
rect 22060 10184 22100 10219
rect 21868 10050 21908 10135
rect 22060 10133 22100 10144
rect 22156 10184 22196 10303
rect 22156 10135 22196 10144
rect 22251 10184 22293 10193
rect 22251 10144 22252 10184
rect 22292 10144 22293 10184
rect 22251 10135 22293 10144
rect 22348 10184 22388 10891
rect 22636 10445 22676 11320
rect 22635 10436 22677 10445
rect 22635 10396 22636 10436
rect 22676 10396 22677 10436
rect 22635 10387 22677 10396
rect 22348 10135 22388 10144
rect 22252 10050 22292 10135
rect 21964 9689 22004 9774
rect 21963 9680 22005 9689
rect 21963 9640 21964 9680
rect 22004 9640 22005 9680
rect 21963 9631 22005 9640
rect 21964 9512 22004 9521
rect 21868 9428 21908 9437
rect 21580 8623 21620 8632
rect 21772 9344 21812 9353
rect 21484 8538 21524 8623
rect 21676 8588 21716 8597
rect 21772 8588 21812 9304
rect 21868 9092 21908 9388
rect 21964 9353 22004 9472
rect 22060 9512 22100 9521
rect 22444 9512 22484 9521
rect 22100 9472 22292 9512
rect 22060 9463 22100 9472
rect 21963 9344 22005 9353
rect 21963 9304 21964 9344
rect 22004 9304 22005 9344
rect 21963 9295 22005 9304
rect 22252 9344 22292 9472
rect 22252 9295 22292 9304
rect 21868 9052 22196 9092
rect 21963 8924 22005 8933
rect 21963 8884 21964 8924
rect 22004 8884 22005 8924
rect 21963 8875 22005 8884
rect 21964 8840 22004 8875
rect 21964 8789 22004 8800
rect 21867 8756 21909 8765
rect 21867 8716 21868 8756
rect 21908 8716 21909 8756
rect 21867 8707 21909 8716
rect 21868 8672 21908 8707
rect 21868 8621 21908 8632
rect 22060 8672 22100 8681
rect 21716 8548 21812 8588
rect 21676 8539 21716 8548
rect 20907 8504 20949 8513
rect 20907 8464 20908 8504
rect 20948 8464 20949 8504
rect 20907 8455 20949 8464
rect 21099 8504 21141 8513
rect 21099 8464 21100 8504
rect 21140 8464 21141 8504
rect 21099 8455 21141 8464
rect 21196 8504 21236 8513
rect 21579 8504 21621 8513
rect 21236 8464 21428 8504
rect 21196 8455 21236 8464
rect 21196 8177 21236 8262
rect 21195 8168 21237 8177
rect 20812 8128 20948 8168
rect 20716 8000 20756 8009
rect 20619 7916 20661 7925
rect 20716 7916 20756 7960
rect 20812 8000 20852 8011
rect 20812 7925 20852 7960
rect 20619 7876 20620 7916
rect 20660 7876 20756 7916
rect 20811 7916 20853 7925
rect 20811 7876 20812 7916
rect 20852 7876 20853 7916
rect 20619 7867 20661 7876
rect 20811 7867 20853 7876
rect 20523 7664 20565 7673
rect 20523 7624 20524 7664
rect 20564 7624 20565 7664
rect 20523 7615 20565 7624
rect 20427 7412 20469 7421
rect 20427 7372 20428 7412
rect 20468 7372 20469 7412
rect 20427 7363 20469 7372
rect 20428 7160 20468 7363
rect 20524 7169 20564 7615
rect 20908 7496 20948 8128
rect 21195 8128 21196 8168
rect 21236 8128 21237 8168
rect 21195 8119 21237 8128
rect 21099 8084 21141 8093
rect 21099 8044 21100 8084
rect 21140 8044 21141 8084
rect 21099 8035 21141 8044
rect 21004 8000 21044 8009
rect 21004 7841 21044 7960
rect 21100 8000 21140 8035
rect 21100 7949 21140 7960
rect 21257 7985 21297 7994
rect 21003 7832 21045 7841
rect 21003 7792 21004 7832
rect 21044 7792 21045 7832
rect 21003 7783 21045 7792
rect 21257 7580 21297 7945
rect 21388 7748 21428 8464
rect 21579 8464 21580 8504
rect 21620 8464 21621 8504
rect 21579 8455 21621 8464
rect 21580 8084 21620 8455
rect 22060 8345 22100 8632
rect 22059 8336 22101 8345
rect 22059 8296 22060 8336
rect 22100 8296 22101 8336
rect 22059 8287 22101 8296
rect 21675 8168 21717 8177
rect 21675 8128 21676 8168
rect 21716 8128 21717 8168
rect 21675 8119 21717 8128
rect 21580 8035 21620 8044
rect 21483 8000 21525 8009
rect 21483 7960 21484 8000
rect 21524 7960 21525 8000
rect 21483 7951 21525 7960
rect 21676 8000 21716 8119
rect 21676 7951 21716 7960
rect 21484 7866 21524 7951
rect 21388 7708 21620 7748
rect 21257 7540 21428 7580
rect 20908 7456 21332 7496
rect 21196 7328 21236 7337
rect 20716 7288 21196 7328
rect 20428 7111 20468 7120
rect 20523 7160 20565 7169
rect 20523 7120 20524 7160
rect 20564 7120 20565 7160
rect 20523 7111 20565 7120
rect 20620 7160 20660 7171
rect 20620 7085 20660 7120
rect 20619 7076 20661 7085
rect 20619 7036 20620 7076
rect 20660 7036 20661 7076
rect 20619 7027 20661 7036
rect 20524 6992 20564 7001
rect 20524 6497 20564 6952
rect 20523 6488 20565 6497
rect 20523 6448 20524 6488
rect 20564 6448 20565 6488
rect 20523 6439 20565 6448
rect 20716 5648 20756 7288
rect 21196 7279 21236 7288
rect 20811 7160 20853 7169
rect 20811 7120 20812 7160
rect 20852 7120 20853 7160
rect 20811 7111 20853 7120
rect 21004 7160 21044 7171
rect 20812 6161 20852 7111
rect 21004 7085 21044 7120
rect 21003 7076 21045 7085
rect 21003 7036 21004 7076
rect 21044 7036 21045 7076
rect 21003 7027 21045 7036
rect 20811 6152 20853 6161
rect 20811 6112 20812 6152
rect 20852 6112 20853 6152
rect 20811 6103 20853 6112
rect 20716 5599 20756 5608
rect 20812 5648 20852 5657
rect 21292 5648 21332 7456
rect 21388 7085 21428 7540
rect 21484 7160 21524 7169
rect 21387 7076 21429 7085
rect 21387 7036 21388 7076
rect 21428 7036 21429 7076
rect 21387 7027 21429 7036
rect 21484 6992 21524 7120
rect 21580 7160 21620 7708
rect 22060 7589 22100 8287
rect 22156 7673 22196 9052
rect 22444 8849 22484 9472
rect 22539 9512 22581 9521
rect 22539 9472 22540 9512
rect 22580 9472 22581 9512
rect 22539 9463 22581 9472
rect 22636 9512 22676 10387
rect 22732 10184 22772 10193
rect 22732 9689 22772 10144
rect 22731 9680 22773 9689
rect 22731 9640 22732 9680
rect 22772 9640 22773 9680
rect 22731 9631 22773 9640
rect 22636 9463 22676 9472
rect 22732 9512 22772 9521
rect 22540 9378 22580 9463
rect 22732 9101 22772 9472
rect 22828 9185 22868 16696
rect 22923 16687 22965 16696
rect 23884 16400 23924 17107
rect 23788 16360 23924 16400
rect 23019 16232 23061 16241
rect 23019 16192 23020 16232
rect 23060 16192 23061 16232
rect 23019 16183 23061 16192
rect 22923 15056 22965 15065
rect 22923 15016 22924 15056
rect 22964 15016 22965 15056
rect 22923 15007 22965 15016
rect 22924 14561 22964 15007
rect 22923 14552 22965 14561
rect 22923 14512 22924 14552
rect 22964 14512 22965 14552
rect 22923 14503 22965 14512
rect 22923 14132 22965 14141
rect 22923 14092 22924 14132
rect 22964 14092 22965 14132
rect 22923 14083 22965 14092
rect 22924 13998 22964 14083
rect 23020 13217 23060 16183
rect 23788 15476 23828 16360
rect 23883 16232 23925 16241
rect 23883 16192 23884 16232
rect 23924 16192 23925 16232
rect 23883 16183 23925 16192
rect 24076 16232 24116 18964
rect 24267 18836 24309 18845
rect 24267 18796 24268 18836
rect 24308 18796 24309 18836
rect 24267 18787 24309 18796
rect 24171 18584 24213 18593
rect 24171 18544 24172 18584
rect 24212 18544 24213 18584
rect 24171 18535 24213 18544
rect 24172 17753 24212 18535
rect 24171 17744 24213 17753
rect 24171 17704 24172 17744
rect 24212 17704 24213 17744
rect 24171 17695 24213 17704
rect 24268 17744 24308 18787
rect 24364 18584 24404 18964
rect 24459 18836 24501 18845
rect 24459 18796 24460 18836
rect 24500 18796 24501 18836
rect 24459 18787 24501 18796
rect 24843 18836 24885 18845
rect 24843 18796 24844 18836
rect 24884 18796 24885 18836
rect 24843 18787 24885 18796
rect 24364 18535 24404 18544
rect 24460 18584 24500 18787
rect 24460 18535 24500 18544
rect 24651 18584 24693 18593
rect 24651 18544 24652 18584
rect 24692 18544 24693 18584
rect 24651 18535 24693 18544
rect 24844 18584 24884 18787
rect 24844 18535 24884 18544
rect 24652 18450 24692 18535
rect 24748 18500 24788 18509
rect 24459 18416 24501 18425
rect 24459 18376 24460 18416
rect 24500 18376 24501 18416
rect 24459 18367 24501 18376
rect 24460 18282 24500 18367
rect 24748 17996 24788 18460
rect 24652 17956 24788 17996
rect 24172 17576 24212 17695
rect 24172 17527 24212 17536
rect 24268 17072 24308 17704
rect 24363 17744 24405 17753
rect 24363 17704 24364 17744
rect 24404 17704 24405 17744
rect 24363 17695 24405 17704
rect 24652 17744 24692 17956
rect 24843 17912 24885 17921
rect 24843 17872 24844 17912
rect 24884 17872 24885 17912
rect 24843 17863 24885 17872
rect 24652 17695 24692 17704
rect 24748 17828 24788 17837
rect 24268 17023 24308 17032
rect 24364 16988 24404 17695
rect 24460 17660 24500 17669
rect 24460 17408 24500 17620
rect 24748 17408 24788 17788
rect 24844 17778 24884 17863
rect 24940 17828 24980 17837
rect 24460 17368 24788 17408
rect 24460 16988 24500 16997
rect 24364 16948 24460 16988
rect 24460 16939 24500 16948
rect 23884 16098 23924 16183
rect 23980 16064 24020 16073
rect 23884 15476 23924 15485
rect 23788 15436 23884 15476
rect 23884 15427 23924 15436
rect 23691 15308 23733 15317
rect 23691 15268 23692 15308
rect 23732 15268 23733 15308
rect 23691 15259 23733 15268
rect 23692 15140 23732 15259
rect 23404 15100 23732 15140
rect 23115 14804 23157 14813
rect 23115 14764 23116 14804
rect 23156 14764 23157 14804
rect 23115 14755 23157 14764
rect 23116 14216 23156 14755
rect 23116 13460 23156 14176
rect 23308 13460 23348 13469
rect 23116 13420 23308 13460
rect 23308 13411 23348 13420
rect 23019 13208 23061 13217
rect 23019 13168 23020 13208
rect 23060 13168 23061 13208
rect 23019 13159 23061 13168
rect 23307 13208 23349 13217
rect 23307 13168 23308 13208
rect 23348 13168 23349 13208
rect 23404 13208 23444 15100
rect 23980 15065 24020 16024
rect 24076 15140 24116 16192
rect 24268 16820 24308 16829
rect 24268 15569 24308 16780
rect 24652 16745 24692 17368
rect 24747 17240 24789 17249
rect 24747 17200 24748 17240
rect 24788 17200 24789 17240
rect 24747 17191 24789 17200
rect 24844 17240 24884 17249
rect 24940 17240 24980 17788
rect 25036 17744 25076 19207
rect 25228 19122 25268 19207
rect 25324 19205 25364 19216
rect 25420 19256 25460 19265
rect 25516 19256 25556 20047
rect 25612 20045 25652 20056
rect 25708 19517 25748 19602
rect 25707 19508 25749 19517
rect 25707 19468 25708 19508
rect 25748 19468 25749 19508
rect 25707 19459 25749 19468
rect 25708 19256 25748 19265
rect 25516 19216 25708 19256
rect 25420 17996 25460 19216
rect 25708 19207 25748 19216
rect 25900 19256 25940 20140
rect 25996 20096 26036 20105
rect 25996 19937 26036 20056
rect 25995 19928 26037 19937
rect 25995 19888 25996 19928
rect 26036 19888 26037 19928
rect 25995 19879 26037 19888
rect 25995 19340 26037 19349
rect 25995 19300 25996 19340
rect 26036 19300 26037 19340
rect 25995 19291 26037 19300
rect 25900 19207 25940 19216
rect 25996 19256 26036 19291
rect 25996 19205 26036 19216
rect 25516 19088 25556 19097
rect 25516 18920 25556 19048
rect 26092 18920 26132 20728
rect 26188 20684 26228 21568
rect 26380 21559 26420 21568
rect 26571 21608 26613 21617
rect 26571 21568 26572 21608
rect 26612 21568 26613 21608
rect 26571 21559 26613 21568
rect 26572 21474 26612 21559
rect 26188 20635 26228 20644
rect 26476 20768 26516 20777
rect 26187 20012 26229 20021
rect 26187 19972 26188 20012
rect 26228 19972 26229 20012
rect 26187 19963 26229 19972
rect 26188 19265 26228 19963
rect 26476 19349 26516 20728
rect 26571 20096 26613 20105
rect 26571 20056 26572 20096
rect 26612 20056 26613 20096
rect 26571 20047 26613 20056
rect 26572 19962 26612 20047
rect 26859 19844 26901 19853
rect 26859 19804 26860 19844
rect 26900 19804 26901 19844
rect 26859 19795 26901 19804
rect 26860 19710 26900 19795
rect 26475 19340 26517 19349
rect 26475 19300 26476 19340
rect 26516 19300 26517 19340
rect 26475 19291 26517 19300
rect 26187 19256 26229 19265
rect 26187 19216 26188 19256
rect 26228 19216 26229 19256
rect 26187 19207 26229 19216
rect 26956 19256 26996 24088
rect 27339 23708 27381 23717
rect 27339 23668 27340 23708
rect 27380 23668 27381 23708
rect 27339 23659 27381 23668
rect 27340 23574 27380 23659
rect 27051 23120 27093 23129
rect 27051 23080 27052 23120
rect 27092 23080 27093 23120
rect 27051 23071 27093 23080
rect 27052 22709 27092 23071
rect 27051 22700 27093 22709
rect 27051 22660 27052 22700
rect 27092 22660 27093 22700
rect 27051 22651 27093 22660
rect 27244 22448 27284 22457
rect 27148 21608 27188 21617
rect 27244 21608 27284 22408
rect 27188 21568 27284 21608
rect 28012 21608 28052 25516
rect 28108 24893 28148 26515
rect 28492 26321 28532 26781
rect 28587 26648 28629 26657
rect 28587 26608 28588 26648
rect 28628 26608 28629 26648
rect 28587 26599 28629 26608
rect 28684 26648 28724 26657
rect 28491 26312 28533 26321
rect 28491 26272 28492 26312
rect 28532 26272 28533 26312
rect 28491 26263 28533 26272
rect 28491 26144 28533 26153
rect 28491 26104 28492 26144
rect 28532 26104 28533 26144
rect 28491 26095 28533 26104
rect 28588 26139 28628 26599
rect 28684 26489 28724 26608
rect 28683 26480 28725 26489
rect 28683 26440 28684 26480
rect 28724 26440 28725 26480
rect 28683 26431 28725 26440
rect 28492 26010 28532 26095
rect 28588 26090 28628 26099
rect 28684 26144 28724 26153
rect 28780 26144 28820 26851
rect 28876 26816 28916 26935
rect 28971 26900 29013 26909
rect 28971 26860 28972 26900
rect 29012 26860 29013 26900
rect 28971 26851 29013 26860
rect 28876 26573 28916 26776
rect 28972 26732 29012 26851
rect 28972 26683 29012 26692
rect 29068 26816 29108 26825
rect 29068 26573 29108 26776
rect 29164 26816 29204 26825
rect 28875 26564 28917 26573
rect 28875 26524 28876 26564
rect 28916 26524 28917 26564
rect 28875 26515 28917 26524
rect 29067 26564 29109 26573
rect 29067 26524 29068 26564
rect 29108 26524 29109 26564
rect 29067 26515 29109 26524
rect 29164 26312 29204 26776
rect 29260 26321 29300 27523
rect 29643 27404 29685 27413
rect 29643 27364 29644 27404
rect 29684 27364 29685 27404
rect 29643 27355 29685 27364
rect 29547 26816 29589 26825
rect 29547 26776 29548 26816
rect 29588 26776 29589 26816
rect 29547 26767 29589 26776
rect 29644 26816 29684 27355
rect 29835 27068 29877 27077
rect 29835 27028 29836 27068
rect 29876 27028 29877 27068
rect 29835 27019 29877 27028
rect 29644 26767 29684 26776
rect 29548 26682 29588 26767
rect 29355 26648 29397 26657
rect 29355 26608 29356 26648
rect 29396 26608 29397 26648
rect 29836 26648 29876 27019
rect 29932 26816 29972 28867
rect 30219 28412 30261 28421
rect 30219 28372 30220 28412
rect 30260 28372 30261 28412
rect 30219 28363 30261 28372
rect 30220 28278 30260 28363
rect 30027 27656 30069 27665
rect 30027 27616 30028 27656
rect 30068 27616 30069 27656
rect 30027 27607 30069 27616
rect 30124 27656 30164 27665
rect 30028 27522 30068 27607
rect 30124 27077 30164 27616
rect 30220 27656 30260 27667
rect 30220 27581 30260 27616
rect 30316 27656 30356 30808
rect 30892 30437 30932 30522
rect 30411 30428 30453 30437
rect 30411 30388 30412 30428
rect 30452 30388 30453 30428
rect 30411 30379 30453 30388
rect 30700 30428 30740 30437
rect 30891 30428 30933 30437
rect 30740 30388 30836 30428
rect 30700 30379 30740 30388
rect 30412 29597 30452 30379
rect 30700 29840 30740 29849
rect 30508 29800 30700 29840
rect 30411 29588 30453 29597
rect 30411 29548 30412 29588
rect 30452 29548 30453 29588
rect 30411 29539 30453 29548
rect 30412 29168 30452 29179
rect 30412 29093 30452 29128
rect 30411 29084 30453 29093
rect 30411 29044 30412 29084
rect 30452 29044 30453 29084
rect 30411 29035 30453 29044
rect 30508 27824 30548 29800
rect 30700 29791 30740 29800
rect 30699 29000 30741 29009
rect 30699 28960 30700 29000
rect 30740 28960 30741 29000
rect 30699 28951 30741 28960
rect 30700 28866 30740 28951
rect 30796 28673 30836 30388
rect 30891 30388 30892 30428
rect 30932 30388 30933 30428
rect 30891 30379 30933 30388
rect 30988 30260 31028 33823
rect 31083 33704 31125 33713
rect 31083 33664 31084 33704
rect 31124 33664 31125 33704
rect 31083 33655 31125 33664
rect 31180 33704 31220 33713
rect 31084 33570 31124 33655
rect 31180 33125 31220 33664
rect 31276 33704 31316 34579
rect 31660 34494 31700 34579
rect 32620 34376 32660 34385
rect 32716 34376 32756 35008
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 35500 34544 35540 34553
rect 37996 34544 38036 34553
rect 35540 34504 35828 34544
rect 35500 34495 35540 34504
rect 32660 34336 32756 34376
rect 33483 34376 33525 34385
rect 33483 34336 33484 34376
rect 33524 34336 33525 34376
rect 32620 34327 32660 34336
rect 33483 34327 33525 34336
rect 33771 34376 33813 34385
rect 33771 34336 33772 34376
rect 33812 34336 33813 34376
rect 33771 34327 33813 34336
rect 34155 34376 34197 34385
rect 34155 34336 34156 34376
rect 34196 34336 34197 34376
rect 34155 34327 34197 34336
rect 32236 34292 32276 34301
rect 32043 33872 32085 33881
rect 32043 33832 32044 33872
rect 32084 33832 32085 33872
rect 32043 33823 32085 33832
rect 32236 33872 32276 34252
rect 33484 34242 33524 34327
rect 32236 33823 32276 33832
rect 31276 33655 31316 33664
rect 31371 33704 31413 33713
rect 31371 33664 31372 33704
rect 31412 33664 31413 33704
rect 31371 33655 31413 33664
rect 31564 33704 31604 33713
rect 31372 33545 31412 33655
rect 31371 33536 31413 33545
rect 31371 33496 31372 33536
rect 31412 33496 31413 33536
rect 31371 33487 31413 33496
rect 31371 33368 31413 33377
rect 31371 33328 31372 33368
rect 31412 33328 31413 33368
rect 31371 33319 31413 33328
rect 31179 33116 31221 33125
rect 31179 33076 31180 33116
rect 31220 33076 31221 33116
rect 31179 33067 31221 33076
rect 31179 32948 31221 32957
rect 31179 32908 31180 32948
rect 31220 32908 31221 32948
rect 31179 32899 31221 32908
rect 31180 32696 31220 32899
rect 31180 32647 31220 32656
rect 30892 30220 31028 30260
rect 31084 32192 31124 32201
rect 30795 28664 30837 28673
rect 30795 28624 30796 28664
rect 30836 28624 30837 28664
rect 30795 28615 30837 28624
rect 30603 28580 30645 28589
rect 30603 28540 30604 28580
rect 30644 28540 30645 28580
rect 30603 28531 30645 28540
rect 30604 28446 30644 28531
rect 30892 28328 30932 30220
rect 31084 29933 31124 32152
rect 31372 32192 31412 33319
rect 31564 32696 31604 33664
rect 31660 33704 31700 33713
rect 31660 33125 31700 33664
rect 31756 33704 31796 33713
rect 31756 33200 31796 33664
rect 31852 33704 31892 33713
rect 32044 33704 32084 33823
rect 32140 33713 32180 33798
rect 31892 33664 31988 33704
rect 31852 33655 31892 33664
rect 31948 33536 31988 33664
rect 32044 33655 32084 33664
rect 32139 33704 32181 33713
rect 32139 33664 32140 33704
rect 32180 33664 32181 33704
rect 32139 33655 32181 33664
rect 32332 33704 32372 33713
rect 32524 33704 32564 33713
rect 32332 33536 32372 33664
rect 31948 33496 32372 33536
rect 32428 33664 32524 33704
rect 31756 33160 31892 33200
rect 31659 33116 31701 33125
rect 31659 33076 31660 33116
rect 31700 33076 31701 33116
rect 31659 33067 31701 33076
rect 31660 32873 31700 32958
rect 31659 32864 31701 32873
rect 31659 32824 31660 32864
rect 31700 32824 31701 32864
rect 31659 32815 31701 32824
rect 31756 32864 31796 32873
rect 31756 32696 31796 32824
rect 31564 32656 31796 32696
rect 31756 32369 31796 32656
rect 31755 32360 31797 32369
rect 31755 32320 31756 32360
rect 31796 32320 31797 32360
rect 31755 32311 31797 32320
rect 31467 32276 31509 32285
rect 31467 32236 31468 32276
rect 31508 32236 31509 32276
rect 31467 32227 31509 32236
rect 31372 32143 31412 32152
rect 31468 32142 31508 32227
rect 31852 32192 31892 33160
rect 31948 33116 31988 33125
rect 32428 33116 32468 33664
rect 32524 33655 32564 33664
rect 32619 33704 32661 33713
rect 32619 33664 32620 33704
rect 32660 33664 32661 33704
rect 32619 33655 32661 33664
rect 32908 33704 32948 33713
rect 33772 33704 33812 34327
rect 32948 33664 33044 33704
rect 32908 33655 32948 33664
rect 31988 33076 32468 33116
rect 31948 33067 31988 33076
rect 32043 32948 32085 32957
rect 32043 32908 32044 32948
rect 32084 32908 32180 32948
rect 32043 32899 32085 32908
rect 31948 32864 31988 32873
rect 31948 32360 31988 32824
rect 32140 32864 32180 32908
rect 32140 32815 32180 32824
rect 32620 32780 32660 33655
rect 33004 33032 33044 33664
rect 33772 33655 33812 33664
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 33771 33116 33813 33125
rect 33771 33076 33772 33116
rect 33812 33076 33813 33116
rect 33771 33067 33813 33076
rect 34156 33116 34196 34327
rect 34636 34208 34676 34217
rect 35692 34208 35732 34217
rect 34676 34168 35060 34208
rect 34636 34159 34676 34168
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 34924 33452 34964 33463
rect 34924 33377 34964 33412
rect 34923 33368 34965 33377
rect 34923 33328 34924 33368
rect 34964 33328 34965 33368
rect 34923 33319 34965 33328
rect 34156 33067 34196 33076
rect 34347 33116 34389 33125
rect 34347 33076 34348 33116
rect 34388 33076 34389 33116
rect 34347 33067 34389 33076
rect 33004 32983 33044 32992
rect 33675 33032 33717 33041
rect 33675 32992 33676 33032
rect 33716 32992 33717 33032
rect 33675 32983 33717 32992
rect 33291 32948 33333 32957
rect 33291 32908 33292 32948
rect 33332 32908 33333 32948
rect 33291 32899 33333 32908
rect 33484 32948 33524 32957
rect 33195 32864 33237 32873
rect 33195 32824 33196 32864
rect 33236 32824 33237 32864
rect 33195 32815 33237 32824
rect 32428 32740 32660 32780
rect 32139 32696 32181 32705
rect 32139 32656 32140 32696
rect 32180 32656 32181 32696
rect 32139 32647 32181 32656
rect 31948 32311 31988 32320
rect 32044 32192 32084 32201
rect 31852 32152 32044 32192
rect 31755 31940 31797 31949
rect 31755 31900 31756 31940
rect 31796 31900 31797 31940
rect 31755 31891 31797 31900
rect 31756 31806 31796 31891
rect 32044 31688 32084 32152
rect 32140 32192 32180 32647
rect 32235 32360 32277 32369
rect 32235 32320 32236 32360
rect 32276 32320 32277 32360
rect 32235 32311 32277 32320
rect 32428 32360 32468 32740
rect 32812 32696 32852 32705
rect 32852 32656 33140 32696
rect 32812 32647 32852 32656
rect 32428 32311 32468 32320
rect 32140 32143 32180 32152
rect 32236 32192 32276 32311
rect 32811 32192 32853 32201
rect 32276 32152 32468 32192
rect 32236 32143 32276 32152
rect 32044 31648 32372 31688
rect 32044 31445 32084 31648
rect 32235 31520 32277 31529
rect 32235 31480 32236 31520
rect 32276 31480 32277 31520
rect 32235 31471 32277 31480
rect 32043 31436 32085 31445
rect 32043 31396 32044 31436
rect 32084 31396 32085 31436
rect 32043 31387 32085 31396
rect 31660 31352 31700 31361
rect 31564 30680 31604 30689
rect 31083 29924 31125 29933
rect 31083 29884 31084 29924
rect 31124 29884 31125 29924
rect 31083 29875 31125 29884
rect 31467 29924 31509 29933
rect 31467 29884 31468 29924
rect 31508 29884 31509 29924
rect 31467 29875 31509 29884
rect 30987 29336 31029 29345
rect 30987 29296 30988 29336
rect 31028 29296 31029 29336
rect 30987 29287 31029 29296
rect 30988 29252 31028 29287
rect 30988 29201 31028 29212
rect 31083 29168 31125 29177
rect 31372 29168 31412 29177
rect 31083 29128 31084 29168
rect 31124 29128 31125 29168
rect 31083 29119 31125 29128
rect 31180 29128 31372 29168
rect 31084 29034 31124 29119
rect 31180 28664 31220 29128
rect 31372 29119 31412 29128
rect 30316 27607 30356 27616
rect 30412 27784 30548 27824
rect 30700 28288 30932 28328
rect 31084 28624 31220 28664
rect 30219 27572 30261 27581
rect 30219 27532 30220 27572
rect 30260 27532 30261 27572
rect 30219 27523 30261 27532
rect 30123 27068 30165 27077
rect 30123 27028 30124 27068
rect 30164 27028 30165 27068
rect 30123 27019 30165 27028
rect 30124 26900 30164 26909
rect 30164 26860 30260 26900
rect 30124 26851 30164 26860
rect 29932 26776 30068 26816
rect 29932 26648 29972 26657
rect 29836 26608 29932 26648
rect 29355 26599 29397 26608
rect 29932 26599 29972 26608
rect 29356 26514 29396 26599
rect 29164 26263 29204 26272
rect 29259 26312 29301 26321
rect 29259 26272 29260 26312
rect 29300 26272 29301 26312
rect 29259 26263 29301 26272
rect 29547 26312 29589 26321
rect 29547 26272 29548 26312
rect 29588 26272 29589 26312
rect 29547 26263 29589 26272
rect 29068 26144 29108 26153
rect 28724 26104 28820 26144
rect 28972 26104 29068 26144
rect 28684 26095 28724 26104
rect 28204 25892 28244 25901
rect 28244 25852 28532 25892
rect 28204 25843 28244 25852
rect 28203 25388 28245 25397
rect 28203 25348 28204 25388
rect 28244 25348 28245 25388
rect 28203 25339 28245 25348
rect 28204 25304 28244 25339
rect 28204 25253 28244 25264
rect 28107 24884 28149 24893
rect 28107 24844 28108 24884
rect 28148 24844 28149 24884
rect 28107 24835 28149 24844
rect 28108 24632 28148 24641
rect 28108 22793 28148 24592
rect 28203 23792 28245 23801
rect 28203 23752 28204 23792
rect 28244 23752 28245 23792
rect 28203 23743 28245 23752
rect 28204 23120 28244 23743
rect 28204 23071 28244 23080
rect 28107 22784 28149 22793
rect 28107 22744 28108 22784
rect 28148 22744 28149 22784
rect 28107 22735 28149 22744
rect 27148 21559 27188 21568
rect 28012 21559 28052 21568
rect 27435 20768 27477 20777
rect 27435 20728 27436 20768
rect 27476 20728 27477 20768
rect 27435 20719 27477 20728
rect 27436 20634 27476 20719
rect 27147 20516 27189 20525
rect 27147 20476 27148 20516
rect 27188 20476 27189 20516
rect 27147 20467 27189 20476
rect 27148 19508 27188 20467
rect 27820 20189 27860 20274
rect 27819 20180 27861 20189
rect 27819 20140 27820 20180
rect 27860 20140 27861 20180
rect 27819 20131 27861 20140
rect 27532 20096 27572 20105
rect 28492 20096 28532 25852
rect 28972 25649 29012 26104
rect 29068 26095 29108 26104
rect 29260 26144 29300 26263
rect 29260 26095 29300 26104
rect 29356 26144 29396 26153
rect 29356 25985 29396 26104
rect 29355 25976 29397 25985
rect 29355 25936 29356 25976
rect 29396 25936 29397 25976
rect 29355 25927 29397 25936
rect 28971 25640 29013 25649
rect 28971 25600 28972 25640
rect 29012 25600 29013 25640
rect 28971 25591 29013 25600
rect 29259 25388 29301 25397
rect 29259 25348 29260 25388
rect 29300 25348 29301 25388
rect 29259 25339 29301 25348
rect 28876 25304 28916 25313
rect 28588 24380 28628 24389
rect 28588 22709 28628 24340
rect 28876 23885 28916 25264
rect 29260 24632 29300 25339
rect 29548 24632 29588 26263
rect 29643 26228 29685 26237
rect 29643 26188 29644 26228
rect 29684 26188 29685 26228
rect 29643 26179 29685 26188
rect 29644 26144 29684 26179
rect 29644 26093 29684 26104
rect 29836 26144 29876 26153
rect 29836 25901 29876 26104
rect 29932 26144 29972 26153
rect 30028 26144 30068 26776
rect 29972 26104 30068 26144
rect 29932 26095 29972 26104
rect 29644 25892 29684 25901
rect 29644 24800 29684 25852
rect 29835 25892 29877 25901
rect 29835 25852 29836 25892
rect 29876 25852 29877 25892
rect 29835 25843 29877 25852
rect 29836 25304 29876 25315
rect 29836 25229 29876 25264
rect 29835 25220 29877 25229
rect 29835 25180 29836 25220
rect 29876 25180 29877 25220
rect 29835 25171 29877 25180
rect 29644 24760 30068 24800
rect 29644 24632 29684 24641
rect 29548 24592 29644 24632
rect 29260 24583 29300 24592
rect 29644 24583 29684 24592
rect 29836 24632 29876 24641
rect 29739 24380 29781 24389
rect 29739 24340 29740 24380
rect 29780 24340 29781 24380
rect 29739 24331 29781 24340
rect 29740 24246 29780 24331
rect 28875 23876 28917 23885
rect 28875 23836 28876 23876
rect 28916 23836 28917 23876
rect 28875 23827 28917 23836
rect 28876 23204 28916 23827
rect 29452 23792 29492 23801
rect 29740 23792 29780 23801
rect 29492 23752 29740 23792
rect 29452 23743 29492 23752
rect 29740 23743 29780 23752
rect 28972 23624 29012 23633
rect 28972 23381 29012 23584
rect 28971 23372 29013 23381
rect 28971 23332 28972 23372
rect 29012 23332 29013 23372
rect 28971 23323 29013 23332
rect 28876 23155 28916 23164
rect 29644 23120 29684 23129
rect 29260 23080 29644 23120
rect 29163 22952 29205 22961
rect 29163 22912 29164 22952
rect 29204 22912 29205 22952
rect 29163 22903 29205 22912
rect 29164 22793 29204 22903
rect 29163 22784 29205 22793
rect 29163 22744 29164 22784
rect 29204 22744 29205 22784
rect 29163 22735 29205 22744
rect 28587 22700 28629 22709
rect 28587 22660 28588 22700
rect 28628 22660 28629 22700
rect 28587 22651 28629 22660
rect 29164 22532 29204 22735
rect 29164 22483 29204 22492
rect 29164 21776 29204 21785
rect 29260 21776 29300 23080
rect 29644 23071 29684 23080
rect 29836 22952 29876 24592
rect 30028 24632 30068 24760
rect 30028 24583 30068 24592
rect 30124 24645 30164 24654
rect 30124 24389 30164 24605
rect 30123 24380 30165 24389
rect 30123 24340 30124 24380
rect 30164 24340 30165 24380
rect 30123 24331 30165 24340
rect 30220 23381 30260 26860
rect 30316 25892 30356 25901
rect 30316 25304 30356 25852
rect 30412 25565 30452 27784
rect 30507 27656 30549 27665
rect 30507 27616 30508 27656
rect 30548 27616 30549 27656
rect 30507 27607 30549 27616
rect 30700 27656 30740 28288
rect 30700 27607 30740 27616
rect 30795 27656 30837 27665
rect 30795 27616 30796 27656
rect 30836 27616 30837 27656
rect 30795 27607 30837 27616
rect 30508 27522 30548 27607
rect 30796 27522 30836 27607
rect 30507 27404 30549 27413
rect 30988 27404 31028 27413
rect 30507 27364 30508 27404
rect 30548 27364 30549 27404
rect 30507 27355 30549 27364
rect 30604 27364 30988 27404
rect 30508 27270 30548 27355
rect 30508 26816 30548 26825
rect 30508 25892 30548 26776
rect 30604 26816 30644 27364
rect 30988 27355 31028 27364
rect 30988 27077 31028 27162
rect 30987 27068 31029 27077
rect 30987 27028 30988 27068
rect 31028 27028 31029 27068
rect 30987 27019 31029 27028
rect 30700 26825 30740 26910
rect 30891 26900 30933 26909
rect 30891 26860 30892 26900
rect 30932 26860 31028 26900
rect 30891 26851 30933 26860
rect 30604 26767 30644 26776
rect 30699 26816 30741 26825
rect 30699 26776 30700 26816
rect 30740 26776 30741 26816
rect 30699 26767 30741 26776
rect 30988 26816 31028 26860
rect 30988 26767 31028 26776
rect 30796 26648 30836 26657
rect 30700 26608 30796 26648
rect 30603 26144 30645 26153
rect 30603 26104 30604 26144
rect 30644 26104 30645 26144
rect 30603 26095 30645 26104
rect 30700 26144 30740 26608
rect 30796 26599 30836 26608
rect 30796 26489 30836 26494
rect 30795 26480 30837 26489
rect 30795 26440 30796 26480
rect 30836 26440 30837 26480
rect 30795 26431 30837 26440
rect 30796 26370 30836 26431
rect 30796 26321 30836 26330
rect 30700 26095 30740 26104
rect 30604 26010 30644 26095
rect 30603 25892 30645 25901
rect 30508 25852 30604 25892
rect 30644 25852 30645 25892
rect 30603 25843 30645 25852
rect 30411 25556 30453 25565
rect 30411 25516 30412 25556
rect 30452 25516 30453 25556
rect 30411 25507 30453 25516
rect 30316 25255 30356 25264
rect 30508 25472 30548 25481
rect 30315 24884 30357 24893
rect 30315 24844 30316 24884
rect 30356 24844 30357 24884
rect 30315 24835 30357 24844
rect 30316 24632 30356 24835
rect 30411 24800 30453 24809
rect 30411 24760 30412 24800
rect 30452 24760 30453 24800
rect 30411 24751 30453 24760
rect 30316 24583 30356 24592
rect 30316 24464 30356 24473
rect 30412 24464 30452 24751
rect 30356 24424 30452 24464
rect 30316 24415 30356 24424
rect 30411 23792 30453 23801
rect 30411 23752 30412 23792
rect 30452 23752 30453 23792
rect 30411 23743 30453 23752
rect 30412 23658 30452 23743
rect 30219 23372 30261 23381
rect 30219 23332 30220 23372
rect 30260 23332 30261 23372
rect 30219 23323 30261 23332
rect 30316 23120 30356 23129
rect 30316 22961 30356 23080
rect 30411 23120 30453 23129
rect 30411 23080 30412 23120
rect 30452 23080 30453 23120
rect 30411 23071 30453 23080
rect 30412 22986 30452 23071
rect 30028 22952 30068 22961
rect 29836 22912 30028 22952
rect 30028 22903 30068 22912
rect 30315 22952 30357 22961
rect 30315 22912 30316 22952
rect 30356 22912 30357 22952
rect 30315 22903 30357 22912
rect 30315 22700 30357 22709
rect 30315 22660 30316 22700
rect 30356 22660 30357 22700
rect 30315 22651 30357 22660
rect 30316 22280 30356 22651
rect 30316 22231 30356 22240
rect 29204 21736 29300 21776
rect 29164 21727 29204 21736
rect 30219 21608 30261 21617
rect 30219 21568 30220 21608
rect 30260 21568 30261 21608
rect 30219 21559 30261 21568
rect 29835 21440 29877 21449
rect 29835 21400 29836 21440
rect 29876 21400 29877 21440
rect 29835 21391 29877 21400
rect 29836 21306 29876 21391
rect 30028 20936 30068 20945
rect 28683 20768 28725 20777
rect 28683 20728 28684 20768
rect 28724 20728 28725 20768
rect 28683 20719 28725 20728
rect 28588 20096 28628 20105
rect 27532 19517 27572 20056
rect 28300 20056 28588 20096
rect 28204 19844 28244 19853
rect 27148 19459 27188 19468
rect 27531 19508 27573 19517
rect 27531 19468 27532 19508
rect 27572 19468 27573 19508
rect 27531 19459 27573 19468
rect 26996 19216 27572 19256
rect 26956 19207 26996 19216
rect 25516 18880 26132 18920
rect 25995 18752 26037 18761
rect 25995 18712 25996 18752
rect 26036 18712 26037 18752
rect 25995 18703 26037 18712
rect 25707 18416 25749 18425
rect 25707 18376 25708 18416
rect 25748 18376 25749 18416
rect 25707 18367 25749 18376
rect 25612 18332 25652 18341
rect 25515 17996 25557 18005
rect 25420 17956 25516 17996
rect 25556 17956 25557 17996
rect 25515 17947 25557 17956
rect 25131 17912 25173 17921
rect 25131 17872 25132 17912
rect 25172 17872 25173 17912
rect 25131 17863 25173 17872
rect 25036 17695 25076 17704
rect 24884 17200 24980 17240
rect 24844 17191 24884 17200
rect 24748 17072 24788 17191
rect 24748 17023 24788 17032
rect 24940 17072 24980 17081
rect 24651 16736 24693 16745
rect 24651 16696 24652 16736
rect 24692 16696 24693 16736
rect 24651 16687 24693 16696
rect 24748 16064 24788 16073
rect 24267 15560 24309 15569
rect 24267 15520 24268 15560
rect 24308 15520 24309 15560
rect 24267 15511 24309 15520
rect 24364 15476 24404 15485
rect 24076 15100 24308 15140
rect 23979 15056 24021 15065
rect 23979 15016 23980 15056
rect 24020 15016 24021 15056
rect 23979 15007 24021 15016
rect 23595 14720 23637 14729
rect 23595 14680 23596 14720
rect 23636 14680 23637 14720
rect 23595 14671 23637 14680
rect 23692 14720 23732 14729
rect 23596 14586 23636 14671
rect 23500 14552 23540 14561
rect 23500 14057 23540 14512
rect 23499 14048 23541 14057
rect 23499 14008 23500 14048
rect 23540 14008 23541 14048
rect 23499 13999 23541 14008
rect 23692 13385 23732 14680
rect 23788 14720 23828 14729
rect 23788 14561 23828 14680
rect 23980 14720 24020 14729
rect 23787 14552 23829 14561
rect 23787 14512 23788 14552
rect 23828 14512 23829 14552
rect 23787 14503 23829 14512
rect 23980 14477 24020 14680
rect 24075 14720 24117 14729
rect 24075 14680 24076 14720
rect 24116 14680 24117 14720
rect 24075 14671 24117 14680
rect 24172 14720 24212 14729
rect 24076 14586 24116 14671
rect 24172 14561 24212 14680
rect 24171 14552 24213 14561
rect 24171 14512 24172 14552
rect 24212 14512 24213 14552
rect 24171 14503 24213 14512
rect 23979 14468 24021 14477
rect 23979 14428 23980 14468
rect 24020 14428 24021 14468
rect 23979 14419 24021 14428
rect 24268 14216 24308 15100
rect 24364 14720 24404 15436
rect 24748 14813 24788 16024
rect 24843 16064 24885 16073
rect 24843 16024 24844 16064
rect 24884 16024 24885 16064
rect 24843 16015 24885 16024
rect 24844 14972 24884 16015
rect 24940 15065 24980 17032
rect 25132 17072 25172 17863
rect 25420 17744 25460 17753
rect 25228 17704 25420 17744
rect 25228 17240 25268 17704
rect 25420 17695 25460 17704
rect 25228 17191 25268 17200
rect 25323 17240 25365 17249
rect 25323 17200 25324 17240
rect 25364 17200 25365 17240
rect 25323 17191 25365 17200
rect 25132 17023 25172 17032
rect 25228 16232 25268 16241
rect 25324 16232 25364 17191
rect 25420 17072 25460 17081
rect 25516 17072 25556 17947
rect 25612 17249 25652 18292
rect 25611 17240 25653 17249
rect 25611 17200 25612 17240
rect 25652 17200 25653 17240
rect 25611 17191 25653 17200
rect 25460 17032 25556 17072
rect 25612 17072 25652 17081
rect 25420 17023 25460 17032
rect 25612 16745 25652 17032
rect 25708 17072 25748 18367
rect 25803 17996 25845 18005
rect 25803 17956 25804 17996
rect 25844 17956 25845 17996
rect 25803 17947 25845 17956
rect 25708 17023 25748 17032
rect 25804 17072 25844 17947
rect 25804 17023 25844 17032
rect 25900 17072 25940 17081
rect 25611 16736 25653 16745
rect 25611 16696 25612 16736
rect 25652 16696 25653 16736
rect 25611 16687 25653 16696
rect 25268 16192 25364 16232
rect 25228 16183 25268 16192
rect 25227 15560 25269 15569
rect 25227 15520 25228 15560
rect 25268 15520 25269 15560
rect 25227 15511 25269 15520
rect 25228 15426 25268 15511
rect 24939 15056 24981 15065
rect 24939 15016 24940 15056
rect 24980 15016 24981 15056
rect 24939 15007 24981 15016
rect 24844 14923 24884 14932
rect 24747 14804 24789 14813
rect 24747 14764 24748 14804
rect 24788 14764 24789 14804
rect 24747 14755 24789 14764
rect 24556 14720 24596 14729
rect 24404 14680 24500 14720
rect 24364 14671 24404 14680
rect 24268 14176 24404 14216
rect 24268 14048 24308 14057
rect 23691 13376 23733 13385
rect 23691 13336 23692 13376
rect 23732 13336 23733 13376
rect 23691 13327 23733 13336
rect 23500 13208 23540 13217
rect 23404 13168 23500 13208
rect 23540 13168 23732 13208
rect 23307 13159 23349 13168
rect 23500 13159 23540 13168
rect 22923 13124 22965 13133
rect 22923 13084 22924 13124
rect 22964 13084 22965 13124
rect 22923 13075 22965 13084
rect 22924 12990 22964 13075
rect 23020 10865 23060 13159
rect 23308 13074 23348 13159
rect 23500 11696 23540 11705
rect 23500 11285 23540 11656
rect 23595 11696 23637 11705
rect 23595 11656 23596 11696
rect 23636 11656 23637 11696
rect 23595 11647 23637 11656
rect 23692 11696 23732 13168
rect 24268 13133 24308 14008
rect 24267 13124 24309 13133
rect 24267 13084 24268 13124
rect 24308 13084 24309 13124
rect 24267 13075 24309 13084
rect 23979 11696 24021 11705
rect 23732 11656 23924 11696
rect 23692 11647 23732 11656
rect 23596 11562 23636 11647
rect 23499 11276 23541 11285
rect 23499 11236 23500 11276
rect 23540 11236 23541 11276
rect 23499 11227 23541 11236
rect 23403 11192 23445 11201
rect 23403 11152 23404 11192
rect 23444 11152 23445 11192
rect 23403 11143 23445 11152
rect 23019 10856 23061 10865
rect 23019 10816 23020 10856
rect 23060 10816 23061 10856
rect 23019 10807 23061 10816
rect 23020 10352 23060 10361
rect 23404 10352 23444 11143
rect 23500 11024 23540 11227
rect 23884 11201 23924 11656
rect 23979 11656 23980 11696
rect 24020 11656 24021 11696
rect 23979 11647 24021 11656
rect 23980 11562 24020 11647
rect 24171 11276 24213 11285
rect 24171 11236 24172 11276
rect 24212 11236 24213 11276
rect 24171 11227 24213 11236
rect 23883 11192 23925 11201
rect 23883 11152 23884 11192
rect 23924 11152 23925 11192
rect 23883 11143 23925 11152
rect 23596 11024 23636 11033
rect 23500 10984 23596 11024
rect 23596 10975 23636 10984
rect 23692 11024 23732 11033
rect 23884 11024 23924 11033
rect 23692 10865 23732 10984
rect 23788 10984 23884 11024
rect 23691 10856 23733 10865
rect 23691 10816 23692 10856
rect 23732 10816 23733 10856
rect 23691 10807 23733 10816
rect 23060 10312 23252 10352
rect 23404 10312 23540 10352
rect 23020 10303 23060 10312
rect 22923 10268 22965 10277
rect 22923 10228 22924 10268
rect 22964 10228 22965 10268
rect 22923 10219 22965 10228
rect 22924 10184 22964 10219
rect 22924 10133 22964 10144
rect 23020 10184 23060 10193
rect 23020 9848 23060 10144
rect 23212 10184 23252 10312
rect 23212 10135 23252 10144
rect 23308 10184 23348 10193
rect 23308 10025 23348 10144
rect 23403 10184 23445 10193
rect 23403 10144 23404 10184
rect 23444 10144 23445 10184
rect 23403 10135 23445 10144
rect 23500 10184 23540 10312
rect 23696 10268 23738 10277
rect 23696 10228 23697 10268
rect 23737 10228 23738 10268
rect 23696 10219 23738 10228
rect 23307 10016 23349 10025
rect 23307 9976 23308 10016
rect 23348 9976 23349 10016
rect 23307 9967 23349 9976
rect 23404 10016 23444 10135
rect 23404 9967 23444 9976
rect 23500 9848 23540 10144
rect 23595 10184 23637 10193
rect 23595 10144 23596 10184
rect 23636 10144 23637 10184
rect 23595 10135 23637 10144
rect 23697 10184 23737 10219
rect 23020 9808 23540 9848
rect 23307 9680 23349 9689
rect 23307 9640 23308 9680
rect 23348 9640 23349 9680
rect 23307 9631 23349 9640
rect 23212 9512 23252 9521
rect 22924 9472 23212 9512
rect 22827 9176 22869 9185
rect 22827 9136 22828 9176
rect 22868 9136 22869 9176
rect 22827 9127 22869 9136
rect 22731 9092 22773 9101
rect 22731 9052 22732 9092
rect 22772 9052 22773 9092
rect 22731 9043 22773 9052
rect 22828 8933 22868 9018
rect 22827 8924 22869 8933
rect 22827 8884 22828 8924
rect 22868 8884 22869 8924
rect 22827 8875 22869 8884
rect 22443 8840 22485 8849
rect 22443 8800 22444 8840
rect 22484 8800 22485 8840
rect 22443 8791 22485 8800
rect 22732 8681 22772 8766
rect 22924 8756 22964 9472
rect 23212 9463 23252 9472
rect 23115 9260 23157 9269
rect 23115 9220 23116 9260
rect 23156 9220 23157 9260
rect 23115 9211 23157 9220
rect 23019 9176 23061 9185
rect 23019 9136 23020 9176
rect 23060 9136 23061 9176
rect 23019 9127 23061 9136
rect 23020 8756 23060 9127
rect 23116 8840 23156 9211
rect 23211 8840 23253 8849
rect 23116 8800 23158 8840
rect 22828 8716 22964 8756
rect 23013 8716 23060 8756
rect 22731 8672 22773 8681
rect 22731 8632 22732 8672
rect 22772 8632 22773 8672
rect 22731 8623 22773 8632
rect 22347 8588 22389 8597
rect 22347 8548 22348 8588
rect 22388 8548 22389 8588
rect 22347 8539 22389 8548
rect 22348 8429 22388 8539
rect 22347 8420 22389 8429
rect 22347 8380 22348 8420
rect 22388 8380 22389 8420
rect 22347 8371 22389 8380
rect 22539 8420 22581 8429
rect 22539 8380 22540 8420
rect 22580 8380 22581 8420
rect 22539 8371 22581 8380
rect 22348 8000 22388 8371
rect 22348 7951 22388 7960
rect 22443 8000 22485 8009
rect 22443 7960 22444 8000
rect 22484 7960 22485 8000
rect 22443 7951 22485 7960
rect 22540 8000 22580 8371
rect 22828 8168 22868 8716
rect 22919 8651 22959 8660
rect 22919 8513 22959 8611
rect 22918 8504 22960 8513
rect 22918 8464 22919 8504
rect 22959 8464 22960 8504
rect 22918 8455 22960 8464
rect 23013 8429 23053 8716
rect 23118 8681 23158 8800
rect 23211 8800 23212 8840
rect 23252 8800 23253 8840
rect 23211 8791 23253 8800
rect 23116 8672 23158 8681
rect 23156 8632 23158 8672
rect 23116 8623 23156 8632
rect 23212 8588 23252 8791
rect 23308 8672 23348 9631
rect 23308 8597 23348 8632
rect 23403 8672 23445 8681
rect 23403 8632 23404 8672
rect 23444 8632 23445 8672
rect 23403 8623 23445 8632
rect 23212 8539 23252 8548
rect 23307 8588 23349 8597
rect 23307 8548 23308 8588
rect 23348 8548 23349 8588
rect 23307 8539 23349 8548
rect 23308 8508 23348 8539
rect 23404 8538 23444 8623
rect 23013 8420 23061 8429
rect 23013 8380 23020 8420
rect 23060 8380 23061 8420
rect 23019 8371 23061 8380
rect 23115 8336 23157 8345
rect 23500 8336 23540 9808
rect 23596 9512 23636 10135
rect 23697 10133 23737 10144
rect 23788 9680 23828 10984
rect 23884 10975 23924 10984
rect 24075 11024 24117 11033
rect 24075 10984 24076 11024
rect 24116 10984 24117 11024
rect 24075 10975 24117 10984
rect 24172 11024 24212 11227
rect 24364 11192 24404 14176
rect 24460 13628 24500 14680
rect 24556 13880 24596 14680
rect 24651 14720 24693 14729
rect 24651 14680 24652 14720
rect 24692 14680 24693 14720
rect 24651 14671 24693 14680
rect 24652 14586 24692 14671
rect 24556 13831 24596 13840
rect 24460 13588 24596 13628
rect 24459 11528 24501 11537
rect 24459 11488 24460 11528
rect 24500 11488 24501 11528
rect 24459 11479 24501 11488
rect 24460 11394 24500 11479
rect 24364 11152 24500 11192
rect 24172 10975 24212 10984
rect 24268 11024 24308 11033
rect 24076 10890 24116 10975
rect 23884 10772 23924 10781
rect 23884 10184 23924 10732
rect 23980 10436 24020 10445
rect 24268 10436 24308 10984
rect 24363 11024 24405 11033
rect 24363 10984 24364 11024
rect 24404 10984 24405 11024
rect 24363 10975 24405 10984
rect 24364 10890 24404 10975
rect 24020 10396 24308 10436
rect 23980 10387 24020 10396
rect 24460 10352 24500 11152
rect 24556 11033 24596 13588
rect 24748 13544 24788 14755
rect 24940 14729 24980 15007
rect 25131 14888 25173 14897
rect 25131 14848 25132 14888
rect 25172 14848 25173 14888
rect 25131 14839 25173 14848
rect 25132 14754 25172 14839
rect 24939 14720 24981 14729
rect 24939 14680 24940 14720
rect 24980 14680 24981 14720
rect 24939 14671 24981 14680
rect 25324 14561 25364 16192
rect 25900 16232 25940 17032
rect 25900 16183 25940 16192
rect 25515 16064 25557 16073
rect 25515 16024 25516 16064
rect 25556 16024 25557 16064
rect 25515 16015 25557 16024
rect 25707 16064 25749 16073
rect 25707 16024 25708 16064
rect 25748 16024 25749 16064
rect 25707 16015 25749 16024
rect 25516 15930 25556 16015
rect 25708 15930 25748 16015
rect 25996 15140 26036 18703
rect 26092 18584 26132 18593
rect 26188 18584 26228 19207
rect 27340 19088 27380 19097
rect 26132 18544 26228 18584
rect 26956 19048 27340 19088
rect 26092 18535 26132 18544
rect 26379 17996 26421 18005
rect 26379 17956 26380 17996
rect 26420 17956 26421 17996
rect 26379 17947 26421 17956
rect 26380 17744 26420 17947
rect 26380 17695 26420 17704
rect 26668 17660 26708 17669
rect 26572 17249 26612 17334
rect 26571 17240 26613 17249
rect 26571 17200 26572 17240
rect 26612 17200 26613 17240
rect 26571 17191 26613 17200
rect 26380 17081 26420 17166
rect 26379 17072 26421 17081
rect 26379 17032 26380 17072
rect 26420 17032 26421 17072
rect 26379 17023 26421 17032
rect 26572 17072 26612 17083
rect 26572 16997 26612 17032
rect 26571 16988 26613 16997
rect 26571 16948 26572 16988
rect 26612 16948 26613 16988
rect 26571 16939 26613 16948
rect 26572 16745 26612 16939
rect 26571 16736 26613 16745
rect 26571 16696 26572 16736
rect 26612 16696 26613 16736
rect 26571 16687 26613 16696
rect 26091 15812 26133 15821
rect 26091 15772 26092 15812
rect 26132 15772 26133 15812
rect 26091 15763 26133 15772
rect 26092 15644 26132 15763
rect 26092 15595 26132 15604
rect 25420 15100 26036 15140
rect 26284 15308 26324 15317
rect 25420 14720 25460 15100
rect 25420 14671 25460 14680
rect 25516 14720 25556 14729
rect 25323 14552 25365 14561
rect 25323 14512 25324 14552
rect 25364 14512 25365 14552
rect 25323 14503 25365 14512
rect 25516 14141 25556 14680
rect 25804 14720 25844 14729
rect 26187 14720 26229 14729
rect 25844 14680 25940 14720
rect 25804 14671 25844 14680
rect 25803 14468 25845 14477
rect 25803 14428 25804 14468
rect 25844 14428 25845 14468
rect 25803 14419 25845 14428
rect 25515 14132 25557 14141
rect 25515 14092 25516 14132
rect 25556 14092 25557 14132
rect 25515 14083 25557 14092
rect 24940 13880 24980 13889
rect 24980 13840 25076 13880
rect 24940 13831 24980 13840
rect 24748 13504 24980 13544
rect 24652 13208 24692 13219
rect 24652 13133 24692 13168
rect 24651 13124 24693 13133
rect 24651 13084 24652 13124
rect 24692 13084 24693 13124
rect 24651 13075 24693 13084
rect 24843 11948 24885 11957
rect 24843 11908 24844 11948
rect 24884 11908 24885 11948
rect 24843 11899 24885 11908
rect 24844 11780 24884 11899
rect 24844 11731 24884 11740
rect 24747 11192 24789 11201
rect 24747 11152 24748 11192
rect 24788 11152 24789 11192
rect 24747 11143 24789 11152
rect 24555 11024 24597 11033
rect 24748 11024 24788 11143
rect 24555 10984 24556 11024
rect 24596 10984 24692 11024
rect 24555 10975 24597 10984
rect 24555 10436 24597 10445
rect 24555 10396 24556 10436
rect 24596 10396 24597 10436
rect 24555 10387 24597 10396
rect 24172 10312 24500 10352
rect 23980 10184 24020 10193
rect 23884 10144 23980 10184
rect 23980 10135 24020 10144
rect 24076 10184 24116 10193
rect 24076 10025 24116 10144
rect 24075 10016 24117 10025
rect 24075 9976 24076 10016
rect 24116 9976 24117 10016
rect 24075 9967 24117 9976
rect 24172 9941 24212 10312
rect 24556 10268 24596 10387
rect 24521 10228 24596 10268
rect 24521 10199 24561 10228
rect 24268 10184 24308 10193
rect 24268 10025 24308 10144
rect 24363 10184 24405 10193
rect 24363 10144 24364 10184
rect 24404 10144 24405 10184
rect 24521 10150 24561 10159
rect 24363 10135 24405 10144
rect 24364 10050 24404 10135
rect 24267 10016 24309 10025
rect 24267 9976 24268 10016
rect 24308 9976 24309 10016
rect 24267 9967 24309 9976
rect 24171 9932 24213 9941
rect 24171 9892 24172 9932
rect 24212 9892 24213 9932
rect 24171 9883 24213 9892
rect 24652 9848 24692 10984
rect 24748 10975 24788 10984
rect 24843 11024 24885 11033
rect 24843 10984 24844 11024
rect 24884 10984 24885 11024
rect 24843 10975 24885 10984
rect 24844 10890 24884 10975
rect 24940 10940 24980 13504
rect 25036 12125 25076 13840
rect 25804 13460 25844 14419
rect 25900 13973 25940 14680
rect 26187 14680 26188 14720
rect 26228 14680 26229 14720
rect 26187 14671 26229 14680
rect 26092 14561 26132 14646
rect 26188 14586 26228 14671
rect 26091 14552 26133 14561
rect 26091 14512 26092 14552
rect 26132 14512 26133 14552
rect 26091 14503 26133 14512
rect 26091 14300 26133 14309
rect 26091 14260 26092 14300
rect 26132 14260 26133 14300
rect 26091 14251 26133 14260
rect 26092 14216 26132 14251
rect 26092 14165 26132 14176
rect 25899 13964 25941 13973
rect 25899 13924 25900 13964
rect 25940 13924 25941 13964
rect 25899 13915 25941 13924
rect 25804 13411 25844 13420
rect 25900 13796 25940 13805
rect 25612 13208 25652 13217
rect 25612 12713 25652 13168
rect 25611 12704 25653 12713
rect 25611 12664 25612 12704
rect 25652 12664 25653 12704
rect 25611 12655 25653 12664
rect 25612 12284 25652 12293
rect 25035 12116 25077 12125
rect 25035 12076 25036 12116
rect 25076 12076 25077 12116
rect 25035 12067 25077 12076
rect 25036 11453 25076 12067
rect 25035 11444 25077 11453
rect 25035 11404 25036 11444
rect 25076 11404 25077 11444
rect 25035 11395 25077 11404
rect 24940 10891 24980 10900
rect 25036 10856 25076 10865
rect 24747 10436 24789 10445
rect 24747 10396 24748 10436
rect 24788 10396 24789 10436
rect 24747 10387 24789 10396
rect 24268 9808 24692 9848
rect 23788 9640 24116 9680
rect 23692 9596 23732 9607
rect 23692 9521 23732 9556
rect 23596 9008 23636 9472
rect 23691 9512 23733 9521
rect 23980 9512 24020 9521
rect 23691 9472 23692 9512
rect 23732 9472 23733 9512
rect 23691 9463 23733 9472
rect 23788 9472 23980 9512
rect 23596 8968 23732 9008
rect 23595 8840 23637 8849
rect 23595 8800 23596 8840
rect 23636 8800 23637 8840
rect 23595 8791 23637 8800
rect 23596 8504 23636 8791
rect 23692 8681 23732 8968
rect 23788 8933 23828 9472
rect 23980 9463 24020 9472
rect 24076 9437 24116 9640
rect 24171 9512 24213 9521
rect 24171 9472 24172 9512
rect 24212 9472 24213 9512
rect 24171 9463 24213 9472
rect 24075 9428 24117 9437
rect 24075 9388 24076 9428
rect 24116 9388 24117 9428
rect 24075 9379 24117 9388
rect 24172 9378 24212 9463
rect 24171 9260 24213 9269
rect 24171 9220 24172 9260
rect 24212 9220 24213 9260
rect 24171 9211 24213 9220
rect 24172 9126 24212 9211
rect 23787 8924 23829 8933
rect 24268 8924 24308 9808
rect 24652 9680 24692 9689
rect 24364 9512 24404 9521
rect 24364 8933 24404 9472
rect 24460 9512 24500 9521
rect 23787 8884 23788 8924
rect 23828 8884 23829 8924
rect 23787 8875 23829 8884
rect 23980 8884 24308 8924
rect 24363 8924 24405 8933
rect 24363 8884 24364 8924
rect 24404 8884 24405 8924
rect 23691 8672 23733 8681
rect 23691 8632 23692 8672
rect 23732 8632 23733 8672
rect 23691 8623 23733 8632
rect 23788 8672 23828 8875
rect 23980 8756 24020 8884
rect 24363 8875 24405 8884
rect 23980 8716 24021 8756
rect 23788 8623 23828 8632
rect 23883 8672 23925 8681
rect 23883 8632 23884 8672
rect 23924 8632 23925 8672
rect 23883 8623 23925 8632
rect 23884 8538 23924 8623
rect 23981 8588 24021 8716
rect 24076 8681 24116 8766
rect 24363 8756 24405 8765
rect 24363 8716 24364 8756
rect 24404 8716 24405 8756
rect 24363 8707 24405 8716
rect 24075 8672 24117 8681
rect 24075 8632 24076 8672
rect 24116 8632 24117 8672
rect 24075 8623 24117 8632
rect 24172 8672 24212 8681
rect 23980 8548 24021 8588
rect 23596 8455 23636 8464
rect 23115 8296 23116 8336
rect 23156 8296 23157 8336
rect 23115 8287 23157 8296
rect 23404 8296 23540 8336
rect 23595 8336 23637 8345
rect 23595 8296 23596 8336
rect 23636 8296 23637 8336
rect 23019 8252 23061 8261
rect 23019 8212 23020 8252
rect 23060 8212 23061 8252
rect 23019 8203 23061 8212
rect 22444 7866 22484 7951
rect 22155 7664 22197 7673
rect 22155 7624 22156 7664
rect 22196 7624 22197 7664
rect 22155 7615 22197 7624
rect 22059 7580 22101 7589
rect 22059 7540 22060 7580
rect 22100 7540 22101 7580
rect 22059 7531 22101 7540
rect 21675 7328 21717 7337
rect 21675 7288 21676 7328
rect 21716 7288 21717 7328
rect 21675 7279 21717 7288
rect 21580 7111 21620 7120
rect 21484 6952 21620 6992
rect 21483 6404 21525 6413
rect 21483 6364 21484 6404
rect 21524 6364 21525 6404
rect 21483 6355 21525 6364
rect 21387 5816 21429 5825
rect 21387 5776 21388 5816
rect 21428 5776 21429 5816
rect 21387 5767 21429 5776
rect 21388 5682 21428 5767
rect 20852 5608 21292 5648
rect 20812 5599 20852 5608
rect 21292 5599 21332 5608
rect 21484 5648 21524 6355
rect 20524 5564 20564 5573
rect 20564 5524 20660 5564
rect 20524 5515 20564 5524
rect 20620 5144 20660 5524
rect 20812 5480 20852 5489
rect 20852 5440 20948 5480
rect 20812 5431 20852 5440
rect 20908 5237 20948 5440
rect 21484 5396 21524 5608
rect 21580 5573 21620 6952
rect 21676 6988 21716 7279
rect 22347 7244 22389 7253
rect 22347 7204 22348 7244
rect 22388 7204 22389 7244
rect 22347 7195 22389 7204
rect 22251 7160 22293 7169
rect 22251 7120 22252 7160
rect 22292 7120 22293 7160
rect 22251 7111 22293 7120
rect 22348 7160 22388 7195
rect 22252 7026 22292 7111
rect 22348 7109 22388 7120
rect 22540 7160 22580 7960
rect 22636 8128 22868 8168
rect 22636 7505 22676 8128
rect 22732 8000 22772 8009
rect 22732 7841 22772 7960
rect 22924 8000 22964 8009
rect 22731 7832 22773 7841
rect 22731 7792 22732 7832
rect 22772 7792 22773 7832
rect 22731 7783 22773 7792
rect 22731 7580 22773 7589
rect 22731 7540 22732 7580
rect 22772 7540 22773 7580
rect 22731 7531 22773 7540
rect 22635 7496 22677 7505
rect 22635 7456 22636 7496
rect 22676 7456 22677 7496
rect 22635 7447 22677 7456
rect 22540 7111 22580 7120
rect 22636 7160 22676 7447
rect 22636 7111 22676 7120
rect 21676 6939 21716 6948
rect 22539 6908 22581 6917
rect 22539 6868 22540 6908
rect 22580 6868 22581 6908
rect 22539 6859 22581 6868
rect 22540 6488 22580 6859
rect 22540 6439 22580 6448
rect 22636 6413 22676 6498
rect 22732 6497 22772 7531
rect 22924 7421 22964 7960
rect 23020 8000 23060 8203
rect 23020 7951 23060 7960
rect 23020 7832 23060 7841
rect 23116 7832 23156 8287
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 23212 8000 23252 8119
rect 23307 8084 23349 8093
rect 23307 8044 23308 8084
rect 23348 8044 23349 8084
rect 23307 8035 23349 8044
rect 23212 7951 23252 7960
rect 23308 8000 23348 8035
rect 23308 7949 23348 7960
rect 23404 7916 23444 8296
rect 23595 8287 23637 8296
rect 23787 8336 23829 8345
rect 23787 8296 23788 8336
rect 23828 8296 23829 8336
rect 23787 8287 23829 8296
rect 23499 8168 23541 8177
rect 23499 8128 23500 8168
rect 23540 8128 23541 8168
rect 23499 8119 23541 8128
rect 23500 8034 23540 8119
rect 23395 7876 23444 7916
rect 23395 7832 23435 7876
rect 23060 7792 23156 7832
rect 23212 7792 23435 7832
rect 23596 7832 23636 8287
rect 23691 8084 23733 8093
rect 23691 8044 23692 8084
rect 23732 8044 23733 8084
rect 23691 8035 23733 8044
rect 23692 8000 23732 8035
rect 23692 7949 23732 7960
rect 23788 8000 23828 8287
rect 23980 8168 24020 8548
rect 24172 8177 24212 8632
rect 24267 8672 24309 8681
rect 24267 8632 24268 8672
rect 24308 8632 24309 8672
rect 24267 8623 24309 8632
rect 24364 8672 24404 8707
rect 24171 8168 24213 8177
rect 23980 8128 24116 8168
rect 23884 8009 23924 8094
rect 23788 7951 23828 7960
rect 23883 8000 23925 8009
rect 23883 7960 23884 8000
rect 23924 7960 23925 8000
rect 23883 7951 23925 7960
rect 23980 8000 24020 8009
rect 23980 7841 24020 7960
rect 23979 7832 24021 7841
rect 23596 7792 23924 7832
rect 23020 7783 23060 7792
rect 23019 7580 23061 7589
rect 23019 7540 23020 7580
rect 23060 7540 23061 7580
rect 23019 7531 23061 7540
rect 22923 7412 22965 7421
rect 22923 7372 22924 7412
rect 22964 7372 22965 7412
rect 22923 7363 22965 7372
rect 23020 7160 23060 7531
rect 23212 7496 23252 7792
rect 23595 7664 23637 7673
rect 23595 7624 23596 7664
rect 23636 7624 23637 7664
rect 23595 7615 23637 7624
rect 23116 7456 23252 7496
rect 23116 7253 23156 7456
rect 23596 7412 23636 7615
rect 23596 7363 23636 7372
rect 23211 7328 23253 7337
rect 23211 7288 23212 7328
rect 23252 7288 23253 7328
rect 23211 7279 23253 7288
rect 23403 7328 23445 7337
rect 23403 7288 23404 7328
rect 23444 7288 23445 7328
rect 23403 7279 23445 7288
rect 23115 7244 23157 7253
rect 23115 7204 23116 7244
rect 23156 7204 23157 7244
rect 23115 7195 23157 7204
rect 23020 7111 23060 7120
rect 22827 6992 22869 7001
rect 22827 6952 22828 6992
rect 22868 6952 22869 6992
rect 22827 6943 22869 6952
rect 22828 6858 22868 6943
rect 23116 6665 23156 7195
rect 23212 7194 23252 7279
rect 23307 7244 23349 7253
rect 23307 7204 23308 7244
rect 23348 7204 23349 7244
rect 23307 7195 23349 7204
rect 23308 7110 23348 7195
rect 23404 7160 23444 7279
rect 23404 7111 23444 7120
rect 23595 7160 23637 7169
rect 23595 7120 23596 7160
rect 23636 7120 23637 7160
rect 23595 7111 23637 7120
rect 23692 7160 23732 7169
rect 23787 7160 23829 7169
rect 23732 7120 23788 7160
rect 23828 7120 23829 7160
rect 23692 7111 23732 7120
rect 23787 7111 23829 7120
rect 23884 7160 23924 7792
rect 23979 7792 23980 7832
rect 24020 7792 24021 7832
rect 23979 7783 24021 7792
rect 23884 7111 23924 7120
rect 23980 7160 24020 7783
rect 24076 7496 24116 8128
rect 24171 8128 24172 8168
rect 24212 8128 24213 8168
rect 24171 8119 24213 8128
rect 24268 7673 24308 8623
rect 24364 8597 24404 8632
rect 24363 8588 24405 8597
rect 24363 8548 24364 8588
rect 24404 8548 24405 8588
rect 24363 8539 24405 8548
rect 24364 8508 24404 8539
rect 24363 8252 24405 8261
rect 24363 8212 24364 8252
rect 24404 8212 24405 8252
rect 24363 8203 24405 8212
rect 24267 7664 24309 7673
rect 24267 7624 24268 7664
rect 24308 7624 24309 7664
rect 24267 7615 24309 7624
rect 24076 7456 24308 7496
rect 24171 7328 24213 7337
rect 24171 7288 24172 7328
rect 24212 7288 24213 7328
rect 24171 7279 24213 7288
rect 23980 7111 24020 7120
rect 24081 7160 24121 7169
rect 23596 7026 23636 7111
rect 24081 7001 24121 7120
rect 24080 6992 24122 7001
rect 24080 6952 24081 6992
rect 24121 6952 24122 6992
rect 24080 6943 24122 6952
rect 23691 6908 23733 6917
rect 23691 6868 23692 6908
rect 23732 6868 23733 6908
rect 23691 6859 23733 6868
rect 23211 6824 23253 6833
rect 23211 6784 23212 6824
rect 23252 6784 23253 6824
rect 23211 6775 23253 6784
rect 23115 6656 23157 6665
rect 23115 6616 23116 6656
rect 23156 6616 23157 6656
rect 23115 6607 23157 6616
rect 22827 6572 22869 6581
rect 22827 6532 22828 6572
rect 22868 6532 22964 6572
rect 22827 6523 22869 6532
rect 22924 6530 22964 6532
rect 22731 6488 22773 6497
rect 22731 6448 22732 6488
rect 22772 6448 22773 6488
rect 22924 6481 22964 6490
rect 23115 6488 23157 6497
rect 22731 6439 22773 6448
rect 23115 6448 23116 6488
rect 23156 6448 23157 6488
rect 23115 6439 23157 6448
rect 22635 6404 22677 6413
rect 22635 6364 22636 6404
rect 22676 6364 22677 6404
rect 22635 6355 22677 6364
rect 22828 6404 22868 6415
rect 22828 6329 22868 6364
rect 23116 6354 23156 6439
rect 23212 6413 23252 6775
rect 23499 6572 23541 6581
rect 23499 6532 23500 6572
rect 23540 6532 23541 6572
rect 23499 6523 23541 6532
rect 23500 6488 23540 6523
rect 23500 6437 23540 6448
rect 23692 6488 23732 6859
rect 23787 6656 23829 6665
rect 23787 6616 23788 6656
rect 23828 6616 23829 6656
rect 23787 6607 23829 6616
rect 23211 6404 23253 6413
rect 23211 6364 23212 6404
rect 23252 6364 23253 6404
rect 23211 6355 23253 6364
rect 23403 6404 23445 6413
rect 23403 6364 23404 6404
rect 23444 6364 23445 6404
rect 23403 6355 23445 6364
rect 22732 6320 22772 6329
rect 22059 6236 22101 6245
rect 22732 6236 22772 6280
rect 22827 6320 22869 6329
rect 22827 6280 22828 6320
rect 22868 6280 22869 6320
rect 22827 6271 22869 6280
rect 23212 6270 23252 6355
rect 23308 6320 23348 6329
rect 22059 6196 22060 6236
rect 22100 6196 22101 6236
rect 22059 6187 22101 6196
rect 22540 6196 22772 6236
rect 23019 6236 23061 6245
rect 23019 6196 23020 6236
rect 23060 6196 23061 6236
rect 22060 5900 22100 6187
rect 22060 5851 22100 5860
rect 22443 5732 22485 5741
rect 22443 5692 22444 5732
rect 22484 5692 22485 5732
rect 22443 5683 22485 5692
rect 22348 5648 22388 5659
rect 22348 5573 22388 5608
rect 22444 5648 22484 5683
rect 22444 5597 22484 5608
rect 21579 5564 21621 5573
rect 21579 5524 21580 5564
rect 21620 5524 21621 5564
rect 21579 5515 21621 5524
rect 22347 5564 22389 5573
rect 22347 5524 22348 5564
rect 22388 5524 22389 5564
rect 22347 5515 22389 5524
rect 22540 5476 22580 6196
rect 23019 6187 23061 6196
rect 22731 5816 22773 5825
rect 22731 5776 22732 5816
rect 22772 5776 22773 5816
rect 22731 5767 22773 5776
rect 22540 5427 22580 5436
rect 21388 5356 22100 5396
rect 20907 5228 20949 5237
rect 20907 5188 20908 5228
rect 20948 5188 20949 5228
rect 20907 5179 20949 5188
rect 20620 5104 20852 5144
rect 20428 4976 20468 4985
rect 20331 4304 20373 4313
rect 20331 4264 20332 4304
rect 20372 4264 20373 4304
rect 20331 4255 20373 4264
rect 20043 4220 20085 4229
rect 20043 4180 20044 4220
rect 20084 4180 20085 4220
rect 20043 4171 20085 4180
rect 19412 4096 19508 4136
rect 20331 4136 20373 4145
rect 20331 4096 20332 4136
rect 20372 4096 20373 4136
rect 19372 3641 19412 4096
rect 20331 4087 20373 4096
rect 20332 4002 20372 4087
rect 20235 3968 20277 3977
rect 20235 3928 20236 3968
rect 20276 3928 20277 3968
rect 20235 3919 20277 3928
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 19947 3716 19989 3725
rect 19947 3676 19948 3716
rect 19988 3676 19989 3716
rect 19947 3667 19989 3676
rect 19371 3632 19413 3641
rect 19371 3592 19372 3632
rect 19412 3592 19413 3632
rect 19371 3583 19413 3592
rect 19275 3464 19317 3473
rect 19275 3424 19276 3464
rect 19316 3424 19317 3464
rect 19372 3464 19412 3583
rect 19755 3548 19797 3557
rect 19755 3508 19756 3548
rect 19796 3508 19797 3548
rect 19755 3499 19797 3508
rect 19564 3464 19604 3473
rect 19372 3424 19564 3464
rect 19275 3415 19317 3424
rect 19564 3415 19604 3424
rect 19179 3380 19221 3389
rect 19179 3340 19180 3380
rect 19220 3340 19221 3380
rect 19179 3331 19221 3340
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 18315 2876 18357 2885
rect 18124 2836 18260 2876
rect 17931 2827 17973 2836
rect 17835 2792 17877 2801
rect 17835 2752 17836 2792
rect 17876 2752 17877 2792
rect 17835 2743 17877 2752
rect 18027 2792 18069 2801
rect 18027 2752 18028 2792
rect 18068 2752 18069 2792
rect 18027 2743 18069 2752
rect 17836 2624 17876 2743
rect 17836 2575 17876 2584
rect 18028 2540 18068 2743
rect 18028 2491 18068 2500
rect 18123 2540 18165 2549
rect 18123 2500 18124 2540
rect 18164 2500 18165 2540
rect 18123 2491 18165 2500
rect 17931 2456 17973 2465
rect 17931 2416 17932 2456
rect 17972 2416 17973 2456
rect 17931 2407 17973 2416
rect 17740 1903 17780 1912
rect 17932 1952 17972 2407
rect 17932 1903 17972 1912
rect 18028 1952 18068 1961
rect 18124 1952 18164 2491
rect 18068 1912 18164 1952
rect 18220 1952 18260 2836
rect 18315 2836 18316 2876
rect 18356 2836 18357 2876
rect 18315 2827 18357 2836
rect 18316 2624 18356 2827
rect 18316 2549 18356 2584
rect 18412 2624 18452 2633
rect 18315 2540 18357 2549
rect 18315 2500 18316 2540
rect 18356 2500 18357 2540
rect 18315 2491 18357 2500
rect 18316 2460 18356 2491
rect 18412 2465 18452 2584
rect 18508 2624 18548 2633
rect 19180 2624 19220 3331
rect 19276 3330 19316 3415
rect 19371 2960 19413 2969
rect 19371 2920 19372 2960
rect 19412 2920 19413 2960
rect 19371 2911 19413 2920
rect 19276 2624 19316 2633
rect 19180 2584 19276 2624
rect 18411 2456 18453 2465
rect 18411 2416 18412 2456
rect 18452 2416 18453 2456
rect 18411 2407 18453 2416
rect 18028 1903 18068 1912
rect 18220 1903 18260 1912
rect 18220 1784 18260 1793
rect 18508 1784 18548 2584
rect 19276 2575 19316 2584
rect 19372 2624 19412 2911
rect 19467 2708 19509 2717
rect 19467 2668 19468 2708
rect 19508 2668 19509 2708
rect 19467 2659 19509 2668
rect 19372 2575 19412 2584
rect 19468 2624 19508 2659
rect 19468 2573 19508 2584
rect 19659 2624 19701 2633
rect 19659 2584 19660 2624
rect 19700 2584 19701 2624
rect 19756 2624 19796 3499
rect 19851 2624 19893 2633
rect 19756 2584 19852 2624
rect 19892 2584 19893 2624
rect 19659 2575 19701 2584
rect 19851 2575 19893 2584
rect 19948 2624 19988 3667
rect 20139 3464 20181 3473
rect 20139 3424 20140 3464
rect 20180 3424 20181 3464
rect 20139 3415 20181 3424
rect 20140 3305 20180 3415
rect 20139 3296 20181 3305
rect 20139 3256 20140 3296
rect 20180 3256 20181 3296
rect 20139 3247 20181 3256
rect 20236 2876 20276 3919
rect 20428 3716 20468 4936
rect 20524 4976 20564 4987
rect 20524 4901 20564 4936
rect 20620 4976 20660 4985
rect 20523 4892 20565 4901
rect 20523 4852 20524 4892
rect 20564 4852 20565 4892
rect 20523 4843 20565 4852
rect 20620 4565 20660 4936
rect 20716 4976 20756 4985
rect 20619 4556 20661 4565
rect 20619 4516 20620 4556
rect 20660 4516 20661 4556
rect 20619 4507 20661 4516
rect 20716 4388 20756 4936
rect 20620 4348 20756 4388
rect 20620 3968 20660 4348
rect 20812 4304 20852 5104
rect 20908 4901 20948 5179
rect 21388 4985 21428 5356
rect 21484 5153 21524 5238
rect 21483 5144 21525 5153
rect 21483 5104 21484 5144
rect 21524 5104 21525 5144
rect 21483 5095 21525 5104
rect 21580 5060 21620 5069
rect 21387 4976 21429 4985
rect 21387 4936 21388 4976
rect 21428 4936 21429 4976
rect 21387 4927 21429 4936
rect 20907 4892 20949 4901
rect 20907 4852 20908 4892
rect 20948 4852 21044 4892
rect 20907 4843 20949 4852
rect 20907 4472 20949 4481
rect 20907 4432 20908 4472
rect 20948 4432 20949 4472
rect 20907 4423 20949 4432
rect 20908 4313 20948 4423
rect 20524 3928 20620 3968
rect 20524 3725 20564 3928
rect 20620 3919 20660 3928
rect 20716 4264 20852 4304
rect 20907 4304 20949 4313
rect 20907 4264 20908 4304
rect 20948 4264 20949 4304
rect 20619 3800 20661 3809
rect 20619 3760 20620 3800
rect 20660 3760 20661 3800
rect 20619 3751 20661 3760
rect 19948 2575 19988 2584
rect 20044 2836 20276 2876
rect 20332 3676 20468 3716
rect 20523 3716 20565 3725
rect 20523 3676 20524 3716
rect 20564 3676 20565 3716
rect 20332 3464 20372 3676
rect 20523 3667 20565 3676
rect 20620 3632 20660 3751
rect 20620 3583 20660 3592
rect 18603 2540 18645 2549
rect 18603 2500 18604 2540
rect 18644 2500 18645 2540
rect 18603 2491 18645 2500
rect 18604 2406 18644 2491
rect 19180 2456 19220 2465
rect 18988 1952 19028 1961
rect 19028 1912 19124 1952
rect 18988 1903 19028 1912
rect 18260 1744 18548 1784
rect 18795 1784 18837 1793
rect 18795 1744 18796 1784
rect 18836 1744 18837 1784
rect 18220 1735 18260 1744
rect 18795 1735 18837 1744
rect 17451 1700 17493 1709
rect 17451 1660 17452 1700
rect 17492 1660 17493 1700
rect 17451 1651 17493 1660
rect 17356 1147 17396 1156
rect 17259 1112 17301 1121
rect 17259 1072 17260 1112
rect 17300 1072 17301 1112
rect 17259 1063 17301 1072
rect 17452 1112 17492 1651
rect 18796 1650 18836 1735
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 17452 1063 17492 1072
rect 17260 978 17300 1063
rect 19084 944 19124 1912
rect 19180 1112 19220 2416
rect 19371 2456 19413 2465
rect 19371 2416 19372 2456
rect 19412 2416 19413 2456
rect 19371 2407 19413 2416
rect 19660 2456 19700 2575
rect 19852 2490 19892 2575
rect 20044 2456 20084 2836
rect 20140 2633 20180 2718
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 20236 2624 20276 2633
rect 20332 2624 20372 3424
rect 20427 3464 20469 3473
rect 20427 3424 20428 3464
rect 20468 3424 20469 3464
rect 20427 3415 20469 3424
rect 20524 3464 20564 3473
rect 20428 3330 20468 3415
rect 20428 2876 20468 2885
rect 20524 2876 20564 3424
rect 20468 2836 20564 2876
rect 20428 2827 20468 2836
rect 20428 2633 20468 2718
rect 20619 2708 20661 2717
rect 20619 2668 20620 2708
rect 20660 2668 20661 2708
rect 20619 2659 20661 2668
rect 20276 2584 20372 2624
rect 20427 2624 20469 2633
rect 20427 2584 20428 2624
rect 20468 2584 20469 2624
rect 20236 2575 20276 2584
rect 20427 2575 20469 2584
rect 20620 2574 20660 2659
rect 20235 2456 20277 2465
rect 20044 2416 20236 2456
rect 20276 2416 20277 2456
rect 19660 2407 19700 2416
rect 20235 2407 20277 2416
rect 19372 2120 19412 2407
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 19372 2080 19508 2120
rect 19372 1952 19412 1961
rect 19372 1793 19412 1912
rect 19371 1784 19413 1793
rect 19371 1744 19372 1784
rect 19412 1744 19413 1784
rect 19371 1735 19413 1744
rect 19276 1112 19316 1121
rect 19180 1072 19276 1112
rect 19276 1063 19316 1072
rect 19468 1112 19508 2080
rect 20236 1952 20276 2407
rect 20236 1903 20276 1912
rect 20716 1121 20756 4264
rect 20907 4255 20949 4264
rect 20811 4136 20853 4145
rect 20811 4096 20812 4136
rect 20852 4096 20853 4136
rect 20811 4087 20853 4096
rect 20908 4136 20948 4255
rect 20908 4087 20948 4096
rect 20812 4002 20852 4087
rect 21004 3968 21044 4852
rect 21099 4556 21141 4565
rect 21099 4516 21100 4556
rect 21140 4516 21141 4556
rect 21099 4507 21141 4516
rect 20908 3928 21044 3968
rect 20908 3557 20948 3928
rect 21100 3641 21140 4507
rect 21195 4388 21237 4397
rect 21195 4348 21196 4388
rect 21236 4348 21237 4388
rect 21195 4339 21237 4348
rect 21099 3632 21141 3641
rect 21099 3592 21100 3632
rect 21140 3592 21141 3632
rect 21099 3583 21141 3592
rect 20907 3548 20949 3557
rect 20907 3508 20908 3548
rect 20948 3508 20949 3548
rect 20907 3499 20949 3508
rect 20812 3464 20852 3473
rect 20812 3305 20852 3424
rect 20908 3464 20948 3499
rect 20811 3296 20853 3305
rect 20811 3256 20812 3296
rect 20852 3256 20853 3296
rect 20811 3247 20853 3256
rect 20812 3053 20852 3247
rect 20811 3044 20853 3053
rect 20811 3004 20812 3044
rect 20852 3004 20853 3044
rect 20811 2995 20853 3004
rect 20908 2969 20948 3424
rect 21004 3464 21044 3475
rect 21004 3389 21044 3424
rect 21099 3464 21141 3473
rect 21099 3424 21100 3464
rect 21140 3424 21141 3464
rect 21099 3415 21141 3424
rect 21003 3380 21045 3389
rect 21003 3340 21004 3380
rect 21044 3340 21045 3380
rect 21003 3331 21045 3340
rect 21100 3330 21140 3415
rect 20907 2960 20949 2969
rect 20907 2920 20908 2960
rect 20948 2920 20949 2960
rect 20907 2911 20949 2920
rect 21196 2633 21236 4339
rect 21580 3809 21620 5020
rect 21676 4985 21716 5066
rect 21670 4976 21716 4985
rect 21670 4936 21671 4976
rect 21670 4927 21716 4936
rect 21771 4976 21813 4985
rect 21771 4936 21772 4976
rect 21812 4936 21813 4976
rect 21771 4927 21813 4936
rect 21772 4842 21812 4927
rect 21676 4724 21716 4733
rect 21716 4684 22004 4724
rect 21676 4675 21716 4684
rect 21579 3800 21621 3809
rect 21579 3760 21580 3800
rect 21620 3760 21621 3800
rect 21579 3751 21621 3760
rect 21387 3548 21429 3557
rect 21387 3508 21388 3548
rect 21428 3508 21429 3548
rect 21387 3499 21429 3508
rect 21292 3464 21332 3473
rect 21292 3305 21332 3424
rect 21388 3464 21428 3499
rect 21388 3413 21428 3424
rect 21484 3464 21524 3475
rect 21484 3389 21524 3424
rect 21580 3464 21620 3473
rect 21483 3380 21525 3389
rect 21483 3340 21484 3380
rect 21524 3340 21525 3380
rect 21483 3331 21525 3340
rect 21291 3296 21333 3305
rect 21291 3256 21292 3296
rect 21332 3256 21333 3296
rect 21291 3247 21333 3256
rect 21291 3128 21333 3137
rect 21291 3088 21292 3128
rect 21332 3088 21333 3128
rect 21291 3079 21333 3088
rect 21195 2624 21237 2633
rect 21195 2584 21196 2624
rect 21236 2584 21237 2624
rect 21195 2575 21237 2584
rect 21292 2624 21332 3079
rect 21292 2540 21332 2584
rect 21292 2500 21524 2540
rect 21484 1952 21524 2500
rect 21580 1961 21620 3424
rect 21675 3464 21717 3473
rect 21675 3424 21676 3464
rect 21716 3424 21717 3464
rect 21675 3415 21717 3424
rect 21484 1903 21524 1912
rect 21579 1952 21621 1961
rect 21579 1912 21580 1952
rect 21620 1912 21621 1952
rect 21579 1903 21621 1912
rect 21676 1952 21716 3415
rect 21772 3212 21812 3221
rect 21772 2624 21812 3172
rect 21772 2575 21812 2584
rect 21771 2120 21813 2129
rect 21771 2080 21772 2120
rect 21812 2080 21813 2120
rect 21771 2071 21813 2080
rect 21772 1986 21812 2071
rect 21676 1903 21716 1912
rect 21964 1952 22004 4684
rect 22060 4061 22100 5356
rect 22732 4976 22772 5767
rect 23020 5648 23060 6187
rect 23308 5984 23348 6280
rect 23404 6270 23444 6355
rect 23692 6329 23732 6448
rect 23788 6404 23828 6607
rect 23883 6488 23925 6497
rect 23883 6448 23884 6488
rect 23924 6448 23925 6488
rect 23883 6439 23925 6448
rect 24076 6488 24116 6497
rect 24172 6488 24212 7279
rect 24268 6824 24308 7456
rect 24364 7160 24404 8203
rect 24460 8000 24500 9472
rect 24555 9512 24597 9521
rect 24555 9472 24556 9512
rect 24596 9472 24597 9512
rect 24555 9463 24597 9472
rect 24556 8672 24596 9463
rect 24652 9269 24692 9640
rect 24651 9260 24693 9269
rect 24651 9220 24652 9260
rect 24692 9220 24693 9260
rect 24651 9211 24693 9220
rect 24748 9008 24788 10387
rect 25036 10268 25076 10816
rect 25132 10772 25172 10781
rect 25172 10732 25460 10772
rect 25132 10723 25172 10732
rect 25036 10219 25076 10228
rect 24843 10184 24885 10193
rect 24843 10144 24844 10184
rect 24884 10144 24885 10184
rect 24843 10135 24885 10144
rect 25132 10184 25172 10193
rect 24844 9764 24884 10135
rect 25132 9857 25172 10144
rect 25420 10184 25460 10732
rect 25612 10361 25652 12244
rect 25900 11360 25940 13756
rect 26188 13208 26228 13217
rect 26091 13124 26133 13133
rect 26091 13084 26092 13124
rect 26132 13084 26133 13124
rect 26091 13075 26133 13084
rect 26092 12990 26132 13075
rect 26188 12293 26228 13168
rect 26284 12536 26324 15268
rect 26380 14552 26420 14561
rect 26420 14512 26516 14552
rect 26380 14503 26420 14512
rect 26476 14048 26516 14512
rect 26668 14132 26708 17620
rect 26763 16316 26805 16325
rect 26763 16276 26764 16316
rect 26804 16276 26805 16316
rect 26763 16267 26805 16276
rect 26764 15317 26804 16267
rect 26859 16064 26901 16073
rect 26859 16024 26860 16064
rect 26900 16024 26901 16064
rect 26859 16015 26901 16024
rect 26860 15737 26900 16015
rect 26859 15728 26901 15737
rect 26859 15688 26860 15728
rect 26900 15688 26901 15728
rect 26859 15679 26901 15688
rect 26860 15560 26900 15679
rect 26860 15511 26900 15520
rect 26763 15308 26805 15317
rect 26763 15268 26764 15308
rect 26804 15268 26805 15308
rect 26763 15259 26805 15268
rect 26764 14720 26804 15259
rect 26956 14897 26996 19048
rect 27340 19039 27380 19048
rect 27532 18500 27572 19216
rect 28108 19088 28148 19097
rect 27820 19048 28108 19088
rect 27723 18584 27765 18593
rect 27723 18544 27724 18584
rect 27764 18544 27765 18584
rect 27723 18535 27765 18544
rect 27532 17744 27572 18460
rect 27724 18416 27764 18535
rect 27724 18367 27764 18376
rect 27723 18248 27765 18257
rect 27723 18208 27724 18248
rect 27764 18208 27765 18248
rect 27723 18199 27765 18208
rect 27532 17695 27572 17704
rect 27339 17240 27381 17249
rect 27339 17200 27340 17240
rect 27380 17200 27381 17240
rect 27339 17191 27381 17200
rect 27531 17240 27573 17249
rect 27531 17200 27532 17240
rect 27572 17200 27573 17240
rect 27531 17191 27573 17200
rect 27244 16400 27284 16409
rect 27147 16316 27189 16325
rect 27147 16276 27148 16316
rect 27188 16276 27189 16316
rect 27147 16267 27189 16276
rect 27052 16232 27092 16241
rect 27052 15653 27092 16192
rect 27148 16182 27188 16267
rect 27244 16073 27284 16360
rect 27340 16325 27380 17191
rect 27532 17072 27572 17191
rect 27724 17081 27764 18199
rect 27532 17023 27572 17032
rect 27723 17072 27765 17081
rect 27723 17032 27724 17072
rect 27764 17032 27765 17072
rect 27723 17023 27765 17032
rect 27628 16988 27668 16997
rect 27628 16829 27668 16948
rect 27820 16988 27860 19048
rect 28108 19039 28148 19048
rect 28204 18920 28244 19804
rect 28300 19256 28340 20056
rect 28588 20047 28628 20056
rect 28300 19207 28340 19216
rect 28588 19256 28628 19265
rect 28588 19181 28628 19216
rect 28587 19172 28629 19181
rect 28587 19132 28588 19172
rect 28628 19132 28629 19172
rect 28587 19123 28629 19132
rect 28588 18920 28628 19123
rect 28012 18880 28244 18920
rect 28492 18880 28628 18920
rect 27915 18752 27957 18761
rect 27915 18712 27916 18752
rect 27956 18712 27957 18752
rect 27915 18703 27957 18712
rect 27916 18618 27956 18703
rect 28012 18584 28052 18880
rect 28492 18761 28532 18880
rect 28491 18752 28533 18761
rect 28684 18752 28724 20719
rect 29068 20264 29108 20273
rect 29068 20180 29108 20224
rect 30028 20180 30068 20896
rect 28972 20140 29108 20180
rect 29932 20140 30068 20180
rect 28780 19256 28820 19265
rect 28972 19256 29012 20140
rect 29164 20096 29204 20105
rect 29164 19265 29204 20056
rect 29548 20096 29588 20105
rect 29356 19844 29396 19853
rect 28820 19216 29012 19256
rect 29163 19256 29205 19265
rect 29163 19216 29164 19256
rect 29204 19216 29205 19256
rect 28780 19013 28820 19216
rect 29163 19207 29205 19216
rect 29164 19122 29204 19207
rect 29259 19088 29301 19097
rect 29259 19048 29260 19088
rect 29300 19048 29301 19088
rect 29259 19039 29301 19048
rect 28779 19004 28821 19013
rect 28779 18964 28780 19004
rect 28820 18964 28821 19004
rect 28779 18955 28821 18964
rect 29260 18954 29300 19039
rect 28491 18712 28492 18752
rect 28532 18712 28533 18752
rect 28491 18703 28533 18712
rect 28588 18712 28724 18752
rect 28203 18668 28245 18677
rect 28203 18628 28204 18668
rect 28244 18628 28245 18668
rect 28203 18619 28245 18628
rect 28012 18257 28052 18544
rect 28107 18584 28149 18593
rect 28107 18544 28108 18584
rect 28148 18544 28149 18584
rect 28107 18535 28149 18544
rect 28011 18248 28053 18257
rect 28011 18208 28012 18248
rect 28052 18208 28053 18248
rect 28011 18199 28053 18208
rect 28012 17921 28052 18006
rect 28011 17912 28053 17921
rect 28011 17872 28012 17912
rect 28052 17872 28053 17912
rect 28011 17863 28053 17872
rect 28011 17744 28053 17753
rect 28011 17704 28012 17744
rect 28052 17704 28053 17744
rect 28011 17695 28053 17704
rect 28012 17610 28052 17695
rect 28108 17408 28148 18535
rect 28204 18534 28244 18619
rect 28395 18500 28437 18509
rect 28395 18460 28396 18500
rect 28436 18460 28437 18500
rect 28395 18451 28437 18460
rect 28204 17585 28244 17670
rect 28203 17576 28245 17585
rect 28203 17536 28204 17576
rect 28244 17536 28245 17576
rect 28203 17527 28245 17536
rect 28108 17368 28340 17408
rect 28203 17240 28245 17249
rect 28203 17200 28204 17240
rect 28244 17200 28245 17240
rect 28108 17165 28148 17196
rect 28203 17191 28245 17200
rect 28107 17156 28149 17165
rect 28107 17116 28108 17156
rect 28148 17116 28149 17156
rect 28107 17107 28149 17116
rect 27915 17072 27957 17081
rect 27915 17032 27916 17072
rect 27956 17032 27957 17072
rect 27915 17023 27957 17032
rect 28108 17072 28148 17107
rect 27820 16939 27860 16948
rect 27724 16904 27764 16913
rect 27435 16820 27477 16829
rect 27435 16780 27436 16820
rect 27476 16780 27477 16820
rect 27435 16771 27477 16780
rect 27627 16820 27669 16829
rect 27627 16780 27628 16820
rect 27668 16780 27669 16820
rect 27627 16771 27669 16780
rect 27339 16316 27381 16325
rect 27339 16276 27340 16316
rect 27380 16276 27381 16316
rect 27339 16267 27381 16276
rect 27243 16064 27285 16073
rect 27243 16024 27244 16064
rect 27284 16024 27285 16064
rect 27243 16015 27285 16024
rect 27340 15896 27380 16267
rect 27436 16232 27476 16771
rect 27724 16493 27764 16864
rect 27916 16820 27956 17023
rect 28108 16829 28148 17032
rect 28204 17072 28244 17191
rect 28204 17023 28244 17032
rect 28300 17072 28340 17368
rect 28396 17333 28436 18451
rect 28492 18332 28532 18341
rect 28492 17921 28532 18292
rect 28491 17912 28533 17921
rect 28491 17872 28492 17912
rect 28532 17872 28533 17912
rect 28491 17863 28533 17872
rect 28588 17417 28628 18712
rect 28684 18584 28724 18595
rect 28684 18509 28724 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 28779 18535 28821 18544
rect 29356 18584 29396 19804
rect 29548 19601 29588 20056
rect 29932 20096 29972 20140
rect 29932 20047 29972 20056
rect 30220 19760 30260 21559
rect 30508 20777 30548 25432
rect 30604 21533 30644 25843
rect 31084 25229 31124 28624
rect 31468 28580 31508 29875
rect 31564 29345 31604 30640
rect 31563 29336 31605 29345
rect 31563 29296 31564 29336
rect 31604 29296 31605 29336
rect 31563 29287 31605 29296
rect 31660 29093 31700 31312
rect 31948 31352 31988 31361
rect 31755 30680 31797 30689
rect 31755 30640 31756 30680
rect 31796 30640 31797 30680
rect 31755 30631 31797 30640
rect 31948 30680 31988 31312
rect 32236 30848 32276 31471
rect 32236 30799 32276 30808
rect 31756 30546 31796 30631
rect 31948 30437 31988 30640
rect 32044 30680 32084 30689
rect 32332 30680 32372 31648
rect 32428 31604 32468 32152
rect 32811 32152 32812 32192
rect 32852 32152 32853 32192
rect 32811 32143 32853 32152
rect 32908 32192 32948 32201
rect 33100 32192 33140 32656
rect 33196 32360 33236 32815
rect 33196 32311 33236 32320
rect 32948 32152 33044 32192
rect 32908 32143 32948 32152
rect 32428 31555 32468 31564
rect 32620 32108 32660 32117
rect 32620 31529 32660 32068
rect 32812 32058 32852 32143
rect 32619 31520 32661 31529
rect 32619 31480 32620 31520
rect 32660 31480 32661 31520
rect 32619 31471 32661 31480
rect 32907 31520 32949 31529
rect 32907 31480 32908 31520
rect 32948 31480 32949 31520
rect 32907 31471 32949 31480
rect 32908 31352 32948 31471
rect 32908 31303 32948 31312
rect 33004 30773 33044 32152
rect 33100 32143 33140 32152
rect 33292 31940 33332 32899
rect 33484 32201 33524 32908
rect 33676 32898 33716 32983
rect 33483 32192 33525 32201
rect 33483 32152 33484 32192
rect 33524 32152 33525 32192
rect 33483 32143 33525 32152
rect 33772 32192 33812 33067
rect 34348 32982 34388 33067
rect 33868 32873 33908 32958
rect 34155 32948 34197 32957
rect 34155 32908 34156 32948
rect 34196 32908 34197 32948
rect 34155 32899 34197 32908
rect 33867 32864 33909 32873
rect 33867 32824 33868 32864
rect 33908 32824 33909 32864
rect 33867 32815 33909 32824
rect 33964 32864 34004 32873
rect 33964 32360 34004 32824
rect 34156 32864 34196 32899
rect 34156 32813 34196 32824
rect 35020 32864 35060 34168
rect 35404 34168 35692 34208
rect 35404 33788 35444 34168
rect 35692 34159 35732 34168
rect 35404 33739 35444 33748
rect 35212 33704 35252 33713
rect 35116 33452 35156 33461
rect 35116 32873 35156 33412
rect 35212 33116 35252 33664
rect 35788 33704 35828 34504
rect 37036 34504 37652 34544
rect 36363 34376 36405 34385
rect 36363 34336 36364 34376
rect 36404 34336 36405 34376
rect 36363 34327 36405 34336
rect 36556 34376 36596 34385
rect 36364 34242 36404 34327
rect 35788 33655 35828 33664
rect 35883 33368 35925 33377
rect 35883 33328 35884 33368
rect 35924 33328 35925 33368
rect 35883 33319 35925 33328
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 33964 32320 34868 32360
rect 33772 32143 33812 32152
rect 33196 31900 33332 31940
rect 33868 31940 33908 31949
rect 33196 31613 33236 31900
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 33195 31604 33237 31613
rect 33195 31564 33196 31604
rect 33236 31564 33237 31604
rect 33195 31555 33237 31564
rect 33387 31604 33429 31613
rect 33387 31564 33388 31604
rect 33428 31564 33429 31604
rect 33387 31555 33429 31564
rect 33388 31352 33428 31555
rect 33292 30848 33332 30857
rect 33388 30848 33428 31312
rect 33332 30808 33428 30848
rect 33772 31184 33812 31193
rect 33292 30799 33332 30808
rect 33003 30764 33045 30773
rect 33003 30724 33004 30764
rect 33044 30724 33045 30764
rect 33003 30715 33045 30724
rect 32084 30640 32276 30680
rect 32044 30631 32084 30640
rect 31756 30428 31796 30437
rect 31756 29252 31796 30388
rect 31947 30428 31989 30437
rect 31947 30388 31948 30428
rect 31988 30388 31989 30428
rect 31947 30379 31989 30388
rect 32236 30176 32276 30640
rect 32332 30605 32372 30640
rect 32428 30680 32468 30689
rect 32331 30596 32373 30605
rect 32331 30556 32332 30596
rect 32372 30556 32373 30596
rect 32331 30547 32373 30556
rect 32236 30136 32372 30176
rect 32235 30008 32277 30017
rect 32235 29968 32236 30008
rect 32276 29968 32277 30008
rect 32235 29959 32277 29968
rect 31852 29672 31892 29681
rect 31852 29513 31892 29632
rect 32043 29672 32085 29681
rect 32043 29632 32044 29672
rect 32084 29632 32085 29672
rect 32043 29623 32085 29632
rect 32044 29538 32084 29623
rect 31851 29504 31893 29513
rect 31851 29464 31852 29504
rect 31892 29464 31893 29504
rect 31851 29455 31893 29464
rect 31852 29252 31892 29261
rect 31756 29212 31852 29252
rect 31852 29203 31892 29212
rect 32236 29168 32276 29959
rect 32332 29336 32372 30136
rect 32428 29513 32468 30640
rect 32524 30680 32564 30689
rect 32524 30437 32564 30640
rect 33195 30680 33237 30689
rect 33195 30640 33196 30680
rect 33236 30640 33237 30680
rect 33195 30631 33237 30640
rect 33676 30680 33716 30689
rect 32811 30596 32853 30605
rect 32811 30556 32812 30596
rect 32852 30556 32853 30596
rect 32811 30547 32853 30556
rect 32523 30428 32565 30437
rect 32523 30388 32524 30428
rect 32564 30388 32565 30428
rect 32523 30379 32565 30388
rect 32716 29840 32756 29849
rect 32716 29513 32756 29800
rect 32812 29765 32852 30547
rect 32907 30428 32949 30437
rect 32907 30388 32908 30428
rect 32948 30388 32949 30428
rect 32907 30379 32949 30388
rect 32908 29840 32948 30379
rect 32908 29791 32948 29800
rect 33003 29840 33045 29849
rect 33003 29800 33004 29840
rect 33044 29800 33045 29840
rect 33003 29791 33045 29800
rect 33100 29840 33140 29851
rect 32811 29756 32853 29765
rect 32811 29716 32812 29756
rect 32852 29716 32853 29756
rect 32811 29707 32853 29716
rect 32427 29504 32469 29513
rect 32427 29464 32428 29504
rect 32468 29464 32469 29504
rect 32427 29455 32469 29464
rect 32715 29504 32757 29513
rect 32715 29464 32716 29504
rect 32756 29464 32757 29504
rect 32715 29455 32757 29464
rect 32332 29296 32564 29336
rect 32236 29119 32276 29128
rect 31659 29084 31701 29093
rect 31659 29044 31660 29084
rect 31700 29044 31701 29084
rect 31659 29035 31701 29044
rect 32427 28664 32469 28673
rect 32427 28624 32428 28664
rect 32468 28624 32469 28664
rect 32427 28615 32469 28624
rect 31180 28540 31508 28580
rect 31180 27665 31220 28540
rect 31563 28496 31605 28505
rect 31563 28456 31564 28496
rect 31604 28456 31605 28496
rect 31563 28447 31605 28456
rect 32235 28496 32277 28505
rect 32235 28456 32236 28496
rect 32276 28456 32277 28496
rect 32235 28447 32277 28456
rect 31275 28412 31317 28421
rect 31275 28372 31276 28412
rect 31316 28372 31317 28412
rect 31275 28363 31317 28372
rect 31276 28328 31316 28363
rect 31276 28277 31316 28288
rect 31468 28328 31508 28337
rect 31468 27749 31508 28288
rect 31564 28328 31604 28447
rect 32044 28337 32084 28422
rect 31564 28279 31604 28288
rect 31756 28328 31796 28337
rect 31948 28328 31988 28337
rect 31796 28288 31948 28328
rect 31756 28279 31796 28288
rect 31948 28279 31988 28288
rect 32043 28328 32085 28337
rect 32043 28288 32044 28328
rect 32084 28288 32085 28328
rect 32043 28279 32085 28288
rect 32140 28328 32180 28337
rect 31659 28160 31701 28169
rect 31659 28120 31660 28160
rect 31700 28120 31701 28160
rect 31659 28111 31701 28120
rect 31660 28026 31700 28111
rect 31275 27740 31317 27749
rect 31275 27700 31276 27740
rect 31316 27700 31317 27740
rect 31275 27691 31317 27700
rect 31467 27740 31509 27749
rect 31467 27700 31468 27740
rect 31508 27700 31509 27740
rect 31467 27691 31509 27700
rect 31179 27656 31221 27665
rect 31179 27616 31180 27656
rect 31220 27616 31221 27656
rect 31179 27607 31221 27616
rect 31276 27606 31316 27691
rect 31372 27656 31412 27665
rect 31372 27413 31412 27616
rect 31659 27656 31701 27665
rect 31659 27616 31660 27656
rect 31700 27616 31701 27656
rect 31659 27607 31701 27616
rect 32043 27656 32085 27665
rect 32043 27616 32044 27656
rect 32084 27616 32085 27656
rect 32043 27607 32085 27616
rect 31660 27522 31700 27607
rect 31371 27404 31413 27413
rect 31371 27364 31372 27404
rect 31412 27364 31413 27404
rect 31371 27355 31413 27364
rect 31948 27404 31988 27413
rect 31180 26816 31220 26825
rect 31180 26237 31220 26776
rect 31276 26816 31316 26825
rect 31276 26489 31316 26776
rect 31467 26816 31509 26825
rect 31467 26776 31468 26816
rect 31508 26776 31509 26816
rect 31467 26767 31509 26776
rect 31852 26816 31892 26825
rect 31948 26816 31988 27364
rect 31892 26776 31988 26816
rect 31852 26767 31892 26776
rect 31275 26480 31317 26489
rect 31468 26480 31508 26767
rect 31275 26440 31276 26480
rect 31316 26440 31317 26480
rect 31275 26431 31317 26440
rect 31372 26440 31508 26480
rect 31755 26480 31797 26489
rect 31755 26440 31756 26480
rect 31796 26440 31797 26480
rect 31179 26228 31221 26237
rect 31179 26188 31180 26228
rect 31220 26188 31221 26228
rect 31372 26228 31412 26440
rect 31755 26431 31797 26440
rect 31372 26188 31508 26228
rect 31179 26179 31221 26188
rect 31180 26133 31220 26179
rect 31372 26133 31412 26142
rect 31180 26093 31372 26133
rect 31180 25817 31220 26093
rect 31372 26084 31412 26093
rect 31372 25976 31412 25985
rect 31468 25976 31508 26188
rect 31412 25936 31508 25976
rect 31564 26144 31604 26153
rect 31372 25927 31412 25936
rect 31564 25901 31604 26104
rect 31660 26144 31700 26153
rect 31756 26144 31796 26431
rect 31700 26104 31796 26144
rect 31852 26144 31892 26153
rect 31660 26095 31700 26104
rect 31563 25892 31605 25901
rect 31563 25852 31564 25892
rect 31604 25852 31605 25892
rect 31563 25843 31605 25852
rect 31179 25808 31221 25817
rect 31179 25768 31180 25808
rect 31220 25768 31221 25808
rect 31179 25759 31221 25768
rect 31852 25397 31892 26104
rect 32044 25556 32084 27607
rect 32140 27077 32180 28288
rect 32236 28328 32276 28447
rect 32236 28253 32276 28288
rect 32428 28328 32468 28615
rect 32524 28580 32564 29296
rect 32524 28531 32564 28540
rect 32812 28337 32852 29707
rect 33004 29336 33044 29791
rect 33100 29765 33140 29800
rect 33196 29840 33236 30631
rect 33676 30521 33716 30640
rect 33772 30605 33812 31144
rect 33868 30689 33908 31900
rect 34060 30857 34100 32320
rect 34155 32192 34197 32201
rect 34155 32152 34156 32192
rect 34196 32152 34197 32192
rect 34155 32143 34197 32152
rect 34539 32192 34581 32201
rect 34539 32152 34540 32192
rect 34580 32152 34581 32192
rect 34539 32143 34581 32152
rect 34156 31529 34196 32143
rect 34540 32058 34580 32143
rect 34252 32024 34292 32033
rect 34252 31688 34292 31984
rect 34828 32024 34868 32320
rect 35020 32285 35060 32824
rect 35115 32864 35157 32873
rect 35115 32824 35116 32864
rect 35156 32824 35157 32864
rect 35115 32815 35157 32824
rect 35212 32705 35252 33076
rect 35884 32864 35924 33319
rect 36556 33284 36596 34336
rect 36651 34376 36693 34385
rect 36651 34336 36652 34376
rect 36692 34336 36693 34376
rect 36651 34327 36693 34336
rect 36748 34376 36788 34385
rect 36652 34242 36692 34327
rect 36651 33704 36693 33713
rect 36651 33664 36652 33704
rect 36692 33664 36693 33704
rect 36651 33655 36693 33664
rect 36652 33570 36692 33655
rect 36364 33244 36596 33284
rect 35979 33032 36021 33041
rect 35979 32992 35980 33032
rect 36020 32992 36021 33032
rect 35979 32983 36021 32992
rect 36267 33032 36309 33041
rect 36364 33032 36404 33244
rect 36267 32992 36268 33032
rect 36308 32992 36404 33032
rect 36460 33032 36500 33041
rect 36500 32992 36692 33032
rect 36267 32983 36309 32992
rect 36460 32983 36500 32992
rect 35884 32815 35924 32824
rect 35211 32696 35253 32705
rect 35211 32656 35212 32696
rect 35252 32656 35253 32696
rect 35211 32647 35253 32656
rect 35787 32360 35829 32369
rect 35787 32320 35788 32360
rect 35828 32320 35829 32360
rect 35787 32311 35829 32320
rect 35019 32276 35061 32285
rect 35019 32236 35020 32276
rect 35060 32236 35061 32276
rect 35019 32227 35061 32236
rect 35788 32226 35828 32311
rect 35211 32192 35253 32201
rect 35211 32152 35212 32192
rect 35252 32152 35253 32192
rect 35211 32143 35253 32152
rect 35691 32192 35733 32201
rect 35691 32152 35692 32192
rect 35732 32152 35733 32192
rect 35691 32143 35733 32152
rect 35980 32192 36020 32983
rect 36172 32864 36212 32873
rect 36172 32369 36212 32824
rect 36268 32864 36308 32983
rect 36268 32815 36308 32824
rect 36460 32864 36500 32873
rect 36171 32360 36213 32369
rect 36171 32320 36172 32360
rect 36212 32320 36213 32360
rect 36171 32311 36213 32320
rect 36268 32360 36308 32369
rect 36460 32360 36500 32824
rect 36652 32864 36692 32992
rect 36652 32815 36692 32824
rect 36748 32780 36788 34336
rect 37036 34376 37076 34504
rect 37036 34327 37076 34336
rect 37228 34376 37268 34385
rect 37132 34292 37172 34301
rect 36844 34208 36884 34217
rect 36844 32957 36884 34168
rect 36843 32948 36885 32957
rect 36843 32908 36844 32948
rect 36884 32908 36885 32948
rect 36843 32899 36885 32908
rect 36748 32740 37076 32780
rect 36651 32528 36693 32537
rect 36651 32488 36652 32528
rect 36692 32488 36693 32528
rect 36651 32479 36693 32488
rect 36308 32320 36500 32360
rect 36268 32311 36308 32320
rect 36556 32285 36596 32316
rect 36555 32276 36597 32285
rect 36555 32236 36556 32276
rect 36596 32236 36597 32276
rect 36555 32227 36597 32236
rect 34828 31975 34868 31984
rect 34252 31648 34868 31688
rect 34155 31520 34197 31529
rect 34155 31480 34156 31520
rect 34196 31480 34197 31520
rect 34155 31471 34197 31480
rect 34059 30848 34101 30857
rect 34059 30808 34060 30848
rect 34100 30808 34101 30848
rect 34059 30799 34101 30808
rect 33867 30680 33909 30689
rect 33867 30640 33868 30680
rect 33908 30640 33909 30680
rect 33867 30631 33909 30640
rect 34060 30680 34100 30689
rect 34156 30680 34196 31471
rect 34732 31277 34772 31362
rect 34828 31352 34868 31648
rect 35116 31352 35156 31361
rect 34828 31312 35116 31352
rect 35116 31303 35156 31312
rect 34731 31268 34773 31277
rect 34731 31228 34732 31268
rect 34772 31228 34773 31268
rect 34731 31219 34773 31228
rect 35212 31184 35252 32143
rect 35692 32058 35732 32143
rect 35980 31856 36020 32152
rect 36076 32192 36116 32201
rect 36076 32033 36116 32152
rect 36172 32192 36212 32201
rect 36075 32024 36117 32033
rect 36075 31984 36076 32024
rect 36116 31984 36117 32024
rect 36075 31975 36117 31984
rect 35692 31816 36020 31856
rect 35595 31268 35637 31277
rect 35595 31228 35596 31268
rect 35636 31228 35637 31268
rect 35595 31219 35637 31228
rect 35116 31144 35252 31184
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 34539 30848 34581 30857
rect 34539 30808 34540 30848
rect 34580 30808 34581 30848
rect 34539 30799 34581 30808
rect 35019 30848 35061 30857
rect 35019 30808 35020 30848
rect 35060 30808 35061 30848
rect 35019 30799 35061 30808
rect 34252 30680 34292 30689
rect 34156 30640 34252 30680
rect 33771 30596 33813 30605
rect 33771 30556 33772 30596
rect 33812 30556 33813 30596
rect 33771 30547 33813 30556
rect 33675 30512 33717 30521
rect 33675 30472 33676 30512
rect 33716 30472 33717 30512
rect 33675 30463 33717 30472
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 33387 30008 33429 30017
rect 33387 29968 33388 30008
rect 33428 29968 33429 30008
rect 33387 29959 33429 29968
rect 33388 29874 33428 29959
rect 33196 29791 33236 29800
rect 33963 29840 34005 29849
rect 33963 29800 33964 29840
rect 34004 29800 34005 29840
rect 33963 29791 34005 29800
rect 33099 29756 33141 29765
rect 33099 29716 33100 29756
rect 33140 29716 33141 29756
rect 33099 29707 33141 29716
rect 33964 29706 34004 29791
rect 33004 29296 33236 29336
rect 33099 29168 33141 29177
rect 33099 29128 33100 29168
rect 33140 29128 33141 29168
rect 33099 29119 33141 29128
rect 33003 29084 33045 29093
rect 33003 29044 33004 29084
rect 33044 29044 33045 29084
rect 33003 29035 33045 29044
rect 32908 28496 32948 28505
rect 32428 28279 32468 28288
rect 32811 28328 32853 28337
rect 32811 28288 32812 28328
rect 32852 28288 32853 28328
rect 32811 28279 32853 28288
rect 32235 28244 32277 28253
rect 32235 28204 32236 28244
rect 32276 28204 32277 28244
rect 32235 28195 32277 28204
rect 32236 28164 32276 28195
rect 32619 28160 32661 28169
rect 32619 28120 32620 28160
rect 32660 28120 32661 28160
rect 32619 28111 32661 28120
rect 32620 27656 32660 28111
rect 32908 27833 32948 28456
rect 32907 27824 32949 27833
rect 32907 27784 32908 27824
rect 32948 27784 32949 27824
rect 32907 27775 32949 27784
rect 32620 27607 32660 27616
rect 32235 27488 32277 27497
rect 32235 27448 32236 27488
rect 32276 27448 32277 27488
rect 32235 27439 32277 27448
rect 32811 27488 32853 27497
rect 32811 27448 32812 27488
rect 32852 27448 32853 27488
rect 32811 27439 32853 27448
rect 32139 27068 32181 27077
rect 32139 27028 32140 27068
rect 32180 27028 32181 27068
rect 32139 27019 32181 27028
rect 32236 26816 32276 27439
rect 32812 27354 32852 27439
rect 32236 26767 32276 26776
rect 32235 26648 32277 26657
rect 32235 26608 32236 26648
rect 32276 26608 32277 26648
rect 32235 26599 32277 26608
rect 32044 25507 32084 25516
rect 31851 25388 31893 25397
rect 31851 25348 31852 25388
rect 31892 25348 31893 25388
rect 31851 25339 31893 25348
rect 32236 25313 32276 26599
rect 32811 26144 32853 26153
rect 32811 26104 32812 26144
rect 32852 26104 32853 26144
rect 33004 26144 33044 29035
rect 33100 29034 33140 29119
rect 33196 28496 33236 29296
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 33388 28496 33428 28505
rect 33196 28456 33332 28496
rect 33196 28328 33236 28339
rect 33100 28313 33140 28322
rect 33100 27413 33140 28273
rect 33196 28253 33236 28288
rect 33195 28244 33237 28253
rect 33195 28204 33196 28244
rect 33236 28204 33237 28244
rect 33195 28195 33237 28204
rect 33292 27656 33332 28456
rect 33428 28456 33620 28496
rect 33388 28447 33428 28456
rect 33388 28328 33428 28337
rect 33580 28328 33620 28456
rect 34060 28421 34100 30640
rect 34252 30631 34292 30640
rect 34540 30680 34580 30799
rect 34540 30631 34580 30640
rect 34636 30680 34676 30689
rect 34155 30512 34197 30521
rect 34155 30472 34156 30512
rect 34196 30472 34197 30512
rect 34155 30463 34197 30472
rect 34156 29000 34196 30463
rect 34636 30353 34676 30640
rect 34732 30680 34772 30691
rect 34732 30605 34772 30640
rect 34828 30680 34868 30689
rect 35020 30680 35060 30799
rect 34868 30640 34964 30680
rect 34828 30631 34868 30640
rect 34731 30596 34773 30605
rect 34731 30556 34732 30596
rect 34772 30556 34773 30596
rect 34731 30547 34773 30556
rect 34635 30344 34677 30353
rect 34635 30304 34636 30344
rect 34676 30304 34677 30344
rect 34635 30295 34677 30304
rect 34636 29840 34676 29849
rect 34252 29800 34636 29840
rect 34924 29840 34964 30640
rect 35020 30344 35060 30640
rect 35116 30680 35156 31144
rect 35596 30848 35636 31219
rect 35596 30799 35636 30808
rect 35116 30631 35156 30640
rect 35212 30680 35252 30689
rect 35212 30521 35252 30640
rect 35308 30680 35348 30689
rect 35500 30680 35540 30689
rect 35348 30640 35500 30680
rect 35308 30631 35348 30640
rect 35500 30631 35540 30640
rect 35692 30680 35732 31816
rect 36076 31520 36116 31975
rect 36172 31949 36212 32152
rect 36460 32192 36500 32203
rect 36460 32117 36500 32152
rect 36556 32192 36596 32227
rect 36459 32108 36501 32117
rect 36459 32068 36460 32108
rect 36500 32068 36501 32108
rect 36459 32059 36501 32068
rect 36171 31940 36213 31949
rect 36171 31900 36172 31940
rect 36212 31900 36213 31940
rect 36171 31891 36213 31900
rect 36172 31613 36212 31891
rect 36171 31604 36213 31613
rect 36171 31564 36172 31604
rect 36212 31564 36213 31604
rect 36171 31555 36213 31564
rect 35884 31480 36116 31520
rect 35692 30631 35732 30640
rect 35787 30680 35829 30689
rect 35787 30640 35788 30680
rect 35828 30640 35829 30680
rect 35787 30631 35829 30640
rect 35788 30546 35828 30631
rect 35211 30512 35253 30521
rect 35211 30472 35212 30512
rect 35252 30472 35253 30512
rect 35211 30463 35253 30472
rect 35020 30304 35252 30344
rect 35020 29840 35060 29849
rect 34924 29800 35020 29840
rect 34252 29336 34292 29800
rect 34636 29791 34676 29800
rect 35020 29791 35060 29800
rect 35212 29840 35252 30304
rect 35691 29924 35733 29933
rect 35691 29884 35692 29924
rect 35732 29884 35733 29924
rect 35691 29875 35733 29884
rect 35212 29791 35252 29800
rect 35308 29840 35348 29849
rect 35115 29672 35157 29681
rect 35115 29632 35116 29672
rect 35156 29632 35157 29672
rect 35115 29623 35157 29632
rect 35116 29538 35156 29623
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 34252 29287 34292 29296
rect 34443 29336 34485 29345
rect 34443 29296 34444 29336
rect 34484 29296 34485 29336
rect 34443 29287 34485 29296
rect 34444 29168 34484 29287
rect 34444 29119 34484 29128
rect 35115 29168 35157 29177
rect 35115 29128 35116 29168
rect 35156 29128 35157 29168
rect 35115 29119 35157 29128
rect 34156 28960 34388 29000
rect 34059 28412 34101 28421
rect 34059 28372 34060 28412
rect 34100 28372 34101 28412
rect 34059 28363 34101 28372
rect 33428 28288 33524 28328
rect 33388 28279 33428 28288
rect 33484 27824 33524 28288
rect 33580 28279 33620 28288
rect 33771 28328 33813 28337
rect 33771 28288 33772 28328
rect 33812 28288 33813 28328
rect 33771 28279 33813 28288
rect 33676 27824 33716 27833
rect 33484 27784 33676 27824
rect 33676 27775 33716 27784
rect 33388 27656 33428 27665
rect 33292 27616 33388 27656
rect 33388 27607 33428 27616
rect 33772 27656 33812 28279
rect 33963 28244 34005 28253
rect 33963 28204 33964 28244
rect 34004 28204 34005 28244
rect 33963 28195 34005 28204
rect 33772 27607 33812 27616
rect 33868 27656 33908 27665
rect 33292 27413 33332 27498
rect 33868 27497 33908 27616
rect 33964 27656 34004 28195
rect 33867 27488 33909 27497
rect 33867 27448 33868 27488
rect 33908 27448 33909 27488
rect 33867 27439 33909 27448
rect 33099 27404 33141 27413
rect 33099 27364 33100 27404
rect 33140 27364 33141 27404
rect 33099 27355 33141 27364
rect 33291 27404 33333 27413
rect 33291 27364 33292 27404
rect 33332 27364 33333 27404
rect 33291 27355 33333 27364
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 33867 27068 33909 27077
rect 33867 27028 33868 27068
rect 33908 27028 33909 27068
rect 33867 27019 33909 27028
rect 33100 26816 33140 26825
rect 33100 26657 33140 26776
rect 33099 26648 33141 26657
rect 33099 26608 33100 26648
rect 33140 26608 33141 26648
rect 33099 26599 33141 26608
rect 33100 26144 33140 26153
rect 33004 26104 33100 26144
rect 32811 26095 32853 26104
rect 33100 26095 33140 26104
rect 32715 25472 32757 25481
rect 32715 25432 32716 25472
rect 32756 25432 32757 25472
rect 32715 25423 32757 25432
rect 32235 25304 32277 25313
rect 32235 25264 32236 25304
rect 32276 25264 32277 25304
rect 32235 25255 32277 25264
rect 32620 25304 32660 25313
rect 31083 25220 31125 25229
rect 31083 25180 31084 25220
rect 31124 25180 31125 25220
rect 31083 25171 31125 25180
rect 31659 25220 31701 25229
rect 31659 25180 31660 25220
rect 31700 25180 31701 25220
rect 31659 25171 31701 25180
rect 31275 24800 31317 24809
rect 31275 24760 31276 24800
rect 31316 24760 31317 24800
rect 31275 24751 31317 24760
rect 31276 24666 31316 24751
rect 30796 24632 30836 24641
rect 30796 24137 30836 24592
rect 31660 24632 31700 25171
rect 31660 24583 31700 24592
rect 32139 24632 32181 24641
rect 32139 24592 32140 24632
rect 32180 24592 32181 24632
rect 32139 24583 32181 24592
rect 32140 24498 32180 24583
rect 30987 24380 31029 24389
rect 30987 24340 30988 24380
rect 31028 24340 31029 24380
rect 30987 24331 31029 24340
rect 32043 24380 32085 24389
rect 32043 24340 32044 24380
rect 32084 24340 32085 24380
rect 32043 24331 32085 24340
rect 30795 24128 30837 24137
rect 30700 24088 30796 24128
rect 30836 24088 30837 24128
rect 30700 23120 30740 24088
rect 30795 24079 30837 24088
rect 30700 23071 30740 23080
rect 30796 23960 30836 23969
rect 30796 23036 30836 23920
rect 30988 23792 31028 24331
rect 32044 24246 32084 24331
rect 31276 23969 31316 24054
rect 31275 23960 31317 23969
rect 31275 23920 31276 23960
rect 31316 23920 31317 23960
rect 31275 23911 31317 23920
rect 32139 23960 32181 23969
rect 32139 23920 32140 23960
rect 32180 23920 32181 23960
rect 32139 23911 32181 23920
rect 30988 23743 31028 23752
rect 31084 23792 31124 23801
rect 31084 23549 31124 23752
rect 31275 23792 31317 23801
rect 31275 23752 31276 23792
rect 31316 23752 31317 23792
rect 31275 23743 31317 23752
rect 32140 23792 32180 23911
rect 32140 23743 32180 23752
rect 31276 23658 31316 23743
rect 32043 23708 32085 23717
rect 32043 23668 32044 23708
rect 32084 23668 32085 23708
rect 32043 23659 32085 23668
rect 31468 23624 31508 23633
rect 31372 23584 31468 23624
rect 31083 23540 31125 23549
rect 31083 23500 31084 23540
rect 31124 23500 31125 23540
rect 31083 23491 31125 23500
rect 31084 23204 31124 23213
rect 31372 23204 31412 23584
rect 31468 23575 31508 23584
rect 31947 23372 31989 23381
rect 31947 23332 31948 23372
rect 31988 23332 31989 23372
rect 31947 23323 31989 23332
rect 31124 23164 31412 23204
rect 31084 23155 31124 23164
rect 31468 23120 31508 23129
rect 31180 23080 31468 23120
rect 31180 23036 31220 23080
rect 31468 23071 31508 23080
rect 30796 22996 31220 23036
rect 31467 22952 31509 22961
rect 31467 22912 31468 22952
rect 31508 22912 31509 22952
rect 31467 22903 31509 22912
rect 30699 22700 30741 22709
rect 30699 22660 30700 22700
rect 30740 22660 30741 22700
rect 30699 22651 30741 22660
rect 30603 21524 30645 21533
rect 30603 21484 30604 21524
rect 30644 21484 30645 21524
rect 30603 21475 30645 21484
rect 30507 20768 30549 20777
rect 30507 20728 30508 20768
rect 30548 20728 30549 20768
rect 30507 20719 30549 20728
rect 30700 20180 30740 22651
rect 31180 22280 31220 22289
rect 30987 21608 31029 21617
rect 30987 21568 30988 21608
rect 31028 21568 31029 21608
rect 30987 21559 31029 21568
rect 31084 21608 31124 21619
rect 30795 21524 30837 21533
rect 30795 21484 30796 21524
rect 30836 21484 30837 21524
rect 30795 21475 30837 21484
rect 30796 20852 30836 21475
rect 30988 21474 31028 21559
rect 31084 21533 31124 21568
rect 31083 21524 31125 21533
rect 31083 21484 31084 21524
rect 31124 21484 31125 21524
rect 31083 21475 31125 21484
rect 31180 21449 31220 22240
rect 31468 22028 31508 22903
rect 31851 22280 31893 22289
rect 31851 22240 31852 22280
rect 31892 22240 31893 22280
rect 31851 22231 31893 22240
rect 31564 22196 31604 22205
rect 31756 22196 31796 22205
rect 31604 22156 31756 22196
rect 31564 22147 31604 22156
rect 31756 22147 31796 22156
rect 31468 21988 31700 22028
rect 31563 21776 31605 21785
rect 31563 21736 31564 21776
rect 31604 21736 31605 21776
rect 31563 21727 31605 21736
rect 31276 21608 31316 21617
rect 31468 21608 31508 21617
rect 31316 21568 31468 21608
rect 31276 21559 31316 21568
rect 31468 21559 31508 21568
rect 31564 21608 31604 21727
rect 31564 21559 31604 21568
rect 31660 21608 31700 21988
rect 31660 21559 31700 21568
rect 31756 21608 31796 21619
rect 31756 21533 31796 21568
rect 31755 21524 31797 21533
rect 31755 21484 31756 21524
rect 31796 21484 31797 21524
rect 31755 21475 31797 21484
rect 31852 21449 31892 22231
rect 31179 21440 31221 21449
rect 31179 21400 31180 21440
rect 31220 21400 31221 21440
rect 31179 21391 31221 21400
rect 31276 21440 31316 21449
rect 31371 21440 31413 21449
rect 31316 21400 31372 21440
rect 31412 21400 31413 21440
rect 31276 21391 31316 21400
rect 31371 21391 31413 21400
rect 31851 21440 31893 21449
rect 31851 21400 31852 21440
rect 31892 21400 31893 21440
rect 31851 21391 31893 21400
rect 31948 20945 31988 23323
rect 31659 20936 31701 20945
rect 31659 20896 31660 20936
rect 31700 20896 31701 20936
rect 31659 20887 31701 20896
rect 31947 20936 31989 20945
rect 31947 20896 31948 20936
rect 31988 20896 31989 20936
rect 31947 20887 31989 20896
rect 30796 20803 30836 20812
rect 31660 20768 31700 20887
rect 32044 20768 32084 23659
rect 32236 23120 32276 25255
rect 32620 24809 32660 25264
rect 32619 24800 32661 24809
rect 32619 24760 32620 24800
rect 32660 24760 32661 24800
rect 32619 24751 32661 24760
rect 32716 24464 32756 25423
rect 32716 24415 32756 24424
rect 32715 23876 32757 23885
rect 32715 23836 32716 23876
rect 32756 23836 32757 23876
rect 32715 23827 32757 23836
rect 32331 23792 32373 23801
rect 32331 23752 32332 23792
rect 32372 23752 32373 23792
rect 32331 23743 32373 23752
rect 32428 23792 32468 23801
rect 32332 23658 32372 23743
rect 32332 23120 32372 23129
rect 32236 23080 32332 23120
rect 32332 23071 32372 23080
rect 32428 22541 32468 23752
rect 32524 23792 32564 23803
rect 32524 23717 32564 23752
rect 32620 23792 32660 23801
rect 32523 23708 32565 23717
rect 32523 23668 32524 23708
rect 32564 23668 32565 23708
rect 32523 23659 32565 23668
rect 32523 23456 32565 23465
rect 32523 23416 32524 23456
rect 32564 23416 32565 23456
rect 32523 23407 32565 23416
rect 32427 22532 32469 22541
rect 32332 22492 32428 22532
rect 32468 22492 32469 22532
rect 32332 21785 32372 22492
rect 32427 22483 32469 22492
rect 32427 22280 32469 22289
rect 32427 22240 32428 22280
rect 32468 22240 32469 22280
rect 32427 22231 32469 22240
rect 32428 22146 32468 22231
rect 32524 21953 32564 23407
rect 32620 22448 32660 23752
rect 32716 23465 32756 23827
rect 32812 23708 32852 26095
rect 33003 25892 33045 25901
rect 33003 25852 33004 25892
rect 33044 25852 33045 25892
rect 33003 25843 33045 25852
rect 33004 25304 33044 25843
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 33387 25472 33429 25481
rect 33387 25432 33388 25472
rect 33428 25432 33429 25472
rect 33387 25423 33429 25432
rect 33004 25255 33044 25264
rect 33388 25304 33428 25423
rect 33388 25255 33428 25264
rect 32907 24800 32949 24809
rect 32907 24760 32908 24800
rect 32948 24760 32949 24800
rect 32907 24751 32949 24760
rect 33004 24760 33236 24800
rect 32908 24632 32948 24751
rect 33004 24716 33044 24760
rect 33004 24667 33044 24676
rect 32908 23969 32948 24592
rect 33100 24632 33140 24641
rect 32907 23960 32949 23969
rect 32907 23920 32908 23960
rect 32948 23920 32949 23960
rect 32907 23911 32949 23920
rect 33004 23885 33044 23970
rect 33003 23876 33045 23885
rect 33003 23836 33004 23876
rect 33044 23836 33045 23876
rect 33003 23827 33045 23836
rect 32812 23668 33044 23708
rect 32715 23456 32757 23465
rect 32715 23416 32716 23456
rect 32756 23416 32757 23456
rect 32715 23407 32757 23416
rect 32620 22408 32852 22448
rect 32620 22280 32660 22289
rect 32523 21944 32565 21953
rect 32523 21904 32524 21944
rect 32564 21904 32565 21944
rect 32523 21895 32565 21904
rect 32331 21776 32373 21785
rect 32620 21776 32660 22240
rect 32812 22280 32852 22408
rect 32907 22364 32949 22373
rect 32907 22324 32908 22364
rect 32948 22324 32949 22364
rect 32907 22315 32949 22324
rect 32715 22196 32757 22205
rect 32715 22156 32716 22196
rect 32756 22156 32757 22196
rect 32715 22147 32757 22156
rect 32716 22062 32756 22147
rect 32812 22112 32852 22240
rect 32908 22280 32948 22315
rect 32908 22229 32948 22240
rect 32812 22072 32948 22112
rect 32715 21944 32757 21953
rect 32715 21904 32716 21944
rect 32756 21904 32757 21944
rect 32715 21895 32757 21904
rect 32331 21736 32332 21776
rect 32372 21736 32564 21776
rect 32331 21727 32373 21736
rect 32235 21608 32277 21617
rect 32235 21568 32236 21608
rect 32276 21568 32277 21608
rect 32235 21559 32277 21568
rect 32332 21608 32372 21619
rect 32139 21440 32181 21449
rect 32139 21400 32140 21440
rect 32180 21400 32181 21440
rect 32139 21391 32181 21400
rect 32140 21306 32180 21391
rect 32236 21020 32276 21559
rect 32332 21533 32372 21568
rect 32427 21608 32469 21617
rect 32427 21568 32428 21608
rect 32468 21568 32469 21608
rect 32427 21559 32469 21568
rect 32524 21608 32564 21736
rect 32620 21727 32660 21736
rect 32524 21559 32564 21568
rect 32331 21524 32373 21533
rect 32331 21484 32332 21524
rect 32372 21484 32373 21524
rect 32331 21475 32373 21484
rect 32428 21474 32468 21559
rect 32236 20971 32276 20980
rect 32332 20768 32372 20777
rect 32044 20728 32332 20768
rect 31660 20719 31700 20728
rect 32332 20719 32372 20728
rect 32716 20768 32756 21895
rect 32811 21692 32853 21701
rect 32811 21652 32812 21692
rect 32852 21652 32853 21692
rect 32811 21643 32853 21652
rect 32812 21558 32852 21643
rect 32908 21533 32948 22072
rect 32907 21524 32949 21533
rect 32907 21484 32908 21524
rect 32948 21484 32949 21524
rect 32907 21475 32949 21484
rect 32716 20719 32756 20728
rect 33004 20180 33044 23668
rect 33100 23297 33140 24592
rect 33196 24044 33236 24760
rect 33291 24632 33333 24641
rect 33291 24592 33292 24632
rect 33332 24592 33333 24632
rect 33868 24632 33908 27019
rect 33964 26312 34004 27616
rect 34060 26900 34100 28363
rect 34252 28160 34292 28169
rect 34156 27740 34196 27749
rect 34252 27740 34292 28120
rect 34196 27700 34292 27740
rect 34156 27691 34196 27700
rect 34251 27068 34293 27077
rect 34251 27028 34252 27068
rect 34292 27028 34293 27068
rect 34251 27019 34293 27028
rect 34252 26934 34292 27019
rect 34155 26900 34197 26909
rect 34060 26860 34156 26900
rect 34196 26860 34197 26900
rect 34155 26851 34197 26860
rect 33964 26272 34100 26312
rect 33963 26144 34005 26153
rect 33963 26104 33964 26144
rect 34004 26104 34005 26144
rect 33963 26095 34005 26104
rect 33964 26010 34004 26095
rect 34060 26069 34100 26272
rect 34059 26060 34101 26069
rect 34059 26020 34060 26060
rect 34100 26020 34101 26060
rect 34059 26011 34101 26020
rect 33964 24632 34004 24641
rect 33868 24592 33964 24632
rect 33291 24583 33333 24592
rect 33964 24583 34004 24592
rect 33292 24498 33332 24583
rect 34060 24464 34100 26011
rect 34156 24632 34196 26851
rect 34348 26237 34388 28960
rect 35116 28580 35156 29119
rect 35308 29009 35348 29800
rect 35692 29840 35732 29875
rect 35692 29429 35732 29800
rect 35884 29840 35924 31480
rect 35979 31352 36021 31361
rect 35979 31312 35980 31352
rect 36020 31312 36021 31352
rect 35979 31303 36021 31312
rect 35980 31218 36020 31303
rect 36363 31016 36405 31025
rect 36363 30976 36364 31016
rect 36404 30976 36405 31016
rect 36363 30967 36405 30976
rect 36075 30764 36117 30773
rect 36075 30724 36076 30764
rect 36116 30724 36117 30764
rect 36075 30715 36117 30724
rect 36076 30092 36116 30715
rect 36171 30512 36213 30521
rect 36171 30472 36172 30512
rect 36212 30472 36213 30512
rect 36171 30463 36213 30472
rect 36172 30378 36212 30463
rect 36076 30043 36116 30052
rect 35884 29791 35924 29800
rect 35788 29756 35828 29765
rect 35691 29420 35733 29429
rect 35691 29380 35692 29420
rect 35732 29380 35733 29420
rect 35691 29371 35733 29380
rect 35788 29261 35828 29716
rect 36364 29429 36404 30967
rect 36460 30680 36500 32059
rect 36556 31025 36596 32152
rect 36652 32192 36692 32479
rect 36652 32143 36692 32152
rect 36748 32192 36788 32201
rect 36939 32192 36981 32201
rect 36788 32152 36884 32192
rect 36748 32143 36788 32152
rect 36555 31016 36597 31025
rect 36555 30976 36556 31016
rect 36596 30976 36597 31016
rect 36555 30967 36597 30976
rect 36555 30848 36597 30857
rect 36555 30808 36556 30848
rect 36596 30808 36597 30848
rect 36555 30799 36597 30808
rect 36460 30631 36500 30640
rect 36556 30680 36596 30799
rect 36651 30764 36693 30773
rect 36651 30724 36652 30764
rect 36692 30724 36693 30764
rect 36651 30715 36693 30724
rect 36556 30631 36596 30640
rect 36652 30630 36692 30715
rect 36747 30680 36789 30689
rect 36747 30640 36748 30680
rect 36788 30640 36789 30680
rect 36747 30631 36789 30640
rect 36748 30546 36788 30631
rect 36555 30512 36597 30521
rect 36555 30472 36556 30512
rect 36596 30472 36597 30512
rect 36555 30463 36597 30472
rect 36363 29420 36405 29429
rect 36363 29380 36364 29420
rect 36404 29380 36405 29420
rect 36363 29371 36405 29380
rect 35787 29252 35829 29261
rect 35787 29212 35788 29252
rect 35828 29212 35829 29252
rect 35787 29203 35829 29212
rect 35691 29168 35733 29177
rect 35691 29128 35692 29168
rect 35732 29128 35733 29168
rect 35691 29119 35733 29128
rect 36556 29168 36596 30463
rect 36748 29933 36788 29964
rect 36747 29924 36789 29933
rect 36747 29884 36748 29924
rect 36788 29884 36789 29924
rect 36747 29875 36789 29884
rect 36748 29840 36788 29875
rect 36748 29345 36788 29800
rect 36747 29336 36789 29345
rect 36747 29296 36748 29336
rect 36788 29296 36789 29336
rect 36747 29287 36789 29296
rect 36556 29119 36596 29128
rect 35692 29034 35732 29119
rect 35307 29000 35349 29009
rect 35307 28960 35308 29000
rect 35348 28960 35349 29000
rect 36844 29000 36884 32152
rect 36939 32152 36940 32192
rect 36980 32152 36981 32192
rect 36939 32143 36981 32152
rect 36940 32058 36980 32143
rect 37036 31949 37076 32740
rect 37132 32537 37172 34252
rect 37131 32528 37173 32537
rect 37131 32488 37132 32528
rect 37172 32488 37173 32528
rect 37131 32479 37173 32488
rect 37228 32285 37268 34336
rect 37324 32780 37364 32789
rect 37516 32780 37556 32789
rect 37364 32740 37516 32780
rect 37324 32731 37364 32740
rect 37516 32731 37556 32740
rect 37227 32276 37269 32285
rect 37227 32236 37228 32276
rect 37268 32236 37269 32276
rect 37227 32227 37269 32236
rect 37612 32192 37652 34504
rect 37900 34504 37996 34544
rect 37803 34376 37845 34385
rect 37803 34336 37804 34376
rect 37844 34336 37845 34376
rect 37803 34327 37845 34336
rect 37804 33872 37844 34327
rect 37804 33823 37844 33832
rect 37900 32864 37940 34504
rect 37996 34495 38036 34504
rect 37995 34376 38037 34385
rect 37995 34336 37996 34376
rect 38036 34336 38037 34376
rect 37995 34327 38037 34336
rect 37996 33704 38036 34327
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 37996 33655 38036 33664
rect 38763 33704 38805 33713
rect 38763 33664 38764 33704
rect 38804 33664 38805 33704
rect 38763 33655 38805 33664
rect 38667 33452 38709 33461
rect 38667 33412 38668 33452
rect 38708 33412 38709 33452
rect 38667 33403 38709 33412
rect 38668 33318 38708 33403
rect 37900 32815 37940 32824
rect 38764 32864 38804 33655
rect 39627 33452 39669 33461
rect 39627 33412 39628 33452
rect 39668 33412 39669 33452
rect 39627 33403 39669 33412
rect 38187 32696 38229 32705
rect 38187 32656 38188 32696
rect 38228 32656 38229 32696
rect 38187 32647 38229 32656
rect 38092 32192 38132 32201
rect 37035 31940 37077 31949
rect 37035 31900 37036 31940
rect 37076 31900 37077 31940
rect 37035 31891 37077 31900
rect 36940 30680 36980 30689
rect 36940 29840 36980 30640
rect 37036 30680 37076 31891
rect 37132 31604 37172 31613
rect 37612 31604 37652 32152
rect 37172 31564 37652 31604
rect 37804 32152 38092 32192
rect 37132 31555 37172 31564
rect 37516 31184 37556 31193
rect 37556 31144 37652 31184
rect 37516 31135 37556 31144
rect 37227 30848 37269 30857
rect 37227 30808 37228 30848
rect 37268 30808 37269 30848
rect 37227 30799 37269 30808
rect 37036 30353 37076 30640
rect 37132 30680 37172 30689
rect 37035 30344 37077 30353
rect 37035 30304 37036 30344
rect 37076 30304 37077 30344
rect 37035 30295 37077 30304
rect 37132 30185 37172 30640
rect 37228 30680 37268 30799
rect 37420 30680 37460 30689
rect 37131 30176 37173 30185
rect 37131 30136 37132 30176
rect 37172 30136 37173 30176
rect 37131 30127 37173 30136
rect 37228 30008 37268 30640
rect 37132 29968 37268 30008
rect 37324 30640 37420 30680
rect 36940 29791 36980 29800
rect 37035 29840 37077 29849
rect 37035 29800 37036 29840
rect 37076 29800 37077 29840
rect 37035 29791 37077 29800
rect 37132 29840 37172 29968
rect 37324 29849 37364 30640
rect 37420 30631 37460 30640
rect 37419 29924 37461 29933
rect 37419 29884 37420 29924
rect 37460 29884 37461 29924
rect 37419 29875 37461 29884
rect 37323 29840 37365 29849
rect 37132 29791 37172 29800
rect 37228 29825 37268 29834
rect 37036 29756 37076 29791
rect 37323 29800 37324 29840
rect 37364 29800 37365 29840
rect 37323 29791 37365 29800
rect 37420 29790 37460 29875
rect 37228 29765 37268 29785
rect 37036 29705 37076 29716
rect 37227 29756 37269 29765
rect 37227 29716 37228 29756
rect 37268 29716 37269 29756
rect 37227 29707 37269 29716
rect 36939 29672 36981 29681
rect 36939 29632 36940 29672
rect 36980 29632 36981 29672
rect 36939 29623 36981 29632
rect 36940 29168 36980 29623
rect 36940 29119 36980 29128
rect 37228 29168 37268 29707
rect 37323 29336 37365 29345
rect 37323 29296 37324 29336
rect 37364 29296 37365 29336
rect 37323 29287 37365 29296
rect 37228 29119 37268 29128
rect 37324 29168 37364 29287
rect 37419 29252 37461 29261
rect 37419 29212 37420 29252
rect 37460 29212 37461 29252
rect 37419 29203 37461 29212
rect 37324 29119 37364 29128
rect 37420 29168 37460 29203
rect 37420 29117 37460 29128
rect 37515 29168 37557 29177
rect 37515 29128 37516 29168
rect 37556 29128 37557 29168
rect 37515 29119 37557 29128
rect 37516 29034 37556 29119
rect 36844 28960 36980 29000
rect 35307 28951 35349 28960
rect 35116 28531 35156 28540
rect 35691 28412 35733 28421
rect 35979 28412 36021 28421
rect 35691 28372 35692 28412
rect 35732 28372 35733 28412
rect 35691 28363 35733 28372
rect 35884 28372 35980 28412
rect 36020 28372 36021 28412
rect 34444 28328 34484 28337
rect 34444 27665 34484 28288
rect 35403 28328 35445 28337
rect 35403 28288 35404 28328
rect 35444 28288 35445 28328
rect 35403 28279 35445 28288
rect 35692 28328 35732 28363
rect 35404 28194 35444 28279
rect 35692 28277 35732 28288
rect 35884 28328 35924 28372
rect 35979 28363 36021 28372
rect 35884 28279 35924 28288
rect 36844 28328 36884 28337
rect 36172 28160 36212 28169
rect 35500 28120 36172 28160
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 34539 27824 34581 27833
rect 34539 27784 34540 27824
rect 34580 27784 34581 27824
rect 34539 27775 34581 27784
rect 34443 27656 34485 27665
rect 34443 27616 34444 27656
rect 34484 27616 34485 27656
rect 34443 27607 34485 27616
rect 34540 27656 34580 27775
rect 34540 27607 34580 27616
rect 35403 27656 35445 27665
rect 35403 27616 35404 27656
rect 35444 27616 35445 27656
rect 35403 27607 35445 27616
rect 34444 26657 34484 27607
rect 35404 27522 35444 27607
rect 34731 26900 34773 26909
rect 34731 26860 34732 26900
rect 34772 26860 34773 26900
rect 34731 26851 34773 26860
rect 34635 26816 34677 26825
rect 34635 26776 34636 26816
rect 34676 26776 34677 26816
rect 34635 26767 34677 26776
rect 34732 26816 34772 26851
rect 34636 26682 34676 26767
rect 34732 26765 34772 26776
rect 34924 26816 34964 26825
rect 35307 26816 35349 26825
rect 34964 26776 35156 26816
rect 34924 26767 34964 26776
rect 34443 26648 34485 26657
rect 34443 26608 34444 26648
rect 34484 26608 34485 26648
rect 34443 26599 34485 26608
rect 34828 26648 34868 26657
rect 34868 26608 35060 26648
rect 34828 26599 34868 26608
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34347 26228 34389 26237
rect 34347 26188 34348 26228
rect 34388 26188 34484 26228
rect 34347 26179 34389 26188
rect 34347 25892 34389 25901
rect 34347 25852 34348 25892
rect 34388 25852 34389 25892
rect 34347 25843 34389 25852
rect 34348 25758 34388 25843
rect 34251 25304 34293 25313
rect 34251 25264 34252 25304
rect 34292 25264 34293 25304
rect 34251 25255 34293 25264
rect 34252 25170 34292 25255
rect 34252 24632 34292 24641
rect 34156 24592 34252 24632
rect 33868 24424 34100 24464
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 33196 24004 33620 24044
rect 33483 23876 33525 23885
rect 33483 23836 33484 23876
rect 33524 23836 33525 23876
rect 33483 23827 33525 23836
rect 33195 23792 33237 23801
rect 33195 23752 33196 23792
rect 33236 23752 33237 23792
rect 33195 23743 33237 23752
rect 33388 23792 33428 23801
rect 33196 23624 33236 23743
rect 33196 23575 33236 23584
rect 33099 23288 33141 23297
rect 33099 23248 33100 23288
rect 33140 23248 33141 23288
rect 33099 23239 33141 23248
rect 33388 22868 33428 23752
rect 33484 23792 33524 23827
rect 33484 23741 33524 23752
rect 33580 23792 33620 24004
rect 33580 23743 33620 23752
rect 33675 23792 33717 23801
rect 33675 23752 33676 23792
rect 33716 23752 33717 23792
rect 33675 23743 33717 23752
rect 33868 23792 33908 24424
rect 34059 24212 34101 24221
rect 34059 24172 34060 24212
rect 34100 24172 34101 24212
rect 34059 24163 34101 24172
rect 33676 23658 33716 23743
rect 33675 23540 33717 23549
rect 33675 23500 33676 23540
rect 33716 23500 33717 23540
rect 33675 23491 33717 23500
rect 33483 23288 33525 23297
rect 33483 23248 33484 23288
rect 33524 23248 33525 23288
rect 33483 23239 33525 23248
rect 33676 23288 33716 23491
rect 33868 23465 33908 23752
rect 33964 23792 34004 23801
rect 33867 23456 33909 23465
rect 33867 23416 33868 23456
rect 33908 23416 33909 23456
rect 33867 23407 33909 23416
rect 33964 23381 34004 23752
rect 34060 23792 34100 24163
rect 34252 24137 34292 24592
rect 34444 24221 34484 26188
rect 35020 26144 35060 26608
rect 35116 26489 35156 26776
rect 35307 26776 35308 26816
rect 35348 26776 35349 26816
rect 35307 26767 35349 26776
rect 35404 26816 35444 26825
rect 35500 26816 35540 28120
rect 36172 28111 36212 28120
rect 35979 27740 36021 27749
rect 35979 27700 35980 27740
rect 36020 27700 36021 27740
rect 35979 27691 36021 27700
rect 35595 27068 35637 27077
rect 35595 27028 35596 27068
rect 35636 27028 35637 27068
rect 35595 27019 35637 27028
rect 35444 26776 35540 26816
rect 35596 26816 35636 27019
rect 35404 26767 35444 26776
rect 35596 26767 35636 26776
rect 35788 26816 35828 26825
rect 35980 26816 36020 27691
rect 36844 27497 36884 28288
rect 36940 27824 36980 28960
rect 37035 28916 37077 28925
rect 37035 28876 37036 28916
rect 37076 28876 37077 28916
rect 37035 28867 37077 28876
rect 37036 28580 37076 28867
rect 37612 28664 37652 31144
rect 37036 28531 37076 28540
rect 37516 28624 37652 28664
rect 37132 28328 37172 28337
rect 37516 28328 37556 28624
rect 37708 28496 37748 28505
rect 37172 28288 37556 28328
rect 37612 28456 37708 28496
rect 37132 28279 37172 28288
rect 36940 27784 37172 27824
rect 36940 27656 36980 27665
rect 36555 27488 36597 27497
rect 36555 27448 36556 27488
rect 36596 27448 36597 27488
rect 36555 27439 36597 27448
rect 36843 27488 36885 27497
rect 36843 27448 36844 27488
rect 36884 27448 36885 27488
rect 36843 27439 36885 27448
rect 36556 27354 36596 27439
rect 35828 26776 36020 26816
rect 35788 26767 35828 26776
rect 35308 26648 35348 26767
rect 35692 26732 35732 26741
rect 35348 26608 35636 26648
rect 35308 26599 35348 26608
rect 35115 26480 35157 26489
rect 35115 26440 35116 26480
rect 35156 26440 35157 26480
rect 35115 26431 35157 26440
rect 35499 26480 35541 26489
rect 35499 26440 35500 26480
rect 35540 26440 35541 26480
rect 35499 26431 35541 26440
rect 35500 26312 35540 26431
rect 35500 26263 35540 26272
rect 35403 26228 35445 26237
rect 35403 26188 35404 26228
rect 35444 26188 35445 26228
rect 35403 26179 35445 26188
rect 35020 26095 35060 26104
rect 35212 26144 35252 26155
rect 35212 26069 35252 26104
rect 35308 26144 35348 26153
rect 35211 26060 35253 26069
rect 35211 26020 35212 26060
rect 35252 26020 35253 26060
rect 35211 26011 35253 26020
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 35212 24632 35252 26011
rect 35308 24800 35348 26104
rect 35404 26144 35444 26179
rect 35404 26093 35444 26104
rect 35596 25304 35636 26608
rect 35692 25640 35732 26692
rect 35692 25600 35828 25640
rect 35596 25255 35636 25264
rect 35692 25304 35732 25315
rect 35692 25229 35732 25264
rect 35788 25304 35828 25600
rect 35788 25255 35828 25264
rect 35883 25304 35925 25313
rect 35883 25264 35884 25304
rect 35924 25264 35925 25304
rect 35883 25255 35925 25264
rect 35691 25220 35733 25229
rect 35691 25180 35692 25220
rect 35732 25180 35733 25220
rect 35691 25171 35733 25180
rect 35884 25170 35924 25255
rect 35980 25229 36020 26776
rect 36940 26489 36980 27616
rect 36939 26480 36981 26489
rect 36939 26440 36940 26480
rect 36980 26440 36981 26480
rect 36939 26431 36981 26440
rect 36555 26312 36597 26321
rect 36555 26272 36556 26312
rect 36596 26272 36597 26312
rect 36555 26263 36597 26272
rect 36556 26178 36596 26263
rect 36172 26144 36212 26153
rect 36172 25556 36212 26104
rect 37036 26144 37076 26153
rect 36267 26060 36309 26069
rect 36267 26020 36268 26060
rect 36308 26020 36309 26060
rect 36267 26011 36309 26020
rect 36172 25507 36212 25516
rect 36268 25304 36308 26011
rect 36651 25808 36693 25817
rect 36651 25768 36652 25808
rect 36692 25768 36693 25808
rect 36651 25759 36693 25768
rect 36459 25388 36501 25397
rect 36459 25348 36460 25388
rect 36500 25348 36501 25388
rect 36459 25339 36501 25348
rect 36268 25255 36308 25264
rect 35979 25220 36021 25229
rect 35979 25180 35980 25220
rect 36020 25180 36021 25220
rect 35979 25171 36021 25180
rect 36460 25220 36500 25339
rect 36460 25171 36500 25180
rect 36652 25318 36692 25759
rect 35404 25136 35444 25145
rect 35444 25096 35636 25136
rect 35404 25087 35444 25096
rect 35404 24800 35444 24809
rect 35308 24760 35404 24800
rect 35404 24751 35444 24760
rect 35596 24632 35636 25096
rect 36076 24632 36116 24641
rect 35596 24592 36076 24632
rect 35212 24583 35252 24592
rect 36076 24583 36116 24592
rect 36555 24464 36597 24473
rect 36555 24424 36556 24464
rect 36596 24424 36597 24464
rect 36555 24415 36597 24424
rect 35404 24380 35444 24389
rect 34443 24212 34485 24221
rect 34443 24172 34444 24212
rect 34484 24172 34485 24212
rect 34443 24163 34485 24172
rect 34251 24128 34293 24137
rect 34251 24088 34252 24128
rect 34292 24088 34293 24128
rect 34251 24079 34293 24088
rect 33963 23372 34005 23381
rect 33963 23332 33964 23372
rect 34004 23332 34005 23372
rect 33963 23323 34005 23332
rect 33676 23239 33716 23248
rect 33484 23154 33524 23239
rect 33196 22828 33428 22868
rect 33196 22373 33236 22828
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 34060 22541 34100 23752
rect 34156 23920 34676 23960
rect 34156 23792 34196 23920
rect 34348 23792 34388 23801
rect 34156 23743 34196 23752
rect 34252 23752 34348 23792
rect 34059 22532 34101 22541
rect 34059 22492 34060 22532
rect 34100 22492 34101 22532
rect 34059 22483 34101 22492
rect 34252 22532 34292 23752
rect 34348 23743 34388 23752
rect 34444 23792 34484 23801
rect 34347 23288 34389 23297
rect 34347 23248 34348 23288
rect 34388 23248 34389 23288
rect 34347 23239 34389 23248
rect 34348 23120 34388 23239
rect 34348 23071 34388 23080
rect 34444 22532 34484 23752
rect 34636 23792 34676 23920
rect 34636 23743 34676 23752
rect 34539 23708 34581 23717
rect 34539 23668 34540 23708
rect 34580 23668 34581 23708
rect 34539 23659 34581 23668
rect 34540 23574 34580 23659
rect 34828 23624 34868 23633
rect 34868 23584 35060 23624
rect 34828 23575 34868 23584
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 34539 23288 34581 23297
rect 34539 23248 34540 23288
rect 34580 23248 34581 23288
rect 34539 23239 34581 23248
rect 34252 22483 34292 22492
rect 34348 22492 34484 22532
rect 34155 22448 34197 22457
rect 34155 22408 34156 22448
rect 34196 22408 34197 22448
rect 34155 22399 34197 22408
rect 33195 22364 33237 22373
rect 33195 22324 33196 22364
rect 33236 22324 33237 22364
rect 33195 22315 33237 22324
rect 33772 22280 33812 22291
rect 33772 22205 33812 22240
rect 34059 22280 34101 22289
rect 34059 22240 34060 22280
rect 34100 22240 34101 22280
rect 34059 22231 34101 22240
rect 34156 22280 34196 22399
rect 33771 22196 33813 22205
rect 33771 22156 33772 22196
rect 33812 22156 33813 22196
rect 33771 22147 33813 22156
rect 33100 22112 33140 22121
rect 33100 21701 33140 22072
rect 33099 21692 33141 21701
rect 33099 21652 33100 21692
rect 33140 21652 33141 21692
rect 33099 21643 33141 21652
rect 33196 21608 33236 21617
rect 33099 21524 33141 21533
rect 33099 21484 33100 21524
rect 33140 21484 33141 21524
rect 33099 21475 33141 21484
rect 33100 21020 33140 21475
rect 33196 21449 33236 21568
rect 34060 21608 34100 22231
rect 34156 21617 34196 22240
rect 34060 21559 34100 21568
rect 34155 21608 34197 21617
rect 34155 21568 34156 21608
rect 34196 21568 34197 21608
rect 34155 21559 34197 21568
rect 34348 21533 34388 22492
rect 34443 22364 34485 22373
rect 34443 22324 34444 22364
rect 34484 22324 34485 22364
rect 34443 22315 34485 22324
rect 34444 22230 34484 22315
rect 34540 22280 34580 23239
rect 34923 23204 34965 23213
rect 34923 23164 34924 23204
rect 34964 23164 34965 23204
rect 34923 23155 34965 23164
rect 34924 23070 34964 23155
rect 34731 22952 34773 22961
rect 34731 22912 34732 22952
rect 34772 22912 34773 22952
rect 34731 22903 34773 22912
rect 34732 22818 34772 22903
rect 34827 22532 34869 22541
rect 34827 22492 34828 22532
rect 34868 22492 34869 22532
rect 34827 22483 34869 22492
rect 34540 22231 34580 22240
rect 34828 22280 34868 22483
rect 35020 22457 35060 23584
rect 35404 23297 35444 24340
rect 35500 23792 35540 23801
rect 35403 23288 35445 23297
rect 35403 23248 35404 23288
rect 35444 23248 35445 23288
rect 35403 23239 35445 23248
rect 35500 23129 35540 23752
rect 36364 23792 36404 23803
rect 36364 23717 36404 23752
rect 36363 23708 36405 23717
rect 36363 23668 36364 23708
rect 36404 23668 36405 23708
rect 36363 23659 36405 23668
rect 36556 23708 36596 24415
rect 36652 23876 36692 25278
rect 37036 25229 37076 26104
rect 37132 25724 37172 27784
rect 37324 27656 37364 27665
rect 37612 27656 37652 28456
rect 37708 28447 37748 28456
rect 37707 28328 37749 28337
rect 37804 28328 37844 32152
rect 38092 32143 38132 32152
rect 38188 32033 38228 32647
rect 38187 32024 38229 32033
rect 38187 31984 38188 32024
rect 38228 31984 38229 32024
rect 38187 31975 38229 31984
rect 38764 32024 38804 32824
rect 39628 32192 39668 33403
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 39915 32696 39957 32705
rect 39915 32656 39916 32696
rect 39956 32656 39957 32696
rect 39915 32647 39957 32656
rect 39916 32562 39956 32647
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 39628 32143 39668 32152
rect 40588 32192 40628 32201
rect 39723 32108 39765 32117
rect 39723 32068 39724 32108
rect 39764 32068 39765 32108
rect 39723 32059 39765 32068
rect 38764 31975 38804 31984
rect 39244 32024 39284 32033
rect 38188 31352 38228 31975
rect 38572 31940 38612 31949
rect 38572 31361 38612 31900
rect 39244 31865 39284 31984
rect 39724 31974 39764 32059
rect 39916 31940 39956 31949
rect 39956 31900 40148 31940
rect 39916 31891 39956 31900
rect 38763 31856 38805 31865
rect 38763 31816 38764 31856
rect 38804 31816 38805 31856
rect 38763 31807 38805 31816
rect 39243 31856 39285 31865
rect 39243 31816 39244 31856
rect 39284 31816 39285 31856
rect 39243 31807 39285 31816
rect 38188 31303 38228 31312
rect 38571 31352 38613 31361
rect 38571 31312 38572 31352
rect 38612 31312 38613 31352
rect 38571 31303 38613 31312
rect 38764 31352 38804 31807
rect 38764 31303 38804 31312
rect 39628 31352 39668 31361
rect 38380 31268 38420 31277
rect 38380 30857 38420 31228
rect 38379 30848 38421 30857
rect 38379 30808 38380 30848
rect 38420 30808 38421 30848
rect 38379 30799 38421 30808
rect 38283 30764 38325 30773
rect 38283 30724 38284 30764
rect 38324 30724 38325 30764
rect 38283 30715 38325 30724
rect 38284 30680 38324 30715
rect 38284 30629 38324 30640
rect 38572 30605 38612 31303
rect 39339 31184 39381 31193
rect 39339 31144 39340 31184
rect 39380 31144 39381 31184
rect 39339 31135 39381 31144
rect 38955 30848 38997 30857
rect 38955 30808 38956 30848
rect 38996 30808 38997 30848
rect 38955 30799 38997 30808
rect 38956 30714 38996 30799
rect 39147 30680 39189 30689
rect 39147 30640 39148 30680
rect 39188 30640 39189 30680
rect 39147 30631 39189 30640
rect 39244 30680 39284 30689
rect 38571 30596 38613 30605
rect 38571 30556 38572 30596
rect 38612 30556 38613 30596
rect 38571 30547 38613 30556
rect 38091 30428 38133 30437
rect 38091 30388 38092 30428
rect 38132 30388 38133 30428
rect 38091 30379 38133 30388
rect 38092 30294 38132 30379
rect 38572 29840 38612 30547
rect 39148 30546 39188 30631
rect 38955 30344 38997 30353
rect 39244 30344 39284 30640
rect 39340 30680 39380 31135
rect 39435 30932 39477 30941
rect 39435 30892 39436 30932
rect 39476 30892 39477 30932
rect 39435 30883 39477 30892
rect 39340 30631 39380 30640
rect 39436 30680 39476 30883
rect 39436 30631 39476 30640
rect 39628 30605 39668 31312
rect 40108 30680 40148 31900
rect 40588 31193 40628 32152
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 41932 31520 41972 31529
rect 40587 31184 40629 31193
rect 40587 31144 40588 31184
rect 40628 31144 40629 31184
rect 40587 31135 40629 31144
rect 40779 31184 40821 31193
rect 40779 31144 40780 31184
rect 40820 31144 40821 31184
rect 40779 31135 40821 31144
rect 40780 31050 40820 31135
rect 40108 30631 40148 30640
rect 41452 30680 41492 30689
rect 41836 30680 41876 30689
rect 41932 30680 41972 31480
rect 43276 31352 43316 31361
rect 43180 31184 43220 31193
rect 42892 31144 43180 31184
rect 41492 30640 41684 30680
rect 41452 30631 41492 30640
rect 39627 30596 39669 30605
rect 39627 30556 39628 30596
rect 39668 30556 39669 30596
rect 39627 30547 39669 30556
rect 39628 30462 39668 30547
rect 39819 30428 39861 30437
rect 39819 30388 39820 30428
rect 39860 30388 39861 30428
rect 39819 30379 39861 30388
rect 40012 30428 40052 30437
rect 38955 30304 38956 30344
rect 38996 30304 39284 30344
rect 38955 30295 38997 30304
rect 37899 29168 37941 29177
rect 37899 29128 37900 29168
rect 37940 29128 37941 29168
rect 37899 29119 37941 29128
rect 37707 28288 37708 28328
rect 37748 28288 37844 28328
rect 37707 28279 37749 28288
rect 37364 27616 37652 27656
rect 37324 27607 37364 27616
rect 37708 27068 37748 28279
rect 37708 27019 37748 27028
rect 37323 26564 37365 26573
rect 37323 26524 37324 26564
rect 37364 26524 37365 26564
rect 37323 26515 37365 26524
rect 37324 26228 37364 26515
rect 37900 26396 37940 29119
rect 38091 29000 38133 29009
rect 38572 29000 38612 29800
rect 38091 28960 38092 29000
rect 38132 28960 38133 29000
rect 38091 28951 38133 28960
rect 38188 28960 38612 29000
rect 38092 28866 38132 28951
rect 38188 27656 38228 28960
rect 38380 28328 38420 28337
rect 38380 27749 38420 28288
rect 38379 27740 38421 27749
rect 38379 27700 38380 27740
rect 38420 27700 38421 27740
rect 38379 27691 38421 27700
rect 38188 27607 38228 27616
rect 38763 27572 38805 27581
rect 38763 27532 38764 27572
rect 38804 27532 38805 27572
rect 38763 27523 38805 27532
rect 38476 26984 38516 26993
rect 38187 26816 38229 26825
rect 38187 26776 38188 26816
rect 38228 26776 38229 26816
rect 38187 26767 38229 26776
rect 37995 26648 38037 26657
rect 37995 26608 37996 26648
rect 38036 26608 38037 26648
rect 37995 26599 38037 26608
rect 37708 26356 37940 26396
rect 37419 26312 37461 26321
rect 37419 26272 37420 26312
rect 37460 26272 37461 26312
rect 37419 26263 37461 26272
rect 37324 26179 37364 26188
rect 37228 26144 37268 26155
rect 37228 26069 37268 26104
rect 37420 26144 37460 26263
rect 37420 26095 37460 26104
rect 37227 26060 37269 26069
rect 37227 26020 37228 26060
rect 37268 26020 37269 26060
rect 37227 26011 37269 26020
rect 37228 25901 37268 26011
rect 37708 25976 37748 26356
rect 37803 26228 37845 26237
rect 37803 26188 37804 26228
rect 37844 26188 37845 26228
rect 37803 26179 37845 26188
rect 37804 26094 37844 26179
rect 37900 26144 37940 26155
rect 37900 26069 37940 26104
rect 37996 26144 38036 26599
rect 38188 26153 38228 26767
rect 38476 26741 38516 26944
rect 38764 26816 38804 27523
rect 38859 27488 38901 27497
rect 38859 27448 38860 27488
rect 38900 27448 38901 27488
rect 38859 27439 38901 27448
rect 38764 26767 38804 26776
rect 38860 26816 38900 27439
rect 38475 26732 38517 26741
rect 38475 26692 38476 26732
rect 38516 26692 38517 26732
rect 38475 26683 38517 26692
rect 38379 26480 38421 26489
rect 38379 26440 38380 26480
rect 38420 26440 38421 26480
rect 38379 26431 38421 26440
rect 38380 26312 38420 26431
rect 38380 26263 38420 26272
rect 38283 26228 38325 26237
rect 38283 26188 38284 26228
rect 38324 26188 38325 26228
rect 38283 26179 38325 26188
rect 38475 26228 38517 26237
rect 38475 26188 38476 26228
rect 38516 26188 38517 26228
rect 38475 26179 38517 26188
rect 37996 26095 38036 26104
rect 38092 26144 38132 26153
rect 37899 26060 37941 26069
rect 37899 26020 37900 26060
rect 37940 26020 37941 26060
rect 37899 26011 37941 26020
rect 37708 25936 37844 25976
rect 37227 25892 37269 25901
rect 37227 25852 37228 25892
rect 37268 25852 37269 25892
rect 37227 25843 37269 25852
rect 37132 25684 37748 25724
rect 37131 25556 37173 25565
rect 37131 25516 37132 25556
rect 37172 25516 37173 25556
rect 37131 25507 37173 25516
rect 37132 25304 37172 25507
rect 37611 25388 37653 25397
rect 37611 25348 37612 25388
rect 37652 25348 37653 25388
rect 37611 25339 37653 25348
rect 37708 25388 37748 25684
rect 37708 25339 37748 25348
rect 37132 25255 37172 25264
rect 37612 25254 37652 25339
rect 37035 25220 37077 25229
rect 37035 25180 37036 25220
rect 37076 25180 37077 25220
rect 37035 25171 37077 25180
rect 37707 25136 37749 25145
rect 37707 25096 37708 25136
rect 37748 25096 37749 25136
rect 37707 25087 37749 25096
rect 37708 24632 37748 25087
rect 37708 24583 37748 24592
rect 37804 23876 37844 25936
rect 38092 25817 38132 26104
rect 38187 26144 38229 26153
rect 38187 26104 38188 26144
rect 38228 26104 38229 26144
rect 38187 26095 38229 26104
rect 38284 26144 38324 26179
rect 38284 26093 38324 26104
rect 38476 26144 38516 26179
rect 38187 25892 38229 25901
rect 38187 25852 38188 25892
rect 38228 25852 38229 25892
rect 38187 25843 38229 25852
rect 38091 25808 38133 25817
rect 38091 25768 38092 25808
rect 38132 25768 38133 25808
rect 38091 25759 38133 25768
rect 38091 25304 38133 25313
rect 38091 25264 38092 25304
rect 38132 25264 38133 25304
rect 38091 25255 38133 25264
rect 38188 25304 38228 25843
rect 38476 25817 38516 26104
rect 38572 26144 38612 26153
rect 38763 26144 38805 26153
rect 38612 26104 38708 26144
rect 38572 26095 38612 26104
rect 38475 25808 38517 25817
rect 38475 25768 38476 25808
rect 38516 25768 38517 25808
rect 38475 25759 38517 25768
rect 38228 25264 38324 25304
rect 38188 25255 38228 25264
rect 38092 25170 38132 25255
rect 36652 23836 36740 23876
rect 36700 23834 36740 23836
rect 37804 23827 37844 23836
rect 36700 23785 36740 23794
rect 37228 23792 37268 23801
rect 37708 23792 37748 23801
rect 36556 23659 36596 23668
rect 35692 23624 35732 23633
rect 35692 23213 35732 23584
rect 35691 23204 35733 23213
rect 35691 23164 35692 23204
rect 35732 23164 35733 23204
rect 35691 23155 35733 23164
rect 35211 23120 35253 23129
rect 35211 23080 35212 23120
rect 35252 23080 35253 23120
rect 35211 23071 35253 23080
rect 35308 23120 35348 23129
rect 35019 22448 35061 22457
rect 35019 22408 35020 22448
rect 35060 22408 35061 22448
rect 35019 22399 35061 22408
rect 34828 22231 34868 22240
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 35212 21776 35252 23071
rect 35308 22961 35348 23080
rect 35499 23120 35541 23129
rect 35499 23080 35500 23120
rect 35540 23080 35541 23120
rect 35499 23071 35541 23080
rect 36172 23120 36212 23129
rect 35307 22952 35349 22961
rect 35307 22912 35308 22952
rect 35348 22912 35349 22952
rect 35307 22903 35349 22912
rect 36172 22289 36212 23080
rect 37228 22961 37268 23752
rect 37612 23752 37708 23792
rect 37323 23372 37365 23381
rect 37323 23332 37324 23372
rect 37364 23332 37365 23372
rect 37323 23323 37365 23332
rect 37324 23288 37364 23323
rect 37324 23237 37364 23248
rect 37227 22952 37269 22961
rect 37227 22912 37228 22952
rect 37268 22912 37269 22952
rect 37227 22903 37269 22912
rect 35212 21727 35252 21736
rect 35692 22280 35732 22289
rect 35596 21617 35636 21702
rect 35595 21608 35637 21617
rect 35595 21568 35596 21608
rect 35636 21568 35637 21608
rect 35595 21559 35637 21568
rect 34347 21524 34389 21533
rect 34347 21484 34348 21524
rect 34388 21484 34389 21524
rect 34347 21475 34389 21484
rect 33195 21440 33237 21449
rect 33195 21400 33196 21440
rect 33236 21400 33237 21440
rect 33195 21391 33237 21400
rect 35595 21440 35637 21449
rect 35595 21400 35596 21440
rect 35636 21400 35637 21440
rect 35595 21391 35637 21400
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 33100 20971 33140 20980
rect 35596 20768 35636 21391
rect 35596 20719 35636 20728
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 30700 20140 30836 20180
rect 30796 20096 30836 20140
rect 32908 20140 33044 20180
rect 30796 20047 30836 20056
rect 32044 20096 32084 20105
rect 30220 19720 30548 19760
rect 29547 19592 29589 19601
rect 29547 19552 29548 19592
rect 29588 19552 29589 19592
rect 29547 19543 29589 19552
rect 30315 19592 30357 19601
rect 30315 19552 30316 19592
rect 30356 19552 30357 19592
rect 30315 19543 30357 19552
rect 30316 19508 30356 19543
rect 30316 19457 30356 19468
rect 30508 19265 30548 19720
rect 29740 19256 29780 19265
rect 29740 19097 29780 19216
rect 29836 19256 29876 19265
rect 30316 19256 30356 19265
rect 29739 19088 29781 19097
rect 29739 19048 29740 19088
rect 29780 19048 29781 19088
rect 29739 19039 29781 19048
rect 29547 18668 29589 18677
rect 29547 18628 29548 18668
rect 29588 18628 29589 18668
rect 29547 18619 29589 18628
rect 29356 18535 29396 18544
rect 29548 18584 29588 18619
rect 28683 18500 28725 18509
rect 28683 18460 28684 18500
rect 28724 18460 28725 18500
rect 28683 18451 28725 18460
rect 28683 18332 28725 18341
rect 28683 18292 28684 18332
rect 28724 18292 28725 18332
rect 28683 18283 28725 18292
rect 28684 17744 28724 18283
rect 28587 17408 28629 17417
rect 28587 17368 28588 17408
rect 28628 17368 28629 17408
rect 28587 17359 28629 17368
rect 28395 17324 28437 17333
rect 28395 17284 28396 17324
rect 28436 17284 28437 17324
rect 28395 17275 28437 17284
rect 28684 17249 28724 17704
rect 28780 17744 28820 18535
rect 29548 18533 29588 18544
rect 29644 18584 29684 18593
rect 29740 18584 29780 19039
rect 29836 18761 29876 19216
rect 30028 19216 30316 19256
rect 29835 18752 29877 18761
rect 29835 18712 29836 18752
rect 29876 18712 29877 18752
rect 30028 18752 30068 19216
rect 30316 19207 30356 19216
rect 30507 19256 30549 19265
rect 30507 19216 30508 19256
rect 30548 19216 30549 19256
rect 30507 19207 30549 19216
rect 30508 19122 30548 19207
rect 30124 19088 30164 19097
rect 30164 19048 30356 19088
rect 30124 19039 30164 19048
rect 30028 18712 30164 18752
rect 29835 18703 29877 18712
rect 29684 18544 29780 18584
rect 29835 18584 29877 18593
rect 29835 18544 29836 18584
rect 29876 18544 29877 18584
rect 29644 18535 29684 18544
rect 29835 18535 29877 18544
rect 30028 18584 30068 18593
rect 29836 18450 29876 18535
rect 30028 18425 30068 18544
rect 30027 18416 30069 18425
rect 30027 18376 30028 18416
rect 30068 18376 30069 18416
rect 30027 18367 30069 18376
rect 29356 18332 29396 18341
rect 29164 18292 29356 18332
rect 28875 17912 28917 17921
rect 28875 17872 28876 17912
rect 28916 17872 28917 17912
rect 28875 17863 28917 17872
rect 28780 17695 28820 17704
rect 28779 17576 28821 17585
rect 28779 17536 28780 17576
rect 28820 17536 28821 17576
rect 28876 17576 28916 17863
rect 28972 17828 29012 17839
rect 28972 17753 29012 17788
rect 28971 17744 29013 17753
rect 28971 17704 28972 17744
rect 29012 17704 29013 17744
rect 28971 17695 29013 17704
rect 29164 17744 29204 18292
rect 29356 18283 29396 18292
rect 29932 18332 29972 18341
rect 29356 17912 29396 17921
rect 29739 17912 29781 17921
rect 29396 17872 29492 17912
rect 29356 17863 29396 17872
rect 29452 17753 29492 17872
rect 29739 17872 29740 17912
rect 29780 17872 29781 17912
rect 29739 17863 29781 17872
rect 29356 17744 29396 17753
rect 29164 17704 29356 17744
rect 28876 17536 29108 17576
rect 28779 17527 28821 17536
rect 28683 17240 28725 17249
rect 28683 17200 28684 17240
rect 28724 17200 28725 17240
rect 28683 17191 28725 17200
rect 28396 17081 28436 17166
rect 28300 17023 28340 17032
rect 28395 17072 28437 17081
rect 28395 17032 28396 17072
rect 28436 17032 28437 17072
rect 28395 17023 28437 17032
rect 28588 17072 28628 17081
rect 27820 16780 27956 16820
rect 28107 16820 28149 16829
rect 28107 16780 28108 16820
rect 28148 16780 28149 16820
rect 27723 16484 27765 16493
rect 27723 16444 27724 16484
rect 27764 16444 27765 16484
rect 27723 16435 27765 16444
rect 27820 16316 27860 16780
rect 28107 16771 28149 16780
rect 28395 16400 28437 16409
rect 28395 16360 28396 16400
rect 28436 16360 28437 16400
rect 28395 16351 28437 16360
rect 27436 16073 27476 16192
rect 27628 16276 27860 16316
rect 27915 16316 27957 16325
rect 27915 16276 27916 16316
rect 27956 16276 27957 16316
rect 27435 16064 27477 16073
rect 27435 16024 27436 16064
rect 27476 16024 27477 16064
rect 27435 16015 27477 16024
rect 27148 15856 27380 15896
rect 27051 15644 27093 15653
rect 27051 15604 27052 15644
rect 27092 15604 27093 15644
rect 27051 15595 27093 15604
rect 27051 14972 27093 14981
rect 27051 14932 27052 14972
rect 27092 14932 27093 14972
rect 27051 14923 27093 14932
rect 26955 14888 26997 14897
rect 26955 14848 26956 14888
rect 26996 14848 26997 14888
rect 26955 14839 26997 14848
rect 26859 14804 26901 14813
rect 26859 14764 26860 14804
rect 26900 14764 26901 14804
rect 26859 14755 26901 14764
rect 26764 14671 26804 14680
rect 26860 14670 26900 14755
rect 26955 14720 26997 14729
rect 26955 14680 26956 14720
rect 26996 14680 26997 14720
rect 26955 14671 26997 14680
rect 26956 14141 26996 14671
rect 26955 14132 26997 14141
rect 26668 14092 26900 14132
rect 26516 14008 26804 14048
rect 26476 13999 26516 14008
rect 26475 13880 26517 13889
rect 26475 13840 26476 13880
rect 26516 13840 26517 13880
rect 26475 13831 26517 13840
rect 26476 13208 26516 13831
rect 26476 13159 26516 13168
rect 26764 13208 26804 14008
rect 26764 13159 26804 13168
rect 26860 12545 26900 14092
rect 26955 14092 26956 14132
rect 26996 14092 26997 14132
rect 26955 14083 26997 14092
rect 27052 13880 27092 14923
rect 27148 14720 27188 15856
rect 27339 15644 27381 15653
rect 27339 15604 27340 15644
rect 27380 15604 27381 15644
rect 27339 15595 27381 15604
rect 27340 15510 27380 15595
rect 27532 15560 27572 15569
rect 27628 15560 27668 16276
rect 27915 16267 27957 16276
rect 27916 16232 27956 16267
rect 27916 16181 27956 16192
rect 28011 16232 28053 16241
rect 28011 16192 28012 16232
rect 28052 16192 28053 16232
rect 28011 16183 28053 16192
rect 28108 16232 28148 16241
rect 28012 16098 28052 16183
rect 27915 16064 27957 16073
rect 27915 16024 27916 16064
rect 27956 16024 27957 16064
rect 27915 16015 27957 16024
rect 27572 15520 27668 15560
rect 27820 15560 27860 15571
rect 27532 15511 27572 15520
rect 27820 15485 27860 15520
rect 27819 15476 27861 15485
rect 27819 15436 27820 15476
rect 27860 15436 27861 15476
rect 27819 15427 27861 15436
rect 27435 15308 27477 15317
rect 27435 15268 27436 15308
rect 27476 15268 27477 15308
rect 27435 15259 27477 15268
rect 27243 15140 27285 15149
rect 27243 15100 27244 15140
rect 27284 15100 27285 15140
rect 27243 15091 27285 15100
rect 27244 14972 27284 15091
rect 27244 14923 27284 14932
rect 27339 14888 27381 14897
rect 27339 14848 27340 14888
rect 27380 14848 27381 14888
rect 27339 14839 27381 14848
rect 27340 14743 27380 14839
rect 27340 14694 27380 14703
rect 27148 14671 27188 14680
rect 27436 14636 27476 15259
rect 27340 14596 27476 14636
rect 27532 14720 27572 14729
rect 27148 13880 27188 13889
rect 27052 13840 27148 13880
rect 27148 13831 27188 13840
rect 27243 13796 27285 13805
rect 27340 13796 27380 14596
rect 27532 14561 27572 14680
rect 27724 14720 27764 14731
rect 27820 14729 27860 15427
rect 27724 14645 27764 14680
rect 27819 14720 27861 14729
rect 27819 14680 27820 14720
rect 27860 14680 27861 14720
rect 27819 14671 27861 14680
rect 27628 14636 27668 14645
rect 27531 14552 27573 14561
rect 27531 14512 27532 14552
rect 27572 14512 27573 14552
rect 27531 14503 27573 14512
rect 27436 14141 27476 14226
rect 27435 14132 27477 14141
rect 27435 14092 27436 14132
rect 27476 14092 27477 14132
rect 27435 14083 27477 14092
rect 27628 14057 27668 14596
rect 27723 14636 27765 14645
rect 27723 14596 27724 14636
rect 27764 14596 27765 14636
rect 27723 14587 27765 14596
rect 27532 14048 27572 14057
rect 27435 13964 27477 13973
rect 27435 13924 27436 13964
rect 27476 13924 27477 13964
rect 27435 13915 27477 13924
rect 27243 13756 27244 13796
rect 27284 13756 27380 13796
rect 27243 13747 27285 13756
rect 26956 13208 26996 13217
rect 26284 12487 26324 12496
rect 26859 12536 26901 12545
rect 26859 12496 26860 12536
rect 26900 12496 26901 12536
rect 26859 12487 26901 12496
rect 26283 12368 26325 12377
rect 26283 12328 26284 12368
rect 26324 12328 26325 12368
rect 26283 12319 26325 12328
rect 26187 12284 26229 12293
rect 26187 12244 26188 12284
rect 26228 12244 26229 12284
rect 26187 12235 26229 12244
rect 26188 11621 26228 12235
rect 26187 11612 26229 11621
rect 26187 11572 26188 11612
rect 26228 11572 26229 11612
rect 26187 11563 26229 11572
rect 25708 11320 25940 11360
rect 25611 10352 25653 10361
rect 25611 10312 25612 10352
rect 25652 10312 25653 10352
rect 25611 10303 25653 10312
rect 25708 10277 25748 11320
rect 26284 10436 26324 12319
rect 26956 12041 26996 13168
rect 27147 12620 27189 12629
rect 27147 12580 27148 12620
rect 27188 12580 27189 12620
rect 27147 12571 27189 12580
rect 26955 12032 26997 12041
rect 26955 11992 26956 12032
rect 26996 11992 26997 12032
rect 26955 11983 26997 11992
rect 27148 11873 27188 12571
rect 27244 12536 27284 13747
rect 27147 11864 27189 11873
rect 27147 11824 27148 11864
rect 27188 11824 27189 11864
rect 27147 11815 27189 11824
rect 26859 11780 26901 11789
rect 26859 11740 26860 11780
rect 26900 11740 26901 11780
rect 26859 11731 26901 11740
rect 26572 11696 26612 11707
rect 26572 11621 26612 11656
rect 26667 11696 26709 11705
rect 26667 11656 26668 11696
rect 26708 11656 26709 11696
rect 26667 11647 26709 11656
rect 26571 11612 26613 11621
rect 26571 11572 26572 11612
rect 26612 11572 26613 11612
rect 26571 11563 26613 11572
rect 26668 11562 26708 11647
rect 26860 11646 26900 11731
rect 27052 11696 27092 11705
rect 26956 11656 27052 11696
rect 26956 11033 26996 11656
rect 27052 11647 27092 11656
rect 27148 11360 27188 11815
rect 27052 11320 27188 11360
rect 27052 11192 27092 11320
rect 27052 11143 27092 11152
rect 26955 11024 26997 11033
rect 26955 10984 26956 11024
rect 26996 10984 26997 11024
rect 26955 10975 26997 10984
rect 26284 10387 26324 10396
rect 26956 10277 26996 10975
rect 27244 10949 27284 12496
rect 27339 12536 27381 12545
rect 27339 12496 27340 12536
rect 27380 12496 27381 12536
rect 27339 12487 27381 12496
rect 27340 11705 27380 12487
rect 27436 11948 27476 13915
rect 27532 13805 27572 14008
rect 27627 14048 27669 14057
rect 27627 14008 27628 14048
rect 27668 14008 27669 14048
rect 27627 13999 27669 14008
rect 27820 14048 27860 14059
rect 27820 13973 27860 14008
rect 27819 13964 27861 13973
rect 27819 13924 27820 13964
rect 27860 13924 27861 13964
rect 27819 13915 27861 13924
rect 27916 13805 27956 16015
rect 28011 14888 28053 14897
rect 28011 14848 28012 14888
rect 28052 14848 28053 14888
rect 28011 14839 28053 14848
rect 27531 13796 27573 13805
rect 27531 13756 27532 13796
rect 27572 13756 27573 13796
rect 27531 13747 27573 13756
rect 27915 13796 27957 13805
rect 27915 13756 27916 13796
rect 27956 13756 27957 13796
rect 27915 13747 27957 13756
rect 27724 13208 27764 13217
rect 27532 13168 27724 13208
rect 27532 12704 27572 13168
rect 27724 13159 27764 13168
rect 27819 13208 27861 13217
rect 27819 13168 27820 13208
rect 27860 13168 27861 13208
rect 27819 13159 27861 13168
rect 27916 13208 27956 13217
rect 27820 13074 27860 13159
rect 27916 12956 27956 13168
rect 28012 13208 28052 14839
rect 28108 14720 28148 16192
rect 28396 15653 28436 16351
rect 28588 16064 28628 17032
rect 28683 17072 28725 17081
rect 28683 17032 28684 17072
rect 28724 17032 28725 17072
rect 28683 17023 28725 17032
rect 28780 17072 28820 17527
rect 28971 17408 29013 17417
rect 28971 17368 28972 17408
rect 29012 17368 29013 17408
rect 28971 17359 29013 17368
rect 28875 17240 28917 17249
rect 28875 17200 28876 17240
rect 28916 17200 28917 17240
rect 28875 17191 28917 17200
rect 28780 17023 28820 17032
rect 28876 17072 28916 17191
rect 28876 17023 28916 17032
rect 28684 16938 28724 17023
rect 28972 16904 29012 17359
rect 29068 17072 29108 17536
rect 29164 17249 29204 17704
rect 29356 17695 29396 17704
rect 29451 17744 29493 17753
rect 29451 17704 29452 17744
rect 29492 17704 29493 17744
rect 29451 17695 29493 17704
rect 29740 17744 29780 17863
rect 29740 17695 29780 17704
rect 29836 17744 29876 17753
rect 29932 17744 29972 18292
rect 30028 17921 30068 18006
rect 30027 17912 30069 17921
rect 30027 17872 30028 17912
rect 30068 17872 30069 17912
rect 30027 17863 30069 17872
rect 30028 17744 30068 17753
rect 29932 17704 30028 17744
rect 29355 17576 29397 17585
rect 29355 17536 29356 17576
rect 29396 17536 29397 17576
rect 29355 17527 29397 17536
rect 29163 17240 29205 17249
rect 29163 17200 29164 17240
rect 29204 17200 29205 17240
rect 29163 17191 29205 17200
rect 29068 17023 29108 17032
rect 29068 16904 29108 16913
rect 28972 16864 29068 16904
rect 29068 16855 29108 16864
rect 29164 16577 29204 17191
rect 29259 17072 29301 17081
rect 29259 17032 29260 17072
rect 29300 17032 29301 17072
rect 29259 17023 29301 17032
rect 29356 17072 29396 17527
rect 29356 17023 29396 17032
rect 29260 16938 29300 17023
rect 29452 16904 29492 17695
rect 29547 17576 29589 17585
rect 29836 17576 29876 17704
rect 29547 17536 29548 17576
rect 29588 17536 29972 17576
rect 29547 17527 29589 17536
rect 29548 17442 29588 17527
rect 29356 16864 29492 16904
rect 29548 17072 29588 17081
rect 29163 16568 29205 16577
rect 29163 16528 29164 16568
rect 29204 16528 29205 16568
rect 29163 16519 29205 16528
rect 29259 16316 29301 16325
rect 29259 16276 29260 16316
rect 29300 16276 29301 16316
rect 29259 16267 29301 16276
rect 29260 16064 29300 16267
rect 29356 16232 29396 16864
rect 29451 16568 29493 16577
rect 29451 16528 29452 16568
rect 29492 16528 29493 16568
rect 29451 16519 29493 16528
rect 29356 16183 29396 16192
rect 29452 16232 29492 16519
rect 29548 16484 29588 17032
rect 29932 17072 29972 17536
rect 30028 17081 30068 17704
rect 29932 17023 29972 17032
rect 30027 17072 30069 17081
rect 30027 17032 30028 17072
rect 30068 17032 30069 17072
rect 30027 17023 30069 17032
rect 29643 16988 29685 16997
rect 29643 16948 29644 16988
rect 29684 16948 29685 16988
rect 29643 16939 29685 16948
rect 29836 16988 29876 16997
rect 29644 16854 29684 16939
rect 29740 16904 29780 16913
rect 29644 16484 29684 16493
rect 29548 16444 29644 16484
rect 29644 16435 29684 16444
rect 29644 16232 29684 16241
rect 29452 16183 29492 16192
rect 29548 16192 29644 16232
rect 29548 16064 29588 16192
rect 29644 16183 29684 16192
rect 29740 16064 29780 16864
rect 29836 16577 29876 16948
rect 29835 16568 29877 16577
rect 29835 16528 29836 16568
rect 29876 16528 29877 16568
rect 29835 16519 29877 16528
rect 29835 16148 29877 16157
rect 29835 16108 29836 16148
rect 29876 16108 29877 16148
rect 29835 16099 29877 16108
rect 28588 16024 28916 16064
rect 29260 16024 29588 16064
rect 29644 16024 29780 16064
rect 28491 15728 28533 15737
rect 28491 15688 28492 15728
rect 28532 15688 28533 15728
rect 28491 15679 28533 15688
rect 28395 15644 28437 15653
rect 28395 15604 28396 15644
rect 28436 15604 28437 15644
rect 28395 15595 28437 15604
rect 28396 15401 28436 15595
rect 28492 15594 28532 15679
rect 28588 15644 28628 15653
rect 28395 15392 28437 15401
rect 28395 15352 28396 15392
rect 28436 15352 28437 15392
rect 28395 15343 28437 15352
rect 28588 14897 28628 15604
rect 28683 15644 28725 15653
rect 28683 15604 28684 15644
rect 28724 15604 28725 15644
rect 28683 15595 28725 15604
rect 28684 15560 28724 15595
rect 28684 15509 28724 15520
rect 28780 15560 28820 15569
rect 28683 15392 28725 15401
rect 28683 15352 28684 15392
rect 28724 15352 28725 15392
rect 28683 15343 28725 15352
rect 28684 15258 28724 15343
rect 28780 14981 28820 15520
rect 28876 15149 28916 16024
rect 29259 15728 29301 15737
rect 29259 15688 29260 15728
rect 29300 15688 29301 15728
rect 29259 15679 29301 15688
rect 29067 15644 29109 15653
rect 29067 15604 29068 15644
rect 29108 15604 29109 15644
rect 29067 15595 29109 15604
rect 28972 15560 29012 15569
rect 28972 15317 29012 15520
rect 29068 15560 29108 15595
rect 29260 15594 29300 15679
rect 29068 15509 29108 15520
rect 29164 15560 29204 15569
rect 29164 15401 29204 15520
rect 29163 15392 29205 15401
rect 29163 15352 29164 15392
rect 29204 15352 29205 15392
rect 29163 15343 29205 15352
rect 28971 15308 29013 15317
rect 28971 15268 28972 15308
rect 29012 15268 29013 15308
rect 28971 15259 29013 15268
rect 28875 15140 28917 15149
rect 29356 15140 29396 16024
rect 29547 15644 29589 15653
rect 29547 15604 29548 15644
rect 29588 15604 29589 15644
rect 29547 15595 29589 15604
rect 28875 15100 28876 15140
rect 28916 15100 28917 15140
rect 28875 15091 28917 15100
rect 28972 15100 29396 15140
rect 29451 15140 29493 15149
rect 29451 15100 29452 15140
rect 29492 15100 29493 15140
rect 28779 14972 28821 14981
rect 28779 14932 28780 14972
rect 28820 14932 28821 14972
rect 28779 14923 28821 14932
rect 28587 14888 28629 14897
rect 28587 14848 28588 14888
rect 28628 14848 28629 14888
rect 28587 14839 28629 14848
rect 28779 14804 28821 14813
rect 28779 14764 28780 14804
rect 28820 14764 28821 14804
rect 28779 14755 28821 14764
rect 28108 14561 28148 14680
rect 28204 14720 28244 14729
rect 28204 14645 28244 14680
rect 28683 14720 28725 14729
rect 28683 14680 28684 14720
rect 28724 14680 28725 14720
rect 28683 14671 28725 14680
rect 28780 14720 28820 14755
rect 28203 14636 28245 14645
rect 28203 14596 28204 14636
rect 28244 14596 28245 14636
rect 28203 14587 28245 14596
rect 28107 14552 28149 14561
rect 28107 14512 28108 14552
rect 28148 14512 28149 14552
rect 28107 14503 28149 14512
rect 28204 14216 28244 14587
rect 28492 14552 28532 14561
rect 28684 14552 28724 14671
rect 28108 14176 28244 14216
rect 28396 14512 28492 14552
rect 28532 14512 28724 14552
rect 28108 13973 28148 14176
rect 28204 14048 28244 14057
rect 28107 13964 28149 13973
rect 28107 13924 28108 13964
rect 28148 13924 28149 13964
rect 28107 13915 28149 13924
rect 28107 13796 28149 13805
rect 28107 13756 28108 13796
rect 28148 13756 28149 13796
rect 28107 13747 28149 13756
rect 28012 13159 28052 13168
rect 27724 12916 27956 12956
rect 27628 12713 27668 12732
rect 27627 12704 27669 12713
rect 27572 12664 27628 12704
rect 27668 12664 27669 12704
rect 27532 12655 27572 12664
rect 27627 12655 27669 12664
rect 27724 12629 27764 12916
rect 28108 12872 28148 13747
rect 28204 13208 28244 14008
rect 28299 14048 28341 14057
rect 28299 14008 28300 14048
rect 28340 14008 28341 14048
rect 28299 13999 28341 14008
rect 28396 14048 28436 14512
rect 28492 14503 28532 14512
rect 28396 13999 28436 14008
rect 28492 14048 28532 14057
rect 28780 14048 28820 14680
rect 28972 14720 29012 15100
rect 29451 15091 29493 15100
rect 29162 14804 29204 14813
rect 29162 14764 29163 14804
rect 29203 14764 29204 14804
rect 29162 14755 29204 14764
rect 29164 14720 29204 14755
rect 29012 14680 29108 14720
rect 28972 14671 29012 14680
rect 28960 14561 29000 14580
rect 28876 14552 28916 14561
rect 28960 14552 29013 14561
rect 28916 14512 28972 14552
rect 29012 14512 29013 14552
rect 28876 14503 28916 14512
rect 28971 14503 29013 14512
rect 28875 14384 28917 14393
rect 29068 14384 29108 14680
rect 29164 14671 29204 14680
rect 29259 14720 29301 14729
rect 29259 14680 29260 14720
rect 29300 14680 29301 14720
rect 29259 14671 29301 14680
rect 29356 14720 29396 14729
rect 29260 14586 29300 14671
rect 29356 14561 29396 14680
rect 29452 14720 29492 15091
rect 29452 14671 29492 14680
rect 29355 14552 29397 14561
rect 29355 14512 29356 14552
rect 29396 14512 29397 14552
rect 29355 14503 29397 14512
rect 28875 14344 28876 14384
rect 28916 14344 28917 14384
rect 28875 14335 28917 14344
rect 28972 14344 29108 14384
rect 28532 14008 28820 14048
rect 28492 13999 28532 14008
rect 28300 13914 28340 13999
rect 28684 13376 28724 13385
rect 28684 13217 28724 13336
rect 28300 13208 28340 13217
rect 28204 13168 28300 13208
rect 27916 12832 28148 12872
rect 28204 12982 28244 12991
rect 27819 12788 27861 12797
rect 27819 12748 27820 12788
rect 27860 12748 27861 12788
rect 27819 12739 27861 12748
rect 27820 12704 27860 12739
rect 27820 12653 27860 12664
rect 27723 12620 27765 12629
rect 27723 12580 27724 12620
rect 27764 12580 27765 12620
rect 27723 12571 27765 12580
rect 27916 12536 27956 12832
rect 27916 12487 27956 12496
rect 28012 12536 28052 12545
rect 27723 12452 27765 12461
rect 27723 12412 27724 12452
rect 27764 12412 27765 12452
rect 27723 12403 27765 12412
rect 27532 11948 27572 11957
rect 27436 11908 27532 11948
rect 27532 11899 27572 11908
rect 27339 11696 27381 11705
rect 27339 11656 27340 11696
rect 27380 11656 27381 11696
rect 27339 11647 27381 11656
rect 27627 11612 27669 11621
rect 27627 11572 27628 11612
rect 27668 11572 27669 11612
rect 27627 11563 27669 11572
rect 27531 11528 27573 11537
rect 27531 11488 27532 11528
rect 27572 11488 27573 11528
rect 27531 11479 27573 11488
rect 27340 11024 27380 11033
rect 27243 10940 27285 10949
rect 27243 10900 27244 10940
rect 27284 10900 27285 10940
rect 27243 10891 27285 10900
rect 25707 10268 25749 10277
rect 25707 10228 25708 10268
rect 25748 10228 25749 10268
rect 25707 10219 25749 10228
rect 26955 10268 26997 10277
rect 26955 10228 26956 10268
rect 26996 10228 26997 10268
rect 26955 10219 26997 10228
rect 25420 10135 25460 10144
rect 25516 10184 25556 10193
rect 25323 10100 25365 10109
rect 25323 10060 25324 10100
rect 25364 10060 25365 10100
rect 25323 10051 25365 10060
rect 25324 9966 25364 10051
rect 25131 9848 25173 9857
rect 25131 9808 25132 9848
rect 25172 9808 25268 9848
rect 25131 9799 25173 9808
rect 24844 9724 24980 9764
rect 24844 9512 24884 9523
rect 24844 9437 24884 9472
rect 24940 9512 24980 9724
rect 25131 9680 25173 9689
rect 25131 9640 25132 9680
rect 25172 9640 25173 9680
rect 25131 9631 25173 9640
rect 25132 9546 25172 9631
rect 24940 9463 24980 9472
rect 25036 9512 25076 9521
rect 24843 9428 24885 9437
rect 24843 9388 24844 9428
rect 24884 9388 24885 9428
rect 24843 9379 24885 9388
rect 24652 8968 24788 9008
rect 24652 8765 24692 8968
rect 24844 8924 24884 9379
rect 25036 9269 25076 9472
rect 25228 9428 25268 9808
rect 25516 9689 25556 10144
rect 25611 10184 25653 10193
rect 25611 10144 25612 10184
rect 25652 10144 25653 10184
rect 25611 10135 25653 10144
rect 25612 10050 25652 10135
rect 25515 9680 25557 9689
rect 25515 9640 25516 9680
rect 25556 9640 25557 9680
rect 25515 9631 25557 9640
rect 25324 9512 25364 9523
rect 25324 9437 25364 9472
rect 25515 9512 25557 9521
rect 25515 9472 25516 9512
rect 25556 9472 25557 9512
rect 25515 9463 25557 9472
rect 25132 9388 25268 9428
rect 25323 9428 25365 9437
rect 25323 9388 25324 9428
rect 25364 9388 25365 9428
rect 25035 9260 25077 9269
rect 25035 9220 25036 9260
rect 25076 9220 25077 9260
rect 25035 9211 25077 9220
rect 24940 8924 24980 8933
rect 24844 8884 24940 8924
rect 24940 8875 24980 8884
rect 24747 8840 24789 8849
rect 24747 8800 24748 8840
rect 24788 8800 24789 8840
rect 24747 8791 24789 8800
rect 24651 8756 24693 8765
rect 24651 8716 24652 8756
rect 24692 8716 24693 8756
rect 24651 8707 24693 8716
rect 24556 8623 24596 8632
rect 24748 8672 24788 8791
rect 24939 8756 24981 8765
rect 24939 8716 24940 8756
rect 24980 8716 24981 8756
rect 24939 8707 24981 8716
rect 24748 8623 24788 8632
rect 24651 8504 24693 8513
rect 24651 8464 24652 8504
rect 24692 8464 24693 8504
rect 24651 8455 24693 8464
rect 24652 8370 24692 8455
rect 24843 8336 24885 8345
rect 24843 8296 24844 8336
rect 24884 8296 24885 8336
rect 24843 8287 24885 8296
rect 24651 8252 24693 8261
rect 24651 8212 24652 8252
rect 24692 8212 24693 8252
rect 24651 8203 24693 8212
rect 24555 8168 24597 8177
rect 24555 8128 24556 8168
rect 24596 8128 24597 8168
rect 24555 8119 24597 8128
rect 24460 7757 24500 7960
rect 24556 8000 24596 8119
rect 24556 7925 24596 7960
rect 24652 8000 24692 8203
rect 24652 7951 24692 7960
rect 24747 8000 24789 8009
rect 24747 7960 24748 8000
rect 24788 7960 24789 8000
rect 24747 7951 24789 7960
rect 24555 7916 24597 7925
rect 24555 7876 24556 7916
rect 24596 7876 24597 7916
rect 24555 7867 24597 7876
rect 24748 7866 24788 7951
rect 24459 7748 24501 7757
rect 24459 7708 24460 7748
rect 24500 7708 24501 7748
rect 24459 7699 24501 7708
rect 24651 7664 24693 7673
rect 24651 7624 24652 7664
rect 24692 7624 24693 7664
rect 24651 7615 24693 7624
rect 24555 7580 24597 7589
rect 24555 7540 24556 7580
rect 24596 7540 24597 7580
rect 24555 7531 24597 7540
rect 24459 7496 24501 7505
rect 24459 7456 24460 7496
rect 24500 7456 24501 7496
rect 24459 7447 24501 7456
rect 24460 7337 24500 7447
rect 24459 7328 24501 7337
rect 24459 7288 24460 7328
rect 24500 7288 24501 7328
rect 24459 7279 24501 7288
rect 24556 7253 24596 7531
rect 24555 7244 24597 7253
rect 24555 7204 24556 7244
rect 24596 7204 24597 7244
rect 24555 7195 24597 7204
rect 24364 7111 24404 7120
rect 24460 7160 24500 7169
rect 24460 7001 24500 7120
rect 24556 7160 24596 7195
rect 24556 7110 24596 7120
rect 24652 7160 24692 7615
rect 24652 7111 24692 7120
rect 24747 7160 24789 7169
rect 24747 7120 24748 7160
rect 24788 7120 24789 7160
rect 24747 7111 24789 7120
rect 24844 7160 24884 8287
rect 24940 8000 24980 8707
rect 24940 7832 24980 7960
rect 25036 8672 25076 8681
rect 25132 8672 25172 9388
rect 25323 9379 25365 9388
rect 25516 9378 25556 9463
rect 25323 9260 25365 9269
rect 25323 9220 25324 9260
rect 25364 9220 25365 9260
rect 25323 9211 25365 9220
rect 25420 9260 25460 9269
rect 25076 8632 25172 8672
rect 25036 8000 25076 8632
rect 25131 8504 25173 8513
rect 25131 8464 25132 8504
rect 25172 8464 25173 8504
rect 25131 8455 25173 8464
rect 25036 7951 25076 7960
rect 24940 7792 24981 7832
rect 24941 7748 24981 7792
rect 24844 7111 24884 7120
rect 24940 7708 24981 7748
rect 24459 6992 24501 7001
rect 24459 6952 24460 6992
rect 24500 6952 24501 6992
rect 24459 6943 24501 6952
rect 24268 6784 24500 6824
rect 24116 6448 24212 6488
rect 24267 6488 24309 6497
rect 24267 6448 24268 6488
rect 24308 6448 24309 6488
rect 24076 6439 24116 6448
rect 24267 6439 24309 6448
rect 24460 6488 24500 6784
rect 23788 6355 23828 6364
rect 23691 6320 23733 6329
rect 23691 6280 23692 6320
rect 23732 6280 23733 6320
rect 23691 6271 23733 6280
rect 23884 6320 23924 6439
rect 23979 6404 24021 6413
rect 23979 6364 23980 6404
rect 24020 6364 24021 6404
rect 23979 6355 24021 6364
rect 23884 6271 23924 6280
rect 23980 6270 24020 6355
rect 24268 6354 24308 6439
rect 24171 6320 24213 6329
rect 24171 6280 24172 6320
rect 24212 6280 24213 6320
rect 24171 6271 24213 6280
rect 23308 5944 23540 5984
rect 23020 5599 23060 5608
rect 23212 5648 23252 5657
rect 23115 5480 23157 5489
rect 23115 5440 23116 5480
rect 23156 5440 23157 5480
rect 23115 5431 23157 5440
rect 23116 5346 23156 5431
rect 23019 5312 23061 5321
rect 23019 5272 23020 5312
rect 23060 5272 23061 5312
rect 23019 5263 23061 5272
rect 22732 4927 22772 4936
rect 22924 4976 22964 4985
rect 23020 4976 23060 5263
rect 22964 4936 23060 4976
rect 23116 4976 23156 4987
rect 22924 4927 22964 4936
rect 23116 4901 23156 4936
rect 23115 4892 23157 4901
rect 23115 4852 23116 4892
rect 23156 4852 23157 4892
rect 23115 4843 23157 4852
rect 23212 4817 23252 5608
rect 23308 5648 23348 5657
rect 23308 5405 23348 5608
rect 23500 5648 23540 5944
rect 23979 5816 24021 5825
rect 23979 5776 23980 5816
rect 24020 5776 24021 5816
rect 23979 5767 24021 5776
rect 23500 5599 23540 5608
rect 23595 5648 23637 5657
rect 23595 5608 23596 5648
rect 23636 5608 23637 5648
rect 23595 5599 23637 5608
rect 23788 5648 23828 5659
rect 23596 5514 23636 5599
rect 23788 5573 23828 5608
rect 23980 5648 24020 5767
rect 23980 5599 24020 5608
rect 24075 5648 24117 5657
rect 24075 5608 24076 5648
rect 24116 5608 24117 5648
rect 24075 5599 24117 5608
rect 24172 5648 24212 6271
rect 24267 6236 24309 6245
rect 24267 6196 24268 6236
rect 24308 6196 24309 6236
rect 24267 6187 24309 6196
rect 24268 6102 24308 6187
rect 24364 5657 24404 5742
rect 24172 5599 24212 5608
rect 24363 5648 24405 5657
rect 24460 5648 24500 6448
rect 24748 6413 24788 7111
rect 24940 6908 24980 7708
rect 25132 7673 25172 8455
rect 25227 8336 25269 8345
rect 25227 8296 25228 8336
rect 25268 8296 25269 8336
rect 25227 8287 25269 8296
rect 25228 8168 25268 8287
rect 25228 8119 25268 8128
rect 25227 7916 25269 7925
rect 25227 7876 25228 7916
rect 25268 7876 25269 7916
rect 25227 7867 25269 7876
rect 25131 7664 25173 7673
rect 25131 7624 25132 7664
rect 25172 7624 25173 7664
rect 25131 7615 25173 7624
rect 25036 7412 25076 7421
rect 25131 7412 25173 7421
rect 25076 7372 25132 7412
rect 25172 7372 25173 7412
rect 25036 7363 25076 7372
rect 25131 7363 25173 7372
rect 25228 7412 25268 7867
rect 25324 7673 25364 9211
rect 25420 8261 25460 9220
rect 25708 8672 25748 10219
rect 26668 10184 26708 10193
rect 26572 10100 26612 10109
rect 26572 8924 26612 10060
rect 26668 9101 26708 10144
rect 26956 10184 26996 10219
rect 27340 10193 27380 10984
rect 27532 11024 27572 11479
rect 27532 10975 27572 10984
rect 27628 10856 27668 11563
rect 27724 11024 27764 12403
rect 28012 12284 28052 12496
rect 28108 12536 28148 12547
rect 28108 12461 28148 12496
rect 28204 12536 28244 12942
rect 28300 12704 28340 13168
rect 28396 13208 28436 13217
rect 28396 12881 28436 13168
rect 28491 13208 28533 13217
rect 28491 13168 28492 13208
rect 28532 13168 28533 13208
rect 28491 13159 28533 13168
rect 28683 13208 28725 13217
rect 28683 13168 28684 13208
rect 28724 13168 28725 13208
rect 28683 13159 28725 13168
rect 28395 12872 28437 12881
rect 28395 12832 28396 12872
rect 28436 12832 28437 12872
rect 28395 12823 28437 12832
rect 28492 12713 28532 13159
rect 28876 12872 28916 14335
rect 28972 13040 29012 14344
rect 29355 13376 29397 13385
rect 29355 13336 29356 13376
rect 29396 13336 29397 13376
rect 29355 13327 29397 13336
rect 29067 13292 29109 13301
rect 29067 13252 29068 13292
rect 29108 13252 29109 13292
rect 29067 13243 29109 13252
rect 29068 13208 29108 13243
rect 29068 13157 29108 13168
rect 29164 13208 29204 13217
rect 29164 13049 29204 13168
rect 29260 13208 29300 13217
rect 29163 13040 29205 13049
rect 28972 13000 29108 13040
rect 28684 12832 28916 12872
rect 28491 12704 28533 12713
rect 28300 12664 28436 12704
rect 28300 12536 28340 12545
rect 28204 12496 28300 12536
rect 28107 12452 28149 12461
rect 28107 12412 28108 12452
rect 28148 12412 28149 12452
rect 28107 12403 28149 12412
rect 28204 12284 28244 12496
rect 28300 12487 28340 12496
rect 28396 12536 28436 12664
rect 28491 12664 28492 12704
rect 28532 12664 28533 12704
rect 28491 12655 28533 12664
rect 28396 12461 28436 12496
rect 28491 12536 28533 12545
rect 28491 12496 28492 12536
rect 28532 12496 28533 12536
rect 28491 12487 28533 12496
rect 28588 12536 28628 12547
rect 28395 12452 28437 12461
rect 28395 12412 28396 12452
rect 28436 12412 28437 12452
rect 28395 12403 28437 12412
rect 28012 12244 28244 12284
rect 28011 11696 28053 11705
rect 28011 11656 28012 11696
rect 28052 11656 28053 11696
rect 28011 11647 28053 11656
rect 28012 11562 28052 11647
rect 27724 10975 27764 10984
rect 28107 11024 28149 11033
rect 28107 10984 28108 11024
rect 28148 10984 28149 11024
rect 28107 10975 28149 10984
rect 28108 10890 28148 10975
rect 28012 10856 28052 10865
rect 27628 10816 27764 10856
rect 27724 10697 27764 10816
rect 27723 10688 27765 10697
rect 27723 10648 27724 10688
rect 27764 10648 27765 10688
rect 27723 10639 27765 10648
rect 26956 10133 26996 10144
rect 27051 10184 27093 10193
rect 27051 10144 27052 10184
rect 27092 10144 27093 10184
rect 27051 10135 27093 10144
rect 27339 10184 27381 10193
rect 27339 10144 27340 10184
rect 27380 10144 27381 10184
rect 27339 10135 27381 10144
rect 27724 10184 27764 10639
rect 28012 10352 28052 10816
rect 28012 10312 28148 10352
rect 27724 10135 27764 10144
rect 28011 10184 28053 10193
rect 28011 10144 28012 10184
rect 28052 10144 28053 10184
rect 28011 10135 28053 10144
rect 26859 10100 26901 10109
rect 26859 10060 26860 10100
rect 26900 10060 26901 10100
rect 26859 10051 26901 10060
rect 26667 9092 26709 9101
rect 26667 9052 26668 9092
rect 26708 9052 26709 9092
rect 26667 9043 26709 9052
rect 26572 8884 26804 8924
rect 25516 8632 25708 8672
rect 25419 8252 25461 8261
rect 25419 8212 25420 8252
rect 25460 8212 25461 8252
rect 25419 8203 25461 8212
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 25420 7866 25460 7951
rect 25323 7664 25365 7673
rect 25323 7624 25324 7664
rect 25364 7624 25365 7664
rect 25323 7615 25365 7624
rect 25516 7505 25556 8632
rect 25708 8623 25748 8632
rect 26284 8672 26324 8681
rect 25803 8504 25845 8513
rect 26188 8504 26228 8513
rect 25803 8464 25804 8504
rect 25844 8464 25845 8504
rect 25803 8455 25845 8464
rect 25900 8464 26188 8504
rect 25804 8370 25844 8455
rect 25900 8252 25940 8464
rect 26188 8455 26228 8464
rect 26284 8345 26324 8632
rect 26380 8672 26420 8681
rect 26283 8336 26325 8345
rect 26283 8296 26284 8336
rect 26324 8296 26325 8336
rect 26283 8287 26325 8296
rect 25708 8212 25940 8252
rect 25995 8252 26037 8261
rect 25995 8212 25996 8252
rect 26036 8212 26037 8252
rect 25612 8000 25652 8009
rect 25515 7496 25557 7505
rect 25515 7456 25516 7496
rect 25556 7456 25557 7496
rect 25515 7447 25557 7456
rect 25612 7412 25652 7960
rect 25708 8000 25748 8212
rect 25995 8203 26037 8212
rect 25996 8009 26036 8203
rect 26380 8168 26420 8632
rect 26476 8680 26516 8681
rect 26476 8672 26612 8680
rect 26516 8640 26612 8672
rect 26516 8632 26519 8640
rect 26476 8623 26516 8632
rect 26572 8597 26612 8640
rect 26571 8588 26613 8597
rect 26571 8548 26572 8588
rect 26612 8548 26613 8588
rect 26571 8539 26613 8548
rect 26475 8504 26517 8513
rect 26475 8464 26476 8504
rect 26516 8464 26517 8504
rect 26475 8455 26517 8464
rect 26284 8128 26420 8168
rect 26092 8009 26132 8094
rect 25708 7951 25748 7960
rect 25991 8000 26036 8009
rect 26031 7960 26036 8000
rect 26091 8000 26133 8009
rect 26091 7960 26092 8000
rect 26132 7960 26133 8000
rect 25991 7951 26031 7960
rect 26091 7951 26133 7960
rect 26188 8000 26228 8009
rect 25708 7832 25748 7841
rect 26188 7832 26228 7960
rect 25748 7792 26228 7832
rect 25708 7783 25748 7792
rect 26284 7589 26324 8128
rect 26379 8000 26421 8009
rect 26379 7960 26380 8000
rect 26420 7960 26421 8000
rect 26379 7951 26421 7960
rect 26476 8000 26516 8455
rect 26572 8093 26612 8539
rect 26667 8336 26709 8345
rect 26667 8296 26668 8336
rect 26708 8296 26709 8336
rect 26667 8287 26709 8296
rect 26571 8084 26613 8093
rect 26571 8044 26572 8084
rect 26612 8044 26613 8084
rect 26571 8035 26613 8044
rect 26476 7951 26516 7960
rect 26380 7866 26420 7951
rect 26668 7916 26708 8287
rect 26572 7876 26708 7916
rect 26476 7748 26516 7757
rect 26385 7708 26476 7748
rect 26385 7673 26425 7708
rect 26476 7699 26516 7708
rect 26380 7664 26425 7673
rect 26380 7624 26381 7664
rect 26421 7624 26425 7664
rect 26380 7615 26422 7624
rect 26283 7580 26325 7589
rect 26283 7540 26284 7580
rect 26324 7540 26325 7580
rect 26283 7531 26325 7540
rect 26380 7412 26420 7421
rect 25612 7372 26380 7412
rect 25228 7363 25268 7372
rect 26380 7363 26420 7372
rect 25035 7160 25077 7169
rect 25035 7120 25036 7160
rect 25076 7120 25077 7160
rect 25035 7111 25077 7120
rect 25323 7160 25365 7169
rect 25323 7120 25324 7160
rect 25364 7120 25365 7160
rect 25323 7111 25365 7120
rect 26379 7160 26421 7169
rect 26379 7120 26380 7160
rect 26420 7120 26421 7160
rect 26379 7111 26421 7120
rect 26572 7160 26612 7876
rect 26764 7832 26804 8884
rect 25036 7026 25076 7111
rect 25324 7026 25364 7111
rect 24940 6868 25076 6908
rect 24939 6656 24981 6665
rect 24939 6616 24940 6656
rect 24980 6616 24981 6656
rect 24939 6607 24981 6616
rect 24747 6404 24789 6413
rect 24747 6364 24748 6404
rect 24788 6364 24789 6404
rect 24747 6355 24789 6364
rect 24555 6320 24597 6329
rect 24555 6280 24556 6320
rect 24596 6280 24597 6320
rect 24555 6271 24597 6280
rect 24363 5608 24364 5648
rect 24404 5608 24500 5648
rect 24556 5648 24596 6271
rect 24363 5599 24405 5608
rect 24556 5599 24596 5608
rect 24748 5648 24788 6355
rect 24843 5732 24885 5741
rect 24843 5692 24844 5732
rect 24884 5692 24885 5732
rect 24843 5683 24885 5692
rect 24748 5599 24788 5608
rect 23787 5564 23829 5573
rect 23787 5524 23788 5564
rect 23828 5524 23829 5564
rect 23787 5515 23829 5524
rect 24076 5514 24116 5599
rect 24844 5598 24884 5683
rect 24940 5648 24980 6607
rect 24940 5599 24980 5608
rect 23692 5480 23732 5489
rect 24460 5480 24500 5489
rect 25036 5480 25076 6868
rect 26380 5909 26420 7111
rect 26572 7085 26612 7120
rect 26668 7792 26804 7832
rect 26571 7076 26613 7085
rect 26571 7036 26572 7076
rect 26612 7036 26613 7076
rect 26571 7027 26613 7036
rect 26572 6996 26612 7027
rect 26668 6572 26708 7792
rect 26763 7664 26805 7673
rect 26763 7624 26764 7664
rect 26804 7624 26805 7664
rect 26763 7615 26805 7624
rect 26476 6532 26708 6572
rect 26379 5900 26421 5909
rect 26379 5860 26380 5900
rect 26420 5860 26421 5900
rect 26379 5851 26421 5860
rect 26476 5648 26516 6532
rect 26571 6404 26613 6413
rect 26571 6364 26572 6404
rect 26612 6364 26613 6404
rect 26571 6355 26613 6364
rect 26285 5633 26325 5642
rect 26285 5564 26325 5593
rect 23307 5396 23349 5405
rect 23307 5356 23308 5396
rect 23348 5356 23349 5396
rect 23307 5347 23349 5356
rect 23595 5396 23637 5405
rect 23595 5356 23596 5396
rect 23636 5356 23637 5396
rect 23595 5347 23637 5356
rect 23298 5060 23340 5069
rect 23403 5060 23445 5069
rect 23298 5020 23299 5060
rect 23339 5020 23348 5060
rect 23298 5011 23348 5020
rect 23403 5020 23404 5060
rect 23444 5020 23445 5060
rect 23403 5011 23445 5020
rect 23308 4976 23348 5011
rect 23211 4808 23253 4817
rect 23211 4768 23212 4808
rect 23252 4768 23253 4808
rect 23211 4759 23253 4768
rect 22732 4724 22772 4733
rect 23116 4724 23156 4733
rect 22252 4304 22292 4313
rect 22156 4264 22252 4304
rect 22059 4052 22101 4061
rect 22059 4012 22060 4052
rect 22100 4012 22101 4052
rect 22059 4003 22101 4012
rect 22156 2624 22196 4264
rect 22252 4255 22292 4264
rect 22732 4229 22772 4684
rect 23020 4684 23116 4724
rect 22923 4388 22965 4397
rect 22923 4348 22924 4388
rect 22964 4348 22965 4388
rect 22923 4339 22965 4348
rect 22731 4220 22773 4229
rect 22731 4180 22732 4220
rect 22772 4180 22773 4220
rect 22731 4171 22773 4180
rect 22924 4220 22964 4339
rect 22924 4171 22964 4180
rect 22156 2575 22196 2584
rect 22444 3464 22484 3473
rect 22444 2129 22484 3424
rect 22636 3464 22676 3473
rect 22636 2801 22676 3424
rect 22731 3464 22773 3473
rect 22731 3424 22732 3464
rect 22772 3424 22773 3464
rect 22731 3415 22773 3424
rect 22924 3464 22964 3473
rect 23020 3464 23060 4684
rect 23116 4675 23156 4684
rect 23308 3809 23348 4936
rect 23404 4976 23444 5011
rect 23596 4976 23636 5347
rect 23692 5321 23732 5440
rect 24172 5440 24460 5480
rect 23691 5312 23733 5321
rect 23691 5272 23692 5312
rect 23732 5272 23733 5312
rect 23691 5263 23733 5272
rect 23883 5060 23925 5069
rect 23883 5020 23884 5060
rect 23924 5020 23925 5060
rect 23883 5011 23925 5020
rect 23692 4976 23732 4985
rect 23596 4936 23692 4976
rect 23404 4925 23444 4936
rect 23692 4927 23732 4936
rect 23788 4976 23828 4985
rect 23788 4733 23828 4936
rect 23884 4926 23924 5011
rect 23980 4976 24020 4985
rect 24172 4976 24212 5440
rect 24460 5431 24500 5440
rect 24940 5440 25076 5480
rect 26284 5524 26325 5564
rect 26373 5634 26516 5648
rect 26373 5594 26380 5634
rect 26420 5608 26516 5634
rect 26572 5648 26612 6355
rect 26764 5984 26804 7615
rect 26572 5599 26612 5608
rect 26668 5944 26804 5984
rect 26373 5580 26420 5594
rect 24020 4936 24212 4976
rect 24268 5144 24308 5153
rect 23980 4927 24020 4936
rect 24268 4901 24308 5104
rect 24364 5060 24404 5069
rect 24267 4892 24309 4901
rect 24267 4852 24268 4892
rect 24308 4852 24309 4892
rect 24267 4843 24309 4852
rect 23787 4724 23829 4733
rect 23787 4684 23788 4724
rect 23828 4684 23829 4724
rect 23787 4675 23829 4684
rect 23499 4640 23541 4649
rect 23499 4600 23500 4640
rect 23540 4600 23541 4640
rect 23499 4591 23541 4600
rect 23500 4388 23540 4591
rect 23595 4556 23637 4565
rect 23595 4516 23596 4556
rect 23636 4516 23637 4556
rect 23595 4507 23637 4516
rect 23500 4339 23540 4348
rect 23596 4313 23636 4507
rect 24364 4388 24404 5020
rect 24459 5060 24501 5069
rect 24651 5060 24693 5069
rect 24459 5020 24460 5060
rect 24500 5020 24501 5060
rect 24459 5011 24501 5020
rect 24556 5020 24652 5060
rect 24692 5020 24693 5060
rect 24460 4976 24500 5011
rect 24460 4925 24500 4936
rect 24556 4976 24596 5020
rect 24651 5011 24693 5020
rect 24843 5060 24885 5069
rect 24843 5020 24844 5060
rect 24884 5020 24885 5060
rect 24843 5011 24885 5020
rect 24556 4927 24596 4936
rect 24748 4976 24788 4985
rect 24460 4808 24500 4817
rect 24748 4808 24788 4936
rect 24500 4768 24788 4808
rect 24460 4759 24500 4768
rect 24556 4388 24596 4397
rect 24364 4348 24556 4388
rect 24556 4339 24596 4348
rect 24844 4313 24884 5011
rect 24940 4565 24980 5440
rect 26284 5405 26324 5524
rect 26373 5489 26413 5580
rect 26373 5480 26421 5489
rect 26373 5440 26380 5480
rect 26420 5440 26421 5480
rect 26379 5431 26421 5440
rect 26476 5480 26516 5489
rect 26668 5480 26708 5944
rect 26860 5900 26900 10051
rect 27052 9680 27092 10135
rect 28012 10050 28052 10135
rect 27052 9631 27092 9640
rect 27916 9596 27956 9605
rect 26956 9512 26996 9523
rect 26956 9437 26996 9472
rect 27244 9512 27284 9521
rect 26955 9428 26997 9437
rect 26955 9388 26956 9428
rect 26996 9388 26997 9428
rect 26955 9379 26997 9388
rect 27244 9008 27284 9472
rect 27435 9512 27477 9521
rect 27435 9472 27436 9512
rect 27476 9472 27477 9512
rect 27435 9463 27477 9472
rect 27820 9512 27860 9521
rect 27436 9378 27476 9463
rect 27244 8968 27572 9008
rect 27238 8840 27280 8849
rect 27238 8800 27239 8840
rect 27279 8800 27280 8840
rect 27238 8791 27280 8800
rect 27239 8672 27279 8791
rect 27340 8672 27380 8681
rect 27279 8632 27284 8672
rect 27239 8623 27284 8632
rect 27244 8168 27284 8623
rect 27340 8345 27380 8632
rect 27435 8672 27477 8681
rect 27435 8632 27436 8672
rect 27476 8632 27477 8672
rect 27435 8623 27477 8632
rect 27436 8538 27476 8623
rect 27532 8504 27572 8968
rect 27723 8840 27765 8849
rect 27820 8840 27860 9472
rect 27916 9437 27956 9556
rect 27915 9428 27957 9437
rect 27915 9388 27916 9428
rect 27956 9388 27957 9428
rect 27915 9379 27957 9388
rect 27723 8800 27724 8840
rect 27764 8800 27860 8840
rect 28011 8840 28053 8849
rect 28108 8840 28148 10312
rect 28204 10100 28244 12244
rect 28299 11780 28341 11789
rect 28299 11740 28300 11780
rect 28340 11740 28341 11780
rect 28299 11731 28341 11740
rect 28300 11696 28340 11731
rect 28300 11645 28340 11656
rect 28492 11696 28532 12487
rect 28588 12461 28628 12496
rect 28587 12452 28629 12461
rect 28587 12412 28588 12452
rect 28628 12412 28629 12452
rect 28587 12403 28629 12412
rect 28492 11647 28532 11656
rect 28395 11528 28437 11537
rect 28395 11488 28396 11528
rect 28436 11488 28437 11528
rect 28395 11479 28437 11488
rect 28396 11394 28436 11479
rect 28204 10051 28244 10060
rect 28395 10100 28437 10109
rect 28395 10060 28396 10100
rect 28436 10060 28437 10100
rect 28395 10051 28437 10060
rect 28299 9428 28341 9437
rect 28299 9388 28300 9428
rect 28340 9388 28341 9428
rect 28299 9379 28341 9388
rect 28396 9428 28436 10051
rect 28396 9379 28436 9388
rect 28492 9512 28532 9521
rect 28203 9344 28245 9353
rect 28203 9304 28204 9344
rect 28244 9304 28245 9344
rect 28203 9295 28245 9304
rect 28300 9344 28340 9379
rect 28204 9210 28244 9295
rect 28300 9293 28340 9304
rect 28492 8840 28532 9472
rect 28587 9512 28629 9521
rect 28587 9472 28588 9512
rect 28628 9472 28629 9512
rect 28587 9463 28629 9472
rect 28588 9378 28628 9463
rect 28011 8800 28012 8840
rect 28052 8800 28148 8840
rect 28300 8800 28532 8840
rect 27723 8791 27765 8800
rect 28011 8791 28053 8800
rect 28300 8756 28340 8800
rect 28211 8716 28340 8756
rect 28492 8756 28532 8800
rect 28588 8765 28628 8796
rect 27628 8672 27668 8681
rect 27628 8513 27668 8632
rect 27723 8672 27765 8681
rect 27723 8632 27724 8672
rect 27764 8632 27765 8672
rect 27723 8623 27765 8632
rect 27916 8668 27956 8677
rect 27724 8538 27764 8623
rect 27532 8455 27572 8464
rect 27627 8504 27669 8513
rect 27627 8464 27628 8504
rect 27668 8464 27669 8504
rect 27627 8455 27669 8464
rect 27339 8336 27381 8345
rect 27339 8296 27340 8336
rect 27380 8296 27381 8336
rect 27339 8287 27381 8296
rect 27531 8168 27573 8177
rect 27244 8128 27476 8168
rect 27436 8009 27476 8128
rect 27531 8128 27532 8168
rect 27572 8128 27573 8168
rect 27531 8119 27573 8128
rect 27051 8000 27093 8009
rect 27051 7960 27052 8000
rect 27092 7960 27093 8000
rect 27051 7951 27093 7960
rect 27148 8000 27188 8009
rect 27052 7866 27092 7951
rect 27148 7421 27188 7960
rect 27243 8000 27285 8009
rect 27243 7960 27244 8000
rect 27284 7960 27285 8000
rect 27243 7951 27285 7960
rect 27340 8000 27380 8009
rect 27244 7866 27284 7951
rect 27147 7412 27189 7421
rect 27147 7372 27148 7412
rect 27188 7372 27189 7412
rect 27147 7363 27189 7372
rect 27340 7244 27380 7960
rect 27435 8000 27477 8009
rect 27435 7960 27436 8000
rect 27476 7960 27477 8000
rect 27435 7951 27477 7960
rect 27532 8000 27572 8119
rect 27532 7951 27572 7960
rect 27628 7580 27668 8455
rect 27916 8345 27956 8628
rect 28011 8672 28053 8681
rect 28211 8677 28251 8716
rect 28492 8707 28532 8716
rect 28587 8756 28629 8765
rect 28587 8716 28588 8756
rect 28628 8716 28629 8756
rect 28587 8707 28629 8716
rect 28011 8632 28012 8672
rect 28052 8632 28053 8672
rect 28011 8623 28053 8632
rect 28115 8668 28155 8677
rect 28211 8628 28251 8637
rect 28396 8672 28436 8681
rect 28012 8538 28052 8623
rect 28115 8504 28155 8628
rect 28396 8513 28436 8632
rect 28588 8672 28628 8707
rect 28588 8597 28628 8632
rect 28587 8588 28629 8597
rect 28587 8548 28588 8588
rect 28628 8548 28629 8588
rect 28587 8539 28629 8548
rect 28108 8464 28155 8504
rect 28395 8504 28437 8513
rect 28395 8464 28396 8504
rect 28436 8464 28437 8504
rect 27915 8336 27957 8345
rect 27915 8296 27916 8336
rect 27956 8296 27957 8336
rect 27915 8287 27957 8296
rect 27819 8000 27861 8009
rect 27819 7960 27820 8000
rect 27860 7960 27861 8000
rect 27819 7951 27861 7960
rect 27820 7757 27860 7951
rect 27819 7748 27861 7757
rect 27819 7708 27820 7748
rect 27860 7708 27861 7748
rect 27819 7699 27861 7708
rect 27340 7195 27380 7204
rect 27532 7540 27668 7580
rect 27819 7580 27861 7589
rect 27819 7540 27820 7580
rect 27860 7540 27861 7580
rect 27147 7160 27189 7169
rect 27147 7120 27148 7160
rect 27188 7120 27189 7160
rect 27147 7111 27189 7120
rect 27435 7160 27477 7169
rect 27435 7120 27436 7160
rect 27476 7120 27477 7160
rect 27532 7160 27572 7540
rect 27819 7531 27861 7540
rect 27627 7412 27669 7421
rect 27724 7412 27764 7421
rect 27627 7372 27628 7412
rect 27668 7372 27724 7412
rect 27627 7363 27669 7372
rect 27724 7363 27764 7372
rect 27628 7160 27668 7169
rect 27532 7120 27628 7160
rect 27435 7111 27477 7120
rect 27628 7111 27668 7120
rect 27820 7160 27860 7531
rect 27148 7026 27188 7111
rect 27243 6992 27285 7001
rect 27243 6952 27244 6992
rect 27284 6952 27285 6992
rect 27243 6943 27285 6952
rect 27244 6488 27284 6943
rect 27436 6656 27476 7111
rect 27820 6917 27860 7120
rect 27819 6908 27861 6917
rect 27819 6868 27820 6908
rect 27860 6868 27861 6908
rect 27819 6859 27861 6868
rect 27244 6439 27284 6448
rect 27340 6616 27476 6656
rect 27340 6404 27380 6616
rect 27627 6572 27669 6581
rect 27627 6532 27628 6572
rect 27668 6532 27669 6572
rect 27627 6523 27669 6532
rect 27531 6488 27573 6497
rect 27531 6448 27532 6488
rect 27572 6448 27573 6488
rect 27531 6439 27573 6448
rect 27628 6488 27668 6523
rect 27340 6355 27380 6364
rect 27532 6404 27572 6439
rect 27628 6437 27668 6448
rect 27916 6404 27956 8287
rect 28108 8177 28148 8464
rect 28395 8455 28437 8464
rect 28107 8168 28149 8177
rect 28107 8128 28108 8168
rect 28148 8128 28149 8168
rect 28107 8119 28149 8128
rect 28203 7244 28245 7253
rect 28203 7204 28204 7244
rect 28244 7204 28245 7244
rect 28203 7195 28245 7204
rect 28204 6497 28244 7195
rect 28395 6740 28437 6749
rect 28395 6700 28396 6740
rect 28436 6700 28437 6740
rect 28395 6691 28437 6700
rect 28203 6488 28245 6497
rect 28203 6448 28204 6488
rect 28244 6448 28245 6488
rect 28203 6439 28245 6448
rect 28396 6488 28436 6691
rect 28684 6656 28724 12832
rect 28779 12704 28821 12713
rect 28779 12664 28780 12704
rect 28820 12664 28821 12704
rect 28779 12655 28821 12664
rect 28780 12536 28820 12655
rect 28971 12620 29013 12629
rect 28971 12580 28972 12620
rect 29012 12580 29013 12620
rect 28971 12571 29013 12580
rect 28780 12487 28820 12496
rect 28875 12536 28917 12545
rect 28875 12496 28876 12536
rect 28916 12496 28917 12536
rect 28875 12487 28917 12496
rect 28876 12402 28916 12487
rect 28972 12486 29012 12571
rect 29068 12545 29108 13000
rect 29163 13000 29164 13040
rect 29204 13000 29205 13040
rect 29163 12991 29205 13000
rect 29260 12704 29300 13168
rect 29356 13208 29396 13327
rect 29548 13208 29588 15595
rect 29644 15560 29684 16024
rect 29836 15980 29876 16099
rect 29644 15511 29684 15520
rect 29740 15940 29876 15980
rect 29740 15560 29780 15940
rect 30124 15737 30164 18712
rect 30316 18584 30356 19048
rect 30316 18535 30356 18544
rect 30508 18584 30548 18593
rect 30315 18332 30357 18341
rect 30315 18292 30316 18332
rect 30356 18292 30357 18332
rect 30315 18283 30357 18292
rect 30316 18198 30356 18283
rect 30508 18005 30548 18544
rect 31563 18332 31605 18341
rect 31563 18292 31564 18332
rect 31604 18292 31605 18332
rect 31563 18283 31605 18292
rect 30507 17996 30549 18005
rect 30507 17956 30508 17996
rect 30548 17956 30549 17996
rect 30507 17947 30549 17956
rect 31179 17996 31221 18005
rect 31179 17956 31180 17996
rect 31220 17956 31221 17996
rect 31179 17947 31221 17956
rect 30699 17912 30741 17921
rect 30988 17912 31028 17921
rect 30699 17872 30700 17912
rect 30740 17872 30741 17912
rect 30699 17863 30741 17872
rect 30796 17872 30988 17912
rect 30508 17744 30548 17753
rect 30316 17704 30508 17744
rect 30219 16820 30261 16829
rect 30219 16780 30220 16820
rect 30260 16780 30261 16820
rect 30219 16771 30261 16780
rect 30220 16325 30260 16771
rect 30219 16316 30261 16325
rect 30219 16276 30220 16316
rect 30260 16276 30261 16316
rect 30219 16267 30261 16276
rect 30316 15905 30356 17704
rect 30508 17695 30548 17704
rect 30700 17744 30740 17863
rect 30700 17695 30740 17704
rect 30796 17744 30836 17872
rect 30988 17863 31028 17872
rect 30796 17695 30836 17704
rect 30987 17744 31029 17753
rect 30987 17704 30988 17744
rect 31028 17704 31029 17744
rect 30987 17695 31029 17704
rect 31180 17744 31220 17947
rect 31180 17695 31220 17704
rect 30988 17610 31028 17695
rect 30604 17576 30644 17585
rect 30412 17536 30604 17576
rect 30412 17072 30452 17536
rect 30604 17527 30644 17536
rect 31564 17156 31604 18283
rect 31851 18080 31893 18089
rect 31851 18040 31852 18080
rect 31892 18040 31893 18080
rect 31851 18031 31893 18040
rect 31852 17744 31892 18031
rect 32044 17828 32084 20056
rect 32908 19517 32948 20140
rect 33004 19928 33044 19937
rect 32907 19508 32949 19517
rect 32907 19468 32908 19508
rect 32948 19468 32949 19508
rect 32907 19459 32949 19468
rect 32332 19424 32372 19433
rect 32372 19384 32564 19424
rect 32332 19375 32372 19384
rect 32139 19256 32181 19265
rect 32139 19216 32140 19256
rect 32180 19216 32181 19256
rect 32139 19207 32181 19216
rect 32332 19256 32372 19265
rect 32140 18668 32180 19207
rect 32332 18761 32372 19216
rect 32524 19256 32564 19384
rect 32524 19207 32564 19216
rect 32908 19256 32948 19265
rect 33004 19256 33044 19888
rect 33772 19928 33812 19937
rect 33812 19888 33908 19928
rect 33772 19879 33812 19888
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 32948 19216 33044 19256
rect 33772 19256 33812 19265
rect 32908 19207 32948 19216
rect 32811 19004 32853 19013
rect 32811 18964 32812 19004
rect 32852 18964 32853 19004
rect 32811 18955 32853 18964
rect 32331 18752 32373 18761
rect 32331 18712 32332 18752
rect 32372 18712 32373 18752
rect 32331 18703 32373 18712
rect 32140 18619 32180 18628
rect 32427 18584 32469 18593
rect 32427 18544 32428 18584
rect 32468 18544 32469 18584
rect 32427 18535 32469 18544
rect 32524 18584 32564 18593
rect 32428 17912 32468 18535
rect 32044 17788 32180 17828
rect 31892 17704 32084 17744
rect 31852 17695 31892 17704
rect 31468 17116 31604 17156
rect 30412 17023 30452 17032
rect 30508 17072 30548 17081
rect 30508 16409 30548 17032
rect 30700 17072 30740 17081
rect 30892 17072 30932 17081
rect 30740 17032 30892 17072
rect 30700 17023 30740 17032
rect 30892 17023 30932 17032
rect 30987 17072 31029 17081
rect 30987 17032 30988 17072
rect 31028 17032 31029 17072
rect 30987 17023 31029 17032
rect 31084 17072 31124 17081
rect 30988 16938 31028 17023
rect 30699 16904 30741 16913
rect 30699 16864 30700 16904
rect 30740 16864 30741 16904
rect 30699 16855 30741 16864
rect 30700 16770 30740 16855
rect 31084 16661 31124 17032
rect 31180 17072 31220 17081
rect 31083 16652 31125 16661
rect 31083 16612 31084 16652
rect 31124 16612 31125 16652
rect 31083 16603 31125 16612
rect 30507 16400 30549 16409
rect 31084 16400 31124 16603
rect 31180 16568 31220 17032
rect 31372 17072 31412 17083
rect 31372 16997 31412 17032
rect 31468 17072 31508 17116
rect 31468 17023 31508 17032
rect 31371 16988 31413 16997
rect 31371 16948 31372 16988
rect 31412 16948 31413 16988
rect 31371 16939 31413 16948
rect 31564 16988 31604 16997
rect 31180 16528 31412 16568
rect 30507 16360 30508 16400
rect 30548 16360 30549 16400
rect 30507 16351 30549 16360
rect 30988 16360 31124 16400
rect 31179 16400 31221 16409
rect 31179 16360 31180 16400
rect 31220 16360 31221 16400
rect 30891 16316 30933 16325
rect 30891 16276 30892 16316
rect 30932 16276 30933 16316
rect 30891 16267 30933 16276
rect 30412 16232 30452 16241
rect 30315 15896 30357 15905
rect 30315 15856 30316 15896
rect 30356 15856 30357 15896
rect 30315 15847 30357 15856
rect 30219 15812 30261 15821
rect 30219 15772 30220 15812
rect 30260 15772 30261 15812
rect 30219 15763 30261 15772
rect 29932 15728 29972 15737
rect 30123 15728 30165 15737
rect 29972 15688 30068 15728
rect 29932 15679 29972 15688
rect 29740 15401 29780 15520
rect 29836 15644 29876 15653
rect 29739 15392 29781 15401
rect 29739 15352 29740 15392
rect 29780 15352 29781 15392
rect 29739 15343 29781 15352
rect 29739 15224 29781 15233
rect 29739 15184 29740 15224
rect 29780 15184 29781 15224
rect 29739 15175 29781 15184
rect 29643 14720 29685 14729
rect 29643 14680 29644 14720
rect 29684 14680 29685 14720
rect 29643 14671 29685 14680
rect 29740 14720 29780 15175
rect 29836 15065 29876 15604
rect 29931 15392 29973 15401
rect 29931 15352 29932 15392
rect 29972 15352 29973 15392
rect 29931 15343 29973 15352
rect 29932 15258 29972 15343
rect 29835 15056 29877 15065
rect 29835 15016 29836 15056
rect 29876 15016 29877 15056
rect 29835 15007 29877 15016
rect 29931 14888 29973 14897
rect 29931 14848 29932 14888
rect 29972 14848 29973 14888
rect 29931 14839 29973 14848
rect 29835 14804 29877 14813
rect 29835 14764 29836 14804
rect 29876 14764 29877 14804
rect 29835 14755 29877 14764
rect 29644 14586 29684 14671
rect 29740 14141 29780 14680
rect 29836 14636 29876 14755
rect 29932 14720 29972 14839
rect 29932 14671 29972 14680
rect 29836 14587 29876 14596
rect 29931 14216 29973 14225
rect 29931 14176 29932 14216
rect 29972 14176 29973 14216
rect 29931 14167 29973 14176
rect 29739 14132 29781 14141
rect 29739 14092 29740 14132
rect 29780 14092 29781 14132
rect 29739 14083 29781 14092
rect 29835 13964 29877 13973
rect 29835 13924 29836 13964
rect 29876 13924 29877 13964
rect 29835 13915 29877 13924
rect 29740 13376 29780 13385
rect 29356 13159 29396 13168
rect 29452 13168 29588 13208
rect 29644 13336 29740 13376
rect 29452 12965 29492 13168
rect 29547 13040 29589 13049
rect 29547 13000 29548 13040
rect 29588 13000 29589 13040
rect 29547 12991 29589 13000
rect 29451 12956 29493 12965
rect 29451 12916 29452 12956
rect 29492 12916 29493 12956
rect 29451 12907 29493 12916
rect 29548 12906 29588 12991
rect 29164 12664 29300 12704
rect 29067 12536 29109 12545
rect 29067 12496 29068 12536
rect 29108 12496 29109 12536
rect 29067 12487 29109 12496
rect 29067 12368 29109 12377
rect 29067 12328 29068 12368
rect 29108 12328 29109 12368
rect 29067 12319 29109 12328
rect 28779 12200 28821 12209
rect 28779 12160 28780 12200
rect 28820 12160 28821 12200
rect 28779 12151 28821 12160
rect 28780 11360 28820 12151
rect 28875 11864 28917 11873
rect 29068 11864 29108 12319
rect 29164 12200 29204 12664
rect 29260 12536 29300 12545
rect 29260 12377 29300 12496
rect 29452 12536 29492 12545
rect 29355 12452 29397 12461
rect 29355 12412 29356 12452
rect 29396 12412 29397 12452
rect 29355 12403 29397 12412
rect 29259 12368 29301 12377
rect 29259 12328 29260 12368
rect 29300 12328 29301 12368
rect 29259 12319 29301 12328
rect 29356 12318 29396 12403
rect 29164 12160 29396 12200
rect 28875 11824 28876 11864
rect 28916 11824 29108 11864
rect 28875 11815 28917 11824
rect 28876 11696 28916 11815
rect 28876 11647 28916 11656
rect 29068 11696 29108 11705
rect 28972 11528 29012 11537
rect 28780 11320 28916 11360
rect 28876 10856 28916 11320
rect 28972 11033 29012 11488
rect 28971 11024 29013 11033
rect 28971 10984 28972 11024
rect 29012 10984 29013 11024
rect 28971 10975 29013 10984
rect 29068 10865 29108 11656
rect 29164 11696 29204 11705
rect 29164 11537 29204 11656
rect 29163 11528 29205 11537
rect 29163 11488 29164 11528
rect 29204 11488 29205 11528
rect 29163 11479 29205 11488
rect 29163 11276 29205 11285
rect 29163 11236 29164 11276
rect 29204 11236 29205 11276
rect 29163 11227 29205 11236
rect 29164 11108 29204 11227
rect 29164 11059 29204 11068
rect 29260 11024 29300 11033
rect 28876 10807 28916 10816
rect 29067 10856 29109 10865
rect 29067 10816 29068 10856
rect 29108 10816 29109 10856
rect 29067 10807 29109 10816
rect 29260 10361 29300 10984
rect 29356 10436 29396 12160
rect 29452 11537 29492 12496
rect 29451 11528 29493 11537
rect 29451 11488 29452 11528
rect 29492 11488 29493 11528
rect 29451 11479 29493 11488
rect 29644 11360 29684 13336
rect 29740 13327 29780 13336
rect 29740 13208 29780 13217
rect 29836 13208 29876 13915
rect 29780 13168 29876 13208
rect 29740 13159 29780 13168
rect 29739 13040 29781 13049
rect 29739 13000 29740 13040
rect 29780 13000 29781 13040
rect 29739 12991 29781 13000
rect 29740 11453 29780 12991
rect 29836 12377 29876 13168
rect 29835 12368 29877 12377
rect 29835 12328 29836 12368
rect 29876 12328 29877 12368
rect 29835 12319 29877 12328
rect 29739 11444 29781 11453
rect 29739 11404 29740 11444
rect 29780 11404 29781 11444
rect 29739 11395 29781 11404
rect 29548 11320 29684 11360
rect 29932 11360 29972 14167
rect 30028 13889 30068 15688
rect 30123 15688 30124 15728
rect 30164 15688 30165 15728
rect 30123 15679 30165 15688
rect 30220 15401 30260 15763
rect 30315 15560 30357 15569
rect 30315 15520 30316 15560
rect 30356 15520 30357 15560
rect 30315 15511 30357 15520
rect 30316 15426 30356 15511
rect 30219 15392 30261 15401
rect 30219 15352 30220 15392
rect 30260 15352 30261 15392
rect 30219 15343 30261 15352
rect 30412 15149 30452 16192
rect 30507 16232 30549 16241
rect 30507 16192 30508 16232
rect 30548 16192 30549 16232
rect 30507 16183 30549 16192
rect 30700 16232 30740 16241
rect 30740 16192 30836 16232
rect 30700 16183 30740 16192
rect 30508 16098 30548 16183
rect 30700 16064 30740 16073
rect 30700 15569 30740 16024
rect 30796 15653 30836 16192
rect 30795 15644 30837 15653
rect 30795 15604 30796 15644
rect 30836 15604 30837 15644
rect 30795 15595 30837 15604
rect 30699 15560 30741 15569
rect 30699 15520 30700 15560
rect 30740 15520 30741 15560
rect 30699 15511 30741 15520
rect 30699 15392 30741 15401
rect 30699 15352 30700 15392
rect 30740 15352 30741 15392
rect 30699 15343 30741 15352
rect 30604 15308 30644 15317
rect 30508 15268 30604 15308
rect 30411 15140 30453 15149
rect 30411 15100 30412 15140
rect 30452 15100 30453 15140
rect 30411 15091 30453 15100
rect 30315 15056 30357 15065
rect 30315 15016 30316 15056
rect 30356 15016 30357 15056
rect 30315 15007 30357 15016
rect 30220 14048 30260 14057
rect 30027 13880 30069 13889
rect 30027 13840 30028 13880
rect 30068 13840 30069 13880
rect 30027 13831 30069 13840
rect 30028 13208 30068 13831
rect 30220 13721 30260 14008
rect 30316 14048 30356 15007
rect 30508 14645 30548 15268
rect 30604 15259 30644 15268
rect 30700 14804 30740 15343
rect 30892 15233 30932 16267
rect 30988 16157 31028 16360
rect 31179 16351 31221 16360
rect 31180 16266 31220 16351
rect 31372 16325 31412 16528
rect 31564 16409 31604 16948
rect 31660 16904 31700 16913
rect 31563 16400 31605 16409
rect 31563 16360 31564 16400
rect 31604 16360 31605 16400
rect 31563 16351 31605 16360
rect 31371 16316 31413 16325
rect 31371 16276 31372 16316
rect 31412 16276 31413 16316
rect 31371 16267 31413 16276
rect 31083 16232 31125 16241
rect 31083 16192 31084 16232
rect 31124 16192 31125 16232
rect 31083 16183 31125 16192
rect 31276 16232 31316 16243
rect 30987 16148 31029 16157
rect 30987 16108 30988 16148
rect 31028 16108 31029 16148
rect 30987 16099 31029 16108
rect 31084 16098 31124 16183
rect 31276 16157 31316 16192
rect 31275 16148 31317 16157
rect 31275 16108 31276 16148
rect 31316 16108 31317 16148
rect 31275 16099 31317 16108
rect 31468 16064 31508 16073
rect 31372 16024 31468 16064
rect 31372 15896 31412 16024
rect 31468 16015 31508 16024
rect 31563 16064 31605 16073
rect 31563 16024 31564 16064
rect 31604 16024 31605 16064
rect 31563 16015 31605 16024
rect 30988 15856 31412 15896
rect 31467 15896 31509 15905
rect 31467 15856 31468 15896
rect 31508 15856 31509 15896
rect 30891 15224 30933 15233
rect 30891 15184 30892 15224
rect 30932 15184 30933 15224
rect 30891 15175 30933 15184
rect 30795 15056 30837 15065
rect 30795 15016 30796 15056
rect 30836 15016 30837 15056
rect 30795 15007 30837 15016
rect 30700 14755 30740 14764
rect 30507 14636 30549 14645
rect 30507 14596 30508 14636
rect 30548 14596 30549 14636
rect 30507 14587 30549 14596
rect 30316 13999 30356 14008
rect 30411 14048 30453 14057
rect 30411 14008 30412 14048
rect 30452 14008 30453 14048
rect 30411 13999 30453 14008
rect 30508 14048 30548 14587
rect 30796 14477 30836 15007
rect 30891 14972 30933 14981
rect 30891 14932 30892 14972
rect 30932 14932 30933 14972
rect 30891 14923 30933 14932
rect 30892 14838 30932 14923
rect 30891 14720 30933 14729
rect 30891 14680 30892 14720
rect 30932 14680 30933 14720
rect 30891 14671 30933 14680
rect 30795 14468 30837 14477
rect 30795 14428 30796 14468
rect 30836 14428 30837 14468
rect 30795 14419 30837 14428
rect 30412 13914 30452 13999
rect 30508 13889 30548 14008
rect 30699 14048 30741 14057
rect 30699 14008 30700 14048
rect 30740 14008 30741 14048
rect 30699 13999 30741 14008
rect 30507 13880 30549 13889
rect 30507 13840 30508 13880
rect 30548 13840 30549 13880
rect 30507 13831 30549 13840
rect 30219 13712 30261 13721
rect 30219 13672 30220 13712
rect 30260 13672 30261 13712
rect 30219 13663 30261 13672
rect 30123 13460 30165 13469
rect 30604 13460 30644 13469
rect 30123 13420 30124 13460
rect 30164 13420 30165 13460
rect 30123 13411 30165 13420
rect 30508 13420 30604 13460
rect 30124 13326 30164 13411
rect 30508 13292 30548 13420
rect 30604 13411 30644 13420
rect 30412 13252 30548 13292
rect 30304 13208 30346 13217
rect 30028 13168 30260 13208
rect 30220 13124 30260 13168
rect 30304 13168 30305 13208
rect 30345 13168 30346 13208
rect 30304 13159 30346 13168
rect 30412 13208 30452 13252
rect 30604 13217 30644 13302
rect 30412 13159 30452 13168
rect 30603 13208 30645 13217
rect 30603 13168 30604 13208
rect 30644 13168 30645 13208
rect 30603 13159 30645 13168
rect 30220 13075 30260 13084
rect 30305 13074 30345 13159
rect 30124 13040 30164 13049
rect 30027 12956 30069 12965
rect 30124 12956 30164 13000
rect 30027 12916 30028 12956
rect 30068 12916 30164 12956
rect 30219 12956 30261 12965
rect 30700 12956 30740 13999
rect 30795 13628 30837 13637
rect 30795 13588 30796 13628
rect 30836 13588 30837 13628
rect 30795 13579 30837 13588
rect 30796 13301 30836 13579
rect 30795 13292 30837 13301
rect 30795 13252 30796 13292
rect 30836 13252 30837 13292
rect 30795 13243 30837 13252
rect 30796 13222 30836 13243
rect 30796 13173 30836 13182
rect 30892 13208 30932 14671
rect 30892 13124 30932 13168
rect 30796 13084 30932 13124
rect 30796 12965 30836 13084
rect 30988 13040 31028 15856
rect 31467 15847 31509 15856
rect 31371 15728 31413 15737
rect 31371 15688 31372 15728
rect 31412 15688 31413 15728
rect 31371 15679 31413 15688
rect 31084 14897 31124 14982
rect 31275 14972 31317 14981
rect 31275 14932 31276 14972
rect 31316 14932 31317 14972
rect 31372 14972 31412 15679
rect 31468 15560 31508 15847
rect 31468 15511 31508 15520
rect 31564 15560 31604 16015
rect 31660 15737 31700 16864
rect 31756 16820 31796 16829
rect 31948 16820 31988 16829
rect 31756 16241 31796 16780
rect 31852 16780 31948 16820
rect 31755 16232 31797 16241
rect 31755 16192 31756 16232
rect 31796 16192 31797 16232
rect 31755 16183 31797 16192
rect 31659 15728 31701 15737
rect 31659 15688 31660 15728
rect 31700 15688 31701 15728
rect 31659 15679 31701 15688
rect 31564 15511 31604 15520
rect 31660 15560 31700 15569
rect 31468 14972 31508 14981
rect 31372 14932 31468 14972
rect 31275 14923 31317 14932
rect 31468 14923 31508 14932
rect 31083 14888 31125 14897
rect 31083 14848 31084 14888
rect 31124 14848 31125 14888
rect 31083 14839 31125 14848
rect 31084 14720 31124 14729
rect 31276 14720 31316 14923
rect 31660 14888 31700 15520
rect 31756 15560 31796 15569
rect 31756 14981 31796 15520
rect 31755 14972 31797 14981
rect 31755 14932 31756 14972
rect 31796 14932 31797 14972
rect 31755 14923 31797 14932
rect 31564 14848 31700 14888
rect 31468 14720 31508 14729
rect 31124 14680 31220 14720
rect 31084 14671 31124 14680
rect 31083 13796 31125 13805
rect 31083 13756 31084 13796
rect 31124 13756 31125 13796
rect 31083 13747 31125 13756
rect 30892 13000 31028 13040
rect 30219 12916 30220 12956
rect 30260 12916 30261 12956
rect 30027 12907 30069 12916
rect 30219 12907 30261 12916
rect 30604 12916 30740 12956
rect 30795 12956 30837 12965
rect 30795 12916 30796 12956
rect 30836 12916 30837 12956
rect 30220 11696 30260 12907
rect 30412 12536 30452 12545
rect 30412 11705 30452 12496
rect 30508 12452 30548 12461
rect 30508 12125 30548 12412
rect 30604 12368 30644 12916
rect 30795 12907 30837 12916
rect 30699 12620 30741 12629
rect 30699 12580 30700 12620
rect 30740 12580 30741 12620
rect 30699 12571 30741 12580
rect 30700 12452 30740 12571
rect 30795 12536 30837 12545
rect 30795 12496 30796 12536
rect 30836 12496 30837 12536
rect 30795 12487 30837 12496
rect 30700 12403 30740 12412
rect 30604 12319 30644 12328
rect 30507 12116 30549 12125
rect 30507 12076 30508 12116
rect 30548 12076 30549 12116
rect 30507 12067 30549 12076
rect 30699 12116 30741 12125
rect 30699 12076 30700 12116
rect 30740 12076 30741 12116
rect 30699 12067 30741 12076
rect 30411 11696 30453 11705
rect 30220 11656 30356 11696
rect 29932 11320 30260 11360
rect 29548 11024 29588 11320
rect 29356 10387 29396 10396
rect 29452 10984 29548 11024
rect 29259 10352 29301 10361
rect 29259 10312 29260 10352
rect 29300 10312 29301 10352
rect 29259 10303 29301 10312
rect 29452 10277 29492 10984
rect 29548 10975 29588 10984
rect 30123 11024 30165 11033
rect 30123 10984 30124 11024
rect 30164 10984 30165 11024
rect 30123 10975 30165 10984
rect 30124 10856 30164 10975
rect 30124 10807 30164 10816
rect 29451 10268 29493 10277
rect 29451 10228 29452 10268
rect 29492 10228 29493 10268
rect 29451 10219 29493 10228
rect 29452 10184 29492 10219
rect 29643 10184 29685 10193
rect 29452 10133 29492 10144
rect 29548 10144 29644 10184
rect 29684 10144 29685 10184
rect 29356 10016 29396 10025
rect 29259 9932 29301 9941
rect 29259 9892 29260 9932
rect 29300 9892 29301 9932
rect 29259 9883 29301 9892
rect 29067 9428 29109 9437
rect 29067 9388 29068 9428
rect 29108 9388 29109 9428
rect 29067 9379 29109 9388
rect 28972 8672 29012 8681
rect 28876 8597 28916 8628
rect 28875 8588 28917 8597
rect 28875 8548 28876 8588
rect 28916 8548 28917 8588
rect 28875 8539 28917 8548
rect 28876 8504 28916 8539
rect 28972 8513 29012 8632
rect 28876 8177 28916 8464
rect 28971 8504 29013 8513
rect 28971 8464 28972 8504
rect 29012 8464 29013 8504
rect 28971 8455 29013 8464
rect 29068 8336 29108 9379
rect 29260 9344 29300 9883
rect 29356 9353 29396 9976
rect 29548 9596 29588 10144
rect 29643 10135 29685 10144
rect 29836 10184 29876 10193
rect 29644 10050 29684 10135
rect 29739 10100 29781 10109
rect 29739 10060 29740 10100
rect 29780 10060 29781 10100
rect 29739 10051 29781 10060
rect 29740 9966 29780 10051
rect 29836 9689 29876 10144
rect 30220 10184 30260 11320
rect 30220 10135 30260 10144
rect 30316 10016 30356 11656
rect 30411 11656 30412 11696
rect 30452 11656 30453 11696
rect 30411 11647 30453 11656
rect 30508 11360 30548 12067
rect 30412 11320 30548 11360
rect 30412 10184 30452 11320
rect 30412 10135 30452 10144
rect 30700 10184 30740 12067
rect 30796 12041 30836 12487
rect 30795 12032 30837 12041
rect 30795 11992 30796 12032
rect 30836 11992 30837 12032
rect 30795 11983 30837 11992
rect 30796 11453 30836 11983
rect 30795 11444 30837 11453
rect 30795 11404 30796 11444
rect 30836 11404 30837 11444
rect 30795 11395 30837 11404
rect 30796 11024 30836 11033
rect 30892 11024 30932 13000
rect 31084 12797 31124 13747
rect 31083 12788 31125 12797
rect 31083 12748 31084 12788
rect 31124 12748 31125 12788
rect 31083 12739 31125 12748
rect 30988 12536 31028 12545
rect 30988 11789 31028 12496
rect 31084 12452 31124 12739
rect 31084 12403 31124 12412
rect 31180 12368 31220 14680
rect 31316 14680 31468 14720
rect 31276 14671 31316 14680
rect 31468 14561 31508 14680
rect 31467 14552 31509 14561
rect 31467 14512 31468 14552
rect 31508 14512 31509 14552
rect 31467 14503 31509 14512
rect 31564 13712 31604 14848
rect 31756 14720 31796 14729
rect 31660 14678 31700 14687
rect 31660 13796 31700 14638
rect 31756 14393 31796 14680
rect 31755 14384 31797 14393
rect 31755 14344 31756 14384
rect 31796 14344 31797 14384
rect 31755 14335 31797 14344
rect 31756 14057 31796 14142
rect 31755 14048 31797 14057
rect 31755 14008 31756 14048
rect 31796 14008 31797 14048
rect 31755 13999 31797 14008
rect 31852 13964 31892 16780
rect 31948 16771 31988 16780
rect 32044 16157 32084 17704
rect 32140 16829 32180 17788
rect 32428 17669 32468 17872
rect 32524 17753 32564 18544
rect 32812 17837 32852 18955
rect 32907 18752 32949 18761
rect 32907 18712 32908 18752
rect 32948 18712 32949 18752
rect 32907 18703 32949 18712
rect 32908 18618 32948 18703
rect 33772 18593 33812 19216
rect 33004 18584 33044 18593
rect 32811 17828 32853 17837
rect 32811 17788 32812 17828
rect 32852 17788 32853 17828
rect 32811 17779 32853 17788
rect 32523 17744 32565 17753
rect 32523 17704 32524 17744
rect 32564 17704 32565 17744
rect 32523 17695 32565 17704
rect 32427 17660 32469 17669
rect 32427 17620 32428 17660
rect 32468 17620 32469 17660
rect 32427 17611 32469 17620
rect 32235 16988 32277 16997
rect 32235 16948 32236 16988
rect 32276 16948 32277 16988
rect 32235 16939 32277 16948
rect 32139 16820 32181 16829
rect 32139 16780 32140 16820
rect 32180 16780 32181 16820
rect 32139 16771 32181 16780
rect 32140 16325 32180 16771
rect 32139 16316 32181 16325
rect 32139 16276 32140 16316
rect 32180 16276 32181 16316
rect 32139 16267 32181 16276
rect 32140 16232 32180 16267
rect 32140 16181 32180 16192
rect 32043 16148 32085 16157
rect 32043 16108 32044 16148
rect 32084 16108 32085 16148
rect 32043 16099 32085 16108
rect 32139 16064 32181 16073
rect 32139 16024 32140 16064
rect 32180 16024 32181 16064
rect 32139 16015 32181 16024
rect 32140 15065 32180 16015
rect 32236 15560 32276 16939
rect 32428 16661 32468 17611
rect 32524 17081 32564 17695
rect 32523 17072 32565 17081
rect 32523 17032 32524 17072
rect 32564 17032 32565 17072
rect 32523 17023 32565 17032
rect 32620 17072 32660 17081
rect 32620 16829 32660 17032
rect 32619 16820 32661 16829
rect 32619 16780 32620 16820
rect 32660 16780 32661 16820
rect 32619 16771 32661 16780
rect 32427 16652 32469 16661
rect 32427 16612 32428 16652
rect 32468 16612 32469 16652
rect 32427 16603 32469 16612
rect 32331 16484 32373 16493
rect 32331 16444 32332 16484
rect 32372 16444 32373 16484
rect 32331 16435 32373 16444
rect 32332 16232 32372 16435
rect 32332 16183 32372 16192
rect 32428 16232 32468 16603
rect 33004 16409 33044 18544
rect 33099 18584 33141 18593
rect 33099 18544 33100 18584
rect 33140 18544 33141 18584
rect 33099 18535 33141 18544
rect 33196 18584 33236 18593
rect 33100 18450 33140 18535
rect 33196 17912 33236 18544
rect 33676 18584 33716 18593
rect 33676 18341 33716 18544
rect 33771 18584 33813 18593
rect 33771 18544 33772 18584
rect 33812 18544 33813 18584
rect 33771 18535 33813 18544
rect 33675 18332 33717 18341
rect 33675 18292 33676 18332
rect 33716 18292 33717 18332
rect 33675 18283 33717 18292
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 33196 17872 33524 17912
rect 33099 17828 33141 17837
rect 33099 17788 33100 17828
rect 33140 17788 33141 17828
rect 33099 17779 33141 17788
rect 33100 17744 33140 17779
rect 32619 16400 32661 16409
rect 32619 16360 32620 16400
rect 32660 16360 32661 16400
rect 32619 16351 32661 16360
rect 33003 16400 33045 16409
rect 33003 16360 33004 16400
rect 33044 16360 33045 16400
rect 33003 16351 33045 16360
rect 32620 16266 32660 16351
rect 32428 16157 32468 16192
rect 32427 16148 32469 16157
rect 32427 16108 32428 16148
rect 32468 16108 32469 16148
rect 32427 16099 32469 16108
rect 32524 16148 32564 16157
rect 32428 16068 32468 16099
rect 32524 15728 32564 16108
rect 32619 16064 32661 16073
rect 32619 16024 32620 16064
rect 32660 16024 32661 16064
rect 32619 16015 32661 16024
rect 32620 15930 32660 16015
rect 32811 15980 32853 15989
rect 32811 15940 32812 15980
rect 32852 15940 32853 15980
rect 32811 15931 32853 15940
rect 32428 15688 32564 15728
rect 32332 15560 32372 15569
rect 32236 15520 32332 15560
rect 32332 15511 32372 15520
rect 32139 15056 32181 15065
rect 32139 15016 32140 15056
rect 32180 15016 32181 15056
rect 32139 15007 32181 15016
rect 32428 14972 32468 15688
rect 32523 15560 32565 15569
rect 32523 15520 32524 15560
rect 32564 15520 32565 15560
rect 32523 15511 32565 15520
rect 32620 15560 32660 15569
rect 32660 15520 32756 15560
rect 32620 15511 32660 15520
rect 32524 15426 32564 15511
rect 32619 15392 32661 15401
rect 32619 15352 32620 15392
rect 32660 15352 32661 15392
rect 32619 15343 32661 15352
rect 32620 15258 32660 15343
rect 32428 14923 32468 14932
rect 32716 14888 32756 15520
rect 32812 15233 32852 15931
rect 33100 15728 33140 17704
rect 33196 17744 33236 17755
rect 33196 17669 33236 17704
rect 33291 17744 33333 17753
rect 33291 17704 33292 17744
rect 33332 17704 33333 17744
rect 33291 17695 33333 17704
rect 33195 17660 33237 17669
rect 33195 17620 33196 17660
rect 33236 17620 33237 17660
rect 33195 17611 33237 17620
rect 33292 17610 33332 17695
rect 33387 17660 33429 17669
rect 33387 17620 33388 17660
rect 33428 17620 33429 17660
rect 33387 17611 33429 17620
rect 33484 17660 33524 17872
rect 33580 17660 33620 17669
rect 33484 17620 33580 17660
rect 33388 17526 33428 17611
rect 33484 17408 33524 17620
rect 33580 17611 33620 17620
rect 33004 15688 33140 15728
rect 33196 17368 33524 17408
rect 32811 15224 32853 15233
rect 32811 15184 32812 15224
rect 32852 15184 32853 15224
rect 32811 15175 32853 15184
rect 32620 14848 32756 14888
rect 32811 14888 32853 14897
rect 32811 14848 32812 14888
rect 32852 14848 32853 14888
rect 31948 14720 31988 14729
rect 31948 14561 31988 14680
rect 32044 14720 32084 14729
rect 31947 14552 31989 14561
rect 31947 14512 31948 14552
rect 31988 14512 31989 14552
rect 31947 14503 31989 14512
rect 31947 14300 31989 14309
rect 31947 14260 31948 14300
rect 31988 14260 31989 14300
rect 31947 14251 31989 14260
rect 31948 14069 31988 14251
rect 31948 14020 31988 14029
rect 32044 13973 32084 14680
rect 32139 14720 32181 14729
rect 32139 14680 32140 14720
rect 32180 14680 32181 14720
rect 32139 14671 32181 14680
rect 32236 14720 32276 14729
rect 32620 14720 32660 14848
rect 32811 14839 32853 14848
rect 32276 14680 32660 14720
rect 32716 14720 32756 14729
rect 32236 14671 32276 14680
rect 32140 14586 32180 14671
rect 32716 14561 32756 14680
rect 32812 14720 32852 14839
rect 32812 14671 32852 14680
rect 32908 14561 32948 14643
rect 32715 14552 32757 14561
rect 32715 14512 32716 14552
rect 32756 14512 32757 14552
rect 32715 14503 32757 14512
rect 32907 14552 32949 14561
rect 32907 14508 32908 14552
rect 32948 14508 32949 14552
rect 32907 14503 32949 14508
rect 32908 14499 32948 14503
rect 32139 14468 32181 14477
rect 32139 14428 32140 14468
rect 32180 14428 32181 14468
rect 32139 14419 32181 14428
rect 32140 14048 32180 14419
rect 33004 14393 33044 15688
rect 33100 15560 33140 15569
rect 33100 14897 33140 15520
rect 33196 15560 33236 17368
rect 33292 17072 33332 17081
rect 33292 16913 33332 17032
rect 33676 17072 33716 17081
rect 33868 17072 33908 19888
rect 35692 19769 35732 22240
rect 36171 22280 36213 22289
rect 36171 22240 36172 22280
rect 36212 22240 36213 22280
rect 36171 22231 36213 22240
rect 36843 22280 36885 22289
rect 36843 22240 36844 22280
rect 36884 22240 36885 22280
rect 36843 22231 36885 22240
rect 36459 21524 36501 21533
rect 36459 21484 36460 21524
rect 36500 21484 36501 21524
rect 36459 21475 36501 21484
rect 36460 21390 36500 21475
rect 36747 21440 36789 21449
rect 36747 21400 36748 21440
rect 36788 21400 36789 21440
rect 36747 21391 36789 21400
rect 36748 21306 36788 21391
rect 35980 20768 36020 20777
rect 35980 20180 36020 20728
rect 36844 20768 36884 22231
rect 37324 22196 37364 22205
rect 37324 21785 37364 22156
rect 37323 21776 37365 21785
rect 37323 21736 37324 21776
rect 37364 21736 37365 21776
rect 37323 21727 37365 21736
rect 36844 20180 36884 20728
rect 37420 21608 37460 21617
rect 35980 20140 36116 20180
rect 36844 20140 36980 20180
rect 36076 19928 36116 20140
rect 36652 20096 36692 20105
rect 36555 20012 36597 20021
rect 36555 19972 36556 20012
rect 36596 19972 36597 20012
rect 36555 19963 36597 19972
rect 36076 19879 36116 19888
rect 36556 19878 36596 19963
rect 36652 19937 36692 20056
rect 36651 19928 36693 19937
rect 36651 19888 36652 19928
rect 36692 19888 36693 19928
rect 36651 19879 36693 19888
rect 36844 19844 36884 19853
rect 36748 19804 36844 19844
rect 35307 19760 35349 19769
rect 35307 19720 35308 19760
rect 35348 19720 35349 19760
rect 35307 19711 35349 19720
rect 35691 19760 35733 19769
rect 35691 19720 35692 19760
rect 35732 19720 35733 19760
rect 35691 19711 35733 19720
rect 35212 19424 35252 19433
rect 35020 19384 35212 19424
rect 34924 19256 34964 19267
rect 34924 19181 34964 19216
rect 34251 19172 34293 19181
rect 34251 19132 34252 19172
rect 34292 19132 34293 19172
rect 34251 19123 34293 19132
rect 34923 19172 34965 19181
rect 34923 19132 34924 19172
rect 34964 19132 34965 19172
rect 34923 19123 34965 19132
rect 34155 18332 34197 18341
rect 34155 18292 34156 18332
rect 34196 18292 34197 18332
rect 34155 18283 34197 18292
rect 34059 17660 34101 17669
rect 34059 17620 34060 17660
rect 34100 17620 34101 17660
rect 34059 17611 34101 17620
rect 33716 17032 33908 17072
rect 33676 17023 33716 17032
rect 33291 16904 33333 16913
rect 33291 16864 33292 16904
rect 33332 16864 33333 16904
rect 33291 16855 33333 16864
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 34060 16232 34100 17611
rect 34156 16316 34196 18283
rect 34252 17744 34292 19123
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 34348 18584 34388 18593
rect 34540 18584 34580 18593
rect 34388 18544 34540 18584
rect 34348 18535 34388 18544
rect 34540 18535 34580 18544
rect 34924 18584 34964 18593
rect 35020 18584 35060 19384
rect 35212 19375 35252 19384
rect 35115 19172 35157 19181
rect 35115 19132 35116 19172
rect 35156 19132 35157 19172
rect 35115 19123 35157 19132
rect 34964 18544 35060 18584
rect 34924 18535 34964 18544
rect 34252 17695 34292 17704
rect 34443 17744 34485 17753
rect 34443 17704 34444 17744
rect 34484 17704 34485 17744
rect 34443 17695 34485 17704
rect 34156 16267 34196 16276
rect 34060 16183 34100 16192
rect 34251 16232 34293 16241
rect 34251 16192 34252 16232
rect 34292 16192 34293 16232
rect 34251 16183 34293 16192
rect 34252 16098 34292 16183
rect 33579 16064 33621 16073
rect 33579 16024 33580 16064
rect 33620 16024 33621 16064
rect 33579 16015 33621 16024
rect 33580 15728 33620 16015
rect 33580 15679 33620 15688
rect 33388 15569 33428 15654
rect 33675 15644 33717 15653
rect 33675 15604 33676 15644
rect 33716 15604 33717 15644
rect 33675 15595 33717 15604
rect 34155 15644 34197 15653
rect 34155 15604 34156 15644
rect 34196 15604 34197 15644
rect 34155 15595 34197 15604
rect 33196 15511 33236 15520
rect 33387 15560 33429 15569
rect 33387 15520 33388 15560
rect 33428 15520 33429 15560
rect 33387 15511 33429 15520
rect 33676 15560 33716 15595
rect 33676 15509 33716 15520
rect 33963 15560 34005 15569
rect 33963 15520 33964 15560
rect 34004 15520 34005 15560
rect 33963 15511 34005 15520
rect 34060 15560 34100 15571
rect 33388 15317 33428 15402
rect 33387 15308 33429 15317
rect 33387 15268 33388 15308
rect 33428 15268 33429 15308
rect 33387 15259 33429 15268
rect 33868 15308 33908 15317
rect 33868 15149 33908 15268
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 33867 15140 33909 15149
rect 33867 15100 33868 15140
rect 33908 15100 33909 15140
rect 33867 15091 33909 15100
rect 33867 14972 33909 14981
rect 33867 14932 33868 14972
rect 33908 14932 33909 14972
rect 33867 14923 33909 14932
rect 33099 14888 33141 14897
rect 33099 14848 33100 14888
rect 33140 14848 33141 14888
rect 33099 14839 33141 14848
rect 33292 14888 33332 14897
rect 33195 14804 33237 14813
rect 33195 14764 33196 14804
rect 33236 14764 33237 14804
rect 33195 14755 33237 14764
rect 33100 14720 33140 14729
rect 32907 14384 32949 14393
rect 32907 14344 32908 14384
rect 32948 14344 32949 14384
rect 33004 14384 33050 14393
rect 33004 14344 33009 14384
rect 33049 14344 33050 14384
rect 32907 14335 32949 14344
rect 33008 14335 33050 14344
rect 32235 14132 32277 14141
rect 32235 14092 32236 14132
rect 32276 14092 32277 14132
rect 32235 14083 32277 14092
rect 32140 13999 32180 14008
rect 32043 13964 32085 13973
rect 31852 13924 31991 13964
rect 31951 13880 31991 13924
rect 32043 13924 32044 13964
rect 32084 13924 32085 13964
rect 32043 13915 32085 13924
rect 32236 13964 32276 14083
rect 32523 14048 32565 14057
rect 32523 14008 32524 14048
rect 32564 14008 32565 14048
rect 32523 13999 32565 14008
rect 32715 14048 32757 14057
rect 32715 14008 32716 14048
rect 32756 14008 32757 14048
rect 32715 13999 32757 14008
rect 31948 13840 31991 13880
rect 31852 13796 31892 13805
rect 31660 13756 31852 13796
rect 31852 13747 31892 13756
rect 31564 13672 31796 13712
rect 31756 13628 31796 13672
rect 31756 13588 31892 13628
rect 31659 13544 31701 13553
rect 31659 13504 31660 13544
rect 31700 13504 31701 13544
rect 31659 13495 31701 13504
rect 31660 13460 31700 13495
rect 31660 13409 31700 13420
rect 31564 13208 31604 13217
rect 31564 12713 31604 13168
rect 31755 13208 31797 13217
rect 31755 13168 31756 13208
rect 31796 13168 31797 13208
rect 31755 13159 31797 13168
rect 31756 13074 31796 13159
rect 31563 12704 31605 12713
rect 31563 12664 31564 12704
rect 31604 12664 31605 12704
rect 31563 12655 31605 12664
rect 31852 12704 31892 13588
rect 31852 12655 31892 12664
rect 31660 12545 31700 12630
rect 31371 12536 31413 12545
rect 31371 12496 31372 12536
rect 31412 12496 31413 12536
rect 31371 12487 31413 12496
rect 31564 12536 31604 12545
rect 31275 12452 31317 12461
rect 31275 12412 31276 12452
rect 31316 12412 31317 12452
rect 31275 12403 31317 12412
rect 31180 12319 31220 12328
rect 31276 12318 31316 12403
rect 31372 12402 31412 12487
rect 31564 12125 31604 12496
rect 31659 12536 31701 12545
rect 31659 12496 31660 12536
rect 31700 12496 31701 12536
rect 31659 12487 31701 12496
rect 31852 12536 31892 12545
rect 31852 12209 31892 12496
rect 31948 12536 31988 13840
rect 32236 13805 32276 13924
rect 32428 13964 32468 13973
rect 32331 13880 32373 13889
rect 32331 13840 32332 13880
rect 32372 13840 32373 13880
rect 32331 13831 32373 13840
rect 32235 13796 32277 13805
rect 32235 13756 32236 13796
rect 32276 13756 32277 13796
rect 32235 13747 32277 13756
rect 32332 13746 32372 13831
rect 32236 13376 32276 13385
rect 32428 13376 32468 13924
rect 32524 13721 32564 13999
rect 32716 13914 32756 13999
rect 32812 13962 32852 13971
rect 32523 13712 32565 13721
rect 32523 13672 32524 13712
rect 32564 13672 32565 13712
rect 32523 13663 32565 13672
rect 32428 13336 32660 13376
rect 32044 13301 32084 13332
rect 32043 13292 32085 13301
rect 32043 13252 32044 13292
rect 32084 13252 32085 13292
rect 32043 13243 32085 13252
rect 32140 13292 32180 13301
rect 32044 13208 32084 13243
rect 32044 12536 32084 13168
rect 32140 12797 32180 13252
rect 32236 13217 32276 13336
rect 32332 13292 32372 13301
rect 32235 13208 32277 13217
rect 32235 13168 32236 13208
rect 32276 13168 32277 13208
rect 32235 13159 32277 13168
rect 32332 13133 32372 13252
rect 32428 13208 32468 13217
rect 32331 13124 32373 13133
rect 32331 13084 32332 13124
rect 32372 13084 32373 13124
rect 32331 13075 32373 13084
rect 32428 12965 32468 13168
rect 32427 12956 32469 12965
rect 32427 12916 32428 12956
rect 32468 12916 32469 12956
rect 32427 12907 32469 12916
rect 32139 12788 32181 12797
rect 32139 12748 32140 12788
rect 32180 12748 32181 12788
rect 32139 12739 32181 12748
rect 32427 12704 32469 12713
rect 32427 12664 32428 12704
rect 32468 12664 32469 12704
rect 32427 12655 32469 12664
rect 32428 12620 32468 12655
rect 32428 12569 32468 12580
rect 32332 12536 32372 12545
rect 32044 12521 32145 12536
rect 32044 12496 32105 12521
rect 31948 12487 31988 12496
rect 32105 12452 32145 12481
rect 32105 12412 32276 12452
rect 31851 12200 31893 12209
rect 31851 12160 31852 12200
rect 31892 12160 31893 12200
rect 31851 12151 31893 12160
rect 31563 12116 31605 12125
rect 31563 12076 31564 12116
rect 31604 12076 31605 12116
rect 31563 12067 31605 12076
rect 32043 12116 32085 12125
rect 32043 12076 32044 12116
rect 32084 12076 32085 12116
rect 32043 12067 32085 12076
rect 31563 11948 31605 11957
rect 31563 11908 31564 11948
rect 31604 11908 31605 11948
rect 31563 11899 31605 11908
rect 30987 11780 31029 11789
rect 30987 11740 30988 11780
rect 31028 11740 31029 11780
rect 30987 11731 31029 11740
rect 31371 11780 31413 11789
rect 31371 11740 31372 11780
rect 31412 11740 31413 11780
rect 31371 11731 31413 11740
rect 31083 11696 31125 11705
rect 31083 11656 31084 11696
rect 31124 11656 31125 11696
rect 31083 11647 31125 11656
rect 31084 11453 31124 11647
rect 31083 11444 31125 11453
rect 31083 11404 31084 11444
rect 31124 11404 31125 11444
rect 31083 11395 31125 11404
rect 31372 11360 31412 11731
rect 31468 11696 31508 11707
rect 31564 11696 31604 11899
rect 31660 11873 31700 11958
rect 31659 11864 31701 11873
rect 31659 11824 31660 11864
rect 31700 11824 31701 11864
rect 31659 11815 31701 11824
rect 31851 11864 31893 11873
rect 31851 11824 31852 11864
rect 31892 11824 31893 11864
rect 31851 11815 31893 11824
rect 32044 11864 32084 12067
rect 32044 11815 32084 11824
rect 31660 11696 31700 11705
rect 31564 11656 31660 11696
rect 31468 11621 31508 11656
rect 31660 11647 31700 11656
rect 31467 11612 31509 11621
rect 31467 11572 31468 11612
rect 31508 11572 31509 11612
rect 31467 11563 31509 11572
rect 31563 11444 31605 11453
rect 31563 11404 31564 11444
rect 31604 11404 31605 11444
rect 31563 11395 31605 11404
rect 31372 11320 31508 11360
rect 30836 10984 30932 11024
rect 31468 11024 31508 11320
rect 31564 11192 31604 11395
rect 31755 11192 31797 11201
rect 31564 11152 31700 11192
rect 30796 10975 30836 10984
rect 31468 10975 31508 10984
rect 31563 11024 31605 11033
rect 31563 10984 31564 11024
rect 31604 10984 31605 11024
rect 31563 10975 31605 10984
rect 31564 10890 31604 10975
rect 31660 10520 31700 11152
rect 31755 11152 31756 11192
rect 31796 11152 31797 11192
rect 31755 11143 31797 11152
rect 31756 11058 31796 11143
rect 31468 10480 31700 10520
rect 31371 10352 31413 10361
rect 31371 10312 31372 10352
rect 31412 10312 31413 10352
rect 31371 10303 31413 10312
rect 31372 10184 31412 10303
rect 31468 10268 31508 10480
rect 31468 10219 31508 10228
rect 31564 10352 31604 10361
rect 31564 10193 31604 10312
rect 31755 10352 31797 10361
rect 31755 10312 31756 10352
rect 31796 10312 31797 10352
rect 31755 10303 31797 10312
rect 31659 10268 31701 10277
rect 31659 10228 31660 10268
rect 31700 10228 31701 10268
rect 31659 10219 31701 10228
rect 30740 10144 31220 10184
rect 30700 10135 30740 10144
rect 30508 10100 30548 10109
rect 30508 10016 30548 10060
rect 30316 9976 30548 10016
rect 29835 9680 29877 9689
rect 29835 9640 29836 9680
rect 29876 9640 29877 9680
rect 30508 9680 30548 9976
rect 30796 9680 30836 9689
rect 30508 9640 30644 9680
rect 29835 9631 29877 9640
rect 29548 9547 29588 9556
rect 30219 9596 30261 9605
rect 30219 9556 30220 9596
rect 30260 9556 30261 9596
rect 30219 9547 30261 9556
rect 29644 9512 29684 9523
rect 29644 9437 29684 9472
rect 29932 9512 29972 9521
rect 29643 9428 29685 9437
rect 29643 9388 29644 9428
rect 29684 9388 29685 9428
rect 29643 9379 29685 9388
rect 29932 9353 29972 9472
rect 30220 9462 30260 9547
rect 30316 9512 30356 9521
rect 29260 9295 29300 9304
rect 29355 9344 29397 9353
rect 29355 9304 29356 9344
rect 29396 9304 29397 9344
rect 29355 9295 29397 9304
rect 29931 9344 29973 9353
rect 29931 9304 29932 9344
rect 29972 9304 29973 9344
rect 29931 9295 29973 9304
rect 30316 8933 30356 9472
rect 30412 9512 30452 9521
rect 30412 9017 30452 9472
rect 30508 9512 30548 9521
rect 30411 9008 30453 9017
rect 30411 8968 30412 9008
rect 30452 8968 30453 9008
rect 30411 8959 30453 8968
rect 30315 8924 30357 8933
rect 30315 8884 30316 8924
rect 30356 8884 30357 8924
rect 30315 8875 30357 8884
rect 29260 8840 29300 8849
rect 30508 8840 30548 9472
rect 30604 9344 30644 9640
rect 30836 9640 31028 9680
rect 30796 9631 30836 9640
rect 30699 9596 30741 9605
rect 30699 9556 30700 9596
rect 30740 9556 30741 9596
rect 30699 9547 30741 9556
rect 30700 9512 30740 9547
rect 30700 9461 30740 9472
rect 30892 9512 30932 9523
rect 30892 9437 30932 9472
rect 30891 9428 30933 9437
rect 30891 9388 30892 9428
rect 30932 9388 30933 9428
rect 30891 9379 30933 9388
rect 30604 9304 30740 9344
rect 30700 8849 30740 9304
rect 29300 8800 29684 8840
rect 29260 8791 29300 8800
rect 29163 8756 29205 8765
rect 29163 8716 29164 8756
rect 29204 8716 29205 8756
rect 29163 8707 29205 8716
rect 29164 8672 29204 8707
rect 29164 8513 29204 8632
rect 29356 8672 29396 8681
rect 29547 8672 29589 8681
rect 29396 8632 29492 8672
rect 29356 8623 29396 8632
rect 29163 8504 29205 8513
rect 29163 8464 29164 8504
rect 29204 8464 29205 8504
rect 29163 8455 29205 8464
rect 29068 8296 29204 8336
rect 28875 8168 28917 8177
rect 28875 8128 28876 8168
rect 28916 8128 28917 8168
rect 28875 8119 28917 8128
rect 29067 7580 29109 7589
rect 29067 7540 29068 7580
rect 29108 7540 29109 7580
rect 29067 7531 29109 7540
rect 28779 7244 28821 7253
rect 28779 7204 28780 7244
rect 28820 7204 28821 7244
rect 28779 7195 28821 7204
rect 28396 6439 28436 6448
rect 28492 6616 28724 6656
rect 27532 6353 27572 6364
rect 27724 6364 27956 6404
rect 27435 6320 27477 6329
rect 27435 6280 27436 6320
rect 27476 6280 27477 6320
rect 27435 6271 27477 6280
rect 27436 6186 27476 6271
rect 27148 5900 27188 5909
rect 26283 5396 26325 5405
rect 26283 5356 26284 5396
rect 26324 5356 26325 5396
rect 26283 5347 26325 5356
rect 26476 4985 26516 5440
rect 26572 5440 26708 5480
rect 26764 5860 27148 5900
rect 25036 4976 25076 4985
rect 26092 4976 26132 4985
rect 25076 4936 25172 4976
rect 25036 4927 25076 4936
rect 25035 4724 25077 4733
rect 25035 4684 25036 4724
rect 25076 4684 25077 4724
rect 25035 4675 25077 4684
rect 25036 4590 25076 4675
rect 24939 4556 24981 4565
rect 24939 4516 24940 4556
rect 24980 4516 24981 4556
rect 24939 4507 24981 4516
rect 23595 4304 23637 4313
rect 23595 4264 23596 4304
rect 23636 4264 23637 4304
rect 23595 4255 23637 4264
rect 24075 4304 24117 4313
rect 24075 4264 24076 4304
rect 24116 4264 24117 4304
rect 24075 4255 24117 4264
rect 24843 4304 24885 4313
rect 24843 4264 24844 4304
rect 24884 4264 24885 4304
rect 24843 4255 24885 4264
rect 23307 3800 23349 3809
rect 23307 3760 23308 3800
rect 23348 3760 23349 3800
rect 23307 3751 23349 3760
rect 23499 3716 23541 3725
rect 23499 3676 23500 3716
rect 23540 3676 23541 3716
rect 23499 3667 23541 3676
rect 22964 3424 23060 3464
rect 23500 3464 23540 3667
rect 22924 3415 22964 3424
rect 23500 3415 23540 3424
rect 23596 3464 23636 4255
rect 23788 4136 23828 4145
rect 23788 3977 23828 4096
rect 23979 4136 24021 4145
rect 23979 4096 23980 4136
rect 24020 4096 24021 4136
rect 23979 4087 24021 4096
rect 23787 3968 23829 3977
rect 23787 3928 23788 3968
rect 23828 3928 23829 3968
rect 23787 3919 23829 3928
rect 23787 3632 23829 3641
rect 23787 3592 23788 3632
rect 23828 3592 23829 3632
rect 23787 3583 23829 3592
rect 23980 3632 24020 4087
rect 24076 3964 24116 4255
rect 24076 3915 24116 3924
rect 24172 4136 24212 4145
rect 24172 3725 24212 4096
rect 24268 4136 24308 4145
rect 24171 3716 24213 3725
rect 24171 3676 24172 3716
rect 24212 3676 24213 3716
rect 24171 3667 24213 3676
rect 24268 3641 24308 4096
rect 25132 4136 25172 4936
rect 25804 4936 26092 4976
rect 25419 4640 25461 4649
rect 25419 4600 25420 4640
rect 25460 4600 25461 4640
rect 25419 4591 25461 4600
rect 25420 4397 25460 4591
rect 25419 4388 25461 4397
rect 25419 4348 25420 4388
rect 25460 4348 25461 4388
rect 25419 4339 25461 4348
rect 25323 4304 25365 4313
rect 25323 4264 25324 4304
rect 25364 4264 25365 4304
rect 25323 4255 25365 4264
rect 25132 4087 25172 4096
rect 25228 4136 25268 4145
rect 24363 4052 24405 4061
rect 24363 4012 24364 4052
rect 24404 4012 24405 4052
rect 24363 4003 24405 4012
rect 23980 3583 24020 3592
rect 24267 3632 24309 3641
rect 24267 3592 24268 3632
rect 24308 3592 24309 3632
rect 24267 3583 24309 3592
rect 23788 3498 23828 3583
rect 24075 3548 24117 3557
rect 24075 3508 24076 3548
rect 24116 3508 24117 3548
rect 24075 3499 24117 3508
rect 23596 3415 23636 3424
rect 23691 3464 23733 3473
rect 23691 3424 23692 3464
rect 23732 3424 23733 3464
rect 23691 3415 23733 3424
rect 24076 3464 24116 3499
rect 22732 3330 22772 3415
rect 23692 3330 23732 3415
rect 24076 3413 24116 3424
rect 24172 3464 24212 3473
rect 24172 3305 24212 3424
rect 24267 3464 24309 3473
rect 24267 3424 24268 3464
rect 24308 3424 24309 3464
rect 24267 3415 24309 3424
rect 24268 3330 24308 3415
rect 24364 3305 24404 4003
rect 25228 3800 25268 4096
rect 25324 4136 25364 4255
rect 25324 4087 25364 4096
rect 25420 4136 25460 4339
rect 25612 4145 25652 4230
rect 25420 4087 25460 4096
rect 25611 4136 25653 4145
rect 25611 4096 25612 4136
rect 25652 4096 25653 4136
rect 25611 4087 25653 4096
rect 25804 4136 25844 4936
rect 26092 4927 26132 4936
rect 26188 4976 26228 4985
rect 26091 4808 26133 4817
rect 26091 4768 26092 4808
rect 26132 4768 26133 4808
rect 26091 4759 26133 4768
rect 25899 4220 25941 4229
rect 25899 4180 25900 4220
rect 25940 4180 25941 4220
rect 25899 4171 25941 4180
rect 25804 4087 25844 4096
rect 25900 4136 25940 4171
rect 26092 4145 26132 4759
rect 26188 4388 26228 4936
rect 26284 4976 26324 4985
rect 26284 4817 26324 4936
rect 26380 4976 26420 4985
rect 26283 4808 26325 4817
rect 26283 4768 26284 4808
rect 26324 4768 26325 4808
rect 26283 4759 26325 4768
rect 26380 4556 26420 4936
rect 26475 4976 26517 4985
rect 26475 4936 26476 4976
rect 26516 4936 26517 4976
rect 26475 4927 26517 4936
rect 26572 4976 26612 5440
rect 26380 4516 26516 4556
rect 26380 4388 26420 4397
rect 26188 4348 26380 4388
rect 26380 4339 26420 4348
rect 26380 4229 26420 4260
rect 26379 4220 26421 4229
rect 26379 4180 26380 4220
rect 26420 4180 26421 4220
rect 26379 4171 26421 4180
rect 25900 4085 25940 4096
rect 26091 4136 26133 4145
rect 26091 4096 26092 4136
rect 26132 4096 26133 4136
rect 26091 4087 26133 4096
rect 26188 4136 26228 4147
rect 26092 4002 26132 4087
rect 26188 4061 26228 4096
rect 26380 4136 26420 4171
rect 26187 4052 26229 4061
rect 26187 4012 26188 4052
rect 26228 4012 26229 4052
rect 26187 4003 26229 4012
rect 26380 3977 26420 4096
rect 26476 4061 26516 4516
rect 26475 4052 26517 4061
rect 26475 4012 26476 4052
rect 26516 4012 26517 4052
rect 26475 4003 26517 4012
rect 25708 3968 25748 3977
rect 25612 3928 25708 3968
rect 25228 3760 25460 3800
rect 25420 3557 25460 3760
rect 25515 3632 25557 3641
rect 25515 3592 25516 3632
rect 25556 3592 25557 3632
rect 25515 3583 25557 3592
rect 25419 3548 25461 3557
rect 25419 3508 25420 3548
rect 25460 3508 25461 3548
rect 25419 3499 25461 3508
rect 24460 3464 24500 3473
rect 24460 3389 24500 3424
rect 25324 3389 25364 3474
rect 24459 3380 24501 3389
rect 24459 3340 24460 3380
rect 24500 3340 24501 3380
rect 24459 3331 24501 3340
rect 25323 3380 25365 3389
rect 25323 3340 25324 3380
rect 25364 3340 25365 3380
rect 25323 3331 25365 3340
rect 24171 3296 24213 3305
rect 24171 3256 24172 3296
rect 24212 3256 24213 3296
rect 24171 3247 24213 3256
rect 24363 3296 24405 3305
rect 24363 3256 24364 3296
rect 24404 3256 24405 3296
rect 24363 3247 24405 3256
rect 22924 3212 22964 3221
rect 22635 2792 22677 2801
rect 22635 2752 22636 2792
rect 22676 2752 22677 2792
rect 22635 2743 22677 2752
rect 22924 2540 22964 3172
rect 24172 2876 24212 2885
rect 24460 2876 24500 3331
rect 25132 3212 25172 3221
rect 25172 3172 25364 3212
rect 25132 3163 25172 3172
rect 25131 2960 25173 2969
rect 25131 2920 25132 2960
rect 25172 2920 25173 2960
rect 25131 2911 25173 2920
rect 24212 2836 24500 2876
rect 25132 2876 25172 2911
rect 24172 2827 24212 2836
rect 25132 2825 25172 2836
rect 22636 2500 22964 2540
rect 23020 2624 23060 2633
rect 22443 2120 22485 2129
rect 22443 2080 22444 2120
rect 22484 2080 22485 2120
rect 22443 2071 22485 2080
rect 22539 2036 22581 2045
rect 22539 1996 22540 2036
rect 22580 1996 22581 2036
rect 22539 1987 22581 1996
rect 21964 1903 22004 1912
rect 22443 1952 22485 1961
rect 22443 1912 22444 1952
rect 22484 1912 22485 1952
rect 22443 1903 22485 1912
rect 22444 1818 22484 1903
rect 22540 1902 22580 1987
rect 22636 1952 22676 2500
rect 23020 2465 23060 2584
rect 25324 2624 25364 3172
rect 25420 2801 25460 3499
rect 25516 3498 25556 3583
rect 25419 2792 25461 2801
rect 25419 2752 25420 2792
rect 25460 2752 25461 2792
rect 25419 2743 25461 2752
rect 25324 2575 25364 2584
rect 23019 2456 23061 2465
rect 23019 2416 23020 2456
rect 23060 2416 23061 2456
rect 23019 2407 23061 2416
rect 24075 2456 24117 2465
rect 24075 2416 24076 2456
rect 24116 2416 24117 2456
rect 24075 2407 24117 2416
rect 22923 2036 22965 2045
rect 22923 1996 22924 2036
rect 22964 1996 22965 2036
rect 22923 1987 22965 1996
rect 22636 1903 22676 1912
rect 22924 1902 22964 1987
rect 23308 1952 23348 1961
rect 24076 1952 24116 2407
rect 24172 1952 24212 1961
rect 23348 1912 23444 1952
rect 24076 1912 24172 1952
rect 23308 1903 23348 1912
rect 23404 1280 23444 1912
rect 24172 1903 24212 1912
rect 25612 1952 25652 3928
rect 25708 3919 25748 3928
rect 26379 3968 26421 3977
rect 26379 3928 26380 3968
rect 26420 3928 26421 3968
rect 26379 3919 26421 3928
rect 26572 3557 26612 4936
rect 26668 4976 26708 4987
rect 26668 4901 26708 4936
rect 26764 4976 26804 5860
rect 27148 5851 27188 5860
rect 26859 5648 26901 5657
rect 26859 5608 26860 5648
rect 26900 5608 26901 5648
rect 26859 5599 26901 5608
rect 26860 5514 26900 5599
rect 27052 5144 27092 5153
rect 27092 5104 27476 5144
rect 27052 5095 27092 5104
rect 26667 4892 26709 4901
rect 26667 4852 26668 4892
rect 26708 4852 26709 4892
rect 26667 4843 26709 4852
rect 26668 4304 26708 4313
rect 26668 4145 26708 4264
rect 26667 4136 26709 4145
rect 26667 4096 26668 4136
rect 26708 4096 26709 4136
rect 26667 4087 26709 4096
rect 26764 4136 26804 4936
rect 26859 4976 26901 4985
rect 26859 4936 26860 4976
rect 26900 4936 26901 4976
rect 26859 4927 26901 4936
rect 27243 4976 27285 4985
rect 27243 4936 27244 4976
rect 27284 4936 27285 4976
rect 27243 4927 27285 4936
rect 27340 4976 27380 4985
rect 27436 4976 27476 5104
rect 27532 4976 27572 4985
rect 27436 4936 27532 4976
rect 26860 4842 26900 4927
rect 27244 4842 27284 4927
rect 27340 4817 27380 4936
rect 27532 4927 27572 4936
rect 27147 4808 27189 4817
rect 27147 4768 27148 4808
rect 27188 4768 27189 4808
rect 27147 4759 27189 4768
rect 27339 4808 27381 4817
rect 27628 4808 27668 4817
rect 27339 4768 27340 4808
rect 27380 4768 27381 4808
rect 27339 4759 27381 4768
rect 27436 4768 27628 4808
rect 26764 3809 26804 4096
rect 26860 4136 26900 4145
rect 26763 3800 26805 3809
rect 26763 3760 26764 3800
rect 26804 3760 26805 3800
rect 26763 3751 26805 3760
rect 26571 3548 26613 3557
rect 26571 3508 26572 3548
rect 26612 3508 26613 3548
rect 26571 3499 26613 3508
rect 26380 3464 26420 3473
rect 25708 3212 25748 3221
rect 25748 3172 25940 3212
rect 25708 3163 25748 3172
rect 25900 2624 25940 3172
rect 25900 2575 25940 2584
rect 26380 2540 26420 3424
rect 26763 3464 26805 3473
rect 26860 3464 26900 4096
rect 26763 3424 26764 3464
rect 26804 3424 26900 3464
rect 26763 3415 26805 3424
rect 26764 3330 26804 3415
rect 26571 3212 26613 3221
rect 26571 3172 26572 3212
rect 26612 3172 26613 3212
rect 26571 3163 26613 3172
rect 26572 2876 26612 3163
rect 27148 3137 27188 4759
rect 27340 4136 27380 4145
rect 27243 3548 27285 3557
rect 27243 3508 27244 3548
rect 27284 3508 27285 3548
rect 27243 3499 27285 3508
rect 27147 3128 27189 3137
rect 27147 3088 27148 3128
rect 27188 3088 27189 3128
rect 27147 3079 27189 3088
rect 27244 3053 27284 3499
rect 27243 3044 27285 3053
rect 27243 3004 27244 3044
rect 27284 3004 27285 3044
rect 27243 2995 27285 3004
rect 26572 2827 26612 2836
rect 27052 2876 27092 2885
rect 27340 2876 27380 4096
rect 27436 3893 27476 4768
rect 27628 4759 27668 4768
rect 27627 4472 27669 4481
rect 27627 4432 27628 4472
rect 27668 4432 27669 4472
rect 27627 4423 27669 4432
rect 27628 4304 27668 4423
rect 27628 4255 27668 4264
rect 27532 4136 27572 4145
rect 27532 3977 27572 4096
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 27628 4002 27668 4087
rect 27531 3968 27573 3977
rect 27531 3928 27532 3968
rect 27572 3928 27573 3968
rect 27531 3919 27573 3928
rect 27435 3884 27477 3893
rect 27435 3844 27436 3884
rect 27476 3844 27477 3884
rect 27435 3835 27477 3844
rect 27627 3884 27669 3893
rect 27627 3844 27628 3884
rect 27668 3844 27669 3884
rect 27627 3835 27669 3844
rect 27531 3800 27573 3809
rect 27531 3760 27532 3800
rect 27572 3760 27573 3800
rect 27531 3751 27573 3760
rect 27435 3548 27477 3557
rect 27435 3508 27436 3548
rect 27476 3508 27477 3548
rect 27435 3499 27477 3508
rect 27436 3464 27476 3499
rect 27436 3413 27476 3424
rect 27435 3212 27477 3221
rect 27435 3172 27436 3212
rect 27476 3172 27477 3212
rect 27435 3163 27477 3172
rect 27092 2836 27380 2876
rect 27052 2827 27092 2836
rect 26284 2500 26420 2540
rect 27148 2624 27188 2633
rect 27148 2540 27188 2584
rect 27436 2540 27476 3163
rect 27532 2624 27572 3751
rect 27628 3464 27668 3835
rect 27628 3415 27668 3424
rect 27628 3212 27668 3221
rect 27628 2885 27668 3172
rect 27627 2876 27669 2885
rect 27627 2836 27628 2876
rect 27668 2836 27669 2876
rect 27627 2827 27669 2836
rect 27532 2575 27572 2584
rect 27148 2500 27436 2540
rect 25612 1903 25652 1912
rect 25996 1952 26036 1961
rect 26036 1912 26132 1952
rect 25996 1903 26036 1912
rect 25324 1700 25364 1709
rect 25324 1289 25364 1660
rect 23404 1231 23444 1240
rect 25323 1280 25365 1289
rect 25323 1240 25324 1280
rect 25364 1240 25365 1280
rect 25323 1231 25365 1240
rect 26092 1280 26132 1912
rect 26284 1289 26324 2500
rect 27436 2491 27476 2500
rect 26859 1952 26901 1961
rect 26859 1912 26860 1952
rect 26900 1912 26901 1952
rect 26859 1903 26901 1912
rect 26860 1818 26900 1903
rect 26092 1231 26132 1240
rect 26283 1280 26325 1289
rect 26283 1240 26284 1280
rect 26324 1240 26325 1280
rect 26283 1231 26325 1240
rect 26667 1280 26709 1289
rect 26667 1240 26668 1280
rect 26708 1240 26709 1280
rect 26667 1231 26709 1240
rect 19468 1063 19508 1072
rect 19563 1112 19605 1121
rect 19563 1072 19564 1112
rect 19604 1072 19605 1112
rect 19563 1063 19605 1072
rect 20715 1112 20757 1121
rect 20715 1072 20716 1112
rect 20756 1072 20757 1112
rect 20715 1063 20757 1072
rect 26668 1112 26708 1231
rect 27724 1121 27764 6364
rect 28204 6354 28244 6439
rect 28204 6236 28244 6245
rect 28108 6196 28204 6236
rect 27820 5648 27860 5657
rect 27820 5489 27860 5608
rect 27915 5648 27957 5657
rect 27915 5608 27916 5648
rect 27956 5608 27957 5648
rect 27915 5599 27957 5608
rect 27819 5480 27861 5489
rect 27819 5440 27820 5480
rect 27860 5440 27861 5480
rect 27819 5431 27861 5440
rect 27916 4976 27956 5599
rect 28108 5153 28148 6196
rect 28204 6187 28244 6196
rect 28492 5657 28532 6616
rect 28587 6488 28629 6497
rect 28587 6448 28588 6488
rect 28628 6448 28629 6488
rect 28587 6439 28629 6448
rect 28780 6488 28820 7195
rect 29068 7160 29108 7531
rect 29068 7111 29108 7120
rect 29164 6497 29204 8296
rect 29452 8009 29492 8632
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 29644 8672 29684 8800
rect 30412 8800 30548 8840
rect 30699 8840 30741 8849
rect 30699 8800 30700 8840
rect 30740 8800 30741 8840
rect 29644 8623 29684 8632
rect 29740 8672 29780 8683
rect 29548 8538 29588 8623
rect 29740 8597 29780 8632
rect 29836 8672 29876 8681
rect 29739 8588 29781 8597
rect 29739 8548 29740 8588
rect 29780 8548 29781 8588
rect 29739 8539 29781 8548
rect 29836 8177 29876 8632
rect 30065 8672 30105 8683
rect 30065 8597 30105 8632
rect 30220 8672 30260 8681
rect 30064 8588 30106 8597
rect 30064 8548 30065 8588
rect 30105 8548 30106 8588
rect 30064 8539 30106 8548
rect 29835 8168 29877 8177
rect 29835 8128 29836 8168
rect 29876 8128 29877 8168
rect 29835 8119 29877 8128
rect 29451 8000 29493 8009
rect 29451 7960 29452 8000
rect 29492 7960 29493 8000
rect 29451 7951 29493 7960
rect 29835 8000 29877 8009
rect 29835 7960 29836 8000
rect 29876 7960 29877 8000
rect 29835 7951 29877 7960
rect 29932 8000 29972 8009
rect 29355 7412 29397 7421
rect 29355 7372 29356 7412
rect 29396 7372 29397 7412
rect 29355 7363 29397 7372
rect 29259 7244 29301 7253
rect 29259 7204 29260 7244
rect 29300 7204 29301 7244
rect 29259 7195 29301 7204
rect 29260 7160 29300 7195
rect 29260 7109 29300 7120
rect 29356 6749 29396 7363
rect 29452 7160 29492 7951
rect 29836 7866 29876 7951
rect 29932 7664 29972 7960
rect 30027 8000 30069 8009
rect 30027 7960 30028 8000
rect 30068 7960 30069 8000
rect 30027 7951 30069 7960
rect 30124 8000 30164 8009
rect 30028 7866 30068 7951
rect 30124 7673 30164 7960
rect 29644 7624 29972 7664
rect 30123 7664 30165 7673
rect 30123 7624 30124 7664
rect 30164 7624 30165 7664
rect 29644 7328 29684 7624
rect 30123 7615 30165 7624
rect 30220 7589 30260 8632
rect 30315 8672 30357 8681
rect 30315 8632 30316 8672
rect 30356 8632 30357 8672
rect 30315 8623 30357 8632
rect 30316 8538 30356 8623
rect 30412 8504 30452 8800
rect 30699 8791 30741 8800
rect 30988 8765 31028 9640
rect 31083 9260 31125 9269
rect 31083 9220 31084 9260
rect 31124 9220 31125 9260
rect 31083 9211 31125 9220
rect 30603 8756 30645 8765
rect 30603 8716 30604 8756
rect 30644 8716 30645 8756
rect 30603 8707 30645 8716
rect 30987 8756 31029 8765
rect 30987 8716 30988 8756
rect 31028 8716 31029 8756
rect 30987 8707 31029 8716
rect 30508 8672 30548 8681
rect 30508 8513 30548 8632
rect 30604 8672 30644 8707
rect 30604 8621 30644 8632
rect 30412 8455 30452 8464
rect 30507 8504 30549 8513
rect 30507 8464 30508 8504
rect 30548 8464 30549 8504
rect 30507 8455 30549 8464
rect 30987 8168 31029 8177
rect 30987 8128 30988 8168
rect 31028 8128 31029 8168
rect 30987 8119 31029 8128
rect 30603 8000 30645 8009
rect 30603 7960 30604 8000
rect 30644 7960 30645 8000
rect 30603 7951 30645 7960
rect 30411 7916 30453 7925
rect 30411 7876 30412 7916
rect 30452 7876 30453 7916
rect 30411 7867 30453 7876
rect 30027 7580 30069 7589
rect 29644 7279 29684 7288
rect 29932 7540 30028 7580
rect 30068 7540 30069 7580
rect 29548 7244 29588 7253
rect 29548 7169 29588 7204
rect 29739 7244 29781 7253
rect 29739 7204 29740 7244
rect 29780 7204 29781 7244
rect 29739 7195 29781 7204
rect 29452 7111 29492 7120
rect 29547 7160 29589 7169
rect 29547 7120 29548 7160
rect 29588 7120 29589 7160
rect 29547 7111 29589 7120
rect 29451 6824 29493 6833
rect 29451 6784 29452 6824
rect 29492 6784 29493 6824
rect 29451 6775 29493 6784
rect 29355 6740 29397 6749
rect 29355 6700 29356 6740
rect 29396 6700 29397 6740
rect 29355 6691 29397 6700
rect 28780 6439 28820 6448
rect 28971 6488 29013 6497
rect 28971 6448 28972 6488
rect 29012 6448 29013 6488
rect 28971 6439 29013 6448
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 29260 6488 29300 6497
rect 29356 6488 29396 6691
rect 29300 6448 29396 6488
rect 29452 6488 29492 6775
rect 29548 6656 29588 7111
rect 29740 7110 29780 7195
rect 29836 7160 29876 7169
rect 29836 6917 29876 7120
rect 29835 6908 29877 6917
rect 29835 6868 29836 6908
rect 29876 6868 29877 6908
rect 29835 6859 29877 6868
rect 29548 6616 29780 6656
rect 29260 6439 29300 6448
rect 29452 6439 29492 6448
rect 29644 6488 29684 6497
rect 28588 6354 28628 6439
rect 28972 6354 29012 6439
rect 29164 6354 29204 6439
rect 29547 6404 29589 6413
rect 29547 6364 29548 6404
rect 29588 6364 29589 6404
rect 29547 6355 29589 6364
rect 29548 6270 29588 6355
rect 29644 6329 29684 6448
rect 29740 6413 29780 6616
rect 29836 6488 29876 6497
rect 29739 6404 29781 6413
rect 29836 6404 29876 6448
rect 29932 6488 29972 7540
rect 30027 7531 30069 7540
rect 30219 7580 30261 7589
rect 30219 7540 30220 7580
rect 30260 7540 30261 7580
rect 30219 7531 30261 7540
rect 30123 7496 30165 7505
rect 30123 7456 30124 7496
rect 30164 7456 30165 7496
rect 30123 7447 30165 7456
rect 30027 7328 30069 7337
rect 30027 7288 30028 7328
rect 30068 7288 30069 7328
rect 30027 7279 30069 7288
rect 30028 7160 30068 7279
rect 30124 7244 30164 7447
rect 30412 7337 30452 7867
rect 30507 7496 30549 7505
rect 30507 7456 30508 7496
rect 30548 7456 30549 7496
rect 30507 7447 30549 7456
rect 30124 7195 30164 7204
rect 30220 7328 30260 7337
rect 30028 7111 30068 7120
rect 30220 6833 30260 7288
rect 30411 7328 30453 7337
rect 30411 7288 30412 7328
rect 30452 7288 30453 7328
rect 30411 7279 30453 7288
rect 30316 7244 30356 7253
rect 30316 6917 30356 7204
rect 30411 7160 30453 7169
rect 30411 7120 30412 7160
rect 30452 7120 30453 7160
rect 30411 7111 30453 7120
rect 30412 7026 30452 7111
rect 30315 6908 30357 6917
rect 30315 6868 30316 6908
rect 30356 6868 30357 6908
rect 30315 6859 30357 6868
rect 30219 6824 30261 6833
rect 30219 6784 30220 6824
rect 30260 6784 30261 6824
rect 30219 6775 30261 6784
rect 30123 6740 30165 6749
rect 30123 6700 30124 6740
rect 30164 6700 30165 6740
rect 30123 6691 30165 6700
rect 30124 6656 30164 6691
rect 30124 6605 30164 6616
rect 29972 6448 30164 6488
rect 29932 6439 29972 6448
rect 29739 6364 29740 6404
rect 29780 6364 29876 6404
rect 29739 6355 29781 6364
rect 29643 6320 29685 6329
rect 29643 6280 29644 6320
rect 29684 6280 29685 6320
rect 29643 6271 29685 6280
rect 28588 6236 28628 6245
rect 28204 5648 28244 5657
rect 28107 5144 28149 5153
rect 28107 5104 28108 5144
rect 28148 5104 28149 5144
rect 28107 5095 28149 5104
rect 27916 4649 27956 4936
rect 28108 4892 28148 4901
rect 27915 4640 27957 4649
rect 27915 4600 27916 4640
rect 27956 4600 27957 4640
rect 27915 4591 27957 4600
rect 28108 4481 28148 4852
rect 28204 4733 28244 5608
rect 28396 5648 28436 5657
rect 28300 5480 28340 5489
rect 28300 5069 28340 5440
rect 28299 5060 28341 5069
rect 28299 5020 28300 5060
rect 28340 5020 28341 5060
rect 28299 5011 28341 5020
rect 28396 4901 28436 5608
rect 28491 5648 28533 5657
rect 28491 5608 28492 5648
rect 28532 5608 28533 5648
rect 28491 5599 28533 5608
rect 28492 5514 28532 5599
rect 28395 4892 28437 4901
rect 28395 4852 28396 4892
rect 28436 4852 28437 4892
rect 28395 4843 28437 4852
rect 28203 4724 28245 4733
rect 28203 4684 28204 4724
rect 28244 4684 28245 4724
rect 28203 4675 28245 4684
rect 28107 4472 28149 4481
rect 28107 4432 28108 4472
rect 28148 4432 28149 4472
rect 28107 4423 28149 4432
rect 28300 4304 28340 4313
rect 28588 4304 28628 6196
rect 28972 6236 29012 6245
rect 29012 6196 29108 6236
rect 28972 6187 29012 6196
rect 28972 5657 29012 5742
rect 28876 5648 28916 5657
rect 28779 5480 28821 5489
rect 28876 5480 28916 5608
rect 28971 5648 29013 5657
rect 28971 5608 28972 5648
rect 29012 5608 29013 5648
rect 28971 5599 29013 5608
rect 28779 5440 28780 5480
rect 28820 5440 28916 5480
rect 28971 5480 29013 5489
rect 28971 5440 28972 5480
rect 29012 5440 29013 5480
rect 28779 5431 28821 5440
rect 28971 5431 29013 5440
rect 28779 5228 28821 5237
rect 28779 5188 28780 5228
rect 28820 5188 28821 5228
rect 28779 5179 28821 5188
rect 28780 5060 28820 5179
rect 28780 5011 28820 5020
rect 28684 4976 28724 4985
rect 28684 4397 28724 4936
rect 28875 4976 28917 4985
rect 28875 4936 28876 4976
rect 28916 4936 28917 4976
rect 28875 4927 28917 4936
rect 28972 4976 29012 5431
rect 28972 4927 29012 4936
rect 28876 4842 28916 4927
rect 29068 4817 29108 6196
rect 29644 5648 29684 5657
rect 29452 5608 29644 5648
rect 29259 5480 29301 5489
rect 29259 5440 29260 5480
rect 29300 5440 29301 5480
rect 29259 5431 29301 5440
rect 29260 5346 29300 5431
rect 29163 5144 29205 5153
rect 29163 5104 29164 5144
rect 29204 5104 29205 5144
rect 29163 5095 29205 5104
rect 29260 5144 29300 5153
rect 29452 5144 29492 5608
rect 29644 5599 29684 5608
rect 29740 5648 29780 5657
rect 29740 5489 29780 5608
rect 29836 5648 29876 5657
rect 29739 5480 29781 5489
rect 29739 5440 29740 5480
rect 29780 5440 29781 5480
rect 29739 5431 29781 5440
rect 29547 5312 29589 5321
rect 29547 5272 29548 5312
rect 29588 5272 29589 5312
rect 29547 5263 29589 5272
rect 29300 5104 29492 5144
rect 29164 4976 29204 5095
rect 29260 4985 29300 5104
rect 29164 4927 29204 4936
rect 29259 4976 29301 4985
rect 29259 4936 29260 4976
rect 29300 4936 29301 4976
rect 29259 4927 29301 4936
rect 29356 4976 29396 4987
rect 29356 4901 29396 4936
rect 29451 4976 29493 4985
rect 29451 4936 29452 4976
rect 29492 4936 29493 4976
rect 29451 4927 29493 4936
rect 29355 4892 29397 4901
rect 29355 4852 29356 4892
rect 29396 4852 29397 4892
rect 29355 4843 29397 4852
rect 29067 4808 29109 4817
rect 29067 4768 29068 4808
rect 29108 4768 29109 4808
rect 29067 4759 29109 4768
rect 28971 4724 29013 4733
rect 28971 4684 28972 4724
rect 29012 4684 29013 4724
rect 28971 4675 29013 4684
rect 28779 4640 28821 4649
rect 28779 4600 28780 4640
rect 28820 4600 28821 4640
rect 28779 4591 28821 4600
rect 28683 4388 28725 4397
rect 28683 4348 28684 4388
rect 28724 4348 28725 4388
rect 28683 4339 28725 4348
rect 27820 4264 28300 4304
rect 27820 4136 27860 4264
rect 27820 4087 27860 4096
rect 27916 4136 27956 4145
rect 27916 3809 27956 4096
rect 28107 4136 28149 4145
rect 28107 4096 28108 4136
rect 28148 4096 28149 4136
rect 28107 4087 28149 4096
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 28012 3918 28052 4003
rect 28108 4002 28148 4087
rect 27915 3800 27957 3809
rect 27915 3760 27916 3800
rect 27956 3760 27957 3800
rect 27915 3751 27957 3760
rect 28108 3473 28148 3558
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 27916 3464 27956 3473
rect 27820 3221 27860 3415
rect 27916 3296 27956 3424
rect 28107 3464 28149 3473
rect 28107 3424 28108 3464
rect 28148 3424 28149 3464
rect 28107 3415 28149 3424
rect 28204 3464 28244 4264
rect 28300 4255 28340 4264
rect 28396 4264 28628 4304
rect 28396 4145 28436 4264
rect 28395 4136 28437 4145
rect 28395 4096 28396 4136
rect 28436 4096 28437 4136
rect 28395 4087 28437 4096
rect 28587 4136 28629 4145
rect 28587 4096 28588 4136
rect 28628 4096 28629 4136
rect 28587 4087 28629 4096
rect 28684 4136 28724 4145
rect 28780 4136 28820 4591
rect 28724 4096 28820 4136
rect 28684 4087 28724 4096
rect 28588 4002 28628 4087
rect 28780 3910 28820 3919
rect 28587 3884 28629 3893
rect 28587 3844 28588 3884
rect 28628 3844 28629 3884
rect 28587 3835 28629 3844
rect 28491 3716 28533 3725
rect 28491 3676 28492 3716
rect 28532 3676 28533 3716
rect 28491 3667 28533 3676
rect 28204 3296 28244 3424
rect 27916 3256 28244 3296
rect 28300 3464 28340 3473
rect 27819 3212 27861 3221
rect 27819 3172 27820 3212
rect 27860 3172 27861 3212
rect 27819 3163 27861 3172
rect 27915 3128 27957 3137
rect 27915 3088 27916 3128
rect 27956 3088 27957 3128
rect 27915 3079 27957 3088
rect 27916 2624 27956 3079
rect 28011 3044 28053 3053
rect 28011 3004 28012 3044
rect 28052 3004 28053 3044
rect 28011 2995 28053 3004
rect 27916 2575 27956 2584
rect 28012 1952 28052 2995
rect 28300 2885 28340 3424
rect 28395 3464 28437 3473
rect 28395 3424 28396 3464
rect 28436 3424 28437 3464
rect 28395 3415 28437 3424
rect 28396 3330 28436 3415
rect 28299 2876 28341 2885
rect 28299 2836 28300 2876
rect 28340 2836 28341 2876
rect 28299 2827 28341 2836
rect 28108 2633 28148 2718
rect 28107 2624 28149 2633
rect 28107 2584 28108 2624
rect 28148 2584 28149 2624
rect 28107 2575 28149 2584
rect 28492 2624 28532 3667
rect 28588 3632 28628 3835
rect 28780 3632 28820 3870
rect 28972 3641 29012 4675
rect 29068 4145 29108 4759
rect 29067 4136 29109 4145
rect 29067 4096 29068 4136
rect 29108 4096 29109 4136
rect 29067 4087 29109 4096
rect 29260 4136 29300 4145
rect 29068 3968 29108 3977
rect 29068 3893 29108 3928
rect 29067 3884 29109 3893
rect 29067 3844 29068 3884
rect 29108 3844 29109 3884
rect 29067 3835 29109 3844
rect 29068 3833 29108 3835
rect 29163 3800 29205 3809
rect 29163 3760 29164 3800
rect 29204 3760 29205 3800
rect 29163 3751 29205 3760
rect 28876 3632 28916 3641
rect 28780 3592 28876 3632
rect 28588 3583 28628 3592
rect 28876 3583 28916 3592
rect 28971 3632 29013 3641
rect 28971 3592 28972 3632
rect 29012 3592 29013 3632
rect 28971 3583 29013 3592
rect 29164 3632 29204 3751
rect 29260 3725 29300 4096
rect 29356 3893 29396 4843
rect 29452 4649 29492 4927
rect 29451 4640 29493 4649
rect 29451 4600 29452 4640
rect 29492 4600 29493 4640
rect 29451 4591 29493 4600
rect 29548 4472 29588 5263
rect 29836 5237 29876 5608
rect 29932 5480 29972 5489
rect 29972 5440 30068 5480
rect 29932 5431 29972 5440
rect 29835 5228 29877 5237
rect 29835 5188 29836 5228
rect 29876 5188 29877 5228
rect 29835 5179 29877 5188
rect 30028 5069 30068 5440
rect 29834 5060 29876 5069
rect 29834 5020 29835 5060
rect 29875 5020 29876 5060
rect 29834 5011 29876 5020
rect 30027 5060 30069 5069
rect 30027 5020 30028 5060
rect 30068 5020 30069 5060
rect 30027 5011 30069 5020
rect 29644 4976 29684 4987
rect 29644 4901 29684 4936
rect 29739 4976 29781 4985
rect 29739 4936 29740 4976
rect 29780 4936 29781 4976
rect 29739 4927 29781 4936
rect 29836 4976 29876 5011
rect 29836 4927 29876 4936
rect 29931 4976 29973 4985
rect 29931 4936 29932 4976
rect 29972 4936 29973 4976
rect 29931 4927 29973 4936
rect 29643 4892 29685 4901
rect 29643 4852 29644 4892
rect 29684 4852 29685 4892
rect 29643 4843 29685 4852
rect 29740 4842 29780 4927
rect 29932 4842 29972 4927
rect 29452 4432 29588 4472
rect 29355 3884 29397 3893
rect 29355 3844 29356 3884
rect 29396 3844 29397 3884
rect 29355 3835 29397 3844
rect 29259 3716 29301 3725
rect 29259 3676 29260 3716
rect 29300 3676 29301 3716
rect 29259 3667 29301 3676
rect 29164 3583 29204 3592
rect 28683 3548 28725 3557
rect 28683 3508 28684 3548
rect 28724 3508 28725 3548
rect 28683 3499 28725 3508
rect 28492 2575 28532 2584
rect 28684 3464 28724 3499
rect 28588 2540 28628 2549
rect 28684 2540 28724 3424
rect 28972 2633 29012 3583
rect 29260 3548 29300 3557
rect 29260 3389 29300 3508
rect 29355 3464 29397 3473
rect 29355 3424 29356 3464
rect 29396 3424 29397 3464
rect 29355 3415 29397 3424
rect 29452 3464 29492 4432
rect 29547 4220 29589 4229
rect 29547 4180 29548 4220
rect 29588 4180 29589 4220
rect 29547 4171 29589 4180
rect 29548 4136 29588 4171
rect 29548 4085 29588 4096
rect 29739 3968 29781 3977
rect 29739 3928 29740 3968
rect 29780 3928 29781 3968
rect 29739 3919 29781 3928
rect 29643 3884 29685 3893
rect 29643 3844 29644 3884
rect 29684 3844 29685 3884
rect 29643 3835 29685 3844
rect 29452 3415 29492 3424
rect 29644 3464 29684 3835
rect 29740 3548 29780 3919
rect 29740 3499 29780 3508
rect 29644 3415 29684 3424
rect 29835 3464 29877 3473
rect 29835 3424 29836 3464
rect 29876 3424 29877 3464
rect 29835 3415 29877 3424
rect 29259 3380 29301 3389
rect 29259 3340 29260 3380
rect 29300 3340 29301 3380
rect 29259 3331 29301 3340
rect 29356 3330 29396 3415
rect 29836 3330 29876 3415
rect 29931 3380 29973 3389
rect 29931 3340 29932 3380
rect 29972 3340 29973 3380
rect 29931 3331 29973 3340
rect 29164 3212 29204 3221
rect 29932 3212 29972 3331
rect 28971 2624 29013 2633
rect 28971 2584 28972 2624
rect 29012 2584 29013 2624
rect 28971 2575 29013 2584
rect 29164 2624 29204 3172
rect 29836 3172 29972 3212
rect 29739 2792 29781 2801
rect 29739 2752 29740 2792
rect 29780 2752 29781 2792
rect 29739 2743 29781 2752
rect 29356 2633 29396 2718
rect 29164 2575 29204 2584
rect 29355 2624 29397 2633
rect 29355 2584 29356 2624
rect 29396 2584 29397 2624
rect 29355 2575 29397 2584
rect 29452 2624 29492 2633
rect 29644 2624 29684 2633
rect 29492 2584 29644 2624
rect 29452 2575 29492 2584
rect 29644 2575 29684 2584
rect 29740 2624 29780 2743
rect 29740 2575 29780 2584
rect 29836 2624 29876 3172
rect 30124 3053 30164 6448
rect 30219 5648 30261 5657
rect 30219 5608 30220 5648
rect 30260 5608 30261 5648
rect 30219 5599 30261 5608
rect 30220 5144 30260 5599
rect 30508 5489 30548 7447
rect 30604 7160 30644 7951
rect 30699 7328 30741 7337
rect 30699 7288 30700 7328
rect 30740 7288 30741 7328
rect 30699 7279 30741 7288
rect 30700 7202 30740 7279
rect 30700 7153 30740 7162
rect 30796 7160 30836 7169
rect 30604 7111 30644 7120
rect 30796 6917 30836 7120
rect 30892 7160 30932 7169
rect 30795 6908 30837 6917
rect 30795 6868 30796 6908
rect 30836 6868 30837 6908
rect 30795 6859 30837 6868
rect 30796 6749 30836 6859
rect 30795 6740 30837 6749
rect 30795 6700 30796 6740
rect 30836 6700 30837 6740
rect 30795 6691 30837 6700
rect 30892 6665 30932 7120
rect 30891 6656 30933 6665
rect 30891 6616 30892 6656
rect 30932 6616 30933 6656
rect 30891 6607 30933 6616
rect 30892 6497 30932 6607
rect 30891 6488 30933 6497
rect 30891 6448 30892 6488
rect 30932 6448 30933 6488
rect 30891 6439 30933 6448
rect 30603 5984 30645 5993
rect 30603 5944 30604 5984
rect 30644 5944 30645 5984
rect 30603 5935 30645 5944
rect 30507 5480 30549 5489
rect 30507 5440 30508 5480
rect 30548 5440 30549 5480
rect 30507 5431 30549 5440
rect 30220 5095 30260 5104
rect 30316 5144 30356 5153
rect 30316 4901 30356 5104
rect 30411 5144 30453 5153
rect 30411 5104 30412 5144
rect 30452 5104 30453 5144
rect 30411 5095 30453 5104
rect 30412 5060 30452 5095
rect 30412 5009 30452 5020
rect 30507 5060 30549 5069
rect 30507 5020 30508 5060
rect 30548 5020 30549 5060
rect 30507 5011 30549 5020
rect 30508 4976 30548 5011
rect 30508 4925 30548 4936
rect 30604 4976 30644 5935
rect 30988 5312 31028 8119
rect 31084 7505 31124 9211
rect 31083 7496 31125 7505
rect 31083 7456 31084 7496
rect 31124 7456 31125 7496
rect 31083 7447 31125 7456
rect 31180 7421 31220 10144
rect 31372 10016 31412 10144
rect 31563 10184 31605 10193
rect 31563 10144 31564 10184
rect 31604 10144 31605 10184
rect 31563 10135 31605 10144
rect 31660 10134 31700 10219
rect 31756 10184 31796 10303
rect 31756 10135 31796 10144
rect 31563 10016 31605 10025
rect 31372 9976 31564 10016
rect 31604 9976 31605 10016
rect 31563 9967 31605 9976
rect 31755 9764 31797 9773
rect 31755 9724 31756 9764
rect 31796 9724 31797 9764
rect 31755 9715 31797 9724
rect 31275 9596 31317 9605
rect 31275 9556 31276 9596
rect 31316 9556 31317 9596
rect 31275 9547 31317 9556
rect 31276 9512 31316 9547
rect 31276 9461 31316 9472
rect 31660 9512 31700 9523
rect 31660 9437 31700 9472
rect 31372 9428 31412 9437
rect 31275 9344 31317 9353
rect 31275 9304 31276 9344
rect 31316 9304 31317 9344
rect 31275 9295 31317 9304
rect 31276 8000 31316 9295
rect 31372 9269 31412 9388
rect 31564 9428 31604 9437
rect 31468 9344 31508 9353
rect 31371 9260 31413 9269
rect 31371 9220 31372 9260
rect 31412 9220 31413 9260
rect 31371 9211 31413 9220
rect 31371 8840 31413 8849
rect 31371 8800 31372 8840
rect 31412 8800 31413 8840
rect 31371 8791 31413 8800
rect 31372 8000 31412 8791
rect 31468 8681 31508 9304
rect 31564 9101 31604 9388
rect 31659 9428 31701 9437
rect 31659 9388 31660 9428
rect 31700 9388 31701 9428
rect 31659 9379 31701 9388
rect 31563 9092 31605 9101
rect 31563 9052 31564 9092
rect 31604 9052 31605 9092
rect 31563 9043 31605 9052
rect 31563 8924 31605 8933
rect 31563 8884 31564 8924
rect 31604 8884 31605 8924
rect 31563 8875 31605 8884
rect 31564 8840 31604 8875
rect 31564 8789 31604 8800
rect 31467 8672 31509 8681
rect 31467 8632 31468 8672
rect 31508 8632 31509 8672
rect 31467 8623 31509 8632
rect 31660 8672 31700 8681
rect 31660 8009 31700 8632
rect 31468 8000 31508 8009
rect 31372 7960 31468 8000
rect 31276 7951 31316 7960
rect 31468 7951 31508 7960
rect 31659 8000 31701 8009
rect 31659 7960 31660 8000
rect 31700 7960 31701 8000
rect 31659 7951 31701 7960
rect 31468 7832 31508 7841
rect 31179 7412 31221 7421
rect 31179 7372 31180 7412
rect 31220 7372 31221 7412
rect 31179 7363 31221 7372
rect 31372 7328 31412 7337
rect 31372 6908 31412 7288
rect 31084 6868 31412 6908
rect 31084 5993 31124 6868
rect 31275 6740 31317 6749
rect 31275 6700 31276 6740
rect 31316 6700 31317 6740
rect 31275 6691 31317 6700
rect 31276 6488 31316 6691
rect 31371 6572 31413 6581
rect 31371 6532 31372 6572
rect 31412 6532 31413 6572
rect 31371 6523 31413 6532
rect 31276 6439 31316 6448
rect 31372 6438 31412 6523
rect 31468 6497 31508 7792
rect 31660 7589 31700 7951
rect 31659 7580 31701 7589
rect 31659 7540 31660 7580
rect 31700 7540 31701 7580
rect 31659 7531 31701 7540
rect 31756 7421 31796 9715
rect 31852 9596 31892 11815
rect 31948 11696 31988 11707
rect 31948 11621 31988 11656
rect 32139 11696 32181 11705
rect 32139 11656 32140 11696
rect 32180 11656 32181 11696
rect 32139 11647 32181 11656
rect 32236 11696 32276 12412
rect 32332 11873 32372 12496
rect 32524 12536 32564 12545
rect 32524 12293 32564 12496
rect 32523 12284 32565 12293
rect 32523 12244 32524 12284
rect 32564 12244 32565 12284
rect 32523 12235 32565 12244
rect 32331 11864 32373 11873
rect 32331 11824 32332 11864
rect 32372 11824 32373 11864
rect 32331 11815 32373 11824
rect 31947 11612 31989 11621
rect 31947 11572 31948 11612
rect 31988 11572 31989 11612
rect 31947 11563 31989 11572
rect 31948 11024 31988 11033
rect 31948 10361 31988 10984
rect 32140 10982 32180 11647
rect 32236 11621 32276 11656
rect 32428 11696 32468 11705
rect 32235 11612 32277 11621
rect 32235 11572 32236 11612
rect 32276 11572 32277 11612
rect 32235 11563 32277 11572
rect 32428 11537 32468 11656
rect 32524 11696 32564 12235
rect 32620 11957 32660 13336
rect 32812 13217 32852 13922
rect 32908 13880 32948 14335
rect 33003 14048 33045 14057
rect 33003 14008 33004 14048
rect 33044 14008 33045 14048
rect 33003 13999 33045 14008
rect 33100 14048 33140 14680
rect 33196 14670 33236 14755
rect 33292 14561 33332 14848
rect 33388 14804 33428 14813
rect 33291 14552 33333 14561
rect 33291 14512 33292 14552
rect 33332 14512 33333 14552
rect 33291 14503 33333 14512
rect 33388 14225 33428 14764
rect 33484 14720 33524 14729
rect 33484 14561 33524 14680
rect 33676 14720 33716 14731
rect 33676 14645 33716 14680
rect 33772 14720 33812 14729
rect 33675 14636 33717 14645
rect 33675 14596 33676 14636
rect 33716 14596 33717 14636
rect 33675 14587 33717 14596
rect 33483 14552 33525 14561
rect 33483 14512 33484 14552
rect 33524 14512 33525 14552
rect 33483 14503 33525 14512
rect 33675 14300 33717 14309
rect 33675 14260 33676 14300
rect 33716 14260 33717 14300
rect 33675 14251 33717 14260
rect 33387 14216 33429 14225
rect 33387 14176 33388 14216
rect 33428 14176 33429 14216
rect 33387 14167 33429 14176
rect 33579 14132 33621 14141
rect 33579 14092 33580 14132
rect 33620 14092 33621 14132
rect 33579 14083 33621 14092
rect 33292 14048 33332 14057
rect 33004 13964 33044 13999
rect 33004 13913 33044 13924
rect 32908 13831 32948 13840
rect 33003 13796 33045 13805
rect 33003 13756 33004 13796
rect 33044 13756 33045 13796
rect 33003 13747 33045 13756
rect 32907 13628 32949 13637
rect 32907 13588 32908 13628
rect 32948 13588 32949 13628
rect 32907 13579 32949 13588
rect 32908 13460 32948 13579
rect 32908 13411 32948 13420
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 33004 13208 33044 13747
rect 33100 13301 33140 14008
rect 33196 14008 33292 14048
rect 33196 13721 33236 14008
rect 33292 13999 33332 14008
rect 33387 14048 33429 14057
rect 33387 14008 33388 14048
rect 33428 14008 33429 14048
rect 33387 13999 33429 14008
rect 33388 13964 33428 13999
rect 33388 13913 33428 13924
rect 33483 13964 33525 13973
rect 33483 13924 33484 13964
rect 33524 13924 33525 13964
rect 33483 13915 33525 13924
rect 33580 13964 33620 14083
rect 33580 13915 33620 13924
rect 33676 14048 33716 14251
rect 33484 13880 33524 13915
rect 33484 13829 33524 13840
rect 33676 13796 33716 14008
rect 33772 13973 33812 14680
rect 33868 14720 33908 14923
rect 33868 14671 33908 14680
rect 33964 14720 34004 15511
rect 34060 15485 34100 15520
rect 34156 15560 34196 15595
rect 34252 15569 34292 15654
rect 34444 15569 34484 17695
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 34539 17072 34581 17081
rect 34539 17032 34540 17072
rect 34580 17032 34581 17072
rect 34539 17023 34581 17032
rect 34540 16938 34580 17023
rect 35116 16064 35156 19123
rect 35308 17837 35348 19711
rect 35596 19256 35636 19265
rect 35596 19013 35636 19216
rect 36556 19256 36596 19265
rect 36748 19256 36788 19804
rect 36844 19795 36884 19804
rect 36596 19216 36788 19256
rect 36556 19207 36596 19216
rect 35595 19004 35637 19013
rect 35595 18964 35596 19004
rect 35636 18964 35637 19004
rect 35595 18955 35637 18964
rect 35787 18584 35829 18593
rect 35787 18544 35788 18584
rect 35828 18544 35829 18584
rect 35787 18535 35829 18544
rect 35788 18450 35828 18535
rect 35980 17912 36020 17921
rect 35788 17872 35980 17912
rect 35307 17828 35349 17837
rect 35307 17788 35308 17828
rect 35348 17788 35349 17828
rect 35307 17779 35349 17788
rect 35308 17744 35348 17779
rect 35308 17694 35348 17704
rect 35691 16988 35733 16997
rect 35691 16948 35692 16988
rect 35732 16948 35733 16988
rect 35691 16939 35733 16948
rect 35692 16854 35732 16939
rect 35595 16400 35637 16409
rect 35595 16360 35596 16400
rect 35636 16360 35637 16400
rect 35595 16351 35637 16360
rect 35211 16316 35253 16325
rect 35211 16276 35212 16316
rect 35252 16276 35253 16316
rect 35211 16267 35253 16276
rect 35212 16182 35252 16267
rect 35020 16024 35156 16064
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 34156 15509 34196 15520
rect 34251 15560 34293 15569
rect 34251 15520 34252 15560
rect 34292 15520 34293 15560
rect 34251 15511 34293 15520
rect 34348 15560 34388 15569
rect 34059 15476 34101 15485
rect 34059 15436 34060 15476
rect 34100 15436 34101 15476
rect 34059 15427 34101 15436
rect 34251 15308 34293 15317
rect 34251 15268 34252 15308
rect 34292 15268 34293 15308
rect 34251 15259 34293 15268
rect 34155 15140 34197 15149
rect 34155 15100 34156 15140
rect 34196 15100 34197 15140
rect 34155 15091 34197 15100
rect 34059 14804 34101 14813
rect 34059 14764 34060 14804
rect 34100 14764 34101 14804
rect 34059 14755 34101 14764
rect 33964 14671 34004 14680
rect 34060 14477 34100 14755
rect 34156 14720 34196 15091
rect 34156 14671 34196 14680
rect 34252 14720 34292 15259
rect 34348 14720 34388 15520
rect 34443 15560 34485 15569
rect 34443 15520 34444 15560
rect 34484 15520 34485 15560
rect 34443 15511 34485 15520
rect 34540 15560 34580 15569
rect 34444 14972 34484 14981
rect 34540 14972 34580 15520
rect 34827 15140 34869 15149
rect 34827 15100 34828 15140
rect 34868 15100 34869 15140
rect 34827 15091 34869 15100
rect 34484 14932 34580 14972
rect 34444 14923 34484 14932
rect 34635 14888 34677 14897
rect 34635 14848 34636 14888
rect 34676 14848 34677 14888
rect 34635 14839 34677 14848
rect 34444 14720 34484 14729
rect 34348 14680 34444 14720
rect 34252 14671 34292 14680
rect 34444 14671 34484 14680
rect 34636 14720 34676 14839
rect 34636 14671 34676 14680
rect 34731 14720 34773 14729
rect 34731 14680 34732 14720
rect 34772 14680 34773 14720
rect 34731 14671 34773 14680
rect 34828 14720 34868 15091
rect 34828 14671 34868 14680
rect 34732 14586 34772 14671
rect 34059 14468 34101 14477
rect 34059 14428 34060 14468
rect 34100 14428 34101 14468
rect 34059 14419 34101 14428
rect 33867 14384 33909 14393
rect 33867 14344 33868 14384
rect 33908 14344 33909 14384
rect 33867 14335 33909 14344
rect 33868 14048 33908 14335
rect 34060 14141 34100 14419
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 34155 14300 34197 14309
rect 34155 14260 34156 14300
rect 34196 14260 34197 14300
rect 34155 14251 34197 14260
rect 34059 14132 34101 14141
rect 34059 14092 34060 14132
rect 34100 14092 34101 14132
rect 34059 14083 34101 14092
rect 33771 13964 33813 13973
rect 33771 13924 33772 13964
rect 33812 13924 33813 13964
rect 33771 13915 33813 13924
rect 33676 13756 33812 13796
rect 33195 13712 33237 13721
rect 33195 13672 33196 13712
rect 33236 13672 33237 13712
rect 33195 13663 33237 13672
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 33099 13292 33141 13301
rect 33099 13252 33100 13292
rect 33140 13252 33141 13292
rect 33099 13243 33141 13252
rect 33004 13159 33044 13168
rect 33579 13208 33621 13217
rect 33579 13168 33580 13208
rect 33620 13168 33621 13208
rect 33579 13159 33621 13168
rect 33676 13208 33716 13217
rect 33772 13208 33812 13756
rect 33868 13217 33908 14008
rect 34156 14048 34196 14251
rect 35020 14216 35060 16024
rect 35212 15560 35252 15569
rect 35404 15560 35444 15569
rect 35252 15520 35404 15560
rect 35212 15511 35252 15520
rect 35404 15511 35444 15520
rect 35115 14384 35157 14393
rect 35115 14344 35116 14384
rect 35156 14344 35157 14384
rect 35115 14335 35157 14344
rect 34828 14176 35060 14216
rect 34251 14132 34293 14141
rect 34251 14092 34252 14132
rect 34292 14092 34293 14132
rect 34251 14083 34293 14092
rect 34156 13999 34196 14008
rect 34060 13964 34100 13973
rect 34060 13376 34100 13924
rect 33964 13336 34100 13376
rect 33716 13168 33812 13208
rect 33867 13208 33909 13217
rect 33867 13168 33868 13208
rect 33908 13168 33909 13208
rect 33676 13159 33716 13168
rect 33867 13159 33909 13168
rect 33580 13074 33620 13159
rect 33867 13040 33909 13049
rect 33867 13000 33868 13040
rect 33908 13000 33909 13040
rect 33964 13040 34004 13336
rect 34060 13208 34100 13217
rect 34252 13208 34292 14083
rect 34443 13544 34485 13553
rect 34443 13504 34444 13544
rect 34484 13504 34485 13544
rect 34443 13495 34485 13504
rect 34444 13385 34484 13495
rect 34443 13376 34485 13385
rect 34443 13336 34444 13376
rect 34484 13336 34485 13376
rect 34443 13327 34485 13336
rect 34348 13217 34388 13302
rect 34100 13168 34292 13208
rect 34347 13208 34389 13217
rect 34347 13168 34348 13208
rect 34388 13168 34389 13208
rect 34060 13159 34100 13168
rect 34347 13159 34389 13168
rect 34156 13040 34196 13049
rect 33964 13000 34100 13040
rect 33867 12991 33909 13000
rect 33868 12906 33908 12991
rect 33195 12536 33237 12545
rect 33195 12496 33196 12536
rect 33236 12496 33237 12536
rect 33195 12487 33237 12496
rect 34060 12536 34100 13000
rect 34060 12487 34100 12496
rect 34156 12536 34196 13000
rect 34347 13040 34389 13049
rect 34347 13000 34348 13040
rect 34388 13000 34389 13040
rect 34347 12991 34389 13000
rect 34251 12620 34293 12629
rect 34251 12580 34252 12620
rect 34292 12580 34293 12620
rect 34251 12571 34293 12580
rect 34156 12487 34196 12496
rect 32619 11948 32661 11957
rect 32619 11908 32620 11948
rect 32660 11908 32661 11948
rect 32619 11899 32661 11908
rect 33003 11864 33045 11873
rect 33003 11824 33004 11864
rect 33044 11824 33045 11864
rect 33003 11815 33045 11824
rect 32427 11528 32469 11537
rect 32427 11488 32428 11528
rect 32468 11488 32469 11528
rect 32427 11479 32469 11488
rect 32524 11453 32564 11656
rect 32620 11696 32660 11705
rect 32523 11444 32565 11453
rect 32523 11404 32524 11444
rect 32564 11404 32567 11444
rect 32523 11395 32567 11404
rect 32527 11360 32567 11395
rect 32620 11360 32660 11656
rect 32907 11696 32949 11705
rect 32907 11656 32908 11696
rect 32948 11656 32949 11696
rect 32907 11647 32949 11656
rect 33004 11696 33044 11815
rect 32715 11612 32757 11621
rect 32715 11572 32716 11612
rect 32756 11572 32757 11612
rect 32715 11563 32757 11572
rect 32716 11478 32756 11563
rect 32908 11562 32948 11647
rect 32811 11528 32853 11537
rect 32811 11488 32812 11528
rect 32852 11488 32853 11528
rect 32811 11479 32853 11488
rect 32527 11320 32574 11360
rect 32620 11320 32756 11360
rect 32331 11276 32373 11285
rect 32331 11236 32332 11276
rect 32372 11236 32373 11276
rect 32534 11276 32574 11320
rect 32534 11236 32660 11276
rect 32331 11227 32373 11236
rect 32332 11024 32372 11227
rect 32427 11192 32469 11201
rect 32427 11152 32428 11192
rect 32468 11152 32469 11192
rect 32427 11143 32469 11152
rect 32222 10982 32262 10991
rect 32043 10940 32085 10949
rect 32140 10942 32222 10982
rect 32332 10975 32372 10984
rect 32043 10900 32044 10940
rect 32084 10900 32085 10940
rect 32222 10933 32262 10942
rect 32043 10891 32085 10900
rect 32044 10806 32084 10891
rect 32140 10814 32180 10823
rect 32140 10529 32180 10774
rect 32428 10772 32468 11143
rect 32523 11024 32565 11033
rect 32523 10984 32524 11024
rect 32564 10984 32565 11024
rect 32523 10975 32565 10984
rect 32524 10890 32564 10975
rect 32620 10940 32660 11236
rect 32716 11201 32756 11320
rect 32715 11192 32757 11201
rect 32715 11152 32716 11192
rect 32756 11152 32757 11192
rect 32715 11143 32757 11152
rect 32715 11024 32757 11033
rect 32715 10984 32716 11024
rect 32756 10984 32757 11024
rect 32715 10975 32757 10984
rect 32620 10891 32660 10900
rect 32716 10856 32756 10975
rect 32716 10807 32756 10816
rect 32812 10940 32852 11479
rect 33004 11360 33044 11656
rect 32908 11320 33044 11360
rect 32908 11024 32948 11320
rect 33196 11285 33236 12487
rect 34252 12368 34292 12571
rect 34348 12536 34388 12991
rect 34444 12629 34484 13327
rect 34828 13217 34868 14176
rect 34924 14048 34964 14057
rect 34924 13805 34964 14008
rect 35020 14048 35060 14176
rect 35020 13999 35060 14008
rect 34923 13796 34965 13805
rect 34923 13756 34924 13796
rect 34964 13756 34965 13796
rect 34923 13747 34965 13756
rect 34827 13208 34869 13217
rect 34827 13168 34828 13208
rect 34868 13168 34869 13208
rect 34827 13159 34869 13168
rect 34924 13208 34964 13219
rect 34924 13133 34964 13168
rect 35020 13208 35060 13217
rect 35116 13208 35156 14335
rect 35212 14216 35252 14225
rect 35212 13889 35252 14176
rect 35403 14048 35445 14057
rect 35403 14008 35404 14048
rect 35444 14008 35445 14048
rect 35403 13999 35445 14008
rect 35404 13914 35444 13999
rect 35211 13880 35253 13889
rect 35211 13840 35212 13880
rect 35252 13840 35253 13880
rect 35211 13831 35253 13840
rect 35596 13376 35636 16351
rect 35788 15560 35828 17872
rect 35980 17863 36020 17872
rect 36555 17072 36597 17081
rect 36555 17032 36556 17072
rect 36596 17032 36597 17072
rect 36555 17023 36597 17032
rect 36652 17072 36692 17083
rect 36459 16988 36501 16997
rect 36459 16948 36460 16988
rect 36500 16948 36501 16988
rect 36459 16939 36501 16948
rect 35980 16820 36020 16829
rect 35980 16232 36020 16780
rect 35980 16183 36020 16192
rect 35788 15511 35828 15520
rect 35979 15224 36021 15233
rect 35979 15184 35980 15224
rect 36020 15184 36021 15224
rect 35979 15175 36021 15184
rect 35980 14300 36020 15175
rect 35692 14260 36020 14300
rect 35692 14048 35732 14260
rect 35884 14057 35924 14142
rect 35692 13999 35732 14008
rect 35883 14048 35925 14057
rect 35883 14008 35884 14048
rect 35924 14008 35925 14048
rect 35883 13999 35925 14008
rect 35980 14048 36020 14260
rect 36172 14216 36212 14225
rect 36172 14057 36212 14176
rect 35980 13999 36020 14008
rect 36171 14048 36213 14057
rect 36364 14048 36404 14057
rect 36171 14008 36172 14048
rect 36212 14008 36213 14048
rect 36171 13999 36213 14008
rect 36268 14008 36364 14048
rect 35692 13880 35732 13889
rect 36268 13880 36308 14008
rect 36364 13999 36404 14008
rect 35732 13840 36308 13880
rect 35692 13831 35732 13840
rect 36364 13796 36404 13805
rect 36268 13756 36364 13796
rect 35596 13336 35828 13376
rect 35060 13168 35156 13208
rect 35020 13159 35060 13168
rect 34923 13124 34965 13133
rect 34923 13084 34924 13124
rect 34964 13084 34965 13124
rect 34923 13075 34965 13084
rect 35019 13040 35061 13049
rect 35019 13000 35020 13040
rect 35060 13000 35061 13040
rect 35019 12991 35061 13000
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 35020 12629 35060 12991
rect 34443 12620 34485 12629
rect 34443 12580 34444 12620
rect 34484 12580 34485 12620
rect 34443 12571 34485 12580
rect 35019 12620 35061 12629
rect 35019 12580 35020 12620
rect 35060 12580 35061 12620
rect 35116 12620 35156 13168
rect 35211 13208 35253 13217
rect 35211 13168 35212 13208
rect 35252 13168 35253 13208
rect 35211 13159 35253 13168
rect 35404 13208 35444 13217
rect 35212 13040 35252 13159
rect 35212 12991 35252 13000
rect 35404 12704 35444 13168
rect 35500 13208 35540 13219
rect 35500 13133 35540 13168
rect 35499 13124 35541 13133
rect 35499 13084 35500 13124
rect 35540 13084 35541 13124
rect 35499 13075 35541 13084
rect 35596 12872 35636 13336
rect 35691 13208 35733 13217
rect 35691 13168 35692 13208
rect 35732 13168 35733 13208
rect 35691 13159 35733 13168
rect 35788 13208 35828 13336
rect 36171 13292 36213 13301
rect 36171 13252 36172 13292
rect 36212 13252 36213 13292
rect 36171 13243 36213 13252
rect 35889 13208 35929 13217
rect 35788 13159 35828 13168
rect 35884 13168 35889 13208
rect 35884 13159 35929 13168
rect 36172 13208 36212 13243
rect 35692 13074 35732 13159
rect 35787 13040 35829 13049
rect 35787 13000 35788 13040
rect 35828 13000 35829 13040
rect 35787 12991 35829 13000
rect 35788 12906 35828 12991
rect 35404 12655 35444 12664
rect 35500 12832 35636 12872
rect 35116 12580 35348 12620
rect 35019 12571 35061 12580
rect 34348 12487 34388 12496
rect 34444 12536 34484 12571
rect 34444 12486 34484 12496
rect 34599 12536 34639 12545
rect 34828 12536 34868 12545
rect 34639 12496 34828 12536
rect 34599 12487 34639 12496
rect 34252 12328 34388 12368
rect 34060 12284 34100 12293
rect 33964 12244 34060 12284
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 33291 11780 33333 11789
rect 33291 11740 33292 11780
rect 33332 11740 33333 11780
rect 33291 11731 33333 11740
rect 33195 11276 33237 11285
rect 33195 11236 33196 11276
rect 33236 11236 33237 11276
rect 33195 11227 33237 11236
rect 32908 10975 32948 10984
rect 33100 11024 33140 11033
rect 32428 10732 32660 10772
rect 32235 10604 32277 10613
rect 32235 10564 32236 10604
rect 32276 10564 32277 10604
rect 32235 10555 32277 10564
rect 32139 10520 32181 10529
rect 32139 10480 32140 10520
rect 32180 10480 32181 10520
rect 32139 10471 32181 10480
rect 31947 10352 31989 10361
rect 31947 10312 31948 10352
rect 31988 10312 31989 10352
rect 31947 10303 31989 10312
rect 31982 10191 32022 10200
rect 31948 10151 31982 10191
rect 31948 10142 32022 10151
rect 32140 10184 32180 10193
rect 31948 9941 31988 10142
rect 32140 10109 32180 10144
rect 32236 10184 32276 10555
rect 32523 10352 32565 10361
rect 32523 10312 32524 10352
rect 32564 10312 32565 10352
rect 32523 10303 32565 10312
rect 32236 10135 32276 10144
rect 32427 10184 32469 10193
rect 32427 10144 32428 10184
rect 32468 10144 32469 10184
rect 32427 10135 32469 10144
rect 32524 10184 32564 10303
rect 32620 10184 32660 10732
rect 32812 10529 32852 10900
rect 32907 10688 32949 10697
rect 32907 10648 32908 10688
rect 32948 10648 32949 10688
rect 32907 10639 32949 10648
rect 32811 10520 32853 10529
rect 32811 10480 32812 10520
rect 32852 10480 32853 10520
rect 32811 10471 32853 10480
rect 32811 10268 32853 10277
rect 32811 10228 32812 10268
rect 32852 10228 32853 10268
rect 32811 10219 32853 10228
rect 32716 10184 32756 10193
rect 32620 10144 32716 10184
rect 32524 10135 32564 10144
rect 32716 10135 32756 10144
rect 32139 10100 32181 10109
rect 32139 10060 32140 10100
rect 32180 10060 32181 10100
rect 32139 10051 32181 10060
rect 32044 10016 32084 10025
rect 31947 9932 31989 9941
rect 31947 9892 31948 9932
rect 31988 9892 31989 9932
rect 31947 9883 31989 9892
rect 31852 9556 31988 9596
rect 31948 9512 31988 9556
rect 32044 9521 32084 9976
rect 32044 9512 32092 9521
rect 32044 9472 32051 9512
rect 32091 9472 32092 9512
rect 31948 9344 31988 9472
rect 32050 9463 32092 9472
rect 31852 9304 31988 9344
rect 32043 9344 32085 9353
rect 32043 9304 32044 9344
rect 32084 9304 32085 9344
rect 31852 8420 31892 9304
rect 32043 9295 32085 9304
rect 31947 8840 31989 8849
rect 31947 8800 31948 8840
rect 31988 8800 31989 8840
rect 31947 8791 31989 8800
rect 31948 8672 31988 8791
rect 32044 8756 32084 9295
rect 32140 8933 32180 10051
rect 32428 10050 32468 10135
rect 32812 10134 32852 10219
rect 32908 10193 32948 10639
rect 33100 10613 33140 10984
rect 33195 11024 33237 11033
rect 33195 10984 33196 11024
rect 33236 10984 33237 11024
rect 33195 10975 33237 10984
rect 33292 11024 33332 11731
rect 33772 11696 33812 11705
rect 33387 11612 33429 11621
rect 33387 11572 33388 11612
rect 33428 11572 33429 11612
rect 33387 11563 33429 11572
rect 33292 10975 33332 10984
rect 33388 11024 33428 11563
rect 33675 11528 33717 11537
rect 33675 11488 33676 11528
rect 33716 11488 33717 11528
rect 33675 11479 33717 11488
rect 33676 11394 33716 11479
rect 33388 10975 33428 10984
rect 33196 10890 33236 10975
rect 33772 10865 33812 11656
rect 33868 11696 33908 11705
rect 33868 11537 33908 11656
rect 33964 11696 34004 12244
rect 34060 12235 34100 12244
rect 34155 12200 34197 12209
rect 34155 12160 34156 12200
rect 34196 12160 34197 12200
rect 34155 12151 34197 12160
rect 33964 11647 34004 11656
rect 34156 11696 34196 12151
rect 34251 11864 34293 11873
rect 34251 11824 34252 11864
rect 34292 11824 34293 11864
rect 34251 11815 34293 11824
rect 33867 11528 33909 11537
rect 33867 11488 33868 11528
rect 33908 11488 33909 11528
rect 33867 11479 33909 11488
rect 33867 11276 33909 11285
rect 33867 11236 33868 11276
rect 33908 11236 33909 11276
rect 33867 11227 33909 11236
rect 33771 10856 33813 10865
rect 33771 10816 33772 10856
rect 33812 10816 33813 10856
rect 33771 10807 33813 10816
rect 33099 10604 33141 10613
rect 33099 10564 33100 10604
rect 33140 10564 33141 10604
rect 33099 10555 33141 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 33003 10436 33045 10445
rect 33003 10396 33004 10436
rect 33044 10396 33045 10436
rect 33003 10387 33045 10396
rect 32907 10184 32949 10193
rect 32907 10144 32908 10184
rect 32948 10144 32949 10184
rect 33004 10184 33044 10387
rect 33100 10361 33140 10446
rect 33483 10436 33525 10445
rect 33483 10396 33484 10436
rect 33524 10396 33525 10436
rect 33483 10387 33525 10396
rect 33099 10352 33141 10361
rect 33099 10312 33100 10352
rect 33140 10312 33141 10352
rect 33099 10303 33141 10312
rect 33484 10302 33524 10387
rect 33100 10184 33140 10193
rect 33004 10144 33100 10184
rect 32907 10135 32949 10144
rect 33100 10135 33140 10144
rect 33292 10184 33332 10195
rect 32908 10050 32948 10135
rect 33292 10109 33332 10144
rect 33580 10184 33620 10193
rect 33291 10100 33333 10109
rect 33291 10060 33292 10100
rect 33332 10060 33333 10100
rect 33291 10051 33333 10060
rect 32619 10016 32661 10025
rect 32619 9976 32620 10016
rect 32660 9976 32661 10016
rect 32619 9967 32661 9976
rect 32235 9848 32277 9857
rect 32235 9808 32236 9848
rect 32276 9808 32277 9848
rect 32235 9799 32277 9808
rect 32236 9344 32276 9799
rect 32236 9295 32276 9304
rect 32428 9260 32468 9269
rect 32468 9220 32564 9260
rect 32428 9211 32468 9220
rect 32235 9008 32277 9017
rect 32235 8968 32236 9008
rect 32276 8968 32277 9008
rect 32235 8959 32277 8968
rect 32139 8924 32181 8933
rect 32139 8884 32140 8924
rect 32180 8884 32181 8924
rect 32139 8875 32181 8884
rect 32236 8840 32276 8959
rect 32044 8716 32180 8756
rect 31948 8623 31988 8632
rect 31852 8380 31988 8420
rect 31851 8252 31893 8261
rect 31851 8212 31852 8252
rect 31892 8212 31893 8252
rect 31851 8203 31893 8212
rect 31852 8000 31892 8203
rect 31852 7951 31892 7960
rect 31948 7916 31988 8380
rect 32140 7925 32180 8716
rect 32236 8000 32276 8800
rect 31948 7867 31988 7876
rect 32139 7916 32181 7925
rect 32139 7876 32140 7916
rect 32180 7876 32181 7916
rect 32139 7867 32181 7876
rect 32044 7832 32084 7841
rect 31755 7412 31797 7421
rect 32044 7412 32084 7792
rect 32140 7782 32180 7867
rect 31755 7372 31756 7412
rect 31796 7372 31797 7412
rect 31755 7363 31797 7372
rect 31852 7372 32084 7412
rect 31659 7328 31701 7337
rect 31659 7288 31660 7328
rect 31700 7288 31701 7328
rect 31659 7279 31701 7288
rect 31660 7160 31700 7279
rect 31564 7120 31660 7160
rect 31467 6488 31509 6497
rect 31467 6448 31468 6488
rect 31508 6448 31509 6488
rect 31467 6439 31509 6448
rect 31468 6354 31508 6439
rect 31564 6329 31604 7120
rect 31660 7111 31700 7120
rect 31756 7160 31796 7169
rect 31756 6581 31796 7120
rect 31852 6988 31892 7372
rect 32139 7328 32181 7337
rect 32139 7288 32140 7328
rect 32180 7288 32181 7328
rect 32139 7279 32181 7288
rect 32043 7160 32085 7169
rect 32043 7120 32044 7160
rect 32084 7120 32085 7160
rect 32043 7111 32085 7120
rect 31852 6939 31892 6948
rect 31755 6572 31797 6581
rect 31947 6572 31989 6581
rect 31755 6532 31756 6572
rect 31796 6532 31797 6572
rect 31755 6523 31797 6532
rect 31852 6532 31948 6572
rect 31988 6532 31989 6572
rect 31660 6488 31700 6497
rect 31563 6320 31605 6329
rect 31563 6280 31564 6320
rect 31604 6280 31605 6320
rect 31563 6271 31605 6280
rect 31564 6068 31604 6271
rect 31660 6245 31700 6448
rect 31852 6488 31892 6532
rect 31947 6523 31989 6532
rect 31852 6439 31892 6448
rect 32044 6488 32084 7111
rect 32044 6439 32084 6448
rect 32140 6404 32180 7279
rect 32236 7169 32276 7960
rect 32524 7589 32564 9220
rect 32523 7580 32565 7589
rect 32523 7540 32524 7580
rect 32564 7540 32565 7580
rect 32523 7531 32565 7540
rect 32523 7412 32565 7421
rect 32523 7372 32524 7412
rect 32564 7372 32565 7412
rect 32523 7363 32565 7372
rect 32331 7328 32373 7337
rect 32331 7288 32332 7328
rect 32372 7288 32373 7328
rect 32331 7279 32373 7288
rect 32428 7328 32468 7337
rect 32332 7244 32372 7279
rect 32332 7193 32372 7204
rect 32235 7160 32277 7169
rect 32235 7120 32236 7160
rect 32276 7120 32277 7160
rect 32235 7111 32277 7120
rect 32236 7026 32276 7111
rect 32428 6656 32468 7288
rect 32524 7244 32564 7363
rect 32524 6833 32564 7204
rect 32620 7160 32660 9967
rect 33580 9269 33620 10144
rect 33868 10184 33908 11227
rect 34156 10949 34196 11656
rect 34252 11696 34292 11815
rect 34252 11647 34292 11656
rect 34155 10940 34197 10949
rect 34155 10900 34156 10940
rect 34196 10900 34197 10940
rect 34155 10891 34197 10900
rect 34348 10865 34388 12328
rect 34444 11740 34772 11780
rect 34444 11528 34484 11740
rect 34732 11696 34772 11740
rect 34732 11647 34772 11656
rect 34828 11696 34868 12496
rect 34924 12536 34964 12545
rect 34924 12293 34964 12496
rect 35308 12536 35348 12580
rect 35308 12487 35348 12496
rect 35211 12452 35253 12461
rect 35211 12412 35212 12452
rect 35252 12412 35253 12452
rect 35211 12403 35253 12412
rect 34923 12284 34965 12293
rect 34923 12244 34924 12284
rect 34964 12244 34965 12284
rect 34923 12235 34965 12244
rect 34828 11647 34868 11656
rect 34923 11696 34965 11705
rect 35212 11696 35252 12403
rect 35500 11705 35540 12832
rect 35595 12620 35637 12629
rect 35595 12580 35596 12620
rect 35636 12580 35637 12620
rect 35595 12571 35637 12580
rect 35596 12536 35636 12571
rect 35596 12485 35636 12496
rect 34923 11656 34924 11696
rect 34964 11656 35060 11696
rect 34923 11647 34965 11656
rect 34636 11537 34676 11622
rect 34924 11562 34964 11647
rect 34444 11479 34484 11488
rect 34635 11528 34677 11537
rect 34635 11488 34636 11528
rect 34676 11488 34677 11528
rect 34635 11479 34677 11488
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 35020 11192 35060 11656
rect 35212 11647 35252 11656
rect 35499 11696 35541 11705
rect 35499 11656 35500 11696
rect 35540 11656 35541 11696
rect 35499 11647 35541 11656
rect 35308 11528 35348 11537
rect 35348 11488 35540 11528
rect 35308 11479 35348 11488
rect 34828 11152 35060 11192
rect 35211 11192 35253 11201
rect 35211 11152 35212 11192
rect 35252 11152 35253 11192
rect 34347 10856 34389 10865
rect 34347 10816 34348 10856
rect 34388 10816 34389 10856
rect 34347 10807 34389 10816
rect 34155 10268 34197 10277
rect 34155 10228 34156 10268
rect 34196 10228 34197 10268
rect 34155 10219 34197 10228
rect 33868 10135 33908 10144
rect 34156 10184 34196 10219
rect 34156 10133 34196 10144
rect 34348 10184 34388 10807
rect 34348 10135 34388 10144
rect 34539 10184 34581 10193
rect 34539 10144 34540 10184
rect 34580 10144 34581 10184
rect 34539 10135 34581 10144
rect 34636 10184 34676 10193
rect 34828 10184 34868 11152
rect 35211 11143 35253 11152
rect 35212 11058 35252 11143
rect 35307 11108 35349 11117
rect 35307 11068 35308 11108
rect 35348 11068 35349 11108
rect 35307 11059 35349 11068
rect 34923 11024 34965 11033
rect 34923 10984 34924 11024
rect 34964 10984 34965 11024
rect 34923 10975 34965 10984
rect 35020 11024 35060 11035
rect 34924 10890 34964 10975
rect 35020 10949 35060 10984
rect 35019 10940 35061 10949
rect 35019 10900 35020 10940
rect 35060 10900 35061 10940
rect 35019 10891 35061 10900
rect 35308 10529 35348 11059
rect 35500 11024 35540 11488
rect 35884 11201 35924 13159
rect 36172 13157 36212 13168
rect 36075 13040 36117 13049
rect 36075 13000 36076 13040
rect 36116 13000 36117 13040
rect 36075 12991 36117 13000
rect 35979 11528 36021 11537
rect 35979 11488 35980 11528
rect 36020 11488 36021 11528
rect 35979 11479 36021 11488
rect 35691 11192 35733 11201
rect 35691 11152 35692 11192
rect 35732 11152 35733 11192
rect 35691 11143 35733 11152
rect 35883 11192 35925 11201
rect 35883 11152 35884 11192
rect 35924 11152 35925 11192
rect 35883 11143 35925 11152
rect 35500 10975 35540 10984
rect 35596 11024 35636 11035
rect 35596 10949 35636 10984
rect 35692 11024 35732 11143
rect 35980 11108 36020 11479
rect 36076 11192 36116 12991
rect 36268 12536 36308 13756
rect 36364 13747 36404 13756
rect 36460 13460 36500 16939
rect 36556 15560 36596 17023
rect 36652 16997 36692 17032
rect 36651 16988 36693 16997
rect 36651 16948 36652 16988
rect 36692 16948 36693 16988
rect 36651 16939 36693 16948
rect 36651 16820 36693 16829
rect 36651 16780 36652 16820
rect 36692 16780 36693 16820
rect 36651 16771 36693 16780
rect 36652 16409 36692 16771
rect 36651 16400 36693 16409
rect 36651 16360 36652 16400
rect 36692 16360 36693 16400
rect 36651 16351 36693 16360
rect 36652 16232 36692 16241
rect 36652 15821 36692 16192
rect 36651 15812 36693 15821
rect 36651 15772 36652 15812
rect 36692 15772 36693 15812
rect 36651 15763 36693 15772
rect 36652 15560 36692 15569
rect 36556 15520 36652 15560
rect 36652 15511 36692 15520
rect 36748 15149 36788 19216
rect 36844 19256 36884 19265
rect 36940 19256 36980 20140
rect 37420 20105 37460 21568
rect 37612 21440 37652 23752
rect 37708 23743 37748 23752
rect 38187 23792 38229 23801
rect 38187 23752 38188 23792
rect 38228 23752 38229 23792
rect 38187 23743 38229 23752
rect 38284 23792 38324 25264
rect 38571 24632 38613 24641
rect 38571 24592 38572 24632
rect 38612 24592 38613 24632
rect 38571 24583 38613 24592
rect 38572 24498 38612 24583
rect 38668 24557 38708 26104
rect 38763 26104 38764 26144
rect 38804 26104 38805 26144
rect 38763 26095 38805 26104
rect 38860 26144 38900 26776
rect 38860 26095 38900 26104
rect 38956 26144 38996 30295
rect 39436 29840 39476 29849
rect 39436 29009 39476 29800
rect 39820 29840 39860 30379
rect 39820 29791 39860 29800
rect 40012 29765 40052 30388
rect 41644 30092 41684 30640
rect 41876 30640 41972 30680
rect 42700 30680 42740 30689
rect 41836 30631 41876 30640
rect 42700 30269 42740 30640
rect 41739 30260 41781 30269
rect 41739 30220 41740 30260
rect 41780 30220 41781 30260
rect 41739 30211 41781 30220
rect 42699 30260 42741 30269
rect 42699 30220 42700 30260
rect 42740 30220 42741 30260
rect 42699 30211 42741 30220
rect 41644 30043 41684 30052
rect 40492 30008 40532 30017
rect 40299 29840 40341 29849
rect 40299 29800 40300 29840
rect 40340 29800 40341 29840
rect 40299 29791 40341 29800
rect 40011 29756 40053 29765
rect 40011 29716 40012 29756
rect 40052 29716 40053 29756
rect 40011 29707 40053 29716
rect 39532 29168 39572 29177
rect 39435 29000 39477 29009
rect 39435 28960 39436 29000
rect 39476 28960 39477 29000
rect 39435 28951 39477 28960
rect 39532 28412 39572 29128
rect 39340 28372 39572 28412
rect 40204 29000 40244 29009
rect 40300 29000 40340 29791
rect 40395 29672 40437 29681
rect 40395 29632 40396 29672
rect 40436 29632 40437 29672
rect 40395 29623 40437 29632
rect 40396 29252 40436 29623
rect 40492 29588 40532 29968
rect 40780 29968 41492 30008
rect 40684 29849 40724 29934
rect 40683 29840 40725 29849
rect 40683 29800 40684 29840
rect 40724 29800 40725 29840
rect 40683 29791 40725 29800
rect 40780 29840 40820 29968
rect 40780 29791 40820 29800
rect 40972 29840 41012 29849
rect 41164 29840 41204 29849
rect 41012 29800 41164 29840
rect 40972 29791 41012 29800
rect 41164 29791 41204 29800
rect 41260 29840 41300 29849
rect 41260 29681 41300 29800
rect 41355 29840 41397 29849
rect 41355 29800 41356 29840
rect 41396 29800 41397 29840
rect 41355 29791 41397 29800
rect 41452 29840 41492 29968
rect 41356 29706 41396 29791
rect 40875 29672 40917 29681
rect 40875 29632 40876 29672
rect 40916 29632 40917 29672
rect 40875 29623 40917 29632
rect 41259 29672 41301 29681
rect 41259 29632 41260 29672
rect 41300 29632 41301 29672
rect 41259 29623 41301 29632
rect 40492 29548 40820 29588
rect 40396 29203 40436 29212
rect 40683 29252 40725 29261
rect 40683 29212 40684 29252
rect 40724 29212 40725 29252
rect 40683 29203 40725 29212
rect 40300 28960 40436 29000
rect 39243 28244 39285 28253
rect 39243 28204 39244 28244
rect 39284 28204 39285 28244
rect 39243 28195 39285 28204
rect 39148 26816 39188 26825
rect 39244 26816 39284 28195
rect 39340 27581 39380 28372
rect 39628 28160 39668 28169
rect 39532 27740 39572 27749
rect 39628 27740 39668 28120
rect 39572 27700 39668 27740
rect 39532 27691 39572 27700
rect 39916 27656 39956 27665
rect 39956 27616 40052 27656
rect 39916 27607 39956 27616
rect 39339 27572 39381 27581
rect 39339 27532 39340 27572
rect 39380 27532 39381 27572
rect 39339 27523 39381 27532
rect 39340 27438 39380 27523
rect 39627 27152 39669 27161
rect 39627 27112 39628 27152
rect 39668 27112 39669 27152
rect 39627 27103 39669 27112
rect 39435 27068 39477 27077
rect 39435 27028 39436 27068
rect 39476 27028 39477 27068
rect 39435 27019 39477 27028
rect 39436 26934 39476 27019
rect 39188 26776 39284 26816
rect 39436 26816 39476 26825
rect 39148 26767 39188 26776
rect 39436 26489 39476 26776
rect 39628 26816 39668 27103
rect 40012 26984 40052 27616
rect 40012 26935 40052 26944
rect 39051 26480 39093 26489
rect 39051 26440 39052 26480
rect 39092 26440 39093 26480
rect 39051 26431 39093 26440
rect 39435 26480 39477 26489
rect 39435 26440 39436 26480
rect 39476 26440 39477 26480
rect 39435 26431 39477 26440
rect 39052 26312 39092 26431
rect 39052 26263 39092 26272
rect 39628 26237 39668 26776
rect 39724 26816 39764 26825
rect 39147 26228 39189 26237
rect 39147 26188 39148 26228
rect 39188 26188 39189 26228
rect 39147 26179 39189 26188
rect 39627 26228 39669 26237
rect 39627 26188 39628 26228
rect 39668 26188 39669 26228
rect 39627 26179 39669 26188
rect 38764 26010 38804 26095
rect 38956 26069 38996 26104
rect 38955 26060 38997 26069
rect 38955 26020 38956 26060
rect 38996 26020 38997 26060
rect 38955 26011 38997 26020
rect 38956 25980 38996 26011
rect 38955 25304 38997 25313
rect 38955 25264 38956 25304
rect 38996 25264 38997 25304
rect 38955 25255 38997 25264
rect 39148 25304 39188 26179
rect 39339 26144 39381 26153
rect 39339 26104 39340 26144
rect 39380 26104 39381 26144
rect 39339 26095 39381 26104
rect 39340 25556 39380 26095
rect 39340 25313 39380 25516
rect 39148 25255 39188 25264
rect 39339 25304 39381 25313
rect 39339 25264 39340 25304
rect 39380 25264 39381 25304
rect 39339 25255 39381 25264
rect 38859 24716 38901 24725
rect 38859 24676 38860 24716
rect 38900 24676 38901 24716
rect 38859 24667 38901 24676
rect 38763 24632 38805 24641
rect 38763 24592 38764 24632
rect 38804 24592 38805 24632
rect 38763 24583 38805 24592
rect 38667 24548 38709 24557
rect 38667 24508 38668 24548
rect 38708 24508 38709 24548
rect 38667 24499 38709 24508
rect 38188 23658 38228 23743
rect 37780 22961 37820 22980
rect 37780 22952 37844 22961
rect 37708 22912 37804 22952
rect 37708 22280 37748 22912
rect 37804 22903 37844 22912
rect 37708 22231 37748 22240
rect 37995 21860 38037 21869
rect 37995 21820 37996 21860
rect 38036 21820 38037 21860
rect 37995 21811 38037 21820
rect 37900 21608 37940 21617
rect 37612 21400 37844 21440
rect 37804 20180 37844 21400
rect 37900 20936 37940 21568
rect 37996 21608 38036 21811
rect 38091 21692 38133 21701
rect 38091 21652 38092 21692
rect 38132 21652 38133 21692
rect 38091 21643 38133 21652
rect 37996 21559 38036 21568
rect 38092 21608 38132 21643
rect 38092 21557 38132 21568
rect 38187 21608 38229 21617
rect 38187 21568 38188 21608
rect 38228 21568 38229 21608
rect 38187 21559 38229 21568
rect 38188 21474 38228 21559
rect 38284 21113 38324 23752
rect 38572 23624 38612 23633
rect 38572 23120 38612 23584
rect 38668 23288 38708 24499
rect 38668 23239 38708 23248
rect 38572 23071 38612 23080
rect 38764 22373 38804 24583
rect 38860 24582 38900 24667
rect 38956 23120 38996 25255
rect 39051 24632 39093 24641
rect 39051 24587 39052 24632
rect 39092 24587 39093 24632
rect 39051 24583 39093 24587
rect 39531 24632 39573 24641
rect 39531 24592 39532 24632
rect 39572 24592 39573 24632
rect 39531 24583 39573 24592
rect 39052 24497 39092 24583
rect 39532 24498 39572 24583
rect 39724 24389 39764 26776
rect 40204 26657 40244 28960
rect 40300 28328 40340 28337
rect 40300 27077 40340 28288
rect 40299 27068 40341 27077
rect 40299 27028 40300 27068
rect 40340 27028 40341 27068
rect 40396 27068 40436 28960
rect 40684 28580 40724 29203
rect 40780 29168 40820 29548
rect 40876 29538 40916 29623
rect 40780 29119 40820 29128
rect 40875 28916 40917 28925
rect 40875 28876 40876 28916
rect 40916 28876 40917 28916
rect 40875 28867 40917 28876
rect 40780 28580 40820 28589
rect 40684 28540 40780 28580
rect 40780 28531 40820 28540
rect 40492 28328 40532 28337
rect 40492 27749 40532 28288
rect 40587 28328 40629 28337
rect 40587 28288 40588 28328
rect 40628 28288 40629 28328
rect 40587 28279 40629 28288
rect 40780 28328 40820 28337
rect 40876 28328 40916 28867
rect 40820 28288 40916 28328
rect 40972 28328 41012 28337
rect 40780 28279 40820 28288
rect 40588 28194 40628 28279
rect 40491 27740 40533 27749
rect 40491 27700 40492 27740
rect 40532 27700 40533 27740
rect 40491 27691 40533 27700
rect 40779 27656 40821 27665
rect 40779 27616 40780 27656
rect 40820 27616 40821 27656
rect 40779 27607 40821 27616
rect 40780 27522 40820 27607
rect 40972 27497 41012 28288
rect 40971 27488 41013 27497
rect 40971 27448 40972 27488
rect 41012 27448 41013 27488
rect 40971 27439 41013 27448
rect 40492 27068 40532 27077
rect 40396 27028 40492 27068
rect 40299 27019 40341 27028
rect 40492 27019 40532 27028
rect 40396 26816 40436 26825
rect 40396 26657 40436 26776
rect 41067 26816 41109 26825
rect 41067 26776 41068 26816
rect 41108 26776 41109 26816
rect 41067 26767 41109 26776
rect 41068 26682 41108 26767
rect 41260 26741 41300 29623
rect 41452 28841 41492 29800
rect 41644 29168 41684 29177
rect 41740 29168 41780 30211
rect 42316 29840 42356 29849
rect 42219 29756 42261 29765
rect 42219 29716 42220 29756
rect 42260 29716 42261 29756
rect 42219 29707 42261 29716
rect 41684 29128 41780 29168
rect 41644 29119 41684 29128
rect 42123 29084 42165 29093
rect 42123 29044 42124 29084
rect 42164 29044 42165 29084
rect 42123 29035 42165 29044
rect 41451 28832 41493 28841
rect 41451 28792 41452 28832
rect 41492 28792 41493 28832
rect 41451 28783 41493 28792
rect 41452 28337 41492 28783
rect 41836 28496 41876 28505
rect 41451 28328 41493 28337
rect 41451 28288 41452 28328
rect 41492 28288 41493 28328
rect 41451 28279 41493 28288
rect 41643 28160 41685 28169
rect 41643 28120 41644 28160
rect 41684 28120 41685 28160
rect 41643 28111 41685 28120
rect 41644 28026 41684 28111
rect 41547 27656 41589 27665
rect 41547 27616 41548 27656
rect 41588 27616 41589 27656
rect 41547 27607 41589 27616
rect 41259 26732 41301 26741
rect 41259 26692 41260 26732
rect 41300 26692 41301 26732
rect 41259 26683 41301 26692
rect 40203 26648 40245 26657
rect 40203 26608 40204 26648
rect 40244 26608 40245 26648
rect 40203 26599 40245 26608
rect 40395 26648 40437 26657
rect 40395 26608 40396 26648
rect 40436 26608 40437 26648
rect 40395 26599 40437 26608
rect 40588 26153 40628 26238
rect 40492 26144 40532 26153
rect 40300 25976 40340 25987
rect 40300 25901 40340 25936
rect 40299 25892 40341 25901
rect 40299 25852 40300 25892
rect 40340 25852 40341 25892
rect 40299 25843 40341 25852
rect 40299 25304 40341 25313
rect 40299 25264 40300 25304
rect 40340 25264 40341 25304
rect 40299 25255 40341 25264
rect 40300 25170 40340 25255
rect 40492 24809 40532 26104
rect 40587 26144 40629 26153
rect 40587 26104 40588 26144
rect 40628 26104 40629 26144
rect 40587 26095 40629 26104
rect 40780 26144 40820 26153
rect 41164 26144 41204 26153
rect 40820 26104 41164 26144
rect 40780 26095 40820 26104
rect 41164 26095 41204 26104
rect 41260 26144 41300 26683
rect 41451 26228 41493 26237
rect 41451 26188 41452 26228
rect 41492 26188 41493 26228
rect 41451 26179 41493 26188
rect 41260 25976 41300 26104
rect 41355 26144 41397 26153
rect 41355 26104 41356 26144
rect 41396 26104 41397 26144
rect 41355 26095 41397 26104
rect 41452 26144 41492 26179
rect 41356 26010 41396 26095
rect 41164 25936 41300 25976
rect 40683 25892 40725 25901
rect 40683 25852 40684 25892
rect 40724 25852 40725 25892
rect 40683 25843 40725 25852
rect 40780 25892 40820 25901
rect 40587 25472 40629 25481
rect 40587 25432 40588 25472
rect 40628 25432 40629 25472
rect 40587 25423 40629 25432
rect 40588 25229 40628 25423
rect 40684 25304 40724 25843
rect 40780 25313 40820 25852
rect 40684 25255 40724 25264
rect 40779 25304 40821 25313
rect 40779 25264 40780 25304
rect 40820 25264 40821 25304
rect 40779 25255 40821 25264
rect 40587 25220 40629 25229
rect 40587 25180 40588 25220
rect 40628 25180 40629 25220
rect 40587 25171 40629 25180
rect 40107 24800 40149 24809
rect 40107 24760 40108 24800
rect 40148 24760 40149 24800
rect 40107 24751 40149 24760
rect 40491 24800 40533 24809
rect 40491 24760 40492 24800
rect 40532 24760 40533 24800
rect 40491 24751 40533 24760
rect 40108 24632 40148 24751
rect 40011 24548 40053 24557
rect 40011 24508 40012 24548
rect 40052 24508 40053 24548
rect 40011 24499 40053 24508
rect 40012 24414 40052 24499
rect 39531 24380 39573 24389
rect 39531 24340 39532 24380
rect 39572 24340 39573 24380
rect 39531 24331 39573 24340
rect 39723 24380 39765 24389
rect 39723 24340 39724 24380
rect 39764 24340 39765 24380
rect 39723 24331 39765 24340
rect 39244 23792 39284 23801
rect 39244 23465 39284 23752
rect 39243 23456 39285 23465
rect 39243 23416 39244 23456
rect 39284 23416 39285 23456
rect 39243 23407 39285 23416
rect 39532 23288 39572 24331
rect 40012 24044 40052 24053
rect 40108 24044 40148 24592
rect 40492 24632 40532 24641
rect 40492 24389 40532 24592
rect 40588 24632 40628 25171
rect 40971 24884 41013 24893
rect 40971 24844 40972 24884
rect 41012 24844 41013 24884
rect 40971 24835 41013 24844
rect 40588 24583 40628 24592
rect 40779 24632 40821 24641
rect 40779 24592 40780 24632
rect 40820 24592 40821 24632
rect 40779 24583 40821 24592
rect 40972 24632 41012 24835
rect 41067 24716 41109 24725
rect 41067 24676 41068 24716
rect 41108 24676 41109 24716
rect 41067 24667 41109 24676
rect 40491 24380 40533 24389
rect 40491 24340 40492 24380
rect 40532 24340 40533 24380
rect 40491 24331 40533 24340
rect 40052 24004 40148 24044
rect 40780 24044 40820 24583
rect 40972 24473 41012 24592
rect 41068 24632 41108 24667
rect 41068 24581 41108 24592
rect 41164 24632 41204 25936
rect 41452 24893 41492 26104
rect 41548 25304 41588 27607
rect 41643 26396 41685 26405
rect 41643 26356 41644 26396
rect 41684 26356 41685 26396
rect 41643 26347 41685 26356
rect 41644 25976 41684 26347
rect 41836 26321 41876 28456
rect 42124 28328 42164 29035
rect 42124 28279 42164 28288
rect 42220 28328 42260 29707
rect 42316 29261 42356 29800
rect 42604 29840 42644 29849
rect 42604 29681 42644 29800
rect 42700 29840 42740 29851
rect 42700 29765 42740 29800
rect 42796 29840 42836 29849
rect 42699 29756 42741 29765
rect 42699 29716 42700 29756
rect 42740 29716 42741 29756
rect 42699 29707 42741 29716
rect 42508 29672 42548 29681
rect 42315 29252 42357 29261
rect 42315 29212 42316 29252
rect 42356 29212 42357 29252
rect 42315 29203 42357 29212
rect 42508 29009 42548 29632
rect 42603 29672 42645 29681
rect 42603 29632 42604 29672
rect 42644 29632 42645 29672
rect 42603 29623 42645 29632
rect 42796 29252 42836 29800
rect 42700 29212 42836 29252
rect 42507 29000 42549 29009
rect 42507 28960 42508 29000
rect 42548 28960 42549 29000
rect 42507 28951 42549 28960
rect 42700 28841 42740 29212
rect 42795 29084 42837 29093
rect 42795 29044 42796 29084
rect 42836 29044 42837 29084
rect 42795 29035 42837 29044
rect 42796 29000 42836 29035
rect 42796 28920 42836 28960
rect 42699 28832 42741 28841
rect 42699 28792 42700 28832
rect 42740 28792 42741 28832
rect 42699 28783 42741 28792
rect 42220 28279 42260 28288
rect 42508 28328 42548 28339
rect 42508 28253 42548 28288
rect 42892 28328 42932 31144
rect 43180 31135 43220 31144
rect 43276 29849 43316 31312
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 44812 30680 44852 30689
rect 44428 30512 44468 30521
rect 43371 30428 43413 30437
rect 43852 30428 43892 30437
rect 43371 30388 43372 30428
rect 43412 30388 43413 30428
rect 43371 30379 43413 30388
rect 43756 30388 43852 30428
rect 43180 29840 43220 29849
rect 43084 29168 43124 29179
rect 43084 29093 43124 29128
rect 43083 29084 43125 29093
rect 43083 29044 43084 29084
rect 43124 29044 43125 29084
rect 43083 29035 43125 29044
rect 42987 28832 43029 28841
rect 42987 28792 42988 28832
rect 43028 28792 43029 28832
rect 42987 28783 43029 28792
rect 42988 28421 43028 28783
rect 43180 28580 43220 29800
rect 43275 29840 43317 29849
rect 43275 29800 43276 29840
rect 43316 29800 43317 29840
rect 43275 29791 43317 29800
rect 43276 29345 43316 29791
rect 43275 29336 43317 29345
rect 43275 29296 43276 29336
rect 43316 29296 43317 29336
rect 43275 29287 43317 29296
rect 43180 28531 43220 28540
rect 42987 28412 43029 28421
rect 42987 28372 42988 28412
rect 43028 28372 43029 28412
rect 42987 28363 43029 28372
rect 42892 28279 42932 28288
rect 42988 28328 43028 28363
rect 42988 28278 43028 28288
rect 43179 28328 43221 28337
rect 43179 28288 43180 28328
rect 43220 28288 43221 28328
rect 43179 28279 43221 28288
rect 43372 28328 43412 30379
rect 43756 30185 43796 30388
rect 43852 30379 43892 30388
rect 43755 30176 43797 30185
rect 43755 30136 43756 30176
rect 43796 30136 43797 30176
rect 43755 30127 43797 30136
rect 43756 29765 43796 30127
rect 44428 29840 44468 30472
rect 44812 30185 44852 30640
rect 45484 30680 45524 30689
rect 45676 30680 45716 30689
rect 45524 30640 45676 30680
rect 45484 30631 45524 30640
rect 45676 30631 45716 30640
rect 45771 30428 45813 30437
rect 45771 30388 45772 30428
rect 45812 30388 45813 30428
rect 45771 30379 45813 30388
rect 45772 30294 45812 30379
rect 45291 30260 45333 30269
rect 45291 30220 45292 30260
rect 45332 30220 45333 30260
rect 45291 30211 45333 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 44811 30176 44853 30185
rect 44811 30136 44812 30176
rect 44852 30136 44853 30176
rect 44811 30127 44853 30136
rect 44428 29791 44468 29800
rect 45292 29840 45332 30211
rect 46251 30008 46293 30017
rect 46251 29968 46252 30008
rect 46292 29968 46293 30008
rect 46251 29959 46293 29968
rect 46635 30008 46677 30017
rect 46635 29968 46636 30008
rect 46676 29968 46677 30008
rect 46635 29959 46677 29968
rect 43755 29756 43797 29765
rect 43755 29716 43756 29756
rect 43796 29716 43797 29756
rect 43755 29707 43797 29716
rect 43852 29756 43892 29765
rect 44044 29756 44084 29765
rect 43892 29716 44044 29756
rect 43852 29707 43892 29716
rect 44044 29707 44084 29716
rect 43756 29345 43796 29430
rect 43755 29336 43797 29345
rect 43755 29296 43756 29336
rect 43796 29296 43797 29336
rect 43755 29287 43797 29296
rect 44235 29336 44277 29345
rect 44235 29296 44236 29336
rect 44276 29296 44277 29336
rect 44235 29287 44277 29296
rect 44044 29168 44084 29177
rect 43660 29128 44044 29168
rect 43467 28412 43509 28421
rect 43467 28372 43468 28412
rect 43508 28372 43509 28412
rect 43467 28363 43509 28372
rect 43372 28279 43412 28288
rect 43468 28328 43508 28363
rect 42315 28244 42357 28253
rect 42315 28204 42316 28244
rect 42356 28204 42357 28244
rect 42315 28195 42357 28204
rect 42507 28244 42549 28253
rect 42507 28204 42508 28244
rect 42548 28204 42549 28244
rect 42507 28195 42549 28204
rect 42123 28160 42165 28169
rect 42123 28120 42124 28160
rect 42164 28120 42165 28160
rect 42123 28111 42165 28120
rect 42124 27656 42164 28111
rect 42219 27740 42261 27749
rect 42219 27700 42220 27740
rect 42260 27700 42261 27740
rect 42219 27691 42261 27700
rect 42124 27607 42164 27616
rect 42220 27606 42260 27691
rect 41931 27488 41973 27497
rect 41931 27448 41932 27488
rect 41972 27448 41973 27488
rect 41931 27439 41973 27448
rect 41932 27354 41972 27439
rect 42027 26816 42069 26825
rect 42027 26776 42028 26816
rect 42068 26776 42069 26816
rect 42027 26767 42069 26776
rect 42028 26682 42068 26767
rect 41835 26312 41877 26321
rect 41835 26272 41836 26312
rect 41876 26272 41877 26312
rect 41835 26263 41877 26272
rect 41931 26228 41973 26237
rect 41931 26188 41932 26228
rect 41972 26188 41973 26228
rect 41931 26179 41973 26188
rect 41644 25927 41684 25936
rect 41451 24884 41493 24893
rect 41451 24844 41452 24884
rect 41492 24844 41493 24884
rect 41451 24835 41493 24844
rect 41548 24809 41588 25264
rect 41643 25304 41685 25313
rect 41643 25264 41644 25304
rect 41684 25264 41685 25304
rect 41643 25255 41685 25264
rect 41547 24800 41589 24809
rect 41547 24760 41548 24800
rect 41588 24760 41589 24800
rect 41547 24751 41589 24760
rect 41644 24800 41684 25255
rect 41644 24751 41684 24760
rect 41932 24800 41972 26179
rect 42028 26144 42068 26153
rect 42028 25817 42068 26104
rect 42316 26144 42356 28195
rect 43180 28194 43220 28279
rect 43468 28277 43508 28288
rect 43660 28328 43700 29128
rect 44044 29119 44084 29128
rect 44140 29168 44180 29177
rect 44140 29000 44180 29128
rect 44236 29168 44276 29287
rect 45292 29177 45332 29800
rect 44236 29119 44276 29128
rect 44332 29168 44372 29177
rect 43948 28960 44180 29000
rect 43755 28496 43797 28505
rect 43755 28456 43756 28496
rect 43796 28456 43797 28496
rect 43755 28447 43797 28456
rect 43660 28279 43700 28288
rect 43563 28244 43605 28253
rect 43563 28204 43564 28244
rect 43604 28204 43605 28244
rect 43563 28195 43605 28204
rect 43564 28110 43604 28195
rect 43756 27656 43796 28447
rect 43851 28328 43893 28337
rect 43851 28288 43852 28328
rect 43892 28288 43893 28328
rect 43851 28279 43893 28288
rect 43948 28328 43988 28960
rect 44140 28421 44180 28468
rect 44332 28421 44372 29128
rect 45291 29168 45333 29177
rect 45291 29128 45292 29168
rect 45332 29128 45333 29168
rect 45291 29119 45333 29128
rect 45484 29168 45524 29177
rect 45196 29000 45236 29009
rect 45292 29000 45332 29119
rect 45484 29000 45524 29128
rect 45868 29168 45908 29177
rect 45236 28960 45428 29000
rect 45484 28960 45812 29000
rect 45196 28951 45236 28960
rect 45195 28496 45237 28505
rect 45195 28456 45196 28496
rect 45236 28456 45237 28496
rect 45195 28447 45237 28456
rect 44139 28412 44181 28421
rect 44139 28363 44140 28412
rect 43852 28194 43892 28279
rect 43948 27824 43988 28288
rect 44043 28328 44085 28337
rect 44043 28288 44044 28328
rect 44084 28288 44085 28328
rect 44180 28363 44181 28412
rect 44331 28412 44373 28421
rect 44331 28372 44332 28412
rect 44372 28372 44373 28412
rect 44331 28363 44373 28372
rect 44140 28324 44180 28333
rect 44332 28328 44372 28363
rect 44043 28279 44085 28288
rect 44044 28194 44084 28279
rect 44332 28277 44372 28288
rect 45196 28328 45236 28447
rect 45196 28279 45236 28288
rect 45099 27824 45141 27833
rect 43948 27784 44276 27824
rect 43756 27607 43796 27616
rect 44140 27656 44180 27665
rect 43564 27404 43604 27413
rect 43564 27161 43604 27364
rect 43563 27152 43605 27161
rect 43563 27112 43564 27152
rect 43604 27112 43605 27152
rect 43563 27103 43605 27112
rect 44140 27077 44180 27616
rect 42987 27068 43029 27077
rect 42987 27028 42988 27068
rect 43028 27028 43029 27068
rect 42987 27019 43029 27028
rect 44139 27068 44181 27077
rect 44139 27028 44140 27068
rect 44180 27028 44181 27068
rect 44139 27019 44181 27028
rect 42795 26984 42837 26993
rect 42795 26944 42796 26984
rect 42836 26944 42837 26984
rect 42795 26935 42837 26944
rect 42700 26816 42740 26825
rect 42700 26312 42740 26776
rect 42796 26816 42836 26935
rect 42988 26934 43028 27019
rect 43467 26984 43509 26993
rect 43467 26944 43468 26984
rect 43508 26944 43509 26984
rect 43467 26935 43509 26944
rect 43755 26984 43797 26993
rect 43755 26944 43756 26984
rect 43796 26944 43797 26984
rect 43755 26935 43797 26944
rect 43371 26900 43413 26909
rect 43371 26860 43372 26900
rect 43412 26860 43413 26900
rect 43371 26851 43413 26860
rect 42796 26767 42836 26776
rect 42988 26816 43028 26825
rect 43180 26816 43220 26825
rect 43028 26776 43180 26816
rect 42988 26767 43028 26776
rect 43180 26767 43220 26776
rect 43276 26816 43316 26827
rect 43276 26741 43316 26776
rect 43372 26816 43412 26851
rect 43372 26765 43412 26776
rect 43468 26816 43508 26935
rect 43468 26767 43508 26776
rect 43660 26816 43700 26825
rect 43275 26732 43317 26741
rect 43275 26692 43276 26732
rect 43316 26692 43317 26732
rect 43275 26683 43317 26692
rect 42796 26312 42836 26321
rect 42700 26272 42796 26312
rect 42796 26263 42836 26272
rect 42316 26069 42356 26104
rect 42891 26144 42933 26153
rect 42891 26104 42892 26144
rect 42932 26104 42933 26144
rect 42891 26095 42933 26104
rect 43083 26144 43125 26153
rect 43083 26104 43084 26144
rect 43124 26104 43125 26144
rect 43083 26095 43125 26104
rect 42315 26060 42357 26069
rect 42315 26020 42316 26060
rect 42356 26020 42357 26060
rect 42315 26011 42357 26020
rect 42316 25980 42356 26011
rect 42892 26010 42932 26095
rect 43084 26010 43124 26095
rect 42027 25808 42069 25817
rect 42027 25768 42028 25808
rect 42068 25768 42069 25808
rect 42027 25759 42069 25768
rect 42699 25808 42741 25817
rect 42699 25768 42700 25808
rect 42740 25768 42741 25808
rect 42699 25759 42741 25768
rect 42700 25556 42740 25759
rect 43660 25556 43700 26776
rect 43756 26816 43796 26935
rect 43756 26767 43796 26776
rect 43948 26816 43988 26825
rect 43851 26648 43893 26657
rect 43851 26608 43852 26648
rect 43892 26608 43893 26648
rect 43851 26599 43893 26608
rect 43852 26514 43892 26599
rect 43948 26489 43988 26776
rect 44236 26741 44276 27784
rect 45099 27784 45100 27824
rect 45140 27784 45141 27824
rect 45099 27775 45141 27784
rect 44524 27656 44564 27665
rect 44564 27616 44948 27656
rect 44524 27607 44564 27616
rect 44620 27112 44852 27152
rect 44235 26732 44277 26741
rect 44235 26692 44236 26732
rect 44276 26692 44277 26732
rect 44235 26683 44277 26692
rect 44427 26732 44469 26741
rect 44427 26692 44428 26732
rect 44468 26692 44469 26732
rect 44427 26683 44469 26692
rect 44140 26648 44180 26657
rect 44044 26608 44140 26648
rect 43947 26480 43989 26489
rect 43947 26440 43948 26480
rect 43988 26440 43989 26480
rect 43947 26431 43989 26440
rect 43756 26144 43796 26153
rect 43756 25817 43796 26104
rect 43947 25976 43989 25985
rect 43947 25936 43948 25976
rect 43988 25936 43989 25976
rect 43947 25927 43989 25936
rect 43948 25842 43988 25927
rect 43755 25808 43797 25817
rect 43755 25768 43756 25808
rect 43796 25768 43797 25808
rect 43755 25759 43797 25768
rect 43756 25556 43796 25565
rect 43660 25516 43756 25556
rect 42700 25507 42740 25516
rect 43756 25507 43796 25516
rect 43371 25388 43413 25397
rect 43371 25348 43372 25388
rect 43412 25348 43413 25388
rect 43371 25339 43413 25348
rect 42891 25304 42933 25313
rect 42891 25264 42892 25304
rect 42932 25264 42933 25304
rect 42891 25255 42933 25264
rect 42892 25170 42932 25255
rect 41164 24583 41204 24592
rect 41259 24632 41301 24641
rect 41259 24592 41260 24632
rect 41300 24592 41301 24632
rect 41259 24583 41301 24592
rect 41452 24632 41492 24643
rect 41740 24641 41780 24726
rect 41932 24725 41972 24760
rect 43083 24800 43125 24809
rect 43083 24760 43084 24800
rect 43124 24760 43125 24800
rect 43083 24751 43125 24760
rect 41931 24716 41973 24725
rect 41931 24676 41932 24716
rect 41972 24676 41973 24716
rect 41931 24667 41973 24676
rect 41260 24498 41300 24583
rect 41452 24557 41492 24592
rect 41548 24632 41588 24641
rect 41451 24548 41493 24557
rect 41451 24508 41452 24548
rect 41492 24508 41493 24548
rect 41451 24499 41493 24508
rect 41548 24473 41588 24592
rect 41739 24632 41781 24641
rect 41932 24636 41972 24667
rect 41739 24592 41740 24632
rect 41780 24592 41781 24632
rect 41739 24583 41781 24592
rect 43084 24632 43124 24751
rect 40971 24464 41013 24473
rect 40971 24424 40972 24464
rect 41012 24424 41013 24464
rect 40971 24415 41013 24424
rect 41547 24464 41589 24473
rect 41547 24424 41548 24464
rect 41588 24424 41589 24464
rect 41547 24415 41589 24424
rect 41931 24464 41973 24473
rect 41931 24424 41932 24464
rect 41972 24424 41973 24464
rect 41931 24415 41973 24424
rect 41259 24380 41301 24389
rect 41259 24340 41260 24380
rect 41300 24340 41301 24380
rect 41259 24331 41301 24340
rect 40012 23995 40052 24004
rect 40780 23995 40820 24004
rect 40492 23960 40532 23969
rect 40532 23920 40628 23960
rect 40492 23911 40532 23920
rect 40107 23792 40149 23801
rect 40107 23752 40108 23792
rect 40148 23752 40149 23792
rect 40107 23743 40149 23752
rect 40108 23658 40148 23743
rect 38956 23071 38996 23080
rect 39052 23248 39380 23288
rect 39052 23120 39092 23248
rect 39052 23071 39092 23080
rect 39148 23120 39188 23129
rect 38763 22364 38805 22373
rect 38763 22324 38764 22364
rect 38804 22324 38805 22364
rect 38763 22315 38805 22324
rect 38571 22280 38613 22289
rect 38571 22240 38572 22280
rect 38612 22240 38613 22280
rect 38571 22231 38613 22240
rect 38572 22146 38612 22231
rect 38667 21860 38709 21869
rect 38667 21820 38668 21860
rect 38708 21820 38709 21860
rect 38667 21811 38709 21820
rect 38379 21692 38421 21701
rect 38379 21652 38380 21692
rect 38420 21652 38421 21692
rect 38379 21643 38421 21652
rect 38380 21558 38420 21643
rect 38475 21524 38517 21533
rect 38475 21484 38476 21524
rect 38516 21484 38517 21524
rect 38475 21475 38517 21484
rect 38283 21104 38325 21113
rect 38283 21064 38284 21104
rect 38324 21064 38420 21104
rect 38283 21055 38325 21064
rect 37900 20896 38324 20936
rect 37995 20768 38037 20777
rect 37995 20728 37996 20768
rect 38036 20728 38037 20768
rect 37995 20719 38037 20728
rect 37996 20600 38036 20719
rect 37996 20551 38036 20560
rect 38187 20600 38229 20609
rect 38187 20560 38188 20600
rect 38228 20560 38229 20600
rect 38187 20551 38229 20560
rect 38188 20466 38228 20551
rect 37995 20348 38037 20357
rect 37995 20308 37996 20348
rect 38036 20308 38037 20348
rect 37995 20299 38037 20308
rect 37804 20131 37844 20140
rect 37419 20096 37461 20105
rect 37419 20056 37420 20096
rect 37460 20056 37461 20096
rect 37419 20047 37461 20056
rect 37516 20096 37556 20105
rect 36884 19216 36980 19256
rect 36844 18593 36884 19216
rect 37516 18752 37556 20056
rect 37900 20096 37940 20107
rect 37900 20021 37940 20056
rect 37996 20096 38036 20299
rect 37996 20047 38036 20056
rect 38091 20096 38133 20105
rect 38091 20056 38092 20096
rect 38132 20056 38133 20096
rect 38091 20047 38133 20056
rect 38284 20096 38324 20896
rect 38380 20782 38420 21064
rect 38380 20733 38420 20742
rect 38380 20189 38420 20274
rect 38379 20180 38421 20189
rect 38379 20140 38380 20180
rect 38420 20140 38421 20180
rect 38379 20131 38421 20140
rect 38284 20047 38324 20056
rect 38476 20096 38516 21475
rect 37899 20012 37941 20021
rect 37899 19972 37900 20012
rect 37940 19972 37941 20012
rect 37899 19963 37941 19972
rect 38092 19962 38132 20047
rect 38476 19853 38516 20056
rect 38571 20096 38613 20105
rect 38571 20056 38572 20096
rect 38612 20056 38613 20096
rect 38571 20047 38613 20056
rect 38572 19962 38612 20047
rect 38475 19844 38517 19853
rect 38475 19804 38476 19844
rect 38516 19804 38517 19844
rect 38475 19795 38517 19804
rect 37900 19636 38228 19676
rect 37804 19256 37844 19265
rect 37804 18845 37844 19216
rect 37803 18836 37845 18845
rect 37803 18796 37804 18836
rect 37844 18796 37845 18836
rect 37803 18787 37845 18796
rect 37036 18712 37556 18752
rect 36843 18584 36885 18593
rect 36843 18544 36844 18584
rect 36884 18544 36885 18584
rect 36843 18535 36885 18544
rect 37036 18584 37076 18712
rect 37900 18668 37940 19636
rect 37995 19508 38037 19517
rect 37995 19468 37996 19508
rect 38036 19468 38037 19508
rect 37995 19459 38037 19468
rect 38188 19508 38228 19636
rect 38188 19459 38228 19468
rect 37900 18619 37940 18628
rect 36843 18416 36885 18425
rect 36843 18376 36844 18416
rect 36884 18376 36885 18416
rect 36843 18367 36885 18376
rect 36844 17744 36884 18367
rect 36844 17695 36884 17704
rect 37036 17156 37076 18544
rect 37419 18584 37461 18593
rect 37419 18544 37420 18584
rect 37460 18544 37461 18584
rect 37419 18535 37461 18544
rect 37420 18500 37460 18535
rect 37420 18449 37460 18460
rect 37996 18416 38036 19459
rect 38668 19433 38708 21811
rect 38764 20357 38804 22315
rect 39148 22280 39188 23080
rect 39052 22240 39188 22280
rect 39244 23120 39284 23129
rect 39340 23120 39380 23248
rect 39532 23239 39572 23248
rect 39436 23120 39476 23129
rect 39724 23120 39764 23129
rect 39340 23080 39436 23120
rect 39476 23080 39724 23120
rect 39052 21869 39092 22240
rect 39147 22112 39189 22121
rect 39147 22072 39148 22112
rect 39188 22072 39189 22112
rect 39147 22063 39189 22072
rect 39051 21860 39093 21869
rect 39051 21820 39052 21860
rect 39092 21820 39093 21860
rect 39051 21811 39093 21820
rect 39052 21608 39092 21617
rect 39052 20777 39092 21568
rect 38860 20768 38900 20777
rect 38860 20609 38900 20728
rect 39051 20768 39093 20777
rect 39051 20728 39052 20768
rect 39092 20728 39093 20768
rect 39051 20719 39093 20728
rect 38859 20600 38901 20609
rect 38859 20560 38860 20600
rect 38900 20560 38901 20600
rect 38859 20551 38901 20560
rect 38763 20348 38805 20357
rect 38763 20308 38764 20348
rect 38804 20308 38805 20348
rect 38763 20299 38805 20308
rect 38764 20096 38804 20299
rect 38764 20047 38804 20056
rect 38956 20096 38996 20105
rect 38859 20012 38901 20021
rect 38859 19972 38860 20012
rect 38900 19972 38901 20012
rect 38859 19963 38901 19972
rect 38860 19878 38900 19963
rect 38956 19517 38996 20056
rect 39148 20012 39188 22063
rect 39244 21608 39284 23080
rect 39436 23071 39476 23080
rect 39724 23071 39764 23080
rect 40396 23120 40436 23129
rect 40396 22709 40436 23080
rect 40491 23120 40533 23129
rect 40491 23080 40492 23120
rect 40532 23080 40533 23120
rect 40491 23071 40533 23080
rect 39723 22700 39765 22709
rect 39723 22660 39724 22700
rect 39764 22660 39765 22700
rect 39723 22651 39765 22660
rect 40395 22700 40437 22709
rect 40395 22660 40396 22700
rect 40436 22660 40437 22700
rect 40395 22651 40437 22660
rect 39724 22532 39764 22651
rect 39724 22483 39764 22492
rect 39915 22364 39957 22373
rect 39915 22324 39916 22364
rect 39956 22324 39957 22364
rect 39915 22315 39957 22324
rect 40396 22364 40436 22373
rect 40492 22364 40532 23071
rect 40588 23036 40628 23920
rect 40876 23792 40916 23803
rect 40876 23717 40916 23752
rect 40875 23708 40917 23717
rect 40875 23668 40876 23708
rect 40916 23668 40917 23708
rect 40875 23659 40917 23668
rect 41068 23624 41108 23633
rect 40972 23584 41068 23624
rect 40684 23204 40724 23213
rect 40972 23204 41012 23584
rect 41068 23575 41108 23584
rect 40724 23164 41012 23204
rect 40684 23155 40724 23164
rect 41068 23120 41108 23129
rect 41068 23036 41108 23080
rect 40588 22996 41108 23036
rect 41067 22448 41109 22457
rect 41067 22408 41068 22448
rect 41108 22408 41109 22448
rect 41067 22399 41109 22408
rect 40436 22324 40532 22364
rect 40779 22364 40821 22373
rect 40779 22324 40780 22364
rect 40820 22324 40821 22364
rect 40396 22315 40436 22324
rect 40779 22315 40821 22324
rect 39339 21776 39381 21785
rect 39339 21736 39340 21776
rect 39380 21736 39381 21776
rect 39339 21727 39381 21736
rect 39340 21642 39380 21727
rect 39244 21559 39284 21568
rect 39435 21608 39477 21617
rect 39435 21568 39436 21608
rect 39476 21568 39477 21608
rect 39435 21559 39477 21568
rect 39532 21608 39572 21617
rect 39436 21474 39476 21559
rect 39339 21020 39381 21029
rect 39339 20980 39340 21020
rect 39380 20980 39381 21020
rect 39339 20971 39381 20980
rect 39340 20852 39380 20971
rect 39340 20803 39380 20812
rect 39435 20768 39477 20777
rect 39435 20728 39436 20768
rect 39476 20728 39477 20768
rect 39435 20719 39477 20728
rect 39436 20634 39476 20719
rect 39532 20264 39572 21568
rect 39819 20852 39861 20861
rect 39819 20812 39820 20852
rect 39860 20812 39861 20852
rect 39819 20803 39861 20812
rect 39820 20768 39860 20803
rect 39820 20717 39860 20728
rect 39916 20768 39956 22315
rect 40204 22280 40244 22289
rect 40107 22196 40149 22205
rect 40107 22156 40108 22196
rect 40148 22156 40149 22196
rect 40107 22147 40149 22156
rect 40108 22062 40148 22147
rect 40204 21617 40244 22240
rect 40780 22280 40820 22315
rect 40780 22229 40820 22240
rect 40875 22280 40917 22289
rect 40875 22240 40876 22280
rect 40916 22240 40917 22280
rect 40875 22231 40917 22240
rect 40972 22280 41012 22289
rect 40876 22146 40916 22231
rect 40972 21869 41012 22240
rect 40971 21860 41013 21869
rect 40971 21820 40972 21860
rect 41012 21820 41013 21860
rect 40971 21811 41013 21820
rect 40491 21776 40533 21785
rect 40491 21736 40492 21776
rect 40532 21736 40533 21776
rect 40491 21727 40533 21736
rect 40299 21692 40341 21701
rect 40299 21652 40300 21692
rect 40340 21652 40341 21692
rect 40299 21643 40341 21652
rect 40203 21608 40245 21617
rect 40203 21568 40204 21608
rect 40244 21568 40245 21608
rect 40203 21559 40245 21568
rect 40300 21608 40340 21643
rect 40107 21440 40149 21449
rect 40107 21400 40108 21440
rect 40148 21400 40149 21440
rect 40107 21391 40149 21400
rect 40108 21306 40148 21391
rect 39916 20719 39956 20728
rect 39244 20224 39572 20264
rect 39244 20180 39284 20224
rect 39244 20131 39284 20140
rect 39340 20096 39380 20105
rect 39340 20012 39380 20056
rect 39148 19972 39380 20012
rect 39628 20096 39668 20105
rect 40300 20096 40340 21568
rect 40395 21608 40437 21617
rect 40395 21568 40396 21608
rect 40436 21568 40437 21608
rect 40395 21559 40437 21568
rect 40492 21608 40532 21727
rect 40971 21692 41013 21701
rect 40971 21652 40972 21692
rect 41012 21652 41013 21692
rect 40971 21643 41013 21652
rect 40492 21559 40532 21568
rect 40588 21608 40628 21617
rect 40780 21608 40820 21617
rect 40628 21568 40780 21608
rect 40588 21559 40628 21568
rect 40780 21559 40820 21568
rect 40972 21608 41012 21643
rect 40396 21474 40436 21559
rect 40972 21557 41012 21568
rect 41068 21608 41108 22399
rect 41164 22280 41204 22291
rect 41164 22205 41204 22240
rect 41260 22280 41300 24331
rect 41355 23792 41397 23801
rect 41740 23792 41780 23801
rect 41355 23752 41356 23792
rect 41396 23752 41397 23792
rect 41355 23743 41397 23752
rect 41452 23752 41740 23792
rect 41260 22231 41300 22240
rect 41163 22196 41205 22205
rect 41163 22156 41164 22196
rect 41204 22156 41205 22196
rect 41163 22147 41205 22156
rect 41163 21860 41205 21869
rect 41163 21820 41164 21860
rect 41204 21820 41205 21860
rect 41163 21811 41205 21820
rect 41068 21559 41108 21568
rect 40875 21440 40917 21449
rect 40875 21400 40876 21440
rect 40916 21400 40917 21440
rect 40875 21391 40917 21400
rect 40780 21356 40820 21365
rect 40492 21316 40780 21356
rect 40492 20768 40532 21316
rect 40780 21307 40820 21316
rect 40492 20719 40532 20728
rect 40876 20768 40916 21391
rect 41164 21197 41204 21811
rect 41260 21776 41300 21785
rect 41356 21776 41396 23743
rect 41452 22532 41492 23752
rect 41740 23743 41780 23752
rect 41932 23792 41972 24415
rect 41932 23743 41972 23752
rect 42027 23792 42069 23801
rect 42027 23752 42028 23792
rect 42068 23752 42069 23792
rect 42027 23743 42069 23752
rect 42124 23792 42164 23801
rect 42028 23658 42068 23743
rect 41547 23624 41589 23633
rect 41547 23584 41548 23624
rect 41588 23584 41589 23624
rect 41547 23575 41589 23584
rect 41452 22483 41492 22492
rect 41452 22280 41492 22289
rect 41548 22280 41588 23575
rect 41931 23120 41973 23129
rect 41931 23080 41932 23120
rect 41972 23080 41973 23120
rect 41931 23071 41973 23080
rect 41932 22986 41972 23071
rect 41643 22952 41685 22961
rect 41643 22912 41644 22952
rect 41684 22912 41685 22952
rect 41643 22903 41685 22912
rect 41492 22240 41588 22280
rect 41644 22280 41684 22903
rect 42124 22625 42164 23752
rect 42603 23708 42645 23717
rect 42603 23668 42604 23708
rect 42644 23668 42645 23708
rect 42603 23659 42645 23668
rect 42219 23624 42261 23633
rect 42219 23584 42220 23624
rect 42260 23584 42261 23624
rect 42219 23575 42261 23584
rect 42220 23490 42260 23575
rect 42604 23574 42644 23659
rect 43084 23129 43124 24592
rect 43275 23792 43317 23801
rect 43275 23752 43276 23792
rect 43316 23752 43317 23792
rect 43275 23743 43317 23752
rect 42603 23120 42645 23129
rect 42603 23080 42604 23120
rect 42644 23080 42645 23120
rect 42603 23071 42645 23080
rect 43083 23120 43125 23129
rect 43083 23080 43084 23120
rect 43124 23080 43125 23120
rect 43083 23071 43125 23080
rect 42123 22616 42165 22625
rect 42123 22576 42124 22616
rect 42164 22576 42165 22616
rect 42123 22567 42165 22576
rect 42507 22616 42549 22625
rect 42507 22576 42508 22616
rect 42548 22576 42549 22616
rect 42507 22567 42549 22576
rect 41931 22448 41973 22457
rect 41931 22408 41932 22448
rect 41972 22408 41973 22448
rect 41931 22399 41973 22408
rect 41835 22364 41877 22373
rect 41835 22324 41836 22364
rect 41876 22324 41877 22364
rect 41835 22315 41877 22324
rect 41452 22231 41492 22240
rect 41644 22231 41684 22240
rect 41739 22280 41781 22289
rect 41739 22240 41740 22280
rect 41780 22240 41781 22280
rect 41739 22231 41781 22240
rect 41836 22280 41876 22315
rect 41740 22146 41780 22231
rect 41836 22229 41876 22240
rect 41932 22280 41972 22399
rect 41932 22231 41972 22240
rect 42123 22112 42165 22121
rect 42123 22072 42124 22112
rect 42164 22072 42165 22112
rect 42123 22063 42165 22072
rect 42124 21978 42164 22063
rect 42508 21785 42548 22567
rect 42507 21776 42549 21785
rect 41300 21736 41396 21776
rect 41932 21736 42356 21776
rect 41260 21727 41300 21736
rect 41932 21608 41972 21736
rect 41932 21559 41972 21568
rect 42124 21608 42164 21617
rect 41259 21524 41301 21533
rect 41259 21484 41260 21524
rect 41300 21484 41301 21524
rect 41259 21475 41301 21484
rect 41163 21188 41205 21197
rect 41163 21148 41164 21188
rect 41204 21148 41205 21188
rect 41163 21139 41205 21148
rect 40876 20719 40916 20728
rect 41067 20768 41109 20777
rect 41067 20728 41068 20768
rect 41108 20728 41109 20768
rect 41067 20719 41109 20728
rect 40396 20096 40436 20105
rect 40300 20056 40396 20096
rect 39532 19844 39572 19853
rect 38955 19508 38997 19517
rect 38955 19468 38956 19508
rect 38996 19468 38997 19508
rect 38955 19459 38997 19468
rect 38667 19424 38709 19433
rect 38667 19384 38668 19424
rect 38708 19384 38709 19424
rect 38667 19375 38709 19384
rect 39148 19424 39188 19433
rect 38379 19340 38421 19349
rect 38379 19300 38380 19340
rect 38420 19300 38421 19340
rect 38379 19291 38421 19300
rect 38188 19256 38228 19265
rect 38188 19088 38228 19216
rect 38380 19256 38420 19291
rect 38476 19265 38516 19350
rect 38380 19205 38420 19216
rect 38475 19256 38517 19265
rect 38475 19216 38476 19256
rect 38516 19216 38517 19256
rect 38668 19256 38708 19375
rect 38956 19349 38996 19380
rect 38955 19340 38997 19349
rect 38955 19300 38956 19340
rect 38996 19300 38997 19340
rect 38955 19291 38997 19300
rect 38764 19256 38804 19265
rect 38668 19216 38764 19256
rect 38475 19207 38517 19216
rect 38764 19207 38804 19216
rect 38860 19256 38900 19267
rect 38860 19181 38900 19216
rect 38956 19256 38996 19291
rect 38859 19172 38901 19181
rect 38859 19132 38860 19172
rect 38900 19132 38901 19172
rect 38859 19123 38901 19132
rect 38668 19088 38708 19097
rect 38188 19048 38668 19088
rect 38668 19039 38708 19048
rect 38956 19013 38996 19216
rect 38955 19004 38997 19013
rect 38955 18964 38956 19004
rect 38996 18964 38997 19004
rect 38955 18955 38997 18964
rect 39148 18929 39188 19384
rect 39532 19265 39572 19804
rect 39628 19685 39668 20056
rect 40396 20047 40436 20056
rect 40684 19844 40724 19853
rect 39627 19676 39669 19685
rect 39627 19636 39628 19676
rect 39668 19636 39669 19676
rect 39627 19627 39669 19636
rect 40107 19424 40149 19433
rect 40107 19384 40108 19424
rect 40148 19384 40149 19424
rect 40107 19375 40149 19384
rect 39531 19256 39573 19265
rect 39531 19216 39532 19256
rect 39572 19216 39573 19256
rect 39531 19207 39573 19216
rect 39628 19256 39668 19267
rect 40012 19265 40052 19350
rect 39628 19181 39668 19216
rect 39916 19256 39956 19265
rect 39627 19172 39669 19181
rect 39627 19132 39628 19172
rect 39668 19132 39669 19172
rect 39627 19123 39669 19132
rect 39724 19088 39764 19097
rect 39764 19048 39860 19088
rect 39724 19039 39764 19048
rect 38283 18920 38325 18929
rect 38283 18880 38284 18920
rect 38324 18880 38325 18920
rect 38283 18871 38325 18880
rect 39147 18920 39189 18929
rect 39147 18880 39148 18920
rect 39188 18880 39189 18920
rect 39147 18871 39189 18880
rect 38284 18584 38324 18871
rect 38475 18836 38517 18845
rect 38475 18796 38476 18836
rect 38516 18796 38517 18836
rect 38475 18787 38517 18796
rect 38284 18535 38324 18544
rect 37900 18376 38036 18416
rect 37707 17744 37749 17753
rect 37707 17704 37708 17744
rect 37748 17704 37749 17744
rect 37707 17695 37749 17704
rect 37708 17610 37748 17695
rect 37324 17576 37364 17585
rect 37364 17536 37460 17576
rect 37324 17527 37364 17536
rect 36940 17116 37076 17156
rect 36844 16829 36884 16914
rect 36843 16820 36885 16829
rect 36843 16780 36844 16820
rect 36884 16780 36885 16820
rect 36843 16771 36885 16780
rect 36940 16652 36980 17116
rect 37324 17072 37364 17081
rect 37132 17032 37324 17072
rect 37035 16988 37077 16997
rect 37035 16948 37036 16988
rect 37076 16948 37077 16988
rect 37035 16939 37077 16948
rect 37036 16854 37076 16939
rect 36844 16612 36980 16652
rect 36844 15233 36884 16612
rect 36940 16484 36980 16493
rect 37132 16484 37172 17032
rect 37324 17023 37364 17032
rect 36980 16444 37172 16484
rect 36940 16435 36980 16444
rect 37420 16400 37460 17536
rect 37036 16360 37460 16400
rect 37708 17072 37748 17081
rect 37708 16400 37748 17032
rect 37804 16400 37844 16409
rect 37708 16360 37804 16400
rect 36940 16232 36980 16241
rect 37036 16232 37076 16360
rect 37804 16351 37844 16360
rect 36940 16073 36980 16192
rect 37035 16211 37076 16232
rect 37324 16232 37364 16241
rect 37132 16211 37172 16220
rect 37035 16171 37132 16211
rect 36939 16064 36981 16073
rect 36939 16024 36940 16064
rect 36980 16024 36981 16064
rect 36939 16015 36981 16024
rect 36939 15476 36981 15485
rect 36939 15436 36940 15476
rect 36980 15436 36981 15476
rect 36939 15427 36981 15436
rect 36843 15224 36885 15233
rect 36843 15184 36844 15224
rect 36884 15184 36885 15224
rect 36843 15175 36885 15184
rect 36747 15140 36789 15149
rect 36747 15100 36748 15140
rect 36788 15100 36789 15140
rect 36747 15091 36789 15100
rect 36940 14897 36980 15427
rect 36939 14888 36981 14897
rect 36939 14848 36940 14888
rect 36980 14848 36981 14888
rect 36939 14839 36981 14848
rect 36556 14048 36596 14057
rect 36556 13889 36596 14008
rect 36651 14048 36693 14057
rect 36651 14008 36652 14048
rect 36692 14008 36693 14048
rect 36651 13999 36693 14008
rect 36843 14048 36885 14057
rect 36843 14008 36844 14048
rect 36884 14008 36885 14048
rect 36843 13999 36885 14008
rect 36940 14048 36980 14839
rect 36652 13914 36692 13999
rect 36844 13914 36884 13999
rect 36555 13880 36597 13889
rect 36555 13840 36556 13880
rect 36596 13840 36597 13880
rect 36555 13831 36597 13840
rect 36651 13796 36693 13805
rect 36651 13756 36652 13796
rect 36692 13756 36693 13796
rect 36651 13747 36693 13756
rect 36460 13420 36596 13460
rect 36460 13217 36500 13302
rect 36459 13208 36501 13217
rect 36459 13168 36460 13208
rect 36500 13168 36501 13208
rect 36459 13159 36501 13168
rect 36363 13124 36405 13133
rect 36363 13084 36364 13124
rect 36404 13084 36405 13124
rect 36363 13075 36405 13084
rect 36364 12990 36404 13075
rect 36556 13040 36596 13420
rect 36460 13000 36596 13040
rect 36268 12496 36404 12536
rect 36268 11696 36308 11705
rect 36268 11537 36308 11656
rect 36172 11528 36212 11537
rect 36172 11369 36212 11488
rect 36267 11528 36309 11537
rect 36267 11488 36268 11528
rect 36308 11488 36309 11528
rect 36267 11479 36309 11488
rect 36171 11360 36213 11369
rect 36171 11320 36172 11360
rect 36212 11320 36213 11360
rect 36171 11311 36213 11320
rect 36364 11201 36404 12496
rect 36460 11276 36500 13000
rect 36652 12125 36692 13747
rect 36940 13217 36980 14008
rect 37036 13385 37076 16171
rect 37132 16162 37172 16171
rect 37228 16211 37268 16220
rect 37364 16192 37556 16232
rect 37324 16183 37364 16192
rect 37228 16157 37268 16171
rect 37227 16148 37269 16157
rect 37227 16108 37228 16148
rect 37268 16108 37269 16148
rect 37227 16099 37269 16108
rect 37228 16076 37268 16099
rect 37419 16064 37461 16073
rect 37419 16024 37420 16064
rect 37460 16024 37461 16064
rect 37419 16015 37461 16024
rect 37420 15930 37460 16015
rect 37419 15560 37461 15569
rect 37419 15520 37420 15560
rect 37460 15520 37461 15560
rect 37419 15511 37461 15520
rect 37132 14216 37172 14225
rect 37035 13376 37077 13385
rect 37035 13336 37036 13376
rect 37076 13336 37077 13376
rect 37035 13327 37077 13336
rect 36939 13208 36981 13217
rect 36939 13168 36940 13208
rect 36980 13168 36981 13208
rect 36939 13159 36981 13168
rect 36651 12116 36693 12125
rect 36651 12076 36652 12116
rect 36692 12076 36693 12116
rect 36651 12067 36693 12076
rect 36940 12041 36980 13159
rect 37036 12536 37076 12545
rect 37132 12536 37172 14176
rect 37324 14048 37364 14057
rect 37324 13469 37364 14008
rect 37323 13460 37365 13469
rect 37323 13420 37324 13460
rect 37364 13420 37365 13460
rect 37323 13411 37365 13420
rect 37323 13208 37365 13217
rect 37323 13168 37324 13208
rect 37364 13168 37365 13208
rect 37323 13159 37365 13168
rect 37420 13208 37460 15511
rect 37516 14813 37556 16192
rect 37804 15308 37844 15317
rect 37804 14981 37844 15268
rect 37900 15140 37940 18376
rect 38188 16400 38228 16409
rect 38228 16360 38420 16400
rect 38188 16351 38228 16360
rect 37996 16232 38036 16241
rect 37996 15401 38036 16192
rect 38188 16232 38228 16241
rect 38092 15728 38132 15737
rect 38188 15728 38228 16192
rect 38380 16232 38420 16360
rect 38380 16183 38420 16192
rect 38132 15688 38228 15728
rect 38092 15679 38132 15688
rect 38188 15560 38228 15569
rect 37995 15392 38037 15401
rect 37995 15352 37996 15392
rect 38036 15352 38037 15392
rect 37995 15343 38037 15352
rect 37900 15100 38036 15140
rect 37611 14972 37653 14981
rect 37611 14932 37612 14972
rect 37652 14932 37653 14972
rect 37611 14923 37653 14932
rect 37803 14972 37845 14981
rect 37803 14932 37804 14972
rect 37844 14932 37845 14972
rect 37803 14923 37845 14932
rect 37515 14804 37557 14813
rect 37515 14764 37516 14804
rect 37556 14764 37557 14804
rect 37515 14755 37557 14764
rect 37420 13159 37460 13168
rect 37516 13208 37556 14755
rect 37612 14720 37652 14923
rect 37899 14888 37941 14897
rect 37899 14848 37900 14888
rect 37940 14848 37941 14888
rect 37899 14839 37941 14848
rect 37900 14754 37940 14839
rect 37612 14561 37652 14680
rect 37611 14552 37653 14561
rect 37611 14512 37612 14552
rect 37652 14512 37653 14552
rect 37611 14503 37653 14512
rect 37996 14141 38036 15100
rect 38188 14813 38228 15520
rect 38283 15560 38325 15569
rect 38283 15520 38284 15560
rect 38324 15520 38325 15560
rect 38283 15511 38325 15520
rect 38380 15560 38420 15569
rect 38284 15426 38324 15511
rect 38380 14897 38420 15520
rect 38379 14888 38421 14897
rect 38379 14848 38380 14888
rect 38420 14848 38421 14888
rect 38379 14839 38421 14848
rect 38187 14804 38229 14813
rect 38187 14764 38188 14804
rect 38228 14764 38229 14804
rect 38187 14755 38229 14764
rect 38283 14216 38325 14225
rect 38283 14176 38284 14216
rect 38324 14176 38325 14216
rect 38283 14167 38325 14176
rect 38380 14216 38420 14225
rect 38476 14216 38516 18787
rect 39147 18584 39189 18593
rect 39147 18544 39148 18584
rect 39188 18544 39189 18584
rect 39147 18535 39189 18544
rect 39148 18450 39188 18535
rect 38859 17744 38901 17753
rect 38859 17704 38860 17744
rect 38900 17704 38901 17744
rect 38859 17695 38901 17704
rect 39532 17744 39572 17753
rect 39820 17744 39860 19048
rect 39916 18929 39956 19216
rect 40011 19256 40053 19265
rect 40011 19216 40012 19256
rect 40052 19216 40053 19256
rect 40011 19207 40053 19216
rect 40108 19256 40148 19375
rect 40108 19207 40148 19216
rect 40491 19256 40533 19265
rect 40491 19216 40492 19256
rect 40532 19216 40533 19256
rect 40491 19207 40533 19216
rect 40395 19172 40437 19181
rect 40395 19132 40396 19172
rect 40436 19132 40437 19172
rect 40395 19123 40437 19132
rect 40204 19088 40244 19097
rect 40244 19048 40340 19088
rect 40204 19039 40244 19048
rect 39915 18920 39957 18929
rect 39915 18880 39916 18920
rect 39956 18880 39957 18920
rect 39915 18871 39957 18880
rect 40203 18920 40245 18929
rect 40203 18880 40204 18920
rect 40244 18880 40245 18920
rect 40203 18871 40245 18880
rect 40204 18080 40244 18871
rect 40300 18500 40340 19048
rect 40396 19038 40436 19123
rect 40492 18752 40532 19207
rect 40684 18929 40724 19804
rect 41068 19256 41108 20719
rect 41260 20096 41300 21475
rect 41740 20768 41780 20777
rect 41644 20728 41740 20768
rect 41644 20105 41684 20728
rect 41740 20719 41780 20728
rect 41739 20348 41781 20357
rect 41739 20308 41740 20348
rect 41780 20308 41781 20348
rect 41739 20299 41781 20308
rect 41260 19853 41300 20056
rect 41643 20096 41685 20105
rect 41643 20056 41644 20096
rect 41684 20056 41685 20096
rect 41643 20047 41685 20056
rect 41740 20096 41780 20299
rect 41932 20273 41972 20358
rect 41931 20264 41973 20273
rect 41931 20224 41932 20264
rect 41972 20224 41973 20264
rect 41931 20215 41973 20224
rect 41740 20047 41780 20056
rect 41836 20096 41876 20105
rect 42028 20096 42068 20105
rect 41259 19844 41301 19853
rect 41259 19804 41260 19844
rect 41300 19804 41301 19844
rect 41259 19795 41301 19804
rect 41836 19769 41876 20056
rect 41932 20056 42028 20096
rect 41835 19760 41877 19769
rect 41835 19720 41836 19760
rect 41876 19720 41877 19760
rect 41835 19711 41877 19720
rect 41932 19265 41972 20056
rect 42028 20047 42068 20056
rect 40683 18920 40725 18929
rect 40683 18880 40684 18920
rect 40724 18880 40725 18920
rect 40683 18871 40725 18880
rect 40492 18703 40532 18712
rect 40300 18460 40436 18500
rect 40299 18332 40341 18341
rect 40299 18292 40300 18332
rect 40340 18292 40341 18332
rect 40299 18283 40341 18292
rect 40300 18198 40340 18283
rect 40204 18040 40340 18080
rect 40204 17744 40244 17753
rect 39820 17704 40204 17744
rect 38860 17610 38900 17695
rect 38571 17072 38613 17081
rect 38571 17032 38572 17072
rect 38612 17032 38613 17072
rect 38571 17023 38613 17032
rect 38572 16938 38612 17023
rect 39532 16997 39572 17704
rect 40204 17695 40244 17704
rect 40300 17744 40340 18040
rect 40396 17744 40436 18460
rect 41068 18341 41108 19216
rect 41931 19256 41973 19265
rect 41931 19216 41932 19256
rect 41972 19216 41973 19256
rect 41931 19207 41973 19216
rect 42124 18593 42164 21568
rect 42219 20600 42261 20609
rect 42219 20560 42220 20600
rect 42260 20560 42261 20600
rect 42219 20551 42261 20560
rect 42220 20012 42260 20551
rect 42220 19963 42260 19972
rect 42316 19433 42356 21736
rect 42507 21736 42508 21776
rect 42548 21736 42549 21776
rect 42507 21727 42549 21736
rect 42604 21776 42644 23071
rect 43084 22952 43124 22961
rect 43276 22952 43316 23743
rect 43372 23288 43412 25339
rect 43852 25304 43892 25313
rect 44044 25304 44084 26608
rect 44140 26599 44180 26608
rect 44331 26396 44373 26405
rect 44331 26356 44332 26396
rect 44372 26356 44373 26396
rect 44331 26347 44373 26356
rect 44235 26228 44277 26237
rect 44235 26188 44236 26228
rect 44276 26188 44277 26228
rect 44235 26179 44277 26188
rect 44236 26094 44276 26179
rect 44332 26144 44372 26347
rect 44332 26095 44372 26104
rect 43892 25264 44084 25304
rect 43852 25255 43892 25264
rect 43563 25220 43605 25229
rect 43563 25180 43564 25220
rect 43604 25180 43605 25220
rect 43563 25171 43605 25180
rect 44331 25220 44373 25229
rect 44331 25180 44332 25220
rect 44372 25180 44373 25220
rect 44331 25171 44373 25180
rect 43564 25086 43604 25171
rect 44332 24716 44372 25171
rect 44428 25136 44468 26683
rect 44523 26480 44565 26489
rect 44523 26440 44524 26480
rect 44564 26440 44565 26480
rect 44523 26431 44565 26440
rect 44524 25304 44564 26431
rect 44620 26321 44660 27112
rect 44715 26984 44757 26993
rect 44715 26944 44716 26984
rect 44756 26944 44757 26984
rect 44715 26935 44757 26944
rect 44716 26648 44756 26935
rect 44812 26816 44852 27112
rect 44812 26767 44852 26776
rect 44716 26608 44852 26648
rect 44715 26480 44757 26489
rect 44715 26440 44716 26480
rect 44756 26440 44757 26480
rect 44715 26431 44757 26440
rect 44619 26312 44661 26321
rect 44619 26272 44620 26312
rect 44660 26272 44661 26312
rect 44619 26263 44661 26272
rect 44620 26144 44660 26155
rect 44620 26069 44660 26104
rect 44619 26060 44661 26069
rect 44619 26020 44620 26060
rect 44660 26020 44661 26060
rect 44619 26011 44661 26020
rect 44524 25255 44564 25264
rect 44620 25304 44660 25313
rect 44620 25136 44660 25264
rect 44716 25304 44756 26431
rect 44716 25255 44756 25264
rect 44812 25304 44852 26608
rect 44908 25472 44948 27616
rect 45100 27068 45140 27775
rect 45388 27665 45428 28960
rect 45580 28496 45620 28505
rect 45484 28456 45580 28496
rect 45387 27656 45429 27665
rect 45387 27616 45388 27656
rect 45428 27616 45429 27656
rect 45387 27607 45429 27616
rect 45388 27522 45428 27607
rect 45291 27404 45333 27413
rect 45291 27364 45292 27404
rect 45332 27364 45333 27404
rect 45291 27355 45333 27364
rect 45100 27019 45140 27028
rect 45003 26900 45045 26909
rect 45003 26860 45004 26900
rect 45044 26860 45045 26900
rect 45003 26851 45045 26860
rect 45004 26816 45044 26851
rect 45004 26765 45044 26776
rect 45292 26816 45332 27355
rect 45387 26984 45429 26993
rect 45387 26944 45388 26984
rect 45428 26944 45429 26984
rect 45387 26935 45429 26944
rect 45292 26767 45332 26776
rect 45388 26816 45428 26935
rect 45388 26767 45428 26776
rect 45003 26648 45045 26657
rect 45484 26648 45524 28456
rect 45580 28447 45620 28456
rect 45579 27236 45621 27245
rect 45579 27196 45580 27236
rect 45620 27196 45621 27236
rect 45579 27187 45621 27196
rect 45580 27068 45620 27187
rect 45580 27019 45620 27028
rect 45003 26608 45004 26648
rect 45044 26608 45045 26648
rect 45003 26599 45045 26608
rect 45388 26608 45524 26648
rect 45580 26816 45620 26825
rect 45772 26816 45812 28960
rect 45868 28253 45908 29128
rect 46252 29168 46292 29959
rect 46636 29874 46676 29959
rect 47884 29840 47924 29849
rect 46444 29672 46484 29681
rect 47788 29672 47828 29681
rect 46484 29632 46580 29672
rect 46444 29623 46484 29632
rect 46252 29119 46292 29128
rect 46540 28337 46580 29632
rect 47115 29168 47157 29177
rect 47115 29128 47116 29168
rect 47156 29128 47157 29168
rect 47115 29119 47157 29128
rect 47116 29034 47156 29119
rect 47403 28496 47445 28505
rect 47403 28456 47404 28496
rect 47444 28456 47445 28496
rect 47403 28447 47445 28456
rect 46156 28328 46196 28337
rect 46444 28328 46484 28337
rect 46196 28288 46444 28328
rect 46156 28279 46196 28288
rect 46444 28279 46484 28288
rect 46539 28328 46581 28337
rect 46539 28288 46540 28328
rect 46580 28288 46581 28328
rect 46539 28279 46581 28288
rect 47115 28328 47157 28337
rect 47115 28288 47116 28328
rect 47156 28288 47157 28328
rect 47115 28279 47157 28288
rect 47404 28328 47444 28447
rect 47404 28279 47444 28288
rect 47500 28328 47540 28337
rect 45867 28244 45909 28253
rect 45867 28204 45868 28244
rect 45908 28204 45909 28244
rect 45867 28195 45909 28204
rect 47116 28194 47156 28279
rect 46060 28160 46100 28169
rect 46100 28120 46196 28160
rect 46060 28111 46100 28120
rect 46059 27236 46101 27245
rect 46059 27196 46060 27236
rect 46100 27196 46101 27236
rect 46059 27187 46101 27196
rect 45963 26984 46005 26993
rect 45963 26944 45964 26984
rect 46004 26944 46005 26984
rect 45963 26935 46005 26944
rect 45867 26816 45909 26825
rect 45772 26776 45868 26816
rect 45908 26776 45909 26816
rect 45004 26228 45044 26599
rect 45004 26179 45044 26188
rect 45388 26144 45428 26608
rect 45580 26573 45620 26776
rect 45867 26767 45909 26776
rect 45868 26682 45908 26767
rect 45964 26741 46004 26935
rect 45963 26732 46005 26741
rect 45963 26692 45964 26732
rect 46004 26692 46005 26732
rect 45963 26683 46005 26692
rect 45579 26564 45621 26573
rect 45579 26524 45580 26564
rect 45620 26524 45621 26564
rect 45579 26515 45621 26524
rect 46060 26321 46100 27187
rect 46059 26312 46101 26321
rect 46059 26272 46060 26312
rect 46100 26272 46101 26312
rect 46059 26263 46101 26272
rect 45388 26095 45428 26104
rect 45963 25976 46005 25985
rect 45963 25936 45964 25976
rect 46004 25936 46005 25976
rect 45963 25927 46005 25936
rect 45579 25892 45621 25901
rect 45579 25852 45580 25892
rect 45620 25852 45621 25892
rect 45579 25843 45621 25852
rect 45100 25472 45140 25481
rect 44908 25432 45100 25472
rect 45100 25423 45140 25432
rect 44812 25255 44852 25264
rect 45580 25304 45620 25843
rect 45580 25255 45620 25264
rect 45964 25318 46004 25927
rect 46156 25397 46196 28120
rect 47500 27749 47540 28288
rect 47596 28328 47636 28337
rect 47499 27740 47541 27749
rect 47499 27700 47500 27740
rect 47540 27700 47541 27740
rect 47499 27691 47541 27700
rect 46251 27656 46293 27665
rect 46251 27616 46252 27656
rect 46292 27616 46293 27656
rect 46251 27607 46293 27616
rect 46828 27656 46868 27665
rect 46252 26144 46292 27607
rect 46540 27404 46580 27413
rect 46444 27364 46540 27404
rect 46444 26405 46484 27364
rect 46540 27355 46580 27364
rect 46731 27404 46773 27413
rect 46731 27364 46732 27404
rect 46772 27364 46773 27404
rect 46731 27355 46773 27364
rect 46732 27270 46772 27355
rect 46539 27068 46581 27077
rect 46539 27028 46540 27068
rect 46580 27028 46581 27068
rect 46539 27019 46581 27028
rect 46540 26934 46580 27019
rect 46731 26984 46773 26993
rect 46731 26944 46732 26984
rect 46772 26944 46773 26984
rect 46731 26935 46773 26944
rect 46443 26396 46485 26405
rect 46443 26356 46444 26396
rect 46484 26356 46485 26396
rect 46443 26347 46485 26356
rect 46252 26095 46292 26104
rect 46251 25556 46293 25565
rect 46251 25516 46252 25556
rect 46292 25516 46293 25556
rect 46251 25507 46293 25516
rect 46155 25388 46197 25397
rect 45964 25229 46004 25278
rect 46060 25348 46156 25388
rect 46196 25348 46197 25388
rect 45771 25220 45813 25229
rect 45771 25180 45772 25220
rect 45812 25180 45813 25220
rect 45771 25171 45813 25180
rect 45963 25220 46005 25229
rect 45963 25180 45964 25220
rect 46004 25180 46005 25220
rect 45963 25171 46005 25180
rect 44428 25096 44660 25136
rect 44332 24667 44372 24676
rect 43948 24632 43988 24641
rect 43660 24592 43948 24632
rect 44620 24632 44660 25096
rect 45483 25136 45525 25145
rect 45483 25096 45484 25136
rect 45524 25096 45525 25136
rect 45483 25087 45525 25096
rect 45484 25002 45524 25087
rect 45772 25086 45812 25171
rect 45964 25154 46004 25171
rect 44716 24632 44756 24641
rect 44620 24592 44716 24632
rect 43660 23960 43700 24592
rect 43948 24583 43988 24592
rect 44716 24583 44756 24592
rect 45676 24632 45716 24641
rect 44908 23960 44948 23969
rect 43660 23911 43700 23920
rect 44812 23920 44908 23960
rect 43372 23239 43412 23248
rect 43564 23248 43796 23288
rect 43124 22912 43316 22952
rect 43468 23120 43508 23129
rect 43084 22903 43124 22912
rect 43468 22700 43508 23080
rect 43564 23120 43604 23248
rect 43564 23071 43604 23080
rect 43660 23120 43700 23129
rect 43563 22868 43605 22877
rect 43563 22828 43564 22868
rect 43604 22828 43605 22868
rect 43563 22819 43605 22828
rect 43084 22660 43508 22700
rect 43084 22532 43124 22660
rect 43564 22532 43604 22819
rect 43660 22793 43700 23080
rect 43659 22784 43701 22793
rect 43659 22744 43660 22784
rect 43700 22744 43701 22784
rect 43659 22735 43701 22744
rect 43084 22483 43124 22492
rect 43372 22492 43604 22532
rect 42987 22364 43029 22373
rect 42987 22324 42988 22364
rect 43028 22324 43029 22364
rect 42987 22315 43029 22324
rect 42604 21727 42644 21736
rect 42796 22280 42836 22289
rect 42411 20600 42453 20609
rect 42411 20560 42412 20600
rect 42452 20560 42453 20600
rect 42411 20551 42453 20560
rect 42315 19424 42357 19433
rect 42315 19384 42316 19424
rect 42356 19384 42357 19424
rect 42315 19375 42357 19384
rect 42219 19256 42261 19265
rect 42219 19216 42220 19256
rect 42260 19216 42261 19256
rect 42219 19207 42261 19216
rect 42316 19256 42356 19265
rect 42220 19122 42260 19207
rect 42316 19088 42356 19216
rect 42412 19256 42452 20551
rect 42508 20180 42548 21727
rect 42796 20609 42836 22240
rect 42988 22280 43028 22315
rect 42988 22229 43028 22240
rect 43180 22280 43220 22289
rect 43180 22121 43220 22240
rect 43372 22280 43412 22492
rect 43756 22373 43796 23248
rect 43947 23120 43989 23129
rect 43947 23080 43948 23120
rect 43988 23080 43989 23120
rect 43947 23071 43989 23080
rect 44236 23120 44276 23129
rect 43948 22986 43988 23071
rect 44236 22961 44276 23080
rect 44428 23120 44468 23129
rect 44235 22952 44277 22961
rect 44235 22912 44236 22952
rect 44276 22912 44277 22952
rect 44235 22903 44277 22912
rect 43852 22868 43892 22877
rect 43852 22457 43892 22828
rect 44139 22868 44181 22877
rect 44139 22828 44140 22868
rect 44180 22828 44181 22868
rect 44139 22819 44181 22828
rect 44140 22734 44180 22819
rect 44428 22709 44468 23080
rect 44812 23120 44852 23920
rect 44908 23911 44948 23920
rect 45676 23885 45716 24592
rect 45675 23876 45717 23885
rect 45388 23836 45676 23876
rect 45716 23836 45717 23876
rect 45195 23792 45237 23801
rect 45195 23752 45196 23792
rect 45236 23752 45237 23792
rect 45195 23743 45237 23752
rect 44812 23071 44852 23080
rect 44427 22700 44469 22709
rect 44427 22660 44428 22700
rect 44468 22660 44469 22700
rect 44427 22651 44469 22660
rect 45196 22625 45236 23743
rect 45195 22616 45237 22625
rect 45195 22576 45196 22616
rect 45236 22576 45237 22616
rect 45195 22567 45237 22576
rect 43851 22448 43893 22457
rect 43851 22408 43852 22448
rect 43892 22408 43893 22448
rect 43851 22399 43893 22408
rect 44043 22448 44085 22457
rect 44043 22408 44044 22448
rect 44084 22408 44085 22448
rect 44043 22399 44085 22408
rect 44523 22448 44565 22457
rect 44523 22408 44524 22448
rect 44564 22408 44565 22448
rect 44523 22399 44565 22408
rect 45003 22448 45045 22457
rect 45003 22408 45004 22448
rect 45044 22408 45045 22448
rect 45003 22399 45045 22408
rect 43755 22364 43797 22373
rect 43755 22324 43756 22364
rect 43796 22324 43797 22364
rect 43755 22315 43797 22324
rect 43372 22231 43412 22240
rect 43468 22280 43508 22289
rect 43468 22205 43508 22240
rect 43659 22280 43701 22289
rect 43659 22240 43660 22280
rect 43700 22240 43701 22280
rect 43659 22231 43701 22240
rect 43852 22280 43892 22291
rect 43467 22196 43509 22205
rect 43467 22156 43468 22196
rect 43508 22156 43509 22196
rect 43467 22147 43509 22156
rect 43179 22112 43221 22121
rect 43179 22072 43180 22112
rect 43220 22072 43221 22112
rect 43179 22063 43221 22072
rect 43084 21608 43124 21617
rect 43371 21608 43413 21617
rect 43124 21568 43316 21608
rect 43084 21559 43124 21568
rect 42891 21440 42933 21449
rect 42891 21400 42892 21440
rect 42932 21400 42933 21440
rect 42891 21391 42933 21400
rect 42892 21029 42932 21391
rect 42891 21020 42933 21029
rect 42891 20980 42892 21020
rect 42932 20980 42933 21020
rect 42891 20971 42933 20980
rect 42892 20886 42932 20971
rect 43276 20777 43316 21568
rect 43371 21568 43372 21608
rect 43412 21568 43413 21608
rect 43371 21559 43413 21568
rect 43372 21474 43412 21559
rect 43468 21533 43508 22147
rect 43660 22146 43700 22231
rect 43852 22205 43892 22240
rect 43948 22280 43988 22289
rect 43851 22196 43893 22205
rect 43851 22156 43852 22196
rect 43892 22156 43893 22196
rect 43851 22147 43893 22156
rect 43564 22112 43604 22121
rect 43467 21524 43509 21533
rect 43467 21484 43468 21524
rect 43508 21484 43509 21524
rect 43467 21475 43509 21484
rect 43084 20768 43124 20777
rect 42795 20600 42837 20609
rect 42795 20560 42796 20600
rect 42836 20560 42837 20600
rect 42795 20551 42837 20560
rect 43084 20273 43124 20728
rect 43275 20768 43317 20777
rect 43275 20728 43276 20768
rect 43316 20728 43317 20768
rect 43275 20719 43317 20728
rect 43083 20264 43125 20273
rect 43083 20224 43084 20264
rect 43124 20224 43125 20264
rect 43083 20215 43125 20224
rect 42508 20140 42644 20180
rect 42507 19760 42549 19769
rect 42507 19720 42508 19760
rect 42548 19720 42549 19760
rect 42507 19711 42549 19720
rect 42412 19207 42452 19216
rect 42508 19256 42548 19711
rect 42508 19207 42548 19216
rect 42604 19088 42644 20140
rect 43179 19676 43221 19685
rect 43179 19636 43180 19676
rect 43220 19636 43221 19676
rect 43179 19627 43221 19636
rect 43180 19508 43220 19627
rect 43180 19459 43220 19468
rect 42891 19424 42933 19433
rect 42891 19384 42892 19424
rect 42932 19384 42933 19424
rect 42891 19375 42933 19384
rect 42892 19290 42932 19375
rect 42316 19048 42644 19088
rect 41643 18584 41685 18593
rect 41643 18544 41644 18584
rect 41684 18544 41685 18584
rect 41643 18535 41685 18544
rect 42123 18584 42165 18593
rect 42508 18584 42548 18593
rect 42123 18544 42124 18584
rect 42164 18544 42165 18584
rect 42123 18535 42165 18544
rect 42220 18544 42508 18584
rect 41644 18450 41684 18535
rect 41067 18332 41109 18341
rect 41067 18292 41068 18332
rect 41108 18292 41109 18332
rect 41067 18283 41109 18292
rect 40492 17912 40532 17921
rect 41740 17912 41780 17921
rect 42220 17912 42260 18544
rect 42508 18535 42548 18544
rect 42892 18584 42932 18593
rect 40532 17872 40724 17912
rect 40492 17863 40532 17872
rect 40492 17744 40532 17753
rect 40396 17704 40492 17744
rect 40300 17695 40340 17704
rect 40492 17695 40532 17704
rect 40684 17744 40724 17872
rect 41780 17872 42260 17912
rect 41740 17863 41780 17872
rect 42892 17753 42932 18544
rect 40684 17695 40724 17704
rect 41355 17744 41397 17753
rect 41355 17704 41356 17744
rect 41396 17704 41397 17744
rect 41355 17695 41397 17704
rect 42891 17744 42933 17753
rect 42891 17704 42892 17744
rect 42932 17704 42933 17744
rect 42891 17695 42933 17704
rect 41356 17610 41396 17695
rect 42987 17660 43029 17669
rect 42987 17620 42988 17660
rect 43028 17620 43029 17660
rect 42987 17611 43029 17620
rect 40299 17072 40341 17081
rect 40299 17032 40300 17072
rect 40340 17032 40341 17072
rect 40299 17023 40341 17032
rect 42892 17072 42932 17081
rect 42988 17072 43028 17611
rect 43276 17156 43316 20719
rect 43371 20096 43413 20105
rect 43371 20056 43372 20096
rect 43412 20056 43413 20096
rect 43371 20047 43413 20056
rect 43372 19962 43412 20047
rect 43564 19004 43604 22072
rect 43948 21188 43988 22240
rect 44044 22280 44084 22399
rect 44044 22231 44084 22240
rect 44139 22280 44181 22289
rect 44139 22240 44140 22280
rect 44180 22240 44181 22280
rect 44139 22231 44181 22240
rect 44332 22280 44372 22289
rect 44140 22146 44180 22231
rect 44044 21608 44084 21617
rect 44044 21449 44084 21568
rect 44235 21608 44277 21617
rect 44235 21568 44236 21608
rect 44276 21568 44277 21608
rect 44235 21559 44277 21568
rect 44332 21608 44372 22240
rect 44236 21474 44276 21559
rect 44332 21533 44372 21568
rect 44428 22280 44468 22289
rect 44331 21524 44373 21533
rect 44331 21484 44332 21524
rect 44372 21484 44373 21524
rect 44331 21475 44373 21484
rect 44043 21440 44085 21449
rect 44043 21400 44044 21440
rect 44084 21400 44085 21440
rect 44043 21391 44085 21400
rect 43852 21148 43988 21188
rect 43755 20600 43797 20609
rect 43755 20560 43756 20600
rect 43796 20560 43797 20600
rect 43755 20551 43797 20560
rect 43756 20466 43796 20551
rect 43852 19685 43892 21148
rect 44236 21020 44276 21029
rect 44428 21020 44468 22240
rect 44524 22280 44564 22399
rect 44812 22280 44852 22289
rect 44524 22231 44564 22240
rect 44716 22240 44812 22280
rect 44620 22112 44660 22121
rect 44524 21608 44564 21617
rect 44620 21608 44660 22072
rect 44564 21568 44660 21608
rect 44524 21559 44564 21568
rect 44523 21440 44565 21449
rect 44523 21400 44524 21440
rect 44564 21400 44565 21440
rect 44523 21391 44565 21400
rect 44524 21306 44564 21391
rect 44044 20980 44236 21020
rect 44276 20980 44468 21020
rect 44044 20768 44084 20980
rect 44236 20971 44276 20980
rect 44044 20719 44084 20728
rect 43948 20600 43988 20609
rect 43948 20357 43988 20560
rect 44619 20600 44661 20609
rect 44619 20560 44620 20600
rect 44660 20560 44661 20600
rect 44619 20551 44661 20560
rect 43947 20348 43989 20357
rect 43947 20308 43948 20348
rect 43988 20308 43989 20348
rect 43947 20299 43989 20308
rect 44620 20180 44660 20551
rect 44620 20131 44660 20140
rect 44236 20096 44276 20105
rect 43851 19676 43893 19685
rect 43851 19636 43852 19676
rect 43892 19636 43893 19676
rect 43851 19627 43893 19636
rect 43851 19508 43893 19517
rect 43851 19468 43852 19508
rect 43892 19468 43893 19508
rect 43851 19459 43893 19468
rect 43852 19265 43892 19459
rect 44236 19433 44276 20056
rect 44235 19424 44277 19433
rect 44235 19384 44236 19424
rect 44276 19384 44277 19424
rect 44235 19375 44277 19384
rect 43851 19256 43893 19265
rect 43851 19216 43852 19256
rect 43892 19216 43893 19256
rect 43851 19207 43893 19216
rect 44044 19256 44084 19265
rect 43852 19122 43892 19207
rect 44044 19004 44084 19216
rect 44235 19256 44277 19265
rect 44716 19256 44756 22240
rect 44812 22231 44852 22240
rect 45004 22280 45044 22399
rect 45004 21701 45044 22240
rect 45196 21776 45236 22567
rect 45388 22457 45428 23836
rect 45675 23827 45717 23836
rect 45772 23801 45812 23886
rect 45771 23792 45813 23801
rect 45771 23752 45772 23792
rect 45812 23752 45813 23792
rect 45771 23743 45813 23752
rect 45868 23792 45908 23801
rect 45676 23624 45716 23633
rect 45716 23584 45812 23624
rect 45676 23575 45716 23584
rect 45676 23120 45716 23129
rect 45484 23080 45676 23120
rect 45387 22448 45429 22457
rect 45387 22408 45388 22448
rect 45428 22408 45429 22448
rect 45387 22399 45429 22408
rect 45388 22280 45428 22291
rect 45388 22205 45428 22240
rect 45387 22196 45429 22205
rect 45387 22156 45388 22196
rect 45428 22156 45429 22196
rect 45387 22147 45429 22156
rect 45196 21727 45236 21736
rect 45292 22112 45332 22121
rect 45003 21692 45045 21701
rect 45003 21652 45004 21692
rect 45044 21652 45045 21692
rect 45003 21643 45045 21652
rect 45292 21617 45332 22072
rect 45291 21608 45333 21617
rect 45291 21568 45292 21608
rect 45332 21568 45333 21608
rect 45291 21559 45333 21568
rect 44907 21188 44949 21197
rect 44907 21148 44908 21188
rect 44948 21148 44949 21188
rect 44907 21139 44949 21148
rect 44908 20768 44948 21139
rect 45387 20768 45429 20777
rect 44948 20728 45236 20768
rect 44908 20719 44948 20728
rect 45196 20264 45236 20728
rect 45387 20728 45388 20768
rect 45428 20728 45429 20768
rect 45387 20719 45429 20728
rect 45388 20634 45428 20719
rect 45196 20215 45236 20224
rect 45484 20105 45524 23080
rect 45676 23071 45716 23080
rect 45772 22952 45812 23584
rect 45868 23549 45908 23752
rect 45963 23792 46005 23801
rect 45963 23752 45964 23792
rect 46004 23752 46005 23792
rect 45963 23743 46005 23752
rect 45964 23658 46004 23743
rect 45867 23540 45909 23549
rect 45867 23500 45868 23540
rect 45908 23500 45909 23540
rect 45867 23491 45909 23500
rect 45580 22912 45812 22952
rect 45580 22280 45620 22912
rect 46060 22868 46100 25348
rect 46155 25339 46197 25348
rect 46155 25220 46197 25229
rect 46155 25180 46156 25220
rect 46196 25180 46197 25220
rect 46155 25171 46197 25180
rect 46156 23792 46196 25171
rect 46252 24800 46292 25507
rect 46443 25304 46485 25313
rect 46443 25264 46444 25304
rect 46484 25264 46485 25304
rect 46443 25255 46485 25264
rect 46347 25220 46389 25229
rect 46347 25180 46348 25220
rect 46388 25180 46389 25220
rect 46347 25171 46389 25180
rect 46348 25052 46388 25171
rect 46444 25170 46484 25255
rect 46539 25136 46581 25145
rect 46539 25096 46540 25136
rect 46580 25096 46581 25136
rect 46539 25087 46581 25096
rect 46348 25012 46484 25052
rect 46252 24751 46292 24760
rect 46348 24632 46388 24641
rect 46252 24044 46292 24053
rect 46348 24044 46388 24592
rect 46444 24632 46484 25012
rect 46540 24641 46580 25087
rect 46732 24725 46772 26935
rect 46828 26489 46868 27616
rect 47020 27404 47060 27413
rect 47020 26909 47060 27364
rect 47019 26900 47061 26909
rect 47019 26860 47020 26900
rect 47060 26860 47061 26900
rect 47019 26851 47061 26860
rect 47212 26648 47252 26657
rect 47212 26489 47252 26608
rect 46827 26480 46869 26489
rect 46827 26440 46828 26480
rect 46868 26440 46869 26480
rect 46827 26431 46869 26440
rect 47211 26480 47253 26489
rect 47211 26440 47212 26480
rect 47252 26440 47253 26480
rect 47211 26431 47253 26440
rect 47403 26480 47445 26489
rect 47403 26440 47404 26480
rect 47444 26440 47445 26480
rect 47403 26431 47445 26440
rect 47404 26312 47444 26431
rect 47404 26237 47444 26272
rect 47403 26228 47445 26237
rect 47403 26188 47404 26228
rect 47444 26188 47445 26228
rect 47403 26179 47445 26188
rect 47115 26144 47157 26153
rect 47115 26104 47116 26144
rect 47156 26104 47157 26144
rect 47115 26095 47157 26104
rect 47019 25556 47061 25565
rect 47019 25516 47020 25556
rect 47060 25516 47061 25556
rect 47019 25507 47061 25516
rect 46923 25388 46965 25397
rect 46923 25348 46924 25388
rect 46964 25348 46965 25388
rect 46923 25339 46965 25348
rect 47020 25388 47060 25507
rect 47020 25339 47060 25348
rect 46924 25254 46964 25339
rect 46827 25220 46869 25229
rect 47116 25220 47156 26095
rect 47403 25724 47445 25733
rect 47403 25684 47404 25724
rect 47444 25684 47445 25724
rect 47403 25675 47445 25684
rect 47211 25640 47253 25649
rect 47211 25600 47212 25640
rect 47252 25600 47253 25640
rect 47211 25591 47253 25600
rect 46827 25180 46828 25220
rect 46868 25180 46869 25220
rect 46827 25171 46869 25180
rect 47020 25180 47156 25220
rect 46731 24716 46773 24725
rect 46731 24676 46732 24716
rect 46772 24676 46773 24716
rect 46731 24667 46773 24676
rect 46444 24583 46484 24592
rect 46539 24632 46581 24641
rect 46539 24592 46540 24632
rect 46580 24592 46581 24632
rect 46539 24583 46581 24592
rect 46732 24632 46772 24667
rect 46540 24498 46580 24583
rect 46732 24582 46772 24592
rect 46828 24632 46868 25171
rect 47020 24800 47060 25180
rect 47212 24800 47252 25591
rect 47404 25304 47444 25675
rect 47596 25649 47636 28288
rect 47691 28328 47733 28337
rect 47691 28288 47692 28328
rect 47732 28288 47733 28328
rect 47691 28279 47733 28288
rect 47692 28194 47732 28279
rect 47692 27656 47732 27665
rect 47692 26405 47732 27616
rect 47691 26396 47733 26405
rect 47691 26356 47692 26396
rect 47732 26356 47733 26396
rect 47691 26347 47733 26356
rect 47788 26144 47828 29632
rect 47884 29345 47924 29800
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 47883 29336 47925 29345
rect 47883 29296 47884 29336
rect 47924 29296 47925 29336
rect 47883 29287 47925 29296
rect 48459 29336 48501 29345
rect 48459 29296 48460 29336
rect 48500 29296 48501 29336
rect 48459 29287 48501 29296
rect 48460 29202 48500 29287
rect 49132 29168 49172 29177
rect 49036 29128 49132 29168
rect 48268 29084 48308 29093
rect 49036 29084 49076 29128
rect 49132 29119 49172 29128
rect 48308 29044 49076 29084
rect 48268 29035 48308 29044
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 48267 28496 48309 28505
rect 48748 28496 48788 28505
rect 48267 28456 48268 28496
rect 48308 28456 48309 28496
rect 48267 28447 48309 28456
rect 48556 28456 48748 28496
rect 47884 28160 47924 28169
rect 47884 27740 47924 28120
rect 47884 27691 47924 27700
rect 48268 27656 48308 28447
rect 48556 28328 48596 28456
rect 48748 28447 48788 28456
rect 49227 28496 49269 28505
rect 49227 28456 49228 28496
rect 49268 28456 49269 28496
rect 49227 28447 49269 28456
rect 48939 28412 48981 28421
rect 48939 28372 48940 28412
rect 48980 28372 48981 28412
rect 48939 28363 48981 28372
rect 48556 28279 48596 28288
rect 48747 28328 48789 28337
rect 48747 28288 48748 28328
rect 48788 28288 48789 28328
rect 48747 28279 48789 28288
rect 48940 28328 48980 28363
rect 49228 28362 49268 28447
rect 48748 28194 48788 28279
rect 48940 28277 48980 28288
rect 49036 28328 49076 28337
rect 49036 27833 49076 28288
rect 50283 28328 50325 28337
rect 50283 28288 50284 28328
rect 50324 28288 50325 28328
rect 50283 28279 50325 28288
rect 50571 28328 50613 28337
rect 50571 28288 50572 28328
rect 50612 28288 50613 28328
rect 50571 28279 50613 28288
rect 49900 28160 49940 28169
rect 49228 28120 49900 28160
rect 49035 27824 49077 27833
rect 49035 27784 49036 27824
rect 49076 27784 49077 27824
rect 49035 27775 49077 27784
rect 48268 27607 48308 27616
rect 49132 27656 49172 27665
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 49132 27077 49172 27616
rect 49131 27068 49173 27077
rect 49131 27028 49132 27068
rect 49172 27028 49173 27068
rect 49131 27019 49173 27028
rect 48171 26984 48213 26993
rect 48171 26944 48172 26984
rect 48212 26944 48213 26984
rect 48171 26935 48213 26944
rect 47884 26816 47924 26825
rect 47884 26489 47924 26776
rect 48172 26816 48212 26935
rect 48172 26767 48212 26776
rect 47979 26732 48021 26741
rect 47979 26692 47980 26732
rect 48020 26692 48021 26732
rect 47979 26683 48021 26692
rect 48939 26732 48981 26741
rect 48939 26692 48940 26732
rect 48980 26692 48981 26732
rect 48939 26683 48981 26692
rect 49036 26732 49076 26741
rect 47883 26480 47925 26489
rect 47883 26440 47884 26480
rect 47924 26440 47925 26480
rect 47883 26431 47925 26440
rect 47788 25733 47828 26104
rect 47884 26130 47924 26139
rect 47884 26069 47924 26090
rect 47883 26060 47925 26069
rect 47980 26060 48020 26683
rect 48267 26312 48309 26321
rect 48267 26272 48268 26312
rect 48308 26272 48309 26312
rect 48267 26263 48309 26272
rect 48940 26312 48980 26683
rect 48940 26263 48980 26272
rect 48076 26153 48116 26238
rect 48075 26144 48117 26153
rect 48075 26104 48076 26144
rect 48116 26104 48117 26144
rect 48075 26095 48117 26104
rect 48268 26144 48308 26263
rect 49036 26153 49076 26692
rect 48268 26095 48308 26104
rect 49035 26144 49077 26153
rect 49035 26104 49036 26144
rect 49076 26104 49077 26144
rect 49035 26095 49077 26104
rect 49132 26144 49172 26153
rect 47883 26020 47884 26060
rect 47924 26020 48020 26060
rect 47883 26011 47925 26020
rect 47884 25995 47924 26011
rect 47883 25808 47925 25817
rect 47883 25768 47884 25808
rect 47924 25768 47925 25808
rect 47883 25759 47925 25768
rect 47787 25724 47829 25733
rect 47787 25684 47788 25724
rect 47828 25684 47829 25724
rect 47787 25675 47829 25684
rect 47595 25640 47637 25649
rect 47595 25600 47596 25640
rect 47636 25600 47637 25640
rect 47595 25591 47637 25600
rect 47499 25472 47541 25481
rect 47499 25432 47500 25472
rect 47540 25432 47541 25472
rect 47499 25423 47541 25432
rect 47404 25255 47444 25264
rect 47500 25304 47540 25423
rect 47500 25255 47540 25264
rect 47595 25304 47637 25313
rect 47595 25264 47596 25304
rect 47636 25264 47637 25304
rect 47595 25255 47637 25264
rect 47787 25304 47829 25313
rect 47787 25264 47788 25304
rect 47828 25264 47829 25304
rect 47787 25255 47829 25264
rect 47884 25304 47924 25759
rect 47980 25304 48020 26020
rect 49132 25985 49172 26104
rect 48075 25976 48117 25985
rect 48075 25936 48076 25976
rect 48116 25936 48117 25976
rect 48075 25927 48117 25936
rect 49131 25976 49173 25985
rect 49131 25936 49132 25976
rect 49172 25936 49173 25976
rect 49131 25927 49173 25936
rect 48076 25842 48116 25927
rect 49228 25808 49268 28120
rect 49900 28111 49940 28120
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 50284 27749 50324 28279
rect 50572 28194 50612 28279
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 50283 27740 50325 27749
rect 50283 27700 50284 27740
rect 50324 27700 50325 27740
rect 50283 27691 50325 27700
rect 50284 27572 50324 27691
rect 50284 27523 50324 27532
rect 51148 27656 51188 27665
rect 50476 27404 50516 27413
rect 49707 26816 49749 26825
rect 49707 26776 49708 26816
rect 49748 26776 49749 26816
rect 49707 26767 49749 26776
rect 49323 26732 49365 26741
rect 49323 26692 49324 26732
rect 49364 26692 49365 26732
rect 49323 26683 49365 26692
rect 49324 26598 49364 26683
rect 49708 26682 49748 26767
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 49132 25768 49268 25808
rect 49804 25892 49844 25901
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 48267 25640 48309 25649
rect 48267 25600 48268 25640
rect 48308 25600 48309 25640
rect 48267 25591 48309 25600
rect 48268 25481 48308 25591
rect 48843 25556 48885 25565
rect 48843 25516 48844 25556
rect 48884 25516 48885 25556
rect 48843 25507 48885 25516
rect 48267 25472 48309 25481
rect 48267 25432 48268 25472
rect 48308 25432 48309 25472
rect 48267 25423 48309 25432
rect 48076 25304 48116 25313
rect 47980 25264 48076 25304
rect 47884 25255 47924 25264
rect 48076 25255 48116 25264
rect 48172 25304 48212 25313
rect 47020 24751 47060 24760
rect 47116 24760 47252 24800
rect 46828 24583 46868 24592
rect 46924 24632 46964 24641
rect 47116 24632 47156 24760
rect 46964 24592 47156 24632
rect 47211 24632 47253 24641
rect 47211 24592 47212 24632
rect 47252 24592 47253 24632
rect 46292 24004 46388 24044
rect 46732 24044 46772 24053
rect 46924 24044 46964 24592
rect 47211 24583 47253 24592
rect 47308 24632 47348 24641
rect 47500 24632 47540 24641
rect 47212 24498 47252 24583
rect 46772 24004 46964 24044
rect 46252 23995 46292 24004
rect 46732 23995 46772 24004
rect 47308 23885 47348 24592
rect 47404 24592 47500 24632
rect 46539 23876 46581 23885
rect 47307 23876 47349 23885
rect 46539 23836 46540 23876
rect 46580 23836 46581 23876
rect 46539 23827 46581 23836
rect 47212 23836 47308 23876
rect 47348 23836 47349 23876
rect 46156 23743 46196 23752
rect 46348 23792 46388 23801
rect 46155 23624 46197 23633
rect 46155 23584 46156 23624
rect 46196 23584 46197 23624
rect 46155 23575 46197 23584
rect 45964 22828 46100 22868
rect 45675 22700 45717 22709
rect 45675 22660 45676 22700
rect 45716 22660 45717 22700
rect 45675 22651 45717 22660
rect 45580 22231 45620 22240
rect 45676 22196 45716 22651
rect 45771 22616 45813 22625
rect 45964 22616 46004 22828
rect 46059 22700 46101 22709
rect 46059 22660 46060 22700
rect 46100 22660 46101 22700
rect 46059 22651 46101 22660
rect 45771 22576 45772 22616
rect 45812 22576 45813 22616
rect 45771 22567 45813 22576
rect 45872 22576 46004 22616
rect 45772 22280 45812 22567
rect 45872 22532 45912 22576
rect 45868 22492 45912 22532
rect 45868 22448 45908 22492
rect 45867 22408 45908 22448
rect 45867 22364 45907 22408
rect 45867 22324 45908 22364
rect 45772 22231 45812 22240
rect 45868 22280 45908 22324
rect 45868 22231 45908 22240
rect 46060 22280 46100 22651
rect 46060 22231 46100 22240
rect 46156 22280 46196 23575
rect 46348 23297 46388 23752
rect 46540 23742 46580 23827
rect 47212 23717 47252 23836
rect 47307 23827 47349 23836
rect 47211 23708 47253 23717
rect 47211 23668 47212 23708
rect 47252 23668 47253 23708
rect 47211 23659 47253 23668
rect 46924 23624 46964 23633
rect 46539 23540 46581 23549
rect 46539 23500 46540 23540
rect 46580 23500 46581 23540
rect 46539 23491 46581 23500
rect 46347 23288 46389 23297
rect 46347 23248 46348 23288
rect 46388 23248 46389 23288
rect 46347 23239 46389 23248
rect 46251 22364 46293 22373
rect 46251 22324 46252 22364
rect 46292 22324 46293 22364
rect 46251 22315 46293 22324
rect 46156 22231 46196 22240
rect 46252 22280 46292 22315
rect 45676 22147 45716 22156
rect 46252 21785 46292 22240
rect 46347 22280 46389 22289
rect 46347 22240 46348 22280
rect 46388 22240 46389 22280
rect 46347 22231 46389 22240
rect 46348 22146 46388 22231
rect 46540 22205 46580 23491
rect 46827 23288 46869 23297
rect 46827 23248 46828 23288
rect 46868 23248 46869 23288
rect 46827 23239 46869 23248
rect 46828 23154 46868 23239
rect 46924 23129 46964 23584
rect 47019 23372 47061 23381
rect 47019 23332 47020 23372
rect 47060 23332 47061 23372
rect 47019 23323 47061 23332
rect 46923 23120 46965 23129
rect 46923 23080 46924 23120
rect 46964 23080 46965 23120
rect 46923 23071 46965 23080
rect 47020 22289 47060 23323
rect 47115 23288 47157 23297
rect 47115 23248 47116 23288
rect 47156 23248 47157 23288
rect 47115 23239 47157 23248
rect 47019 22280 47061 22289
rect 47019 22240 47020 22280
rect 47060 22240 47061 22280
rect 47116 22280 47156 23239
rect 47212 23120 47252 23659
rect 47404 23381 47444 24592
rect 47500 24583 47540 24592
rect 47499 24464 47541 24473
rect 47499 24424 47500 24464
rect 47540 24424 47541 24464
rect 47499 24415 47541 24424
rect 47500 24330 47540 24415
rect 47596 23960 47636 25255
rect 47788 25170 47828 25255
rect 47692 24632 47732 24641
rect 47692 24473 47732 24592
rect 47691 24464 47733 24473
rect 47691 24424 47692 24464
rect 47732 24424 47733 24464
rect 47691 24415 47733 24424
rect 47787 24380 47829 24389
rect 47787 24340 47788 24380
rect 47828 24340 47829 24380
rect 47787 24331 47829 24340
rect 47596 23920 47732 23960
rect 47596 23792 47636 23801
rect 47596 23633 47636 23752
rect 47595 23624 47637 23633
rect 47595 23584 47596 23624
rect 47636 23584 47637 23624
rect 47595 23575 47637 23584
rect 47403 23372 47445 23381
rect 47403 23332 47404 23372
rect 47444 23332 47445 23372
rect 47403 23323 47445 23332
rect 47212 22709 47252 23080
rect 47308 23120 47348 23129
rect 47308 22961 47348 23080
rect 47404 23120 47444 23129
rect 47307 22952 47349 22961
rect 47307 22912 47308 22952
rect 47348 22912 47349 22952
rect 47307 22903 47349 22912
rect 47211 22700 47253 22709
rect 47211 22660 47212 22700
rect 47252 22660 47253 22700
rect 47211 22651 47253 22660
rect 47212 22280 47252 22289
rect 47116 22240 47212 22280
rect 47019 22231 47061 22240
rect 47212 22231 47252 22240
rect 46539 22196 46581 22205
rect 46539 22156 46540 22196
rect 46580 22156 46581 22196
rect 46539 22147 46581 22156
rect 46540 22062 46580 22147
rect 47404 21785 47444 23080
rect 47500 23120 47540 23129
rect 47500 22793 47540 23080
rect 47595 23120 47637 23129
rect 47595 23080 47596 23120
rect 47636 23080 47637 23120
rect 47595 23071 47637 23080
rect 47499 22784 47541 22793
rect 47499 22744 47500 22784
rect 47540 22744 47541 22784
rect 47499 22735 47541 22744
rect 47499 22616 47541 22625
rect 47499 22576 47500 22616
rect 47540 22576 47541 22616
rect 47499 22567 47541 22576
rect 47500 21860 47540 22567
rect 47596 22448 47636 23071
rect 47596 22399 47636 22408
rect 47692 22280 47732 23920
rect 47788 23204 47828 24331
rect 48172 23969 48212 25264
rect 48268 25304 48308 25423
rect 48268 25255 48308 25264
rect 48556 25304 48596 25313
rect 48596 25264 48692 25304
rect 48556 25255 48596 25264
rect 48364 25136 48404 25145
rect 48404 25096 48596 25136
rect 48364 25087 48404 25096
rect 48556 24632 48596 25096
rect 48652 24800 48692 25264
rect 48652 24751 48692 24760
rect 48844 24800 48884 25507
rect 49036 24800 49076 24809
rect 48844 24760 49036 24800
rect 48747 24716 48789 24725
rect 48747 24676 48748 24716
rect 48788 24676 48789 24716
rect 48747 24667 48789 24676
rect 48556 24583 48596 24592
rect 48748 24632 48788 24667
rect 48363 24380 48405 24389
rect 48363 24340 48364 24380
rect 48404 24340 48405 24380
rect 48748 24380 48788 24592
rect 48844 24632 48884 24760
rect 49036 24751 49076 24760
rect 48844 24583 48884 24592
rect 49132 24632 49172 25768
rect 49419 25556 49461 25565
rect 49419 25516 49420 25556
rect 49460 25516 49461 25556
rect 49419 25507 49461 25516
rect 49420 25388 49460 25507
rect 49420 25229 49460 25348
rect 49804 25313 49844 25852
rect 50091 25892 50133 25901
rect 50091 25852 50092 25892
rect 50132 25852 50133 25892
rect 50091 25843 50133 25852
rect 50092 25758 50132 25843
rect 50476 25817 50516 27364
rect 51148 27077 51188 27616
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 50571 27068 50613 27077
rect 51147 27068 51189 27077
rect 50571 27028 50572 27068
rect 50612 27028 50613 27068
rect 50571 27019 50613 27028
rect 51052 27028 51148 27068
rect 51188 27028 51189 27068
rect 50572 26816 50612 27019
rect 50475 25808 50517 25817
rect 50475 25768 50476 25808
rect 50516 25768 50517 25808
rect 50475 25759 50517 25768
rect 49803 25304 49845 25313
rect 49803 25264 49804 25304
rect 49844 25264 49845 25304
rect 49803 25255 49845 25264
rect 50572 25304 50612 26776
rect 50764 26144 50804 26153
rect 50764 25565 50804 26104
rect 50955 26144 50997 26153
rect 50955 26104 50956 26144
rect 50996 26104 50997 26144
rect 50955 26095 50997 26104
rect 51052 26144 51092 27028
rect 51147 27019 51189 27028
rect 51723 27068 51765 27077
rect 51723 27028 51724 27068
rect 51764 27028 51765 27068
rect 51723 27019 51765 27028
rect 51724 26934 51764 27019
rect 51435 26816 51477 26825
rect 51435 26776 51436 26816
rect 51476 26776 51477 26816
rect 51435 26767 51477 26776
rect 51243 26564 51285 26573
rect 51243 26524 51244 26564
rect 51284 26524 51285 26564
rect 51243 26515 51285 26524
rect 51244 26312 51284 26515
rect 51244 26263 51284 26272
rect 51052 26095 51092 26104
rect 51148 26144 51188 26153
rect 50956 26010 50996 26095
rect 50763 25556 50805 25565
rect 50763 25516 50764 25556
rect 50804 25516 50805 25556
rect 50763 25507 50805 25516
rect 51148 25481 51188 26104
rect 51436 25976 51476 26767
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 51436 25927 51476 25936
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 51147 25472 51189 25481
rect 51147 25432 51148 25472
rect 51188 25432 51189 25472
rect 51147 25423 51189 25432
rect 49419 25220 49461 25229
rect 49419 25180 49420 25220
rect 49460 25180 49461 25220
rect 49419 25171 49461 25180
rect 49228 25136 49268 25145
rect 49228 24716 49268 25096
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 49324 24716 49364 24725
rect 49228 24676 49324 24716
rect 49324 24667 49364 24676
rect 49708 24632 49748 24641
rect 49132 24583 49172 24592
rect 49612 24592 49708 24632
rect 48748 24340 48980 24380
rect 48363 24331 48405 24340
rect 48364 24246 48404 24331
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 48171 23960 48213 23969
rect 48940 23960 48980 24340
rect 48171 23920 48172 23960
rect 48212 23920 48213 23960
rect 48171 23911 48213 23920
rect 48748 23920 48980 23960
rect 49612 23960 49652 24592
rect 49708 24583 49748 24592
rect 50572 24632 50612 25264
rect 47883 23876 47925 23885
rect 47883 23836 47884 23876
rect 47924 23836 47925 23876
rect 47883 23827 47925 23836
rect 47788 23155 47828 23164
rect 47788 22280 47828 22289
rect 47692 22240 47788 22280
rect 47788 22231 47828 22240
rect 47884 22280 47924 23827
rect 48748 23792 48788 23920
rect 49612 23911 49652 23920
rect 50475 23876 50517 23885
rect 50475 23836 50476 23876
rect 50516 23836 50517 23876
rect 50475 23827 50517 23836
rect 48748 23743 48788 23752
rect 49132 23792 49172 23801
rect 49804 23792 49844 23801
rect 49172 23752 49804 23792
rect 49132 23743 49172 23752
rect 49804 23743 49844 23752
rect 50476 23792 50516 23827
rect 50476 23741 50516 23752
rect 49036 23624 49076 23633
rect 48940 23584 49036 23624
rect 48171 23120 48213 23129
rect 48171 23080 48172 23120
rect 48212 23080 48213 23120
rect 48171 23071 48213 23080
rect 48172 22986 48212 23071
rect 48363 22952 48405 22961
rect 48363 22912 48364 22952
rect 48404 22912 48405 22952
rect 48363 22903 48405 22912
rect 48075 22784 48117 22793
rect 48075 22744 48076 22784
rect 48116 22744 48117 22784
rect 48075 22735 48117 22744
rect 47500 21820 47732 21860
rect 46156 21776 46196 21785
rect 46251 21776 46293 21785
rect 46196 21736 46252 21776
rect 46292 21736 46293 21776
rect 46156 21727 46196 21736
rect 46251 21727 46293 21736
rect 47211 21776 47253 21785
rect 47211 21736 47212 21776
rect 47252 21736 47253 21776
rect 47211 21727 47253 21736
rect 47403 21776 47445 21785
rect 47403 21736 47404 21776
rect 47444 21736 47445 21776
rect 47692 21776 47732 21820
rect 47692 21736 47828 21776
rect 47403 21727 47445 21736
rect 45579 21692 45621 21701
rect 45579 21652 45580 21692
rect 45620 21652 45621 21692
rect 45579 21643 45621 21652
rect 45580 21608 45620 21643
rect 46252 21642 46292 21727
rect 46347 21692 46389 21701
rect 46347 21652 46348 21692
rect 46388 21652 46389 21692
rect 46347 21643 46389 21652
rect 45580 21557 45620 21568
rect 46348 21524 46388 21643
rect 47019 21608 47061 21617
rect 47019 21568 47020 21608
rect 47060 21568 47061 21608
rect 47019 21559 47061 21568
rect 47116 21608 47156 21617
rect 46348 21475 46388 21484
rect 47020 21474 47060 21559
rect 46539 21440 46581 21449
rect 46539 21400 46540 21440
rect 46580 21400 46581 21440
rect 46539 21391 46581 21400
rect 46732 21440 46772 21449
rect 46347 20768 46389 20777
rect 46347 20728 46348 20768
rect 46388 20728 46389 20768
rect 46347 20719 46389 20728
rect 46540 20768 46580 21391
rect 46540 20719 46580 20728
rect 46348 20105 46388 20719
rect 45483 20096 45525 20105
rect 45483 20056 45484 20096
rect 45524 20056 45525 20096
rect 45483 20047 45525 20056
rect 46347 20096 46389 20105
rect 46347 20056 46348 20096
rect 46388 20056 46389 20096
rect 46732 20096 46772 21400
rect 47116 20609 47156 21568
rect 47212 21608 47252 21727
rect 47595 21692 47637 21701
rect 47595 21652 47596 21692
rect 47636 21652 47637 21692
rect 47595 21643 47637 21652
rect 47212 21559 47252 21568
rect 47308 21608 47348 21617
rect 47500 21608 47540 21617
rect 47348 21568 47500 21608
rect 47308 21559 47348 21568
rect 47500 21559 47540 21568
rect 47596 21558 47636 21643
rect 47691 21608 47733 21617
rect 47691 21568 47692 21608
rect 47732 21568 47733 21608
rect 47691 21559 47733 21568
rect 47788 21608 47828 21736
rect 47788 21559 47828 21568
rect 47692 21440 47732 21559
rect 47884 21440 47924 22240
rect 48076 22280 48116 22735
rect 48364 22532 48404 22903
rect 48940 22793 48980 23584
rect 49036 23575 49076 23584
rect 50187 23624 50229 23633
rect 50187 23584 50188 23624
rect 50228 23584 50229 23624
rect 50187 23575 50229 23584
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 50188 23288 50228 23575
rect 50188 23239 50228 23248
rect 49035 23120 49077 23129
rect 49035 23080 49036 23120
rect 49076 23080 49077 23120
rect 49035 23071 49077 23080
rect 50475 23120 50517 23129
rect 50572 23120 50612 24592
rect 51436 25304 51476 25313
rect 50860 23960 50900 23969
rect 51436 23960 51476 25264
rect 51819 25304 51861 25313
rect 51819 25264 51820 25304
rect 51860 25264 51861 25304
rect 51819 25255 51861 25264
rect 51820 25170 51860 25255
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 51724 24380 51764 24389
rect 51724 23969 51764 24340
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 50900 23920 51476 23960
rect 51723 23960 51765 23969
rect 51723 23920 51724 23960
rect 51764 23920 51765 23960
rect 50860 23911 50900 23920
rect 51723 23911 51765 23920
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 50475 23080 50476 23120
rect 50516 23080 50612 23120
rect 50475 23071 50517 23080
rect 49036 22986 49076 23071
rect 48939 22784 48981 22793
rect 48939 22744 48940 22784
rect 48980 22744 48981 22784
rect 48939 22735 48981 22744
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 48364 22483 48404 22492
rect 49035 22448 49077 22457
rect 49035 22408 49036 22448
rect 49076 22408 49077 22448
rect 49035 22399 49077 22408
rect 48076 22231 48116 22240
rect 49036 22280 49076 22399
rect 47979 22196 48021 22205
rect 47979 22156 47980 22196
rect 48020 22156 48021 22196
rect 47979 22147 48021 22156
rect 47980 22062 48020 22147
rect 49036 22121 49076 22240
rect 49612 22280 49652 22289
rect 49227 22196 49269 22205
rect 49227 22156 49228 22196
rect 49268 22156 49269 22196
rect 49227 22147 49269 22156
rect 49035 22112 49077 22121
rect 49035 22072 49036 22112
rect 49076 22072 49077 22112
rect 49035 22063 49077 22072
rect 49228 22062 49268 22147
rect 47979 21692 48021 21701
rect 47979 21652 47980 21692
rect 48020 21652 48021 21692
rect 47979 21643 48021 21652
rect 47980 21608 48020 21643
rect 47980 21557 48020 21568
rect 48651 21524 48693 21533
rect 48651 21484 48652 21524
rect 48692 21484 48693 21524
rect 48651 21475 48693 21484
rect 47692 21400 47924 21440
rect 48652 21390 48692 21475
rect 49035 21440 49077 21449
rect 49035 21400 49036 21440
rect 49076 21400 49077 21440
rect 49612 21440 49652 22240
rect 50476 22280 50516 23071
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 51627 22448 51669 22457
rect 51627 22408 51628 22448
rect 51668 22408 51669 22448
rect 51627 22399 51669 22408
rect 51628 22314 51668 22399
rect 50476 22231 50516 22240
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 50283 21524 50325 21533
rect 50283 21484 50284 21524
rect 50324 21484 50325 21524
rect 50283 21475 50325 21484
rect 49708 21440 49748 21449
rect 49612 21400 49708 21440
rect 49035 21391 49077 21400
rect 49708 21391 49748 21400
rect 49899 21440 49941 21449
rect 49899 21400 49900 21440
rect 49940 21400 49941 21440
rect 49899 21391 49941 21400
rect 49036 21306 49076 21391
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 49035 20768 49077 20777
rect 49035 20728 49036 20768
rect 49076 20728 49077 20768
rect 49035 20719 49077 20728
rect 49900 20768 49940 21391
rect 49900 20719 49940 20728
rect 50284 20768 50324 21475
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 50284 20719 50324 20728
rect 49036 20634 49076 20719
rect 47115 20600 47157 20609
rect 47115 20560 47116 20600
rect 47156 20560 47157 20600
rect 47115 20551 47157 20560
rect 47212 20600 47252 20609
rect 47787 20600 47829 20609
rect 47884 20600 47924 20609
rect 47252 20560 47636 20600
rect 47212 20551 47252 20560
rect 47596 20180 47636 20560
rect 47787 20560 47788 20600
rect 47828 20560 47884 20600
rect 47787 20551 47829 20560
rect 47884 20551 47924 20560
rect 47596 20131 47636 20140
rect 47212 20096 47252 20105
rect 46732 20056 47212 20096
rect 46347 20047 46389 20056
rect 47212 20047 47252 20056
rect 45099 19424 45141 19433
rect 45099 19384 45100 19424
rect 45140 19384 45141 19424
rect 45099 19375 45141 19384
rect 45100 19290 45140 19375
rect 44235 19216 44236 19256
rect 44276 19216 44277 19256
rect 44235 19207 44277 19216
rect 44620 19216 44756 19256
rect 43564 18964 44084 19004
rect 44236 18584 44276 19207
rect 44236 18535 44276 18544
rect 44620 17669 44660 19216
rect 44716 19088 44756 19097
rect 44716 18593 44756 19048
rect 44715 18584 44757 18593
rect 44715 18544 44716 18584
rect 44756 18544 44757 18584
rect 44715 18535 44757 18544
rect 45484 18584 45524 20047
rect 46348 19962 46388 20047
rect 47788 19937 47828 20551
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 47787 19928 47829 19937
rect 47787 19888 47788 19928
rect 47828 19888 47829 19928
rect 47787 19879 47829 19888
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 46347 19424 46389 19433
rect 46347 19384 46348 19424
rect 46388 19384 46389 19424
rect 46347 19375 46389 19384
rect 45484 18535 45524 18544
rect 46348 18584 46388 19375
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 46348 18535 46388 18544
rect 46731 18584 46773 18593
rect 46731 18544 46732 18584
rect 46772 18544 46773 18584
rect 46731 18535 46773 18544
rect 46732 18450 46772 18535
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 44619 17660 44661 17669
rect 44619 17620 44620 17660
rect 44660 17620 44661 17660
rect 44619 17611 44661 17620
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 43276 17107 43316 17116
rect 42932 17032 43028 17072
rect 44140 17072 44180 17081
rect 42892 17023 42932 17032
rect 39531 16988 39573 16997
rect 39531 16948 39532 16988
rect 39572 16948 39573 16988
rect 39531 16939 39573 16948
rect 39723 16988 39765 16997
rect 39723 16948 39724 16988
rect 39764 16948 39765 16988
rect 39723 16939 39765 16948
rect 39724 16854 39764 16939
rect 39628 16232 39668 16241
rect 39668 16192 39764 16232
rect 39628 16183 39668 16192
rect 39052 16148 39092 16157
rect 39244 16148 39284 16157
rect 39092 16108 39244 16148
rect 39052 16099 39092 16108
rect 39244 16099 39284 16108
rect 39724 15392 39764 16192
rect 39724 15343 39764 15352
rect 38955 14888 38997 14897
rect 39052 14888 39092 14897
rect 38955 14848 38956 14888
rect 38996 14848 39052 14888
rect 38955 14839 38997 14848
rect 39052 14839 39092 14848
rect 39723 14888 39765 14897
rect 39723 14848 39724 14888
rect 39764 14848 39765 14888
rect 39723 14839 39765 14848
rect 38420 14176 38516 14216
rect 38380 14167 38420 14176
rect 37995 14132 38037 14141
rect 37995 14092 37996 14132
rect 38036 14092 38037 14132
rect 37995 14083 38037 14092
rect 37612 14048 37652 14057
rect 37996 14048 38036 14083
rect 37652 14008 37748 14048
rect 37612 13999 37652 14008
rect 37611 13796 37653 13805
rect 37611 13756 37612 13796
rect 37652 13756 37653 13796
rect 37611 13747 37653 13756
rect 37612 13662 37652 13747
rect 37516 13159 37556 13168
rect 37612 13208 37652 13217
rect 37708 13208 37748 14008
rect 37996 13997 38036 14008
rect 37652 13168 37748 13208
rect 37803 13208 37845 13217
rect 37803 13168 37804 13208
rect 37844 13168 37845 13208
rect 37612 13159 37652 13168
rect 37803 13159 37845 13168
rect 37324 12704 37364 13159
rect 37804 13074 37844 13159
rect 38284 12872 38324 14167
rect 38571 14132 38613 14141
rect 38571 14092 38572 14132
rect 38612 14092 38613 14132
rect 38571 14083 38613 14092
rect 37804 12832 38324 12872
rect 37324 12664 37460 12704
rect 37228 12536 37268 12545
rect 37132 12496 37228 12536
rect 37036 12452 37076 12496
rect 37228 12487 37268 12496
rect 37323 12536 37365 12545
rect 37323 12496 37324 12536
rect 37364 12496 37365 12536
rect 37323 12487 37365 12496
rect 37036 12412 37172 12452
rect 37036 12284 37076 12293
rect 36939 12032 36981 12041
rect 36939 11992 36940 12032
rect 36980 11992 36981 12032
rect 36939 11983 36981 11992
rect 37036 11789 37076 12244
rect 37132 12209 37172 12412
rect 37324 12402 37364 12487
rect 37131 12200 37173 12209
rect 37131 12160 37132 12200
rect 37172 12160 37173 12200
rect 37131 12151 37173 12160
rect 37227 12116 37269 12125
rect 37227 12076 37228 12116
rect 37268 12076 37269 12116
rect 37227 12067 37269 12076
rect 37035 11780 37077 11789
rect 37035 11740 37036 11780
rect 37076 11740 37077 11780
rect 37035 11731 37077 11740
rect 36556 11696 36596 11705
rect 36556 11453 36596 11656
rect 36652 11696 36692 11705
rect 36652 11537 36692 11656
rect 36651 11528 36693 11537
rect 36651 11488 36652 11528
rect 36692 11488 36693 11528
rect 36651 11479 36693 11488
rect 36844 11528 36884 11537
rect 36555 11444 36597 11453
rect 36555 11404 36556 11444
rect 36596 11404 36597 11444
rect 36555 11395 36597 11404
rect 36651 11276 36693 11285
rect 36460 11236 36652 11276
rect 36692 11236 36693 11276
rect 36651 11227 36693 11236
rect 36171 11192 36213 11201
rect 36076 11152 36172 11192
rect 36212 11152 36213 11192
rect 36171 11143 36213 11152
rect 36363 11192 36405 11201
rect 36363 11152 36364 11192
rect 36404 11152 36405 11192
rect 36363 11143 36405 11152
rect 35980 11068 36116 11108
rect 35595 10940 35637 10949
rect 35595 10900 35596 10940
rect 35636 10900 35637 10940
rect 35595 10891 35637 10900
rect 35692 10772 35732 10984
rect 35788 11024 35828 11033
rect 35828 10984 35924 11024
rect 35788 10975 35828 10984
rect 35596 10732 35732 10772
rect 34923 10520 34965 10529
rect 34923 10480 34924 10520
rect 34964 10480 34965 10520
rect 34923 10471 34965 10480
rect 35307 10520 35349 10529
rect 35307 10480 35308 10520
rect 35348 10480 35349 10520
rect 35307 10471 35349 10480
rect 34676 10144 34828 10184
rect 34636 10135 34676 10144
rect 34828 10135 34868 10144
rect 34924 10184 34964 10471
rect 35019 10352 35061 10361
rect 35019 10312 35020 10352
rect 35060 10312 35061 10352
rect 35019 10303 35061 10312
rect 34924 10135 34964 10144
rect 35020 10184 35060 10303
rect 35596 10199 35636 10732
rect 35020 10135 35060 10144
rect 35308 10184 35348 10195
rect 34059 10100 34101 10109
rect 34059 10060 34060 10100
rect 34100 10060 34101 10100
rect 34059 10051 34101 10060
rect 34060 9966 34100 10051
rect 34540 10050 34580 10135
rect 35308 10109 35348 10144
rect 35403 10184 35445 10193
rect 35403 10144 35404 10184
rect 35444 10144 35445 10184
rect 35692 10193 35732 10278
rect 35596 10150 35636 10159
rect 35691 10184 35733 10193
rect 35403 10135 35445 10144
rect 35691 10144 35692 10184
rect 35732 10144 35733 10184
rect 35691 10135 35733 10144
rect 35792 10184 35834 10193
rect 35792 10144 35793 10184
rect 35833 10144 35834 10184
rect 35792 10135 35834 10144
rect 35307 10100 35349 10109
rect 35307 10060 35308 10100
rect 35348 10060 35349 10100
rect 35307 10051 35349 10060
rect 35404 10050 35444 10135
rect 35793 10050 35833 10135
rect 35116 10016 35156 10025
rect 35596 10016 35636 10025
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 35116 9521 35156 9976
rect 35500 9976 35596 10016
rect 34156 9512 34196 9521
rect 34444 9512 34484 9521
rect 33579 9260 33621 9269
rect 33579 9220 33580 9260
rect 33620 9220 33621 9260
rect 33579 9211 33621 9220
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 33579 8840 33621 8849
rect 33579 8800 33580 8840
rect 33620 8800 33621 8840
rect 33579 8791 33621 8800
rect 34059 8840 34101 8849
rect 34059 8800 34060 8840
rect 34100 8800 34101 8840
rect 34059 8791 34101 8800
rect 33580 8672 33620 8791
rect 33771 8756 33813 8765
rect 33771 8716 33772 8756
rect 33812 8716 33813 8756
rect 33771 8707 33813 8716
rect 32811 8336 32853 8345
rect 32811 8296 32812 8336
rect 32852 8296 32853 8336
rect 32811 8287 32853 8296
rect 32523 6824 32565 6833
rect 32523 6784 32524 6824
rect 32564 6784 32565 6824
rect 32523 6775 32565 6784
rect 32428 6616 32564 6656
rect 32331 6572 32373 6581
rect 32331 6532 32332 6572
rect 32372 6532 32468 6572
rect 32331 6523 32373 6532
rect 32428 6488 32468 6532
rect 32428 6439 32468 6448
rect 32140 6355 32180 6364
rect 32332 6404 32372 6413
rect 32042 6320 32084 6329
rect 32042 6280 32043 6320
rect 32083 6280 32084 6320
rect 32042 6271 32084 6280
rect 31659 6236 31701 6245
rect 31659 6196 31660 6236
rect 31700 6196 31701 6236
rect 31659 6187 31701 6196
rect 31756 6236 31796 6245
rect 32044 6236 32084 6271
rect 32236 6278 32276 6287
rect 32236 6236 32276 6238
rect 31796 6196 31988 6236
rect 32044 6196 32276 6236
rect 31756 6187 31796 6196
rect 31564 6028 31892 6068
rect 31083 5984 31125 5993
rect 31083 5944 31084 5984
rect 31124 5944 31125 5984
rect 31083 5935 31125 5944
rect 31852 5825 31892 6028
rect 31948 5993 31988 6196
rect 32043 6068 32085 6077
rect 32043 6028 32044 6068
rect 32084 6028 32085 6068
rect 32043 6019 32085 6028
rect 31947 5984 31989 5993
rect 31947 5944 31948 5984
rect 31988 5944 31989 5984
rect 31947 5935 31989 5944
rect 31179 5816 31221 5825
rect 31179 5776 31180 5816
rect 31220 5776 31221 5816
rect 31179 5767 31221 5776
rect 31563 5816 31605 5825
rect 31563 5776 31564 5816
rect 31604 5776 31605 5816
rect 31563 5767 31605 5776
rect 31851 5816 31893 5825
rect 31851 5776 31852 5816
rect 31892 5776 31893 5816
rect 31851 5767 31893 5776
rect 31083 5648 31125 5657
rect 31083 5608 31084 5648
rect 31124 5608 31125 5648
rect 31083 5599 31125 5608
rect 31084 5514 31124 5599
rect 30604 4927 30644 4936
rect 30796 5272 31028 5312
rect 30315 4892 30357 4901
rect 30315 4852 30316 4892
rect 30356 4852 30357 4892
rect 30315 4843 30357 4852
rect 30796 3725 30836 5272
rect 30892 5144 30932 5153
rect 30892 4817 30932 5104
rect 30987 5060 31029 5069
rect 30987 5020 30988 5060
rect 31028 5020 31029 5060
rect 30987 5011 31029 5020
rect 30988 4926 31028 5011
rect 31083 4976 31125 4985
rect 31083 4936 31084 4976
rect 31124 4936 31125 4976
rect 31083 4927 31125 4936
rect 31180 4976 31220 5767
rect 31564 5682 31604 5767
rect 31372 5648 31412 5657
rect 31180 4927 31220 4936
rect 31276 5480 31316 5489
rect 31084 4842 31124 4927
rect 30891 4808 30933 4817
rect 30891 4768 30892 4808
rect 30932 4768 30933 4808
rect 30891 4759 30933 4768
rect 31084 4724 31124 4733
rect 30987 4220 31029 4229
rect 30987 4180 30988 4220
rect 31028 4180 31029 4220
rect 30987 4171 31029 4180
rect 30795 3716 30837 3725
rect 30795 3676 30796 3716
rect 30836 3676 30837 3716
rect 30795 3667 30837 3676
rect 30988 3473 31028 4171
rect 31084 3809 31124 4684
rect 31276 3893 31316 5440
rect 31372 4136 31412 5608
rect 31852 5648 31892 5767
rect 31852 5599 31892 5608
rect 31947 5648 31989 5657
rect 31947 5608 31948 5648
rect 31988 5608 31989 5648
rect 31947 5599 31989 5608
rect 31948 5514 31988 5599
rect 32044 5476 32084 6019
rect 32236 5816 32276 5825
rect 32139 5564 32181 5573
rect 32139 5524 32140 5564
rect 32180 5524 32181 5564
rect 32139 5515 32181 5524
rect 32044 5427 32084 5436
rect 31563 4976 31605 4985
rect 31563 4936 31564 4976
rect 31604 4936 31605 4976
rect 31563 4927 31605 4936
rect 31467 4892 31509 4901
rect 31467 4852 31468 4892
rect 31508 4852 31509 4892
rect 31467 4843 31509 4852
rect 31372 4087 31412 4096
rect 31468 4136 31508 4843
rect 31468 4087 31508 4096
rect 31564 4136 31604 4927
rect 31948 4724 31988 4733
rect 31851 4556 31893 4565
rect 31851 4516 31852 4556
rect 31892 4516 31893 4556
rect 31851 4507 31893 4516
rect 31564 4087 31604 4096
rect 31659 4136 31701 4145
rect 31659 4096 31660 4136
rect 31700 4096 31701 4136
rect 31659 4087 31701 4096
rect 31852 4136 31892 4507
rect 31852 4087 31892 4096
rect 31660 4002 31700 4087
rect 31467 3968 31509 3977
rect 31467 3928 31468 3968
rect 31508 3928 31509 3968
rect 31467 3919 31509 3928
rect 31275 3884 31317 3893
rect 31275 3844 31276 3884
rect 31316 3844 31317 3884
rect 31275 3835 31317 3844
rect 31083 3800 31125 3809
rect 31083 3760 31084 3800
rect 31124 3760 31125 3800
rect 31083 3751 31125 3760
rect 31179 3716 31221 3725
rect 31179 3676 31180 3716
rect 31220 3676 31221 3716
rect 31179 3667 31221 3676
rect 31371 3716 31413 3725
rect 31371 3676 31372 3716
rect 31412 3676 31413 3716
rect 31371 3667 31413 3676
rect 30987 3464 31029 3473
rect 30987 3424 30988 3464
rect 31028 3424 31029 3464
rect 30987 3415 31029 3424
rect 29931 3044 29973 3053
rect 29931 3004 29932 3044
rect 29972 3004 29973 3044
rect 29931 2995 29973 3004
rect 30123 3044 30165 3053
rect 30123 3004 30124 3044
rect 30164 3004 30165 3044
rect 30123 2995 30165 3004
rect 30315 3044 30357 3053
rect 30315 3004 30316 3044
rect 30356 3004 30357 3044
rect 30315 2995 30357 3004
rect 29836 2575 29876 2584
rect 29932 2624 29972 2995
rect 29932 2575 29972 2584
rect 30316 2624 30356 2995
rect 31180 2633 31220 3667
rect 31275 3464 31317 3473
rect 31275 3424 31276 3464
rect 31316 3424 31317 3464
rect 31275 3415 31317 3424
rect 31372 3464 31412 3667
rect 31276 3330 31316 3415
rect 31372 3389 31412 3424
rect 31468 3464 31508 3919
rect 31659 3884 31701 3893
rect 31659 3844 31660 3884
rect 31700 3844 31701 3884
rect 31659 3835 31701 3844
rect 31371 3380 31413 3389
rect 31371 3340 31372 3380
rect 31412 3340 31413 3380
rect 31371 3331 31413 3340
rect 31372 3300 31412 3331
rect 31468 2801 31508 3424
rect 31563 3464 31605 3473
rect 31563 3424 31564 3464
rect 31604 3424 31605 3464
rect 31563 3415 31605 3424
rect 31564 3330 31604 3415
rect 31467 2792 31509 2801
rect 31467 2752 31468 2792
rect 31508 2752 31509 2792
rect 31467 2743 31509 2752
rect 30316 2575 30356 2584
rect 31179 2624 31221 2633
rect 31179 2584 31180 2624
rect 31220 2584 31221 2624
rect 31179 2575 31221 2584
rect 31276 2624 31316 2633
rect 31564 2624 31604 2633
rect 31316 2584 31564 2624
rect 31276 2575 31316 2584
rect 31564 2575 31604 2584
rect 28628 2500 28724 2540
rect 28875 2540 28917 2549
rect 28875 2500 28876 2540
rect 28916 2500 28917 2540
rect 28588 2491 28628 2500
rect 28875 2491 28917 2500
rect 28012 1903 28052 1912
rect 28876 1952 28916 2491
rect 28876 1903 28916 1912
rect 29260 1952 29300 1961
rect 29260 1280 29300 1912
rect 30123 1952 30165 1961
rect 30123 1912 30124 1952
rect 30164 1912 30165 1952
rect 31180 1952 31220 2575
rect 31276 1952 31316 1961
rect 31180 1912 31276 1952
rect 30123 1903 30165 1912
rect 31276 1903 31316 1912
rect 31564 1952 31604 1961
rect 31660 1952 31700 3835
rect 31948 3809 31988 4684
rect 31755 3800 31797 3809
rect 31755 3760 31756 3800
rect 31796 3760 31797 3800
rect 31755 3751 31797 3760
rect 31947 3800 31989 3809
rect 31947 3760 31948 3800
rect 31988 3760 31989 3800
rect 31947 3751 31989 3760
rect 31756 3464 31796 3751
rect 31756 3415 31796 3424
rect 32043 3464 32085 3473
rect 32043 3424 32044 3464
rect 32084 3424 32085 3464
rect 32043 3415 32085 3424
rect 32044 3330 32084 3415
rect 32044 3212 32084 3221
rect 32044 2969 32084 3172
rect 32140 3053 32180 5515
rect 32236 5321 32276 5776
rect 32332 5489 32372 6364
rect 32427 6152 32469 6161
rect 32524 6152 32564 6616
rect 32620 6161 32660 7120
rect 32812 7160 32852 8287
rect 33580 7841 33620 8632
rect 33772 8622 33812 8707
rect 34060 8706 34100 8791
rect 33868 8672 33908 8681
rect 33868 8588 33908 8632
rect 34156 8588 34196 9472
rect 34348 9472 34444 9512
rect 34348 8933 34388 9472
rect 34444 9463 34484 9472
rect 34828 9512 34868 9521
rect 34444 9344 34484 9353
rect 34828 9344 34868 9472
rect 34484 9304 34868 9344
rect 34924 9512 34964 9521
rect 34444 9295 34484 9304
rect 34731 9008 34773 9017
rect 34731 8968 34732 9008
rect 34772 8968 34773 9008
rect 34731 8959 34773 8968
rect 34347 8924 34389 8933
rect 34347 8884 34348 8924
rect 34388 8884 34389 8924
rect 34347 8875 34389 8884
rect 34251 8756 34293 8765
rect 34251 8716 34252 8756
rect 34292 8716 34293 8756
rect 34251 8707 34293 8716
rect 33868 8548 34196 8588
rect 33868 8261 33908 8548
rect 34059 8420 34101 8429
rect 34059 8380 34060 8420
rect 34100 8380 34101 8420
rect 34059 8371 34101 8380
rect 33867 8252 33909 8261
rect 33867 8212 33868 8252
rect 33908 8212 33909 8252
rect 33867 8203 33909 8212
rect 34060 8000 34100 8371
rect 34252 8168 34292 8707
rect 34348 8672 34388 8681
rect 34348 8252 34388 8632
rect 34444 8672 34484 8681
rect 34444 8513 34484 8632
rect 34732 8672 34772 8959
rect 34924 8765 34964 9472
rect 35115 9512 35157 9521
rect 35115 9472 35116 9512
rect 35156 9472 35157 9512
rect 35115 9463 35157 9472
rect 35404 9512 35444 9521
rect 35020 9428 35060 9439
rect 35020 9353 35060 9388
rect 35019 9344 35061 9353
rect 35019 9304 35020 9344
rect 35060 9304 35061 9344
rect 35019 9295 35061 9304
rect 35116 9344 35156 9353
rect 34923 8756 34965 8765
rect 34923 8716 34924 8756
rect 34964 8716 34965 8756
rect 34923 8707 34965 8716
rect 35020 8681 35060 8766
rect 34732 8623 34772 8632
rect 35019 8672 35061 8681
rect 35019 8632 35020 8672
rect 35060 8632 35061 8672
rect 35019 8623 35061 8632
rect 34443 8504 34485 8513
rect 34443 8464 34444 8504
rect 34484 8464 34485 8504
rect 34443 8455 34485 8464
rect 34540 8504 34580 8509
rect 35116 8504 35156 9304
rect 35212 9260 35252 9269
rect 35212 8681 35252 9220
rect 35211 8672 35253 8681
rect 35211 8632 35212 8672
rect 35252 8632 35253 8672
rect 35211 8623 35253 8632
rect 35212 8504 35252 8513
rect 34540 8500 35060 8504
rect 34580 8464 35060 8500
rect 35116 8464 35212 8504
rect 34540 8451 34580 8460
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 34348 8212 34484 8252
rect 34252 8128 34388 8168
rect 34060 7951 34100 7960
rect 34252 8000 34292 8009
rect 33579 7832 33621 7841
rect 33579 7792 33580 7832
rect 33620 7792 33621 7832
rect 33579 7783 33621 7792
rect 34059 7832 34101 7841
rect 34059 7792 34060 7832
rect 34100 7792 34101 7832
rect 34059 7783 34101 7792
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 33004 7328 33044 7337
rect 32812 6917 32852 7120
rect 32908 7244 32948 7253
rect 32811 6908 32853 6917
rect 32811 6868 32812 6908
rect 32852 6868 32853 6908
rect 32811 6859 32853 6868
rect 32716 6497 32756 6582
rect 32715 6488 32757 6497
rect 32908 6488 32948 7204
rect 32715 6448 32716 6488
rect 32756 6448 32948 6488
rect 32715 6439 32757 6448
rect 33004 6404 33044 7288
rect 32812 6364 33044 6404
rect 33100 7244 33140 7253
rect 32812 6320 32852 6364
rect 32716 6280 32852 6320
rect 32427 6112 32428 6152
rect 32468 6112 32564 6152
rect 32619 6152 32661 6161
rect 32619 6112 32620 6152
rect 32660 6112 32661 6152
rect 32427 6103 32469 6112
rect 32619 6103 32661 6112
rect 32619 5984 32661 5993
rect 32619 5944 32620 5984
rect 32660 5944 32661 5984
rect 32619 5935 32661 5944
rect 32523 5816 32565 5825
rect 32523 5776 32524 5816
rect 32564 5776 32565 5816
rect 32523 5767 32565 5776
rect 32524 5648 32564 5767
rect 32524 5599 32564 5608
rect 32620 5648 32660 5935
rect 32620 5599 32660 5608
rect 32331 5480 32373 5489
rect 32331 5440 32332 5480
rect 32372 5440 32373 5480
rect 32331 5431 32373 5440
rect 32716 5476 32756 6280
rect 33003 6236 33045 6245
rect 33003 6196 33004 6236
rect 33044 6196 33045 6236
rect 33003 6187 33045 6196
rect 32811 6152 32853 6161
rect 32811 6112 32812 6152
rect 32852 6112 32853 6152
rect 32811 6103 32853 6112
rect 32716 5427 32756 5436
rect 32619 5396 32661 5405
rect 32619 5356 32620 5396
rect 32660 5356 32661 5396
rect 32619 5347 32661 5356
rect 32235 5312 32277 5321
rect 32235 5272 32236 5312
rect 32276 5272 32277 5312
rect 32235 5263 32277 5272
rect 32620 4976 32660 5347
rect 32715 5060 32757 5069
rect 32715 5020 32716 5060
rect 32756 5020 32757 5060
rect 32715 5011 32757 5020
rect 32620 4927 32660 4936
rect 32716 4976 32756 5011
rect 32716 4229 32756 4936
rect 32812 4817 32852 6103
rect 32907 6068 32949 6077
rect 32907 6028 32908 6068
rect 32948 6028 32949 6068
rect 32907 6019 32949 6028
rect 32908 5648 32948 6019
rect 33004 5984 33044 6187
rect 33100 6161 33140 7204
rect 33195 7160 33237 7169
rect 33195 7120 33196 7160
rect 33236 7120 33237 7160
rect 33195 7111 33237 7120
rect 33196 7026 33236 7111
rect 34060 7076 34100 7783
rect 34252 7589 34292 7960
rect 34348 8000 34388 8128
rect 34348 7951 34388 7960
rect 34347 7832 34389 7841
rect 34347 7792 34348 7832
rect 34388 7792 34389 7832
rect 34347 7783 34389 7792
rect 34348 7698 34388 7783
rect 34251 7580 34293 7589
rect 34251 7540 34252 7580
rect 34292 7540 34293 7580
rect 34251 7531 34293 7540
rect 34252 7412 34292 7531
rect 34252 7363 34292 7372
rect 34347 7412 34389 7421
rect 34347 7372 34348 7412
rect 34388 7372 34389 7412
rect 34347 7363 34389 7372
rect 34444 7412 34484 8212
rect 34827 8168 34869 8177
rect 34827 8128 34828 8168
rect 34868 8128 34869 8168
rect 34827 8119 34869 8128
rect 34924 8168 34964 8177
rect 35020 8168 35060 8464
rect 35212 8455 35252 8464
rect 34964 8128 35060 8168
rect 35307 8168 35349 8177
rect 35307 8128 35308 8168
rect 35348 8128 35349 8168
rect 34924 8119 34964 8128
rect 35307 8119 35349 8128
rect 34828 8009 34868 8119
rect 35308 8013 35348 8119
rect 34732 8000 34772 8009
rect 34574 7985 34614 7994
rect 34540 7945 34574 7985
rect 34540 7936 34614 7945
rect 34540 7421 34580 7936
rect 34444 7363 34484 7372
rect 34539 7412 34581 7421
rect 34539 7372 34540 7412
rect 34580 7372 34581 7412
rect 34539 7363 34581 7372
rect 34155 7160 34197 7169
rect 34155 7120 34156 7160
rect 34196 7120 34197 7160
rect 34155 7111 34197 7120
rect 34348 7160 34388 7363
rect 34636 7253 34676 7338
rect 34635 7244 34677 7253
rect 34732 7244 34772 7960
rect 34827 8000 34869 8009
rect 35020 8000 35060 8009
rect 34827 7960 34828 8000
rect 34868 7960 34869 8000
rect 34827 7951 34869 7960
rect 34924 7960 35020 8000
rect 34828 7866 34868 7951
rect 34635 7204 34636 7244
rect 34676 7204 34772 7244
rect 34635 7195 34677 7204
rect 34444 7160 34484 7169
rect 34348 7120 34444 7160
rect 33964 7036 34100 7076
rect 33195 6824 33237 6833
rect 33195 6784 33196 6824
rect 33236 6784 33237 6824
rect 33195 6775 33237 6784
rect 33196 6656 33236 6775
rect 33196 6607 33236 6616
rect 33868 6488 33908 6497
rect 33964 6488 34004 7036
rect 34156 7026 34196 7111
rect 34059 6908 34101 6917
rect 34059 6868 34060 6908
rect 34100 6868 34101 6908
rect 34059 6859 34101 6868
rect 34060 6656 34100 6859
rect 34348 6833 34388 7120
rect 34444 7111 34484 7120
rect 34539 7160 34581 7169
rect 34539 7120 34540 7160
rect 34580 7120 34581 7160
rect 34539 7111 34581 7120
rect 34636 7160 34676 7195
rect 34636 7111 34676 7120
rect 34924 7160 34964 7960
rect 35020 7951 35060 7960
rect 35116 8000 35156 8009
rect 35308 7964 35348 7973
rect 35116 7841 35156 7960
rect 35404 7916 35444 9472
rect 35500 9512 35540 9976
rect 35596 9967 35636 9976
rect 35884 9932 35924 10984
rect 36076 10520 36116 11068
rect 36171 11024 36213 11033
rect 36171 10984 36172 11024
rect 36212 10984 36213 11024
rect 36171 10975 36213 10984
rect 36268 11024 36308 11033
rect 36172 10890 36212 10975
rect 36268 10865 36308 10984
rect 36363 11024 36405 11033
rect 36363 10984 36364 11024
rect 36404 10984 36405 11024
rect 36363 10975 36405 10984
rect 36460 11024 36500 11033
rect 36267 10856 36309 10865
rect 36267 10816 36268 10856
rect 36308 10816 36309 10856
rect 36267 10807 36309 10816
rect 36076 10480 36308 10520
rect 36075 10352 36117 10361
rect 36075 10312 36076 10352
rect 36116 10312 36117 10352
rect 36075 10303 36117 10312
rect 35979 10184 36021 10193
rect 35979 10144 35980 10184
rect 36020 10144 36021 10184
rect 35979 10135 36021 10144
rect 35692 9892 35924 9932
rect 35595 9848 35637 9857
rect 35595 9808 35596 9848
rect 35636 9808 35637 9848
rect 35595 9799 35637 9808
rect 35500 9463 35540 9472
rect 35596 9512 35636 9799
rect 35596 9463 35636 9472
rect 35692 9512 35732 9892
rect 35883 9680 35925 9689
rect 35883 9640 35884 9680
rect 35924 9640 35925 9680
rect 35883 9631 35925 9640
rect 35692 9463 35732 9472
rect 35787 9512 35829 9521
rect 35787 9472 35788 9512
rect 35828 9472 35829 9512
rect 35787 9463 35829 9472
rect 35884 9512 35924 9631
rect 35884 9463 35924 9472
rect 35788 9344 35828 9463
rect 35692 9304 35828 9344
rect 35883 9344 35925 9353
rect 35883 9304 35884 9344
rect 35924 9304 35925 9344
rect 35595 8672 35637 8681
rect 35595 8632 35596 8672
rect 35636 8632 35637 8672
rect 35595 8623 35637 8632
rect 35692 8672 35732 9304
rect 35883 9295 35925 9304
rect 35884 9210 35924 9295
rect 35787 9176 35829 9185
rect 35787 9136 35788 9176
rect 35828 9136 35829 9176
rect 35787 9127 35829 9136
rect 35692 8623 35732 8632
rect 35788 8672 35828 9127
rect 35980 9092 36020 10135
rect 36076 10016 36116 10303
rect 36076 9967 36116 9976
rect 36268 10184 36308 10480
rect 36364 10361 36404 10975
rect 36460 10772 36500 10984
rect 36652 11024 36692 11035
rect 36844 11033 36884 11488
rect 37132 11528 37172 11537
rect 37035 11276 37077 11285
rect 37035 11236 37036 11276
rect 37076 11236 37077 11276
rect 37035 11227 37077 11236
rect 36939 11108 36981 11117
rect 36939 11068 36940 11108
rect 36980 11068 36981 11108
rect 36939 11059 36981 11068
rect 36652 10949 36692 10984
rect 36843 11024 36885 11033
rect 36843 10984 36844 11024
rect 36884 10984 36885 11024
rect 36843 10975 36885 10984
rect 36651 10940 36693 10949
rect 36651 10900 36652 10940
rect 36692 10900 36693 10940
rect 36651 10891 36693 10900
rect 36748 10940 36788 10951
rect 36748 10865 36788 10900
rect 36940 10940 36980 11059
rect 37036 11024 37076 11227
rect 37132 11117 37172 11488
rect 37131 11108 37173 11117
rect 37131 11068 37132 11108
rect 37172 11068 37173 11108
rect 37131 11059 37173 11068
rect 37036 10975 37076 10984
rect 37228 11024 37268 12067
rect 37323 12032 37365 12041
rect 37323 11992 37324 12032
rect 37364 11992 37365 12032
rect 37323 11983 37365 11992
rect 37228 10975 37268 10984
rect 37324 11024 37364 11983
rect 37324 10975 37364 10984
rect 37420 11696 37460 12664
rect 37516 12629 37556 12660
rect 37515 12620 37557 12629
rect 37515 12580 37516 12620
rect 37556 12580 37557 12620
rect 37515 12571 37557 12580
rect 37516 12536 37556 12571
rect 37516 12461 37556 12496
rect 37804 12536 37844 12832
rect 37996 12704 38036 12713
rect 37996 12545 38036 12664
rect 38187 12620 38229 12629
rect 38187 12580 38188 12620
rect 38228 12580 38229 12620
rect 38187 12571 38229 12580
rect 37804 12487 37844 12496
rect 37995 12536 38037 12545
rect 37995 12496 37996 12536
rect 38036 12496 38037 12536
rect 37995 12487 38037 12496
rect 38188 12536 38228 12571
rect 38188 12485 38228 12496
rect 38284 12536 38324 12832
rect 38284 12487 38324 12496
rect 38476 12704 38516 12713
rect 37515 12452 37557 12461
rect 37515 12412 37516 12452
rect 37556 12412 37557 12452
rect 37515 12403 37557 12412
rect 37612 12452 37652 12461
rect 37612 12209 37652 12412
rect 38187 12284 38229 12293
rect 38187 12244 38188 12284
rect 38228 12244 38229 12284
rect 38187 12235 38229 12244
rect 37611 12200 37653 12209
rect 37611 12160 37612 12200
rect 37652 12160 37653 12200
rect 37611 12151 37653 12160
rect 36940 10891 36980 10900
rect 36747 10856 36789 10865
rect 36747 10816 36748 10856
rect 36788 10816 36789 10856
rect 36747 10807 36789 10816
rect 36844 10856 36884 10865
rect 36460 10732 36596 10772
rect 36556 10445 36596 10732
rect 36844 10520 36884 10816
rect 37227 10772 37269 10781
rect 37227 10732 37228 10772
rect 37268 10732 37269 10772
rect 37227 10723 37269 10732
rect 36844 10480 37172 10520
rect 36555 10436 36597 10445
rect 36555 10396 36556 10436
rect 36596 10396 36597 10436
rect 36555 10387 36597 10396
rect 36363 10352 36405 10361
rect 36363 10312 36364 10352
rect 36404 10312 36405 10352
rect 36363 10303 36405 10312
rect 36843 10352 36885 10361
rect 36843 10312 36844 10352
rect 36884 10312 36885 10352
rect 36843 10303 36885 10312
rect 36555 10268 36597 10277
rect 36555 10228 36556 10268
rect 36596 10228 36597 10268
rect 36555 10219 36597 10228
rect 36268 9689 36308 10144
rect 36363 10184 36405 10193
rect 36363 10144 36364 10184
rect 36404 10144 36405 10184
rect 36363 10135 36405 10144
rect 36556 10184 36596 10219
rect 36748 10193 36788 10278
rect 36267 9680 36309 9689
rect 36267 9640 36268 9680
rect 36308 9640 36309 9680
rect 36267 9631 36309 9640
rect 36172 9512 36212 9521
rect 36364 9512 36404 10135
rect 36556 10133 36596 10144
rect 36747 10184 36789 10193
rect 36747 10144 36748 10184
rect 36788 10144 36789 10184
rect 36747 10135 36789 10144
rect 36844 10184 36884 10303
rect 36844 10135 36884 10144
rect 37132 10184 37172 10480
rect 37132 10135 37172 10144
rect 37228 10184 37268 10723
rect 37323 10436 37365 10445
rect 37323 10396 37324 10436
rect 37364 10396 37365 10436
rect 37323 10387 37365 10396
rect 37228 10135 37268 10144
rect 37324 10184 37364 10387
rect 37420 10361 37460 11656
rect 37899 11696 37941 11705
rect 37899 11656 37900 11696
rect 37940 11656 37941 11696
rect 37899 11647 37941 11656
rect 37611 11276 37653 11285
rect 37611 11236 37612 11276
rect 37652 11236 37653 11276
rect 37611 11227 37653 11236
rect 37516 11192 37556 11201
rect 37516 11033 37556 11152
rect 37515 11024 37557 11033
rect 37515 10984 37516 11024
rect 37556 10984 37557 11024
rect 37515 10975 37557 10984
rect 37515 10688 37557 10697
rect 37515 10648 37516 10688
rect 37556 10648 37557 10688
rect 37515 10639 37557 10648
rect 37419 10352 37461 10361
rect 37419 10312 37420 10352
rect 37460 10312 37461 10352
rect 37419 10303 37461 10312
rect 37324 10135 37364 10144
rect 37419 10184 37461 10193
rect 37419 10144 37420 10184
rect 37460 10144 37461 10184
rect 37419 10135 37461 10144
rect 37516 10184 37556 10639
rect 37612 10613 37652 11227
rect 37804 11108 37844 11117
rect 37708 11024 37748 11033
rect 37708 10865 37748 10984
rect 37707 10856 37749 10865
rect 37707 10816 37708 10856
rect 37748 10816 37749 10856
rect 37707 10807 37749 10816
rect 37611 10604 37653 10613
rect 37611 10564 37612 10604
rect 37652 10564 37653 10604
rect 37611 10555 37653 10564
rect 37708 10445 37748 10807
rect 37707 10436 37749 10445
rect 37516 10135 37556 10144
rect 37612 10396 37708 10436
rect 37748 10396 37749 10436
rect 36651 10016 36693 10025
rect 37036 10016 37076 10025
rect 36651 9976 36652 10016
rect 36692 9976 36693 10016
rect 36651 9967 36693 9976
rect 36748 9976 37036 10016
rect 36652 9882 36692 9967
rect 36212 9472 36404 9512
rect 36172 9463 36212 9472
rect 35788 8623 35828 8632
rect 35884 9052 36020 9092
rect 35596 8538 35636 8623
rect 35499 8504 35541 8513
rect 35499 8464 35500 8504
rect 35540 8464 35541 8504
rect 35499 8455 35541 8464
rect 35500 8370 35540 8455
rect 35787 8336 35829 8345
rect 35884 8336 35924 9052
rect 36748 9008 36788 9976
rect 37036 9967 37076 9976
rect 37227 10016 37269 10025
rect 37227 9976 37228 10016
rect 37268 9976 37269 10016
rect 37227 9967 37269 9976
rect 36652 8968 36788 9008
rect 35787 8296 35788 8336
rect 35828 8296 35924 8336
rect 35980 8672 36020 8681
rect 35787 8287 35829 8296
rect 35595 8168 35637 8177
rect 35595 8128 35596 8168
rect 35636 8128 35637 8168
rect 35595 8119 35637 8128
rect 35308 7876 35444 7916
rect 35500 8000 35540 8009
rect 35115 7832 35157 7841
rect 35115 7792 35116 7832
rect 35156 7792 35157 7832
rect 35115 7783 35157 7792
rect 35115 7664 35157 7673
rect 35115 7624 35116 7664
rect 35156 7624 35157 7664
rect 35115 7615 35157 7624
rect 35116 7328 35156 7615
rect 35308 7580 35348 7876
rect 35116 7279 35156 7288
rect 35212 7540 35348 7580
rect 35404 7748 35444 7757
rect 35019 7244 35061 7253
rect 35019 7204 35020 7244
rect 35060 7204 35061 7244
rect 35019 7195 35061 7204
rect 35212 7244 35252 7540
rect 35212 7195 35252 7204
rect 34540 6992 34580 7111
rect 34444 6952 34580 6992
rect 34924 6992 34964 7120
rect 35020 7110 35060 7195
rect 35308 7169 35348 7254
rect 35404 7253 35444 7708
rect 35403 7244 35445 7253
rect 35403 7204 35404 7244
rect 35444 7204 35445 7244
rect 35403 7195 35445 7204
rect 35307 7160 35349 7169
rect 35307 7120 35308 7160
rect 35348 7120 35349 7160
rect 35307 7111 35349 7120
rect 35115 7076 35157 7085
rect 35115 7036 35116 7076
rect 35156 7036 35157 7076
rect 35115 7027 35157 7036
rect 34924 6952 35060 6992
rect 34155 6824 34197 6833
rect 34155 6784 34156 6824
rect 34196 6784 34197 6824
rect 34155 6775 34197 6784
rect 34347 6824 34389 6833
rect 34347 6784 34348 6824
rect 34388 6784 34389 6824
rect 34347 6775 34389 6784
rect 34060 6607 34100 6616
rect 34156 6488 34196 6775
rect 33964 6448 34100 6488
rect 33868 6329 33908 6448
rect 33195 6320 33237 6329
rect 33195 6280 33196 6320
rect 33236 6280 33237 6320
rect 33195 6271 33237 6280
rect 33867 6320 33909 6329
rect 33867 6280 33868 6320
rect 33908 6280 33909 6320
rect 34060 6320 34100 6448
rect 34156 6439 34196 6448
rect 34348 6488 34388 6497
rect 34348 6320 34388 6448
rect 34060 6280 34388 6320
rect 33867 6271 33909 6280
rect 33099 6152 33141 6161
rect 33099 6112 33100 6152
rect 33140 6112 33141 6152
rect 33099 6103 33141 6112
rect 33004 5944 33140 5984
rect 32908 5599 32948 5608
rect 33003 5648 33045 5657
rect 33003 5608 33004 5648
rect 33044 5608 33045 5648
rect 33003 5599 33045 5608
rect 33100 5648 33140 5944
rect 33196 5648 33236 6271
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 33483 5816 33525 5825
rect 33483 5776 33484 5816
rect 33524 5776 33525 5816
rect 33483 5767 33525 5776
rect 33292 5648 33332 5657
rect 33196 5608 33292 5648
rect 33100 5599 33140 5608
rect 33292 5599 33332 5608
rect 33484 5648 33524 5767
rect 33484 5599 33524 5608
rect 33004 5514 33044 5599
rect 34348 5564 34388 6280
rect 34444 5648 34484 6952
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 35020 6665 35060 6952
rect 34635 6656 34677 6665
rect 34635 6616 34636 6656
rect 34676 6616 34677 6656
rect 34635 6607 34677 6616
rect 35019 6656 35061 6665
rect 35019 6616 35020 6656
rect 35060 6616 35061 6656
rect 35019 6607 35061 6616
rect 34636 6522 34676 6607
rect 34731 6572 34773 6581
rect 34731 6532 34732 6572
rect 34772 6532 34773 6572
rect 34731 6523 34773 6532
rect 34539 5984 34581 5993
rect 34539 5944 34540 5984
rect 34580 5944 34581 5984
rect 34539 5935 34581 5944
rect 34540 5900 34580 5935
rect 34540 5849 34580 5860
rect 34444 5599 34484 5608
rect 34732 5648 34772 6523
rect 35019 6488 35061 6497
rect 35019 6448 35020 6488
rect 35060 6448 35061 6488
rect 35019 6439 35061 6448
rect 35116 6488 35156 7027
rect 35307 6992 35349 7001
rect 35307 6952 35308 6992
rect 35348 6952 35349 6992
rect 35307 6943 35349 6952
rect 35308 6824 35348 6943
rect 35020 6354 35060 6439
rect 34827 5984 34869 5993
rect 34827 5944 34828 5984
rect 34868 5944 34869 5984
rect 34827 5935 34869 5944
rect 34156 5524 34388 5564
rect 33388 5480 33428 5489
rect 33100 5440 33388 5480
rect 32908 4976 32948 4985
rect 33100 4976 33140 5440
rect 33388 5431 33428 5440
rect 32948 4936 33140 4976
rect 32908 4927 32948 4936
rect 33676 4817 33716 4902
rect 33868 4892 33908 4901
rect 32811 4808 32853 4817
rect 32811 4768 32812 4808
rect 32852 4768 32853 4808
rect 32811 4759 32853 4768
rect 33675 4808 33717 4817
rect 33675 4768 33676 4808
rect 33716 4768 33717 4808
rect 33675 4759 33717 4768
rect 32907 4724 32949 4733
rect 32907 4684 32908 4724
rect 32948 4684 32949 4724
rect 32907 4675 32949 4684
rect 32908 4590 32948 4675
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 33868 4397 33908 4852
rect 33867 4388 33909 4397
rect 33867 4348 33868 4388
rect 33908 4348 33909 4388
rect 33867 4339 33909 4348
rect 32715 4220 32757 4229
rect 32715 4180 32716 4220
rect 32756 4180 32757 4220
rect 32715 4171 32757 4180
rect 32236 4136 32276 4145
rect 32907 4136 32949 4145
rect 32276 4096 32372 4136
rect 32236 4087 32276 4096
rect 32332 3296 32372 4096
rect 32907 4096 32908 4136
rect 32948 4096 32949 4136
rect 32907 4087 32949 4096
rect 33100 4136 33140 4145
rect 32908 3632 32948 4087
rect 32908 3583 32948 3592
rect 32332 3247 32372 3256
rect 32139 3044 32181 3053
rect 32139 3004 32140 3044
rect 32180 3004 32181 3044
rect 32139 2995 32181 3004
rect 32043 2960 32085 2969
rect 32043 2920 32044 2960
rect 32084 2920 32085 2960
rect 32043 2911 32085 2920
rect 32140 2836 32468 2876
rect 32140 2540 32180 2836
rect 32428 2792 32468 2836
rect 32428 2743 32468 2752
rect 32236 2591 32276 2635
rect 33100 2633 33140 4096
rect 33579 3632 33621 3641
rect 33579 3592 33580 3632
rect 33620 3592 33621 3632
rect 33579 3583 33621 3592
rect 34059 3632 34101 3641
rect 34156 3632 34196 5524
rect 34732 5480 34772 5608
rect 34828 5648 34868 5935
rect 34828 5599 34868 5608
rect 34923 5648 34965 5657
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 34924 5514 34964 5599
rect 34444 5440 34772 5480
rect 35019 5480 35061 5489
rect 35019 5440 35020 5480
rect 35060 5440 35061 5480
rect 34444 5144 34484 5440
rect 35019 5431 35061 5440
rect 35020 5346 35060 5431
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 35116 5228 35156 6448
rect 35212 6784 35348 6824
rect 35212 6152 35252 6784
rect 35308 6656 35348 6665
rect 35308 6329 35348 6616
rect 35404 6488 35444 6497
rect 35307 6320 35349 6329
rect 35307 6280 35308 6320
rect 35348 6280 35349 6320
rect 35307 6271 35349 6280
rect 35404 6245 35444 6448
rect 35403 6236 35445 6245
rect 35403 6196 35404 6236
rect 35444 6196 35445 6236
rect 35403 6187 35445 6196
rect 35212 6112 35348 6152
rect 35211 5648 35253 5657
rect 35211 5608 35212 5648
rect 35252 5608 35253 5648
rect 35211 5599 35253 5608
rect 35212 5480 35252 5599
rect 35212 5431 35252 5440
rect 35020 5188 35156 5228
rect 34444 5104 34580 5144
rect 34251 4976 34293 4985
rect 34251 4936 34252 4976
rect 34292 4936 34293 4976
rect 34251 4927 34293 4936
rect 34252 4842 34292 4927
rect 34444 4724 34484 4733
rect 34251 4388 34293 4397
rect 34251 4348 34252 4388
rect 34292 4348 34293 4388
rect 34251 4339 34293 4348
rect 34252 4254 34292 4339
rect 34444 3977 34484 4684
rect 34540 4481 34580 5104
rect 34923 5060 34965 5069
rect 35020 5060 35060 5188
rect 34923 5020 34924 5060
rect 34964 5020 35060 5060
rect 35115 5060 35157 5069
rect 35115 5020 35116 5060
rect 35156 5020 35157 5060
rect 34923 5011 34965 5020
rect 35115 5011 35157 5020
rect 34539 4472 34581 4481
rect 34539 4432 34540 4472
rect 34580 4432 34581 4472
rect 34539 4423 34581 4432
rect 34540 4220 34580 4423
rect 34540 4171 34580 4180
rect 34924 3977 34964 5011
rect 35116 4976 35156 5011
rect 35116 4925 35156 4936
rect 35308 4976 35348 6112
rect 35404 5825 35444 6187
rect 35403 5816 35445 5825
rect 35403 5776 35404 5816
rect 35444 5776 35445 5816
rect 35500 5816 35540 7960
rect 35596 6740 35636 8119
rect 35692 8000 35732 8009
rect 35692 7589 35732 7960
rect 35788 8000 35828 8287
rect 35980 8252 36020 8632
rect 36076 8672 36116 8681
rect 36076 8429 36116 8632
rect 36268 8504 36308 8513
rect 36075 8420 36117 8429
rect 36075 8380 36076 8420
rect 36116 8380 36117 8420
rect 36075 8371 36117 8380
rect 36268 8252 36308 8464
rect 36555 8420 36597 8429
rect 36555 8380 36556 8420
rect 36596 8380 36597 8420
rect 36555 8371 36597 8380
rect 35980 8212 36116 8252
rect 35883 8168 35925 8177
rect 35883 8128 35884 8168
rect 35924 8128 35925 8168
rect 35883 8119 35925 8128
rect 35884 8021 35924 8119
rect 35884 7972 35924 7981
rect 35979 8000 36021 8009
rect 35691 7580 35733 7589
rect 35691 7540 35692 7580
rect 35732 7540 35733 7580
rect 35691 7531 35733 7540
rect 35788 7337 35828 7960
rect 35979 7960 35980 8000
rect 36020 7960 36021 8000
rect 35979 7951 36021 7960
rect 35883 7916 35925 7925
rect 35883 7876 35884 7916
rect 35924 7876 35925 7916
rect 35883 7867 35925 7876
rect 35884 7673 35924 7867
rect 35980 7866 36020 7951
rect 35883 7664 35925 7673
rect 35883 7624 35884 7664
rect 35924 7624 35925 7664
rect 35883 7615 35925 7624
rect 35787 7328 35829 7337
rect 35787 7288 35788 7328
rect 35828 7288 35829 7328
rect 35787 7279 35829 7288
rect 35692 7244 35732 7253
rect 35692 7160 35732 7204
rect 35884 7160 35924 7169
rect 35692 7120 35884 7160
rect 35884 7111 35924 7120
rect 35979 7076 36021 7085
rect 36076 7076 36116 8212
rect 36236 8212 36308 8252
rect 36236 8177 36276 8212
rect 36364 8177 36404 8262
rect 36211 8168 36276 8177
rect 36211 8128 36212 8168
rect 36252 8128 36276 8168
rect 36363 8168 36405 8177
rect 36363 8128 36364 8168
rect 36404 8128 36405 8168
rect 36211 8119 36253 8128
rect 36363 8119 36405 8128
rect 36212 8000 36252 8119
rect 36212 7951 36252 7960
rect 36364 8000 36404 8009
rect 36364 7925 36404 7960
rect 36460 8000 36500 8009
rect 36363 7916 36405 7925
rect 36363 7876 36364 7916
rect 36404 7876 36405 7916
rect 36363 7867 36405 7876
rect 36364 7160 36404 7867
rect 36460 7841 36500 7960
rect 36459 7832 36501 7841
rect 36459 7792 36460 7832
rect 36500 7792 36501 7832
rect 36459 7783 36501 7792
rect 36556 7757 36596 8371
rect 36652 8000 36692 8968
rect 36940 8009 36980 8094
rect 36652 7951 36692 7960
rect 36748 8000 36788 8009
rect 36555 7748 36597 7757
rect 36555 7708 36556 7748
rect 36596 7708 36597 7748
rect 36555 7699 36597 7708
rect 35979 7036 35980 7076
rect 36020 7036 36116 7076
rect 36172 7120 36404 7160
rect 35979 7027 36021 7036
rect 35980 6833 36020 7027
rect 35979 6824 36021 6833
rect 35979 6784 35980 6824
rect 36020 6784 36021 6824
rect 35979 6775 36021 6784
rect 35596 6700 35732 6740
rect 35595 6572 35637 6581
rect 35595 6532 35596 6572
rect 35636 6532 35637 6572
rect 35595 6523 35637 6532
rect 35596 6438 35636 6523
rect 35692 5993 35732 6700
rect 35787 6572 35829 6581
rect 35787 6532 35788 6572
rect 35828 6532 35829 6572
rect 35787 6523 35829 6532
rect 35788 6488 35828 6523
rect 35788 6437 35828 6448
rect 35883 6488 35925 6497
rect 35883 6448 35884 6488
rect 35924 6448 35925 6488
rect 35883 6439 35925 6448
rect 35884 6354 35924 6439
rect 35787 6320 35829 6329
rect 35787 6280 35788 6320
rect 35828 6280 35829 6320
rect 35787 6271 35829 6280
rect 35691 5984 35733 5993
rect 35691 5944 35692 5984
rect 35732 5944 35733 5984
rect 35691 5935 35733 5944
rect 35500 5776 35732 5816
rect 35403 5767 35445 5776
rect 35403 5648 35445 5657
rect 35403 5608 35404 5648
rect 35444 5608 35445 5648
rect 35403 5599 35445 5608
rect 35500 5648 35540 5659
rect 35404 5514 35444 5599
rect 35500 5573 35540 5608
rect 35499 5564 35541 5573
rect 35499 5524 35500 5564
rect 35540 5524 35541 5564
rect 35499 5515 35541 5524
rect 35308 4927 35348 4936
rect 35308 4136 35348 4145
rect 35020 4096 35308 4136
rect 34252 3968 34292 3977
rect 34443 3968 34485 3977
rect 34292 3928 34388 3968
rect 34252 3919 34292 3928
rect 34059 3592 34060 3632
rect 34100 3592 34196 3632
rect 34059 3583 34101 3592
rect 33580 3464 33620 3583
rect 33580 3415 33620 3424
rect 33772 3296 33812 3305
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 33291 2876 33333 2885
rect 33291 2836 33292 2876
rect 33332 2836 33333 2876
rect 33291 2827 33333 2836
rect 32811 2624 32853 2633
rect 32811 2584 32812 2624
rect 32852 2584 32853 2624
rect 32811 2575 32853 2584
rect 33099 2624 33141 2633
rect 33099 2584 33100 2624
rect 33140 2584 33141 2624
rect 33099 2575 33141 2584
rect 33292 2624 33332 2827
rect 33292 2575 33332 2584
rect 33676 2624 33716 2633
rect 33772 2624 33812 3256
rect 33716 2584 33812 2624
rect 33676 2575 33716 2584
rect 32236 2549 32276 2551
rect 31604 1912 31700 1952
rect 31948 2500 32180 2540
rect 32235 2540 32277 2549
rect 32235 2500 32236 2540
rect 32276 2500 32277 2540
rect 31948 1952 31988 2500
rect 32235 2491 32277 2500
rect 32812 1961 32852 2575
rect 31564 1903 31604 1912
rect 31948 1903 31988 1912
rect 32811 1952 32853 1961
rect 32811 1912 32812 1952
rect 32852 1912 32853 1952
rect 32811 1903 32853 1912
rect 34060 1952 34100 3583
rect 34348 3464 34388 3928
rect 34443 3928 34444 3968
rect 34484 3928 34485 3968
rect 34443 3919 34485 3928
rect 34923 3968 34965 3977
rect 34923 3928 34924 3968
rect 34964 3928 34965 3968
rect 34923 3919 34965 3928
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 35020 3632 35060 4096
rect 35308 4087 35348 4096
rect 35307 3968 35349 3977
rect 35307 3928 35308 3968
rect 35348 3928 35349 3968
rect 35307 3919 35349 3928
rect 35020 3583 35060 3592
rect 35308 3548 35348 3919
rect 35308 3499 35348 3508
rect 34348 3415 34388 3424
rect 35692 2876 35732 5776
rect 35788 5732 35828 6271
rect 35788 5683 35828 5692
rect 35980 5657 36020 6775
rect 36076 6665 36116 6750
rect 36075 6656 36117 6665
rect 36075 6616 36076 6656
rect 36116 6616 36117 6656
rect 36075 6607 36117 6616
rect 36076 6488 36116 6497
rect 36076 6329 36116 6448
rect 36075 6320 36117 6329
rect 36075 6280 36076 6320
rect 36116 6280 36117 6320
rect 36075 6271 36117 6280
rect 35979 5648 36021 5657
rect 35979 5608 35980 5648
rect 36020 5608 36021 5648
rect 35979 5599 36021 5608
rect 36172 5489 36212 7120
rect 36267 6992 36309 7001
rect 36267 6952 36268 6992
rect 36308 6952 36309 6992
rect 36267 6943 36309 6952
rect 36364 6992 36404 7001
rect 36404 6952 36500 6992
rect 36364 6943 36404 6952
rect 36268 6488 36308 6943
rect 36268 6439 36308 6448
rect 36363 5816 36405 5825
rect 36363 5776 36364 5816
rect 36404 5776 36405 5816
rect 36363 5767 36405 5776
rect 36364 5682 36404 5767
rect 36171 5480 36213 5489
rect 36171 5440 36172 5480
rect 36212 5440 36213 5480
rect 36171 5431 36213 5440
rect 36363 4976 36405 4985
rect 36363 4936 36364 4976
rect 36404 4936 36405 4976
rect 36363 4927 36405 4936
rect 36460 4976 36500 6952
rect 36748 6917 36788 7960
rect 36939 8000 36981 8009
rect 36939 7960 36940 8000
rect 36980 7960 36981 8000
rect 36939 7951 36981 7960
rect 37036 8000 37076 8011
rect 37036 7925 37076 7960
rect 37228 8000 37268 9967
rect 37324 9680 37364 9689
rect 37420 9680 37460 10135
rect 37364 9640 37460 9680
rect 37324 9631 37364 9640
rect 37420 9512 37460 9521
rect 37612 9512 37652 10396
rect 37707 10387 37749 10396
rect 37707 10268 37749 10277
rect 37707 10228 37708 10268
rect 37748 10228 37749 10268
rect 37707 10219 37749 10228
rect 37708 10134 37748 10219
rect 37804 10184 37844 11068
rect 37900 11024 37940 11647
rect 38092 11528 38132 11537
rect 37995 11108 38037 11117
rect 37995 11068 37996 11108
rect 38036 11068 38037 11108
rect 37995 11059 38037 11068
rect 37900 10975 37940 10984
rect 37996 11024 38036 11059
rect 37996 10973 38036 10984
rect 37804 10135 37844 10144
rect 37996 10184 38036 10193
rect 37460 9472 37652 9512
rect 37420 9463 37460 9472
rect 37803 9428 37845 9437
rect 37803 9388 37804 9428
rect 37844 9388 37845 9428
rect 37803 9379 37845 9388
rect 37228 7951 37268 7960
rect 37612 8672 37652 8681
rect 37035 7916 37077 7925
rect 37035 7876 37036 7916
rect 37076 7876 37077 7916
rect 37035 7867 37077 7876
rect 36939 7832 36981 7841
rect 36939 7792 36940 7832
rect 36980 7792 36981 7832
rect 36939 7783 36981 7792
rect 36940 7698 36980 7783
rect 37516 7748 37556 7757
rect 37323 7412 37365 7421
rect 37323 7372 37324 7412
rect 37364 7372 37365 7412
rect 37323 7363 37365 7372
rect 36843 7160 36885 7169
rect 36843 7120 36844 7160
rect 36884 7120 36885 7160
rect 36843 7111 36885 7120
rect 37324 7160 37364 7363
rect 37419 7328 37461 7337
rect 37419 7288 37420 7328
rect 37460 7288 37461 7328
rect 37419 7279 37461 7288
rect 37324 7111 37364 7120
rect 37420 7160 37460 7279
rect 37420 7111 37460 7120
rect 36844 7026 36884 7111
rect 36747 6908 36789 6917
rect 36747 6868 36748 6908
rect 36788 6868 36789 6908
rect 36747 6859 36789 6868
rect 36747 6656 36789 6665
rect 36747 6616 36748 6656
rect 36788 6616 36789 6656
rect 36747 6607 36789 6616
rect 36652 5648 36692 5659
rect 36652 5573 36692 5608
rect 36651 5564 36693 5573
rect 36651 5524 36652 5564
rect 36692 5524 36693 5564
rect 36651 5515 36693 5524
rect 36556 4976 36596 4985
rect 36460 4936 36556 4976
rect 35883 4136 35925 4145
rect 35883 4096 35884 4136
rect 35924 4096 35925 4136
rect 35883 4087 35925 4096
rect 36268 4136 36308 4145
rect 35884 4002 35924 4087
rect 36268 3977 36308 4096
rect 36364 4052 36404 4927
rect 36364 4003 36404 4012
rect 36267 3968 36309 3977
rect 36267 3928 36268 3968
rect 36308 3928 36309 3968
rect 36267 3919 36309 3928
rect 36171 3464 36213 3473
rect 36171 3424 36172 3464
rect 36212 3424 36213 3464
rect 36171 3415 36213 3424
rect 36172 3330 36212 3415
rect 35732 2836 36020 2876
rect 35692 2827 35732 2836
rect 34540 2633 34580 2718
rect 34539 2624 34581 2633
rect 34539 2584 34540 2624
rect 34580 2584 34581 2624
rect 34539 2575 34581 2584
rect 35980 2624 36020 2836
rect 36460 2633 36500 4936
rect 36556 4927 36596 4936
rect 36651 4136 36693 4145
rect 36651 4096 36652 4136
rect 36692 4096 36693 4136
rect 36651 4087 36693 4096
rect 36652 4002 36692 4087
rect 36651 3464 36693 3473
rect 36651 3424 36652 3464
rect 36692 3424 36693 3464
rect 36651 3415 36693 3424
rect 36652 2876 36692 3415
rect 36652 2827 36692 2836
rect 35980 2575 36020 2584
rect 36459 2624 36501 2633
rect 36459 2584 36460 2624
rect 36500 2584 36501 2624
rect 36748 2624 36788 6607
rect 37516 6581 37556 7708
rect 37612 7412 37652 8632
rect 37804 8420 37844 9379
rect 37996 9353 38036 10144
rect 37995 9344 38037 9353
rect 37995 9304 37996 9344
rect 38036 9304 38037 9344
rect 37995 9295 38037 9304
rect 37900 8849 37940 8934
rect 37899 8840 37941 8849
rect 37899 8800 37900 8840
rect 37940 8800 37941 8840
rect 37899 8791 37941 8800
rect 37900 8672 37940 8681
rect 38092 8672 38132 11488
rect 38188 11024 38228 12235
rect 38188 10975 38228 10984
rect 38379 11024 38421 11033
rect 38379 10984 38380 11024
rect 38420 10984 38421 11024
rect 38379 10975 38421 10984
rect 38476 11024 38516 12664
rect 38572 11696 38612 14083
rect 38859 14048 38901 14057
rect 38859 14008 38860 14048
rect 38900 14008 38901 14048
rect 38859 13999 38901 14008
rect 38667 13964 38709 13973
rect 38667 13924 38668 13964
rect 38708 13924 38709 13964
rect 38667 13915 38709 13924
rect 38668 13040 38708 13915
rect 38860 13914 38900 13999
rect 38764 13208 38804 13217
rect 38804 13168 38900 13208
rect 38764 13159 38804 13168
rect 38668 13000 38804 13040
rect 38667 12620 38709 12629
rect 38667 12580 38668 12620
rect 38708 12580 38709 12620
rect 38667 12571 38709 12580
rect 38668 12536 38708 12571
rect 38764 12545 38804 13000
rect 38860 12629 38900 13168
rect 38956 12713 38996 14839
rect 39724 14720 39764 14839
rect 39724 14393 39764 14680
rect 39723 14384 39765 14393
rect 39723 14344 39724 14384
rect 39764 14344 39765 14384
rect 39723 14335 39765 14344
rect 39627 14048 39669 14057
rect 39627 14008 39628 14048
rect 39668 14008 39669 14048
rect 39627 13999 39669 14008
rect 39532 13880 39572 13889
rect 39051 13796 39093 13805
rect 39051 13756 39052 13796
rect 39092 13756 39093 13796
rect 39051 13747 39093 13756
rect 39052 13208 39092 13747
rect 39052 13159 39092 13168
rect 39436 13208 39476 13217
rect 39532 13208 39572 13840
rect 39476 13168 39572 13208
rect 39436 13159 39476 13168
rect 38955 12704 38997 12713
rect 38955 12664 38956 12704
rect 38996 12664 38997 12704
rect 38955 12655 38997 12664
rect 38859 12620 38901 12629
rect 38859 12580 38860 12620
rect 38900 12580 38901 12620
rect 38859 12571 38901 12580
rect 38668 12485 38708 12496
rect 38763 12536 38805 12545
rect 38763 12496 38764 12536
rect 38804 12496 38805 12536
rect 38763 12487 38805 12496
rect 38956 12536 38996 12655
rect 38956 12487 38996 12496
rect 39243 12536 39285 12545
rect 39243 12496 39244 12536
rect 39284 12496 39285 12536
rect 39243 12487 39285 12496
rect 39628 12536 39668 13999
rect 39628 12487 39668 12496
rect 40300 13208 40340 17023
rect 42604 16820 42644 16829
rect 41644 16316 41684 16325
rect 40492 16232 40532 16241
rect 41644 16232 41684 16276
rect 41836 16232 41876 16241
rect 41644 16192 41836 16232
rect 40492 14729 40532 16192
rect 41836 16183 41876 16192
rect 42508 16064 42548 16073
rect 41932 16024 42508 16064
rect 40972 15560 41012 15569
rect 40972 14897 41012 15520
rect 41643 15560 41685 15569
rect 41643 15520 41644 15560
rect 41684 15520 41685 15560
rect 41643 15511 41685 15520
rect 41932 15560 41972 16024
rect 42508 16015 42548 16024
rect 42604 15569 42644 16780
rect 41932 15511 41972 15520
rect 42603 15560 42645 15569
rect 42603 15520 42604 15560
rect 42644 15520 42645 15560
rect 42603 15511 42645 15520
rect 43947 15560 43989 15569
rect 43947 15520 43948 15560
rect 43988 15520 43989 15560
rect 43947 15511 43989 15520
rect 40971 14888 41013 14897
rect 40971 14848 40972 14888
rect 41012 14848 41013 14888
rect 40971 14839 41013 14848
rect 41356 14888 41396 14897
rect 41259 14804 41301 14813
rect 41259 14764 41260 14804
rect 41300 14764 41301 14804
rect 41259 14755 41301 14764
rect 40491 14720 40533 14729
rect 40491 14680 40492 14720
rect 40532 14680 40533 14720
rect 40491 14671 40533 14680
rect 40972 14720 41012 14729
rect 40683 14552 40725 14561
rect 40683 14512 40684 14552
rect 40724 14512 40725 14552
rect 40683 14503 40725 14512
rect 40875 14552 40917 14561
rect 40875 14508 40876 14552
rect 40916 14508 40917 14552
rect 40875 14503 40917 14508
rect 40684 14048 40724 14503
rect 40876 14417 40916 14503
rect 40684 13999 40724 14008
rect 40972 13973 41012 14680
rect 41068 14720 41108 14729
rect 41068 14225 41108 14680
rect 41067 14216 41109 14225
rect 41067 14176 41068 14216
rect 41108 14176 41109 14216
rect 41067 14167 41109 14176
rect 40971 13964 41013 13973
rect 40971 13924 40972 13964
rect 41012 13924 41013 13964
rect 40971 13915 41013 13924
rect 38764 12402 38804 12487
rect 39244 12293 39284 12487
rect 39435 12368 39477 12377
rect 39435 12328 39436 12368
rect 39476 12328 39477 12368
rect 39435 12319 39477 12328
rect 38955 12284 38997 12293
rect 38955 12244 38956 12284
rect 38996 12244 38997 12284
rect 38955 12235 38997 12244
rect 39243 12284 39285 12293
rect 39243 12244 39244 12284
rect 39284 12244 39285 12284
rect 39243 12235 39285 12244
rect 38956 12150 38996 12235
rect 39436 11705 39476 12319
rect 40204 12284 40244 12293
rect 40300 12284 40340 13168
rect 40683 12620 40725 12629
rect 40683 12580 40684 12620
rect 40724 12580 40725 12620
rect 40683 12571 40725 12580
rect 40684 12486 40724 12571
rect 40395 12452 40437 12461
rect 40395 12412 40396 12452
rect 40436 12412 40437 12452
rect 40395 12403 40437 12412
rect 40244 12244 40340 12284
rect 40204 12235 40244 12244
rect 40300 11705 40340 12244
rect 38572 11647 38612 11656
rect 38763 11696 38805 11705
rect 38763 11656 38764 11696
rect 38804 11656 38805 11696
rect 38763 11647 38805 11656
rect 39244 11696 39284 11705
rect 38571 11108 38613 11117
rect 38571 11068 38572 11108
rect 38612 11068 38708 11108
rect 38571 11059 38613 11068
rect 38476 10975 38516 10984
rect 38668 11024 38708 11068
rect 38380 10890 38420 10975
rect 38187 10772 38229 10781
rect 38187 10732 38188 10772
rect 38228 10732 38229 10772
rect 38187 10723 38229 10732
rect 38188 10638 38228 10723
rect 38187 10520 38229 10529
rect 38187 10480 38188 10520
rect 38228 10480 38229 10520
rect 38187 10471 38229 10480
rect 38188 10193 38228 10471
rect 38668 10268 38708 10984
rect 38764 11024 38804 11647
rect 38955 11192 38997 11201
rect 38955 11152 38956 11192
rect 38996 11152 38997 11192
rect 38955 11143 38997 11152
rect 38764 10975 38804 10984
rect 38956 11024 38996 11143
rect 38956 10975 38996 10984
rect 38764 10772 38804 10783
rect 39148 10772 39188 10781
rect 38764 10697 38804 10732
rect 38860 10732 39148 10772
rect 38763 10688 38805 10697
rect 38763 10648 38764 10688
rect 38804 10648 38805 10688
rect 38763 10639 38805 10648
rect 38668 10228 38804 10268
rect 38187 10184 38229 10193
rect 38187 10144 38188 10184
rect 38228 10144 38229 10184
rect 38187 10135 38229 10144
rect 38188 9512 38228 10135
rect 38667 10100 38709 10109
rect 38667 10060 38668 10100
rect 38708 10060 38709 10100
rect 38667 10051 38709 10060
rect 38668 9966 38708 10051
rect 38188 9463 38228 9472
rect 38284 9512 38324 9521
rect 38476 9512 38516 9521
rect 38324 9472 38476 9512
rect 38284 9463 38324 9472
rect 38476 9463 38516 9472
rect 38571 9428 38613 9437
rect 38571 9388 38572 9428
rect 38612 9388 38613 9428
rect 38571 9379 38613 9388
rect 38764 9428 38804 10228
rect 38860 9512 38900 10732
rect 39148 10723 39188 10732
rect 39147 10436 39189 10445
rect 39147 10396 39148 10436
rect 39188 10396 39189 10436
rect 39147 10387 39189 10396
rect 39148 10302 39188 10387
rect 39051 10100 39093 10109
rect 39051 10060 39052 10100
rect 39092 10060 39093 10100
rect 39051 10051 39093 10060
rect 38860 9463 38900 9472
rect 39052 9512 39092 10051
rect 39052 9463 39092 9472
rect 39244 9437 39284 11656
rect 39435 11696 39477 11705
rect 39435 11656 39436 11696
rect 39476 11656 39477 11696
rect 39435 11647 39477 11656
rect 39532 11696 39572 11705
rect 40299 11696 40341 11705
rect 39572 11656 39668 11696
rect 39532 11647 39572 11656
rect 39436 11562 39476 11647
rect 39532 11528 39572 11537
rect 39532 11201 39572 11488
rect 39531 11192 39573 11201
rect 39531 11152 39532 11192
rect 39572 11152 39573 11192
rect 39531 11143 39573 11152
rect 39628 10193 39668 11656
rect 40299 11656 40300 11696
rect 40340 11656 40341 11696
rect 40299 11647 40341 11656
rect 40396 11696 40436 12403
rect 40396 11647 40436 11656
rect 40492 11696 40532 11707
rect 39723 11612 39765 11621
rect 39723 11572 39724 11612
rect 39764 11572 39765 11612
rect 39723 11563 39765 11572
rect 39627 10184 39669 10193
rect 39627 10144 39628 10184
rect 39668 10144 39669 10184
rect 39627 10135 39669 10144
rect 39436 9512 39476 9521
rect 38572 9294 38612 9379
rect 38667 9344 38709 9353
rect 38667 9304 38668 9344
rect 38708 9304 38709 9344
rect 38667 9295 38709 9304
rect 38668 9210 38708 9295
rect 38764 8840 38804 9388
rect 39243 9428 39285 9437
rect 39243 9388 39244 9428
rect 39284 9388 39285 9428
rect 39243 9379 39285 9388
rect 38955 8840 38997 8849
rect 38764 8800 38900 8840
rect 38764 8672 38804 8681
rect 38092 8632 38228 8672
rect 37900 8504 37940 8632
rect 38092 8504 38132 8513
rect 37900 8464 38092 8504
rect 38092 8455 38132 8464
rect 37804 8380 38036 8420
rect 37804 8168 37844 8177
rect 37612 7363 37652 7372
rect 37708 8000 37748 8009
rect 37610 7244 37652 7253
rect 37610 7204 37611 7244
rect 37651 7204 37652 7244
rect 37610 7195 37652 7204
rect 37612 7160 37652 7195
rect 37708 7160 37748 7960
rect 37804 7589 37844 8128
rect 37899 8000 37941 8009
rect 37899 7960 37900 8000
rect 37940 7960 37941 8000
rect 37899 7951 37941 7960
rect 37996 8000 38036 8380
rect 37803 7580 37845 7589
rect 37803 7540 37804 7580
rect 37844 7540 37845 7580
rect 37803 7531 37845 7540
rect 37900 7253 37940 7951
rect 37996 7421 38036 7960
rect 38092 8000 38132 8009
rect 38092 7589 38132 7960
rect 38091 7580 38133 7589
rect 38091 7540 38092 7580
rect 38132 7540 38133 7580
rect 38091 7531 38133 7540
rect 37995 7412 38037 7421
rect 37995 7372 37996 7412
rect 38036 7372 38037 7412
rect 37995 7363 38037 7372
rect 37899 7244 37941 7253
rect 37899 7204 37900 7244
rect 37940 7204 37941 7244
rect 37899 7195 37941 7204
rect 37804 7160 37844 7169
rect 37708 7120 37804 7160
rect 37612 7111 37652 7120
rect 37611 6992 37653 7001
rect 37611 6952 37612 6992
rect 37652 6952 37653 6992
rect 37611 6943 37653 6952
rect 37612 6858 37652 6943
rect 37323 6572 37365 6581
rect 37323 6532 37324 6572
rect 37364 6532 37365 6572
rect 37323 6523 37365 6532
rect 37515 6572 37557 6581
rect 37515 6532 37516 6572
rect 37556 6532 37557 6572
rect 37515 6523 37557 6532
rect 36843 6488 36885 6497
rect 37132 6488 37172 6497
rect 36843 6448 36844 6488
rect 36884 6448 36885 6488
rect 36843 6439 36885 6448
rect 36940 6448 37132 6488
rect 36844 5480 36884 6439
rect 36940 6245 36980 6448
rect 37132 6439 37172 6448
rect 36939 6236 36981 6245
rect 37228 6236 37268 6245
rect 36939 6196 36940 6236
rect 36980 6196 36981 6236
rect 36939 6187 36981 6196
rect 37036 6196 37228 6236
rect 36940 6102 36980 6187
rect 37036 5900 37076 6196
rect 37228 6187 37268 6196
rect 37324 5984 37364 6523
rect 37611 6488 37653 6497
rect 37708 6488 37748 6497
rect 37611 6448 37612 6488
rect 37652 6448 37708 6488
rect 37611 6439 37653 6448
rect 37708 6439 37748 6448
rect 37804 6488 37844 7120
rect 37900 6992 37940 7195
rect 37996 7160 38036 7363
rect 38091 7244 38133 7253
rect 38091 7204 38092 7244
rect 38132 7204 38133 7244
rect 38091 7195 38133 7204
rect 37996 7111 38036 7120
rect 38092 7160 38132 7195
rect 38188 7169 38228 8632
rect 38380 8632 38764 8672
rect 38283 8504 38325 8513
rect 38283 8464 38284 8504
rect 38324 8464 38325 8504
rect 38283 8455 38325 8464
rect 38284 8009 38324 8455
rect 38283 8000 38325 8009
rect 38283 7960 38284 8000
rect 38324 7960 38325 8000
rect 38283 7951 38325 7960
rect 38284 7832 38324 7841
rect 38380 7832 38420 8632
rect 38764 8623 38804 8632
rect 38860 8504 38900 8800
rect 38955 8800 38956 8840
rect 38996 8800 38997 8840
rect 38955 8791 38997 8800
rect 38956 8672 38996 8791
rect 38956 8623 38996 8632
rect 38324 7792 38420 7832
rect 38572 8464 38900 8504
rect 38572 8000 38612 8464
rect 38955 8336 38997 8345
rect 38955 8296 38956 8336
rect 38996 8296 38997 8336
rect 38955 8287 38997 8296
rect 38763 8252 38805 8261
rect 38763 8212 38764 8252
rect 38804 8212 38805 8252
rect 38763 8203 38805 8212
rect 38284 7783 38324 7792
rect 38572 7589 38612 7960
rect 38764 8000 38804 8203
rect 38571 7580 38613 7589
rect 38571 7540 38572 7580
rect 38612 7540 38613 7580
rect 38571 7531 38613 7540
rect 38092 7109 38132 7120
rect 38187 7160 38229 7169
rect 38187 7120 38188 7160
rect 38228 7120 38229 7160
rect 38187 7111 38229 7120
rect 38476 7160 38516 7169
rect 38092 6992 38132 7001
rect 37900 6952 38092 6992
rect 38092 6943 38132 6952
rect 37899 6740 37941 6749
rect 37899 6700 37900 6740
rect 37940 6700 37941 6740
rect 37899 6691 37941 6700
rect 37804 6413 37844 6448
rect 37900 6488 37940 6691
rect 37803 6404 37845 6413
rect 37803 6364 37804 6404
rect 37844 6364 37845 6404
rect 37803 6355 37845 6364
rect 37516 6236 37556 6245
rect 37556 6196 37748 6236
rect 37516 6187 37556 6196
rect 36940 5860 37076 5900
rect 37228 5944 37364 5984
rect 36940 5648 36980 5860
rect 37132 5816 37172 5825
rect 36940 5599 36980 5608
rect 37036 5732 37076 5741
rect 37036 5480 37076 5692
rect 37132 5657 37172 5776
rect 37228 5732 37268 5944
rect 37228 5683 37268 5692
rect 37131 5648 37173 5657
rect 37131 5608 37132 5648
rect 37172 5608 37173 5648
rect 37131 5599 37173 5608
rect 37324 5648 37364 5657
rect 36844 5440 37076 5480
rect 37227 4304 37269 4313
rect 37227 4264 37228 4304
rect 37268 4264 37269 4304
rect 37324 4304 37364 5608
rect 37611 5648 37653 5657
rect 37611 5608 37612 5648
rect 37652 5608 37653 5648
rect 37611 5599 37653 5608
rect 37612 5514 37652 5599
rect 37419 5060 37461 5069
rect 37419 5020 37420 5060
rect 37460 5020 37461 5060
rect 37419 5011 37461 5020
rect 37420 4976 37460 5011
rect 37420 4925 37460 4936
rect 37708 4808 37748 6196
rect 37804 5312 37844 6355
rect 37900 6245 37940 6448
rect 37996 6488 38036 6497
rect 37996 6320 38036 6448
rect 38284 6488 38324 6497
rect 38284 6320 38324 6448
rect 37996 6280 38132 6320
rect 38284 6280 38420 6320
rect 37899 6236 37941 6245
rect 37899 6196 37900 6236
rect 37940 6196 37941 6236
rect 37899 6187 37941 6196
rect 37900 5396 37940 6187
rect 38092 5648 38132 6280
rect 38380 5825 38420 6280
rect 38379 5816 38421 5825
rect 38379 5776 38380 5816
rect 38420 5776 38421 5816
rect 38379 5767 38421 5776
rect 38092 5608 38228 5648
rect 38188 5405 38228 5608
rect 38380 5564 38420 5767
rect 38476 5741 38516 7120
rect 38572 6749 38612 7531
rect 38764 7337 38804 7960
rect 38956 8000 38996 8287
rect 39436 8177 39476 9472
rect 39724 8672 39764 11563
rect 40011 11192 40053 11201
rect 40011 11152 40012 11192
rect 40052 11152 40053 11192
rect 40011 11143 40053 11152
rect 40012 11058 40052 11143
rect 39820 11024 39860 11033
rect 39820 10697 39860 10984
rect 40203 11024 40245 11033
rect 40203 10984 40204 11024
rect 40244 10984 40245 11024
rect 40203 10975 40245 10984
rect 40012 10772 40052 10781
rect 39819 10688 39861 10697
rect 39819 10648 39820 10688
rect 39860 10648 39861 10688
rect 39819 10639 39861 10648
rect 39820 10184 39860 10193
rect 40012 10184 40052 10732
rect 40204 10436 40244 10975
rect 40204 10387 40244 10396
rect 39860 10144 40052 10184
rect 39820 10135 39860 10144
rect 40300 9512 40340 11647
rect 40492 11621 40532 11656
rect 41260 11696 41300 14755
rect 41356 14057 41396 14848
rect 41355 14048 41397 14057
rect 41355 14008 41356 14048
rect 41396 14008 41397 14048
rect 41355 13999 41397 14008
rect 41548 14048 41588 14057
rect 41452 13208 41492 13217
rect 41452 12965 41492 13168
rect 41451 12956 41493 12965
rect 41356 12916 41452 12956
rect 41492 12916 41493 12956
rect 41356 12536 41396 12916
rect 41451 12907 41493 12916
rect 41356 12487 41396 12496
rect 41451 12536 41493 12545
rect 41451 12496 41452 12536
rect 41492 12496 41493 12536
rect 41451 12487 41493 12496
rect 41260 11647 41300 11656
rect 40491 11612 40533 11621
rect 40491 11572 40492 11612
rect 40532 11572 40533 11612
rect 40491 11563 40533 11572
rect 40876 11612 40916 11621
rect 40683 11528 40725 11537
rect 40683 11488 40684 11528
rect 40724 11488 40725 11528
rect 40683 11479 40725 11488
rect 40684 11394 40724 11479
rect 40876 11192 40916 11572
rect 40876 11143 40916 11152
rect 40683 11024 40725 11033
rect 40683 10984 40684 11024
rect 40724 10984 40725 11024
rect 40683 10975 40725 10984
rect 40684 10890 40724 10975
rect 41356 10184 41396 10193
rect 41260 10144 41356 10184
rect 41067 9932 41109 9941
rect 41067 9892 41068 9932
rect 41108 9892 41109 9932
rect 41067 9883 41109 9892
rect 40300 9463 40340 9472
rect 41068 8840 41108 9883
rect 41068 8791 41108 8800
rect 41163 8840 41205 8849
rect 41163 8800 41164 8840
rect 41204 8800 41205 8840
rect 41163 8791 41205 8800
rect 39820 8672 39860 8681
rect 39724 8632 39820 8672
rect 39820 8623 39860 8632
rect 40011 8672 40053 8681
rect 40011 8632 40012 8672
rect 40052 8632 40053 8672
rect 40011 8623 40053 8632
rect 40876 8672 40916 8681
rect 40012 8538 40052 8623
rect 39628 8504 39668 8513
rect 39435 8168 39477 8177
rect 39435 8128 39436 8168
rect 39476 8128 39572 8168
rect 39435 8119 39477 8128
rect 38956 7951 38996 7960
rect 38763 7328 38805 7337
rect 38763 7288 38764 7328
rect 38804 7288 38805 7328
rect 38763 7279 38805 7288
rect 38667 7244 38709 7253
rect 38667 7204 38668 7244
rect 38708 7204 38709 7244
rect 38667 7195 38709 7204
rect 38571 6740 38613 6749
rect 38571 6700 38572 6740
rect 38612 6700 38613 6740
rect 38571 6691 38613 6700
rect 38572 6497 38612 6582
rect 38571 6488 38613 6497
rect 38571 6448 38572 6488
rect 38612 6448 38613 6488
rect 38571 6439 38613 6448
rect 38668 6320 38708 7195
rect 39435 7160 39477 7169
rect 39435 7120 39436 7160
rect 39476 7120 39477 7160
rect 39435 7111 39477 7120
rect 39436 7026 39476 7111
rect 39148 6992 39188 7001
rect 38572 6280 38708 6320
rect 38764 6572 38804 6581
rect 38475 5732 38517 5741
rect 38475 5692 38476 5732
rect 38516 5692 38517 5732
rect 38475 5683 38517 5692
rect 38572 5648 38612 6280
rect 38572 5599 38612 5608
rect 38667 5648 38709 5657
rect 38667 5608 38668 5648
rect 38708 5608 38709 5648
rect 38667 5599 38709 5608
rect 38380 5524 38516 5564
rect 38284 5480 38324 5489
rect 38187 5396 38229 5405
rect 37900 5356 38036 5396
rect 37804 5272 37940 5312
rect 37803 5144 37845 5153
rect 37803 5104 37804 5144
rect 37844 5104 37845 5144
rect 37803 5095 37845 5104
rect 37804 4976 37844 5095
rect 37804 4927 37844 4936
rect 37708 4768 37844 4808
rect 37324 4264 37460 4304
rect 37227 4255 37269 4264
rect 37228 4136 37268 4255
rect 37324 4136 37364 4145
rect 37228 4096 37324 4136
rect 37228 3464 37268 4096
rect 37324 4087 37364 4096
rect 37228 3415 37268 3424
rect 37420 2885 37460 4264
rect 37516 4136 37556 4145
rect 37556 4096 37748 4136
rect 37516 4087 37556 4096
rect 37611 3800 37653 3809
rect 37611 3760 37612 3800
rect 37652 3760 37653 3800
rect 37611 3751 37653 3760
rect 37419 2876 37461 2885
rect 37419 2836 37420 2876
rect 37460 2836 37461 2876
rect 37419 2827 37461 2836
rect 37516 2624 37556 2633
rect 36748 2584 37516 2624
rect 36459 2575 36501 2584
rect 37516 2575 37556 2584
rect 37612 2624 37652 3751
rect 37612 2575 37652 2584
rect 37708 2540 37748 4096
rect 37804 4061 37844 4768
rect 37803 4052 37845 4061
rect 37803 4012 37804 4052
rect 37844 4012 37845 4052
rect 37803 4003 37845 4012
rect 37804 2624 37844 4003
rect 37900 3893 37940 5272
rect 37899 3884 37941 3893
rect 37899 3844 37900 3884
rect 37940 3844 37941 3884
rect 37899 3835 37941 3844
rect 37996 3548 38036 5356
rect 38187 5356 38188 5396
rect 38228 5356 38229 5396
rect 38187 5347 38229 5356
rect 38188 4976 38228 5347
rect 38284 5153 38324 5440
rect 38283 5144 38325 5153
rect 38283 5104 38284 5144
rect 38324 5104 38325 5144
rect 38283 5095 38325 5104
rect 38188 4927 38228 4936
rect 38379 4976 38421 4985
rect 38379 4936 38380 4976
rect 38420 4936 38421 4976
rect 38379 4927 38421 4936
rect 38380 4842 38420 4927
rect 38092 4724 38132 4733
rect 38092 3809 38132 4684
rect 38188 4136 38228 4145
rect 38380 4136 38420 4145
rect 38228 4096 38380 4136
rect 38188 4087 38228 4096
rect 38380 4087 38420 4096
rect 38379 3968 38421 3977
rect 38379 3928 38380 3968
rect 38420 3928 38421 3968
rect 38379 3919 38421 3928
rect 38283 3884 38325 3893
rect 38283 3844 38284 3884
rect 38324 3844 38325 3884
rect 38283 3835 38325 3844
rect 38091 3800 38133 3809
rect 38091 3760 38092 3800
rect 38132 3760 38133 3800
rect 38091 3751 38133 3760
rect 37996 3508 38132 3548
rect 37996 2885 38036 2970
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 37804 2575 37844 2584
rect 37995 2624 38037 2633
rect 37995 2584 37996 2624
rect 38036 2584 38037 2624
rect 38092 2624 38132 3508
rect 38188 2624 38228 2633
rect 38092 2584 38188 2624
rect 37995 2575 38037 2584
rect 38188 2575 38228 2584
rect 38284 2624 38324 3835
rect 38380 3464 38420 3919
rect 38380 3415 38420 3424
rect 38476 2633 38516 5524
rect 38668 5514 38708 5599
rect 38667 5060 38709 5069
rect 38667 5020 38668 5060
rect 38708 5020 38709 5060
rect 38667 5011 38709 5020
rect 38668 4136 38708 5011
rect 38764 4985 38804 6532
rect 39148 6488 39188 6952
rect 39244 6488 39284 6497
rect 39148 6448 39244 6488
rect 39532 6488 39572 8128
rect 39628 8093 39668 8464
rect 39916 8504 39956 8513
rect 39627 8084 39669 8093
rect 39627 8044 39628 8084
rect 39668 8044 39669 8084
rect 39627 8035 39669 8044
rect 39628 6488 39668 6497
rect 39532 6448 39628 6488
rect 39244 6439 39284 6448
rect 39628 6439 39668 6448
rect 39916 6077 39956 8464
rect 40203 8504 40245 8513
rect 40203 8464 40204 8504
rect 40244 8464 40245 8504
rect 40203 8455 40245 8464
rect 40204 8370 40244 8455
rect 40876 8345 40916 8632
rect 41164 8672 41204 8791
rect 41164 8623 41204 8632
rect 40875 8336 40917 8345
rect 40875 8296 40876 8336
rect 40916 8296 40917 8336
rect 40875 8287 40917 8296
rect 41067 8336 41109 8345
rect 41067 8296 41068 8336
rect 41108 8296 41109 8336
rect 41067 8287 41109 8296
rect 41068 8177 41108 8287
rect 41067 8168 41109 8177
rect 41067 8128 41068 8168
rect 41108 8128 41109 8168
rect 41067 8119 41109 8128
rect 40203 8000 40245 8009
rect 40203 7960 40204 8000
rect 40244 7960 40245 8000
rect 40203 7951 40245 7960
rect 41068 8000 41108 8119
rect 41260 8009 41300 10144
rect 41356 10135 41396 10144
rect 41355 10016 41397 10025
rect 41355 9976 41356 10016
rect 41396 9976 41397 10016
rect 41355 9967 41397 9976
rect 41356 9848 41396 9967
rect 41452 9932 41492 12487
rect 41548 12377 41588 14008
rect 41547 12368 41589 12377
rect 41547 12328 41548 12368
rect 41588 12328 41589 12368
rect 41547 12319 41589 12328
rect 41547 11528 41589 11537
rect 41547 11488 41548 11528
rect 41588 11488 41589 11528
rect 41547 11479 41589 11488
rect 41548 11024 41588 11479
rect 41644 11117 41684 15511
rect 43948 15426 43988 15511
rect 44140 15140 44180 17032
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 44428 15308 44468 15317
rect 44140 15100 44276 15140
rect 42123 14804 42165 14813
rect 42123 14764 42124 14804
rect 42164 14764 42165 14804
rect 42123 14755 42165 14764
rect 41740 14720 41780 14729
rect 41740 14216 41780 14680
rect 42124 14720 42164 14755
rect 42124 14669 42164 14680
rect 42987 14720 43029 14729
rect 42987 14680 42988 14720
rect 43028 14680 43029 14720
rect 42987 14671 43029 14680
rect 44140 14720 44180 14729
rect 41740 14167 41780 14176
rect 41835 14216 41877 14225
rect 41835 14176 41836 14216
rect 41876 14176 41877 14216
rect 41835 14167 41877 14176
rect 42028 14216 42068 14225
rect 42068 14176 42164 14216
rect 42028 14167 42068 14176
rect 41739 13964 41781 13973
rect 41739 13924 41740 13964
rect 41780 13924 41781 13964
rect 41739 13915 41781 13924
rect 41740 13208 41780 13915
rect 41836 13712 41876 14167
rect 41931 14048 41973 14057
rect 41931 14008 41932 14048
rect 41972 14008 41973 14048
rect 41931 13999 41973 14008
rect 41932 13914 41972 13999
rect 42027 13880 42069 13889
rect 42027 13840 42028 13880
rect 42068 13840 42069 13880
rect 42027 13831 42069 13840
rect 42028 13712 42068 13831
rect 41836 13672 42068 13712
rect 41932 13208 41972 13672
rect 42028 13217 42068 13302
rect 41780 13168 41876 13208
rect 41740 13159 41780 13168
rect 41739 13040 41781 13049
rect 41739 13000 41740 13040
rect 41780 13000 41781 13040
rect 41836 13040 41876 13168
rect 41932 13159 41972 13168
rect 42027 13208 42069 13217
rect 42027 13168 42028 13208
rect 42068 13168 42069 13208
rect 42027 13159 42069 13168
rect 42124 13049 42164 14176
rect 42508 14048 42548 14057
rect 42508 13889 42548 14008
rect 42507 13880 42549 13889
rect 42507 13840 42508 13880
rect 42548 13840 42549 13880
rect 42507 13831 42549 13840
rect 42795 13880 42837 13889
rect 42795 13840 42796 13880
rect 42836 13840 42837 13880
rect 42795 13831 42837 13840
rect 42411 13376 42453 13385
rect 42411 13336 42412 13376
rect 42452 13336 42453 13376
rect 42411 13327 42453 13336
rect 42316 13292 42356 13301
rect 42220 13208 42260 13217
rect 42123 13040 42165 13049
rect 41836 13000 41972 13040
rect 41739 12991 41781 13000
rect 41740 11621 41780 12991
rect 41932 12788 41972 13000
rect 42123 13000 42124 13040
rect 42164 13000 42165 13040
rect 42123 12991 42165 13000
rect 41932 12748 42164 12788
rect 42124 12704 42164 12748
rect 42124 12655 42164 12664
rect 41835 12620 41877 12629
rect 41835 12580 41836 12620
rect 41876 12580 41877 12620
rect 41835 12571 41877 12580
rect 42028 12620 42068 12629
rect 41836 12536 41876 12571
rect 41836 12377 41876 12496
rect 41932 12536 41972 12547
rect 41932 12461 41972 12496
rect 41931 12452 41973 12461
rect 41931 12412 41932 12452
rect 41972 12412 41973 12452
rect 41931 12403 41973 12412
rect 41835 12368 41877 12377
rect 41835 12328 41836 12368
rect 41876 12328 41877 12368
rect 41835 12319 41877 12328
rect 41932 12284 41972 12293
rect 41739 11612 41781 11621
rect 41739 11572 41740 11612
rect 41780 11572 41781 11612
rect 41739 11563 41781 11572
rect 41643 11108 41685 11117
rect 41643 11068 41644 11108
rect 41684 11068 41685 11108
rect 41643 11059 41685 11068
rect 41548 10975 41588 10984
rect 41644 10361 41684 11059
rect 41740 11024 41780 11033
rect 41643 10352 41685 10361
rect 41643 10312 41644 10352
rect 41684 10312 41685 10352
rect 41643 10303 41685 10312
rect 41740 9941 41780 10984
rect 41932 11024 41972 12244
rect 42028 12125 42068 12580
rect 42220 12452 42260 13168
rect 42316 12452 42356 13252
rect 42412 13242 42452 13327
rect 42508 13292 42548 13301
rect 42508 13217 42548 13252
rect 42507 13208 42549 13217
rect 42507 13168 42508 13208
rect 42548 13168 42549 13208
rect 42507 13159 42549 13168
rect 42604 13208 42644 13217
rect 42508 12713 42548 13159
rect 42507 12704 42549 12713
rect 42507 12664 42508 12704
rect 42548 12664 42549 12704
rect 42604 12704 42644 13168
rect 42796 13208 42836 13831
rect 42796 13159 42836 13168
rect 42604 12664 42836 12704
rect 42507 12655 42549 12664
rect 42604 12536 42644 12545
rect 42220 12412 42265 12452
rect 42316 12412 42452 12452
rect 42123 12368 42165 12377
rect 42123 12328 42124 12368
rect 42164 12328 42165 12368
rect 42123 12319 42165 12328
rect 42124 12234 42164 12319
rect 42225 12284 42265 12412
rect 42220 12244 42265 12284
rect 42027 12116 42069 12125
rect 42027 12076 42028 12116
rect 42068 12076 42069 12116
rect 42027 12067 42069 12076
rect 42220 11957 42260 12244
rect 42412 12041 42452 12412
rect 42604 12377 42644 12496
rect 42699 12536 42741 12545
rect 42699 12496 42700 12536
rect 42740 12496 42741 12536
rect 42699 12487 42741 12496
rect 42603 12368 42645 12377
rect 42603 12328 42604 12368
rect 42644 12328 42645 12368
rect 42603 12319 42645 12328
rect 42700 12293 42740 12487
rect 42507 12284 42549 12293
rect 42507 12244 42508 12284
rect 42548 12244 42549 12284
rect 42507 12235 42549 12244
rect 42699 12284 42741 12293
rect 42699 12244 42700 12284
rect 42740 12244 42741 12284
rect 42699 12235 42741 12244
rect 42411 12032 42453 12041
rect 42411 11992 42412 12032
rect 42452 11992 42453 12032
rect 42411 11983 42453 11992
rect 42027 11948 42069 11957
rect 42027 11908 42028 11948
rect 42068 11908 42069 11948
rect 42027 11899 42069 11908
rect 42219 11948 42261 11957
rect 42219 11908 42220 11948
rect 42260 11908 42261 11948
rect 42219 11899 42261 11908
rect 42028 11444 42068 11899
rect 42508 11789 42548 12235
rect 42699 12032 42741 12041
rect 42699 11992 42700 12032
rect 42740 11992 42741 12032
rect 42699 11983 42741 11992
rect 42507 11780 42549 11789
rect 42507 11740 42508 11780
rect 42548 11740 42549 11780
rect 42507 11731 42549 11740
rect 42123 11696 42165 11705
rect 42123 11656 42124 11696
rect 42164 11656 42165 11696
rect 42123 11647 42165 11656
rect 42124 11562 42164 11647
rect 42219 11444 42261 11453
rect 42028 11404 42220 11444
rect 42260 11404 42261 11444
rect 42219 11395 42261 11404
rect 42123 11276 42165 11285
rect 42123 11236 42124 11276
rect 42164 11236 42165 11276
rect 42123 11227 42165 11236
rect 41932 10975 41972 10984
rect 42124 11024 42164 11227
rect 42124 10975 42164 10984
rect 42220 11024 42260 11395
rect 42508 11369 42548 11731
rect 42507 11360 42549 11369
rect 42507 11320 42508 11360
rect 42548 11320 42549 11360
rect 42507 11311 42549 11320
rect 42412 11192 42452 11201
rect 42452 11152 42548 11192
rect 42412 11143 42452 11152
rect 42220 10975 42260 10984
rect 42316 11108 42356 11117
rect 41836 10940 41876 10949
rect 41739 9932 41781 9941
rect 41452 9892 41588 9932
rect 41356 9808 41492 9848
rect 41452 9512 41492 9808
rect 41452 9463 41492 9472
rect 41355 9428 41397 9437
rect 41355 9388 41356 9428
rect 41396 9388 41397 9428
rect 41355 9379 41397 9388
rect 41356 8681 41396 9379
rect 41548 8849 41588 9892
rect 41739 9892 41740 9932
rect 41780 9892 41781 9932
rect 41739 9883 41781 9892
rect 41739 9680 41781 9689
rect 41739 9640 41740 9680
rect 41780 9640 41781 9680
rect 41739 9631 41781 9640
rect 41740 9428 41780 9631
rect 41740 9379 41780 9388
rect 41547 8840 41589 8849
rect 41547 8800 41548 8840
rect 41588 8800 41589 8840
rect 41547 8791 41589 8800
rect 41451 8756 41493 8765
rect 41451 8716 41452 8756
rect 41492 8716 41493 8756
rect 41451 8707 41493 8716
rect 41355 8672 41397 8681
rect 41355 8632 41356 8672
rect 41396 8632 41397 8672
rect 41355 8623 41397 8632
rect 41356 8504 41396 8623
rect 41356 8455 41396 8464
rect 41452 8504 41492 8707
rect 41548 8588 41588 8791
rect 41548 8539 41588 8548
rect 41644 8672 41684 8681
rect 41452 8455 41492 8464
rect 41451 8084 41493 8093
rect 41451 8044 41452 8084
rect 41492 8044 41493 8084
rect 41451 8035 41493 8044
rect 41068 7951 41108 7960
rect 41259 8000 41301 8009
rect 41259 7960 41260 8000
rect 41300 7960 41301 8000
rect 41259 7951 41301 7960
rect 41452 8000 41492 8035
rect 40108 7412 40148 7421
rect 40204 7412 40244 7951
rect 41452 7949 41492 7960
rect 40148 7372 40244 7412
rect 40108 7363 40148 7372
rect 41644 7337 41684 8632
rect 41740 8672 41780 8681
rect 41740 8513 41780 8632
rect 41739 8504 41781 8513
rect 41739 8464 41740 8504
rect 41780 8464 41781 8504
rect 41739 8455 41781 8464
rect 41643 7328 41685 7337
rect 41643 7288 41644 7328
rect 41684 7288 41685 7328
rect 41643 7279 41685 7288
rect 40587 7244 40629 7253
rect 40587 7204 40588 7244
rect 40628 7204 40629 7244
rect 40587 7195 40629 7204
rect 40396 7160 40436 7169
rect 40396 6488 40436 7120
rect 40588 7110 40628 7195
rect 41260 7160 41300 7169
rect 41260 7085 41300 7120
rect 41452 7160 41492 7169
rect 41644 7160 41684 7279
rect 41492 7120 41684 7160
rect 41836 7160 41876 10900
rect 42219 10352 42261 10361
rect 42219 10312 42220 10352
rect 42260 10312 42261 10352
rect 42219 10303 42261 10312
rect 42220 10184 42260 10303
rect 42316 10277 42356 11068
rect 42412 10772 42452 10781
rect 42315 10268 42357 10277
rect 42315 10228 42316 10268
rect 42356 10228 42357 10268
rect 42315 10219 42357 10228
rect 42220 10135 42260 10144
rect 42412 9521 42452 10732
rect 42124 9512 42164 9521
rect 42411 9512 42453 9521
rect 42164 9472 42356 9512
rect 42124 9463 42164 9472
rect 41932 8504 41972 8513
rect 41972 8464 42260 8504
rect 41932 8455 41972 8464
rect 41931 8000 41973 8009
rect 41931 7960 41932 8000
rect 41972 7960 41973 8000
rect 41931 7951 41973 7960
rect 41932 7866 41972 7951
rect 42220 7412 42260 8464
rect 42316 7916 42356 9472
rect 42411 9472 42412 9512
rect 42452 9472 42453 9512
rect 42411 9463 42453 9472
rect 42508 8429 42548 11152
rect 42603 10184 42645 10193
rect 42603 10144 42604 10184
rect 42644 10144 42645 10184
rect 42603 10135 42645 10144
rect 42604 10050 42644 10135
rect 42700 9353 42740 11983
rect 42796 11369 42836 12664
rect 42988 12545 43028 14671
rect 44140 14216 44180 14680
rect 44236 14720 44276 15100
rect 44428 14897 44468 15268
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 44427 14888 44469 14897
rect 44427 14848 44428 14888
rect 44468 14848 44469 14888
rect 44427 14839 44469 14848
rect 46924 14888 46964 14897
rect 44619 14804 44661 14813
rect 46924 14804 46964 14848
rect 44619 14764 44620 14804
rect 44660 14764 44661 14804
rect 44619 14755 44661 14764
rect 46540 14764 46964 14804
rect 44524 14720 44564 14729
rect 44236 14680 44524 14720
rect 44236 14393 44276 14680
rect 44524 14671 44564 14680
rect 44235 14384 44277 14393
rect 44235 14344 44236 14384
rect 44276 14344 44277 14384
rect 44235 14335 44277 14344
rect 44140 14176 44372 14216
rect 43275 14048 43317 14057
rect 43275 14008 43276 14048
rect 43316 14008 43317 14048
rect 43275 13999 43317 14008
rect 43468 14048 43508 14057
rect 43179 13376 43221 13385
rect 43179 13336 43180 13376
rect 43220 13336 43221 13376
rect 43179 13327 43221 13336
rect 43084 13208 43124 13217
rect 43084 12629 43124 13168
rect 43083 12620 43125 12629
rect 43083 12580 43084 12620
rect 43124 12580 43125 12620
rect 43083 12571 43125 12580
rect 42987 12536 43029 12545
rect 42987 12496 42988 12536
rect 43028 12496 43029 12536
rect 42987 12487 43029 12496
rect 42891 12368 42933 12377
rect 42891 12328 42892 12368
rect 42932 12328 42933 12368
rect 42891 12319 42933 12328
rect 42892 12234 42932 12319
rect 42891 12116 42933 12125
rect 42891 12076 42892 12116
rect 42932 12076 42933 12116
rect 42891 12067 42933 12076
rect 42795 11360 42837 11369
rect 42795 11320 42796 11360
rect 42836 11320 42837 11360
rect 42795 11311 42837 11320
rect 42892 10781 42932 12067
rect 42988 10856 43028 12487
rect 43084 12125 43124 12571
rect 43180 12536 43220 13327
rect 43276 13124 43316 13999
rect 43276 13075 43316 13084
rect 43468 12629 43508 14008
rect 44139 14048 44181 14057
rect 44139 14008 44140 14048
rect 44180 14008 44181 14048
rect 44139 13999 44181 14008
rect 44140 13914 44180 13999
rect 43564 13208 43604 13217
rect 43467 12620 43509 12629
rect 43467 12580 43468 12620
rect 43508 12580 43509 12620
rect 43467 12571 43509 12580
rect 43180 12487 43220 12496
rect 43467 12452 43509 12461
rect 43467 12412 43468 12452
rect 43508 12412 43509 12452
rect 43467 12403 43509 12412
rect 43083 12116 43125 12125
rect 43083 12076 43084 12116
rect 43124 12076 43125 12116
rect 43083 12067 43125 12076
rect 43468 11696 43508 12403
rect 43564 12377 43604 13168
rect 43851 13208 43893 13217
rect 43851 13168 43852 13208
rect 43892 13168 43893 13208
rect 43851 13159 43893 13168
rect 43852 12620 43892 13159
rect 44236 13040 44276 13049
rect 43852 12571 43892 12580
rect 44044 13000 44236 13040
rect 44044 12536 44084 13000
rect 44236 12991 44276 13000
rect 44235 12620 44277 12629
rect 44235 12580 44236 12620
rect 44276 12580 44277 12620
rect 44235 12571 44277 12580
rect 44044 12487 44084 12496
rect 43563 12368 43605 12377
rect 43563 12328 43564 12368
rect 43604 12328 43605 12368
rect 43563 12319 43605 12328
rect 43947 12116 43989 12125
rect 43947 12076 43948 12116
rect 43988 12076 43989 12116
rect 43947 12067 43989 12076
rect 43468 11647 43508 11656
rect 43276 11528 43316 11537
rect 43316 11488 43508 11528
rect 43276 11479 43316 11488
rect 42891 10772 42933 10781
rect 42891 10732 42892 10772
rect 42932 10732 42933 10772
rect 42891 10723 42933 10732
rect 42891 10436 42933 10445
rect 42891 10396 42892 10436
rect 42932 10396 42933 10436
rect 42891 10387 42933 10396
rect 42892 10302 42932 10387
rect 42988 9689 43028 10816
rect 43179 10352 43221 10361
rect 43179 10312 43180 10352
rect 43220 10312 43221 10352
rect 43179 10303 43221 10312
rect 43180 10184 43220 10303
rect 43180 10135 43220 10144
rect 43276 10184 43316 10193
rect 43468 10184 43508 11488
rect 43659 11024 43701 11033
rect 43659 10984 43660 11024
rect 43700 10984 43701 11024
rect 43659 10975 43701 10984
rect 43948 11024 43988 12067
rect 44236 11192 44276 12571
rect 44332 12368 44372 14176
rect 44524 14048 44564 14057
rect 44620 14048 44660 14755
rect 45676 14720 45716 14729
rect 45004 14552 45044 14561
rect 44564 14008 44852 14048
rect 44427 13208 44469 13217
rect 44427 13168 44428 13208
rect 44468 13168 44469 13208
rect 44427 13159 44469 13168
rect 44428 13074 44468 13159
rect 44428 12536 44468 12545
rect 44524 12536 44564 14008
rect 44812 13208 44852 14008
rect 44812 13159 44852 13168
rect 44468 12496 44564 12536
rect 44428 12487 44468 12496
rect 44332 12328 44468 12368
rect 44236 11143 44276 11152
rect 44332 11696 44372 11705
rect 43948 10975 43988 10984
rect 43660 10890 43700 10975
rect 43659 10772 43701 10781
rect 43659 10732 43660 10772
rect 43700 10732 43701 10772
rect 43659 10723 43701 10732
rect 44044 10772 44084 10781
rect 43563 10184 43605 10193
rect 43468 10144 43564 10184
rect 43604 10144 43605 10184
rect 43083 10100 43125 10109
rect 43083 10060 43084 10100
rect 43124 10060 43125 10100
rect 43083 10051 43125 10060
rect 42987 9680 43029 9689
rect 42892 9640 42988 9680
rect 43028 9640 43029 9680
rect 42699 9344 42741 9353
rect 42699 9304 42700 9344
rect 42740 9304 42741 9344
rect 42699 9295 42741 9304
rect 42604 8672 42644 8681
rect 42507 8420 42549 8429
rect 42507 8380 42508 8420
rect 42548 8380 42549 8420
rect 42507 8371 42549 8380
rect 42316 7876 42548 7916
rect 42220 7372 42452 7412
rect 41452 7111 41492 7120
rect 41259 7076 41301 7085
rect 41259 7036 41260 7076
rect 41300 7036 41301 7076
rect 41259 7027 41301 7036
rect 40971 6992 41013 7001
rect 40971 6952 40972 6992
rect 41012 6952 41013 6992
rect 40971 6943 41013 6952
rect 40492 6488 40532 6497
rect 40396 6448 40492 6488
rect 39915 6068 39957 6077
rect 39915 6028 39916 6068
rect 39956 6028 39957 6068
rect 39915 6019 39957 6028
rect 39531 5900 39573 5909
rect 39531 5860 39532 5900
rect 39572 5860 39573 5900
rect 39531 5851 39573 5860
rect 39532 5648 39572 5851
rect 39532 5599 39572 5608
rect 38859 5564 38901 5573
rect 38859 5524 38860 5564
rect 38900 5524 38901 5564
rect 38859 5515 38901 5524
rect 38860 5430 38900 5515
rect 39820 5480 39860 5491
rect 39820 5405 39860 5440
rect 39819 5396 39861 5405
rect 39819 5356 39820 5396
rect 39860 5356 39861 5396
rect 39819 5347 39861 5356
rect 39627 5060 39669 5069
rect 39627 5020 39628 5060
rect 39668 5020 39669 5060
rect 39627 5011 39669 5020
rect 38763 4976 38805 4985
rect 38763 4936 38764 4976
rect 38804 4936 38805 4976
rect 38763 4927 38805 4936
rect 39243 4976 39285 4985
rect 39243 4936 39244 4976
rect 39284 4936 39285 4976
rect 39243 4927 39285 4936
rect 39628 4976 39668 5011
rect 40396 4976 40436 6448
rect 40492 6439 40532 6448
rect 40683 6488 40725 6497
rect 40683 6448 40684 6488
rect 40724 6448 40725 6488
rect 40683 6439 40725 6448
rect 40492 5648 40532 5657
rect 40492 5489 40532 5608
rect 40684 5648 40724 6439
rect 40779 5732 40821 5741
rect 40779 5692 40780 5732
rect 40820 5692 40821 5732
rect 40779 5683 40821 5692
rect 40684 5599 40724 5608
rect 40780 5564 40820 5683
rect 40875 5648 40917 5657
rect 40875 5608 40876 5648
rect 40916 5608 40917 5648
rect 40875 5599 40917 5608
rect 40972 5648 41012 6943
rect 41260 6497 41300 7027
rect 41259 6488 41301 6497
rect 41259 6448 41260 6488
rect 41300 6448 41301 6488
rect 41259 6439 41301 6448
rect 41643 6488 41685 6497
rect 41643 6448 41644 6488
rect 41684 6448 41685 6488
rect 41643 6439 41685 6448
rect 41644 6354 41684 6439
rect 41643 5900 41685 5909
rect 41643 5860 41644 5900
rect 41684 5860 41685 5900
rect 41643 5851 41685 5860
rect 40972 5599 41012 5608
rect 40780 5515 40820 5524
rect 40876 5514 40916 5599
rect 40491 5480 40533 5489
rect 40491 5440 40492 5480
rect 40532 5440 40533 5480
rect 40491 5431 40533 5440
rect 40779 5396 40821 5405
rect 40779 5356 40780 5396
rect 40820 5356 40821 5396
rect 40779 5347 40821 5356
rect 40492 4976 40532 4985
rect 40396 4936 40492 4976
rect 39244 4842 39284 4927
rect 39628 4925 39668 4936
rect 39052 4724 39092 4733
rect 39092 4684 39572 4724
rect 39052 4675 39092 4684
rect 38763 4136 38805 4145
rect 38668 4096 38764 4136
rect 38804 4096 38805 4136
rect 38763 4087 38805 4096
rect 39243 4136 39285 4145
rect 39243 4096 39244 4136
rect 39284 4096 39285 4136
rect 39243 4087 39285 4096
rect 38764 4002 38804 4087
rect 39244 3464 39284 4087
rect 39532 3464 39572 4684
rect 39628 4136 39668 4145
rect 39628 3977 39668 4096
rect 40492 3977 40532 4936
rect 40780 4388 40820 5347
rect 41644 4976 41684 5851
rect 41836 5657 41876 7120
rect 41931 7160 41973 7169
rect 41931 7120 41932 7160
rect 41972 7120 41973 7160
rect 41931 7111 41973 7120
rect 42220 7160 42260 7169
rect 41932 7076 41972 7111
rect 41932 7025 41972 7036
rect 42028 6413 42068 6498
rect 42220 6413 42260 7120
rect 42027 6404 42069 6413
rect 42027 6364 42028 6404
rect 42068 6364 42069 6404
rect 42027 6355 42069 6364
rect 42219 6404 42261 6413
rect 42219 6364 42220 6404
rect 42260 6364 42261 6404
rect 42219 6355 42261 6364
rect 42219 6068 42261 6077
rect 42219 6028 42220 6068
rect 42260 6028 42261 6068
rect 42219 6019 42261 6028
rect 41835 5648 41877 5657
rect 41835 5608 41836 5648
rect 41876 5608 41877 5648
rect 41835 5599 41877 5608
rect 42220 5648 42260 6019
rect 42220 5599 42260 5608
rect 42412 5648 42452 7372
rect 42412 5599 42452 5608
rect 42316 5480 42356 5489
rect 42508 5480 42548 7876
rect 42604 7496 42644 8632
rect 42700 8261 42740 9295
rect 42796 9260 42836 9269
rect 42796 8849 42836 9220
rect 42795 8840 42837 8849
rect 42795 8800 42796 8840
rect 42836 8800 42837 8840
rect 42795 8791 42837 8800
rect 42796 8672 42836 8681
rect 42699 8252 42741 8261
rect 42699 8212 42700 8252
rect 42740 8212 42741 8252
rect 42699 8203 42741 8212
rect 42796 8009 42836 8632
rect 42795 8000 42837 8009
rect 42795 7960 42796 8000
rect 42836 7960 42837 8000
rect 42892 8000 42932 9640
rect 42987 9631 43029 9640
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43084 9512 43124 10051
rect 43276 9680 43316 10144
rect 43563 10135 43605 10144
rect 43564 10050 43604 10135
rect 43371 10016 43413 10025
rect 43371 9972 43372 10016
rect 43412 9972 43413 10016
rect 43371 9967 43413 9972
rect 43372 9881 43412 9967
rect 43660 9932 43700 10723
rect 43564 9892 43700 9932
rect 43276 9640 43412 9680
rect 42988 9378 43028 9463
rect 43084 8924 43124 9472
rect 43276 9512 43316 9523
rect 43276 9437 43316 9472
rect 43275 9428 43317 9437
rect 43275 9388 43276 9428
rect 43316 9388 43317 9428
rect 43275 9379 43317 9388
rect 43179 9344 43221 9353
rect 43179 9304 43180 9344
rect 43220 9304 43221 9344
rect 43179 9295 43221 9304
rect 43180 9210 43220 9295
rect 43084 8884 43316 8924
rect 43084 8000 43124 8009
rect 42892 7960 43084 8000
rect 42795 7951 42837 7960
rect 42987 7832 43029 7841
rect 42987 7792 42988 7832
rect 43028 7792 43029 7832
rect 42987 7783 43029 7792
rect 42604 7456 42836 7496
rect 42699 7328 42741 7337
rect 42699 7288 42700 7328
rect 42740 7288 42741 7328
rect 42699 7279 42741 7288
rect 42603 5648 42645 5657
rect 42603 5608 42604 5648
rect 42644 5608 42645 5648
rect 42603 5599 42645 5608
rect 42700 5648 42740 7279
rect 42700 5599 42740 5608
rect 42604 5514 42644 5599
rect 42796 5564 42836 7456
rect 42891 7328 42933 7337
rect 42891 7288 42892 7328
rect 42932 7288 42933 7328
rect 42891 7279 42933 7288
rect 42892 7194 42932 7279
rect 42988 6320 43028 7783
rect 43084 6488 43124 7960
rect 43276 7412 43316 8884
rect 43372 8681 43412 9640
rect 43468 9260 43508 9269
rect 43468 8765 43508 9220
rect 43467 8756 43509 8765
rect 43467 8716 43468 8756
rect 43508 8716 43509 8756
rect 43467 8707 43509 8716
rect 43371 8672 43413 8681
rect 43371 8632 43372 8672
rect 43412 8632 43413 8672
rect 43371 8623 43413 8632
rect 43467 8504 43509 8513
rect 43467 8464 43468 8504
rect 43508 8464 43509 8504
rect 43467 8455 43509 8464
rect 43468 7841 43508 8455
rect 43467 7832 43509 7841
rect 43467 7792 43468 7832
rect 43508 7792 43509 7832
rect 43467 7783 43509 7792
rect 43564 7664 43604 9892
rect 44044 9521 44084 10732
rect 44236 10436 44276 10445
rect 44332 10436 44372 11656
rect 44428 10781 44468 12328
rect 44715 11948 44757 11957
rect 44715 11908 44716 11948
rect 44756 11908 44757 11948
rect 44715 11899 44757 11908
rect 44716 11814 44756 11899
rect 44811 11780 44853 11789
rect 44811 11740 44812 11780
rect 44852 11740 44853 11780
rect 44811 11731 44853 11740
rect 44812 11696 44852 11731
rect 44812 11645 44852 11656
rect 45004 11033 45044 14512
rect 45388 14048 45428 14057
rect 45291 12536 45333 12545
rect 45291 12496 45292 12536
rect 45332 12496 45333 12536
rect 45291 12487 45333 12496
rect 45292 12402 45332 12487
rect 45099 12284 45141 12293
rect 45099 12244 45100 12284
rect 45140 12244 45141 12284
rect 45099 12235 45141 12244
rect 45100 11948 45140 12235
rect 45100 11899 45140 11908
rect 45099 11360 45141 11369
rect 45099 11320 45100 11360
rect 45140 11320 45141 11360
rect 45099 11311 45141 11320
rect 45100 11192 45140 11311
rect 45388 11201 45428 14008
rect 45676 13889 45716 14680
rect 46540 14720 46580 14764
rect 47596 14720 47636 14729
rect 46540 14671 46580 14680
rect 46636 14680 47596 14720
rect 46636 14048 46676 14680
rect 47596 14671 47636 14680
rect 46636 13999 46676 14008
rect 46924 14552 46964 14561
rect 45675 13880 45717 13889
rect 45675 13840 45676 13880
rect 45716 13840 45717 13880
rect 45675 13831 45717 13840
rect 45676 13208 45716 13217
rect 46828 13208 46868 13217
rect 45676 12545 45716 13168
rect 46636 13168 46828 13208
rect 45675 12536 45717 12545
rect 45675 12496 45676 12536
rect 45716 12496 45717 12536
rect 45675 12487 45717 12496
rect 46444 12284 46484 12293
rect 46444 11873 46484 12244
rect 45771 11864 45813 11873
rect 45771 11824 45772 11864
rect 45812 11824 45813 11864
rect 45771 11815 45813 11824
rect 46443 11864 46485 11873
rect 46443 11824 46444 11864
rect 46484 11824 46485 11864
rect 46443 11815 46485 11824
rect 45772 11696 45812 11815
rect 46636 11789 46676 13168
rect 46828 13159 46868 13168
rect 46924 13040 46964 14512
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 47116 13208 47156 13217
rect 47308 13208 47348 13217
rect 46828 13000 46964 13040
rect 47020 13168 47116 13208
rect 46731 12536 46773 12545
rect 46731 12496 46732 12536
rect 46772 12496 46773 12536
rect 46731 12487 46773 12496
rect 46635 11780 46677 11789
rect 46635 11740 46636 11780
rect 46676 11740 46677 11780
rect 46635 11731 46677 11740
rect 46732 11780 46772 12487
rect 46732 11731 46772 11740
rect 45772 11647 45812 11656
rect 46444 11696 46484 11705
rect 46444 11453 46484 11656
rect 46539 11696 46581 11705
rect 46539 11656 46540 11696
rect 46580 11656 46581 11696
rect 46539 11647 46581 11656
rect 46540 11562 46580 11647
rect 46443 11444 46485 11453
rect 46443 11404 46444 11444
rect 46484 11404 46485 11444
rect 46443 11395 46485 11404
rect 45100 11143 45140 11152
rect 45387 11192 45429 11201
rect 45387 11152 45388 11192
rect 45428 11152 45429 11192
rect 45387 11143 45429 11152
rect 45963 11192 46005 11201
rect 45963 11152 45964 11192
rect 46004 11152 46005 11192
rect 45963 11143 46005 11152
rect 46635 11192 46677 11201
rect 46635 11152 46636 11192
rect 46676 11152 46677 11192
rect 46635 11143 46677 11152
rect 44908 11024 44948 11033
rect 44908 10781 44948 10984
rect 45003 11024 45045 11033
rect 45003 10984 45004 11024
rect 45044 10984 45045 11024
rect 45003 10975 45045 10984
rect 45772 11024 45812 11033
rect 45772 10865 45812 10984
rect 45771 10856 45813 10865
rect 45771 10816 45772 10856
rect 45812 10816 45813 10856
rect 45771 10807 45813 10816
rect 44427 10772 44469 10781
rect 44427 10732 44428 10772
rect 44468 10732 44469 10772
rect 44427 10723 44469 10732
rect 44907 10772 44949 10781
rect 44907 10732 44908 10772
rect 44948 10732 44949 10772
rect 44907 10723 44949 10732
rect 44276 10396 44372 10436
rect 44236 10387 44276 10396
rect 45292 10352 45332 10361
rect 45196 10312 45292 10352
rect 44139 10184 44181 10193
rect 44139 10144 44140 10184
rect 44180 10144 44181 10184
rect 44139 10135 44181 10144
rect 44427 10184 44469 10193
rect 44427 10144 44428 10184
rect 44468 10144 44469 10184
rect 44427 10135 44469 10144
rect 44043 9512 44085 9521
rect 44043 9472 44044 9512
rect 44084 9472 44085 9512
rect 44043 9463 44085 9472
rect 44140 9512 44180 10135
rect 44428 10050 44468 10135
rect 44715 10100 44757 10109
rect 44715 10060 44716 10100
rect 44756 10060 44757 10100
rect 44715 10051 44757 10060
rect 44716 9680 44756 10051
rect 45100 10016 45140 10025
rect 44716 9631 44756 9640
rect 44908 9976 45100 10016
rect 44140 9463 44180 9472
rect 44427 9512 44469 9521
rect 44427 9472 44428 9512
rect 44468 9472 44469 9512
rect 44427 9463 44469 9472
rect 44620 9512 44660 9523
rect 44428 9378 44468 9463
rect 44620 9437 44660 9472
rect 44908 9512 44948 9976
rect 45100 9967 45140 9976
rect 44908 9463 44948 9472
rect 45196 9512 45236 10312
rect 45292 10303 45332 10312
rect 45675 10352 45717 10361
rect 45675 10312 45676 10352
rect 45716 10312 45717 10352
rect 45675 10303 45717 10312
rect 45196 9463 45236 9472
rect 45292 10184 45332 10193
rect 44619 9428 44661 9437
rect 44619 9388 44620 9428
rect 44660 9388 44661 9428
rect 44619 9379 44661 9388
rect 45292 9260 45332 10144
rect 45484 10184 45524 10195
rect 45484 10109 45524 10144
rect 45676 10184 45716 10303
rect 45676 10135 45716 10144
rect 45483 10100 45525 10109
rect 45483 10060 45484 10100
rect 45524 10060 45525 10100
rect 45483 10051 45525 10060
rect 45964 9344 46004 11143
rect 46636 11058 46676 11143
rect 46155 11024 46197 11033
rect 46155 10984 46156 11024
rect 46196 10984 46197 11024
rect 46155 10975 46197 10984
rect 46156 10890 46196 10975
rect 46347 10604 46389 10613
rect 46347 10564 46348 10604
rect 46388 10564 46389 10604
rect 46347 10555 46389 10564
rect 46348 10436 46388 10555
rect 46348 10387 46388 10396
rect 46635 10268 46677 10277
rect 46635 10228 46636 10268
rect 46676 10228 46677 10268
rect 46635 10219 46677 10228
rect 46636 10184 46676 10219
rect 46636 10133 46676 10144
rect 46060 9512 46100 9521
rect 46100 9472 46580 9512
rect 46060 9463 46100 9472
rect 45964 9304 46100 9344
rect 44332 9220 45332 9260
rect 45867 9260 45909 9269
rect 45867 9220 45868 9260
rect 45908 9220 45909 9260
rect 44235 8840 44277 8849
rect 44235 8800 44236 8840
rect 44276 8800 44277 8840
rect 44235 8791 44277 8800
rect 44332 8840 44372 9220
rect 45867 9211 45909 9220
rect 45868 9126 45908 9211
rect 44332 8791 44372 8800
rect 45772 8840 45812 8849
rect 43276 7363 43316 7372
rect 43372 7624 43604 7664
rect 43660 8672 43700 8681
rect 43180 7160 43220 7171
rect 43180 7085 43220 7120
rect 43276 7160 43316 7169
rect 43179 7076 43221 7085
rect 43179 7036 43180 7076
rect 43220 7036 43221 7076
rect 43179 7027 43221 7036
rect 43180 6488 43220 6497
rect 43084 6448 43180 6488
rect 43180 6439 43220 6448
rect 42892 6280 43028 6320
rect 42892 5648 42932 6280
rect 43276 5657 43316 7120
rect 43372 7076 43412 7624
rect 43372 7027 43412 7036
rect 43467 6992 43509 7001
rect 43467 6952 43468 6992
rect 43508 6952 43509 6992
rect 43467 6943 43509 6952
rect 43468 6858 43508 6943
rect 42892 5599 42932 5608
rect 43275 5648 43317 5657
rect 43275 5608 43276 5648
rect 43316 5608 43317 5648
rect 43275 5599 43317 5608
rect 43660 5573 43700 8632
rect 43947 8336 43989 8345
rect 43947 8296 43948 8336
rect 43988 8296 43989 8336
rect 43947 8287 43989 8296
rect 43948 8000 43988 8287
rect 44236 8000 44276 8791
rect 45196 8672 45236 8683
rect 45196 8597 45236 8632
rect 45483 8672 45525 8681
rect 45483 8632 45484 8672
rect 45524 8632 45525 8672
rect 45483 8623 45525 8632
rect 44811 8588 44853 8597
rect 44811 8548 44812 8588
rect 44852 8548 44853 8588
rect 44811 8539 44853 8548
rect 45195 8588 45237 8597
rect 45195 8548 45196 8588
rect 45236 8548 45237 8588
rect 45195 8539 45237 8548
rect 44524 8504 44564 8513
rect 44332 8000 44372 8009
rect 43988 7960 44084 8000
rect 44236 7960 44332 8000
rect 43948 7951 43988 7960
rect 44044 7589 44084 7960
rect 44332 7951 44372 7960
rect 44043 7580 44085 7589
rect 44043 7540 44044 7580
rect 44084 7540 44085 7580
rect 44043 7531 44085 7540
rect 43755 7160 43797 7169
rect 43755 7120 43756 7160
rect 43796 7120 43797 7160
rect 43755 7111 43797 7120
rect 43756 7026 43796 7111
rect 44044 6488 44084 7531
rect 44044 6439 44084 6448
rect 44428 6992 44468 7001
rect 44428 6488 44468 6952
rect 44524 6497 44564 8464
rect 44812 8000 44852 8539
rect 45484 8538 45524 8623
rect 45772 8429 45812 8800
rect 45771 8420 45813 8429
rect 45771 8380 45772 8420
rect 45812 8380 45813 8420
rect 45771 8371 45813 8380
rect 46060 8000 46100 9304
rect 46443 8840 46485 8849
rect 46443 8800 46444 8840
rect 46484 8800 46485 8840
rect 46443 8791 46485 8800
rect 46444 8672 46484 8791
rect 46444 8623 46484 8632
rect 44812 7951 44852 7960
rect 45868 7960 46060 8000
rect 44620 7160 44660 7169
rect 44428 6439 44468 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44620 6320 44660 7120
rect 45292 6992 45332 7001
rect 44716 6497 44756 6582
rect 45292 6497 45332 6952
rect 45580 6992 45620 7001
rect 44715 6488 44757 6497
rect 44715 6448 44716 6488
rect 44756 6448 44757 6488
rect 44715 6439 44757 6448
rect 45291 6488 45333 6497
rect 45291 6448 45292 6488
rect 45332 6448 45333 6488
rect 45291 6439 45333 6448
rect 44524 6280 44660 6320
rect 44715 6320 44757 6329
rect 44715 6280 44716 6320
rect 44756 6280 44757 6320
rect 44235 6068 44277 6077
rect 44235 6028 44236 6068
rect 44276 6028 44277 6068
rect 44235 6019 44277 6028
rect 43947 5648 43989 5657
rect 43947 5608 43948 5648
rect 43988 5608 43989 5648
rect 43947 5599 43989 5608
rect 44236 5648 44276 6019
rect 44236 5599 44276 5608
rect 42796 5515 42836 5524
rect 43659 5564 43701 5573
rect 43659 5524 43660 5564
rect 43700 5524 43701 5564
rect 43659 5515 43701 5524
rect 43948 5514 43988 5599
rect 44428 5564 44468 5573
rect 44524 5564 44564 6280
rect 44715 6271 44757 6280
rect 44716 5648 44756 6271
rect 45003 6068 45045 6077
rect 45003 6028 45004 6068
rect 45044 6028 45045 6068
rect 45003 6019 45045 6028
rect 44716 5599 44756 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45004 5648 45044 6019
rect 45580 5657 45620 6952
rect 45868 6488 45908 7960
rect 46060 7951 46100 7960
rect 46252 7160 46292 7169
rect 46252 6581 46292 7120
rect 46540 7076 46580 9472
rect 46732 9260 46772 9269
rect 46636 8672 46676 8681
rect 46732 8672 46772 9220
rect 46676 8632 46772 8672
rect 46636 8623 46676 8632
rect 46635 8168 46677 8177
rect 46635 8128 46636 8168
rect 46676 8128 46677 8168
rect 46635 8119 46677 8128
rect 46636 7160 46676 8119
rect 46731 7580 46773 7589
rect 46731 7540 46732 7580
rect 46772 7540 46773 7580
rect 46731 7531 46773 7540
rect 46636 7111 46676 7120
rect 46540 7027 46580 7036
rect 46251 6572 46293 6581
rect 46251 6532 46252 6572
rect 46292 6532 46293 6572
rect 46251 6523 46293 6532
rect 45868 6439 45908 6448
rect 46732 6488 46772 7531
rect 46828 7001 46868 13000
rect 46924 12284 46964 12293
rect 46924 11696 46964 12244
rect 46924 11647 46964 11656
rect 47020 10604 47060 13168
rect 47116 13159 47156 13168
rect 47212 13168 47308 13208
rect 47116 13040 47156 13049
rect 47116 11705 47156 13000
rect 47115 11696 47157 11705
rect 47115 11656 47116 11696
rect 47156 11656 47157 11696
rect 47115 11647 47157 11656
rect 47212 10613 47252 13168
rect 47308 13159 47348 13168
rect 47404 13208 47444 13217
rect 47444 13168 47732 13208
rect 47404 13159 47444 13168
rect 47595 12536 47637 12545
rect 47595 12496 47596 12536
rect 47636 12496 47637 12536
rect 47595 12487 47637 12496
rect 47596 12402 47636 12487
rect 47308 11696 47348 11705
rect 47308 11117 47348 11656
rect 47307 11108 47349 11117
rect 47307 11068 47308 11108
rect 47348 11068 47349 11108
rect 47307 11059 47349 11068
rect 47692 11033 47732 13168
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 48652 12536 48692 12545
rect 48652 12293 48692 12496
rect 47980 12284 48020 12293
rect 47980 11453 48020 12244
rect 48651 12284 48693 12293
rect 48651 12244 48652 12284
rect 48692 12244 48693 12284
rect 48651 12235 48693 12244
rect 49323 12200 49365 12209
rect 49323 12160 49324 12200
rect 49364 12160 49365 12200
rect 49323 12151 49365 12160
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 49324 11948 49364 12151
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 49324 11899 49364 11908
rect 48172 11696 48212 11705
rect 47979 11444 48021 11453
rect 47979 11404 47980 11444
rect 48020 11404 48021 11444
rect 47979 11395 48021 11404
rect 48172 11201 48212 11656
rect 48843 11696 48885 11705
rect 48843 11656 48844 11696
rect 48884 11656 48885 11696
rect 48843 11647 48885 11656
rect 48363 11444 48405 11453
rect 48363 11404 48364 11444
rect 48404 11404 48405 11444
rect 48363 11395 48405 11404
rect 48171 11192 48213 11201
rect 48171 11152 48172 11192
rect 48212 11152 48213 11192
rect 48171 11143 48213 11152
rect 47787 11108 47829 11117
rect 47787 11068 47788 11108
rect 47828 11068 47829 11108
rect 47787 11059 47829 11068
rect 48075 11108 48117 11117
rect 48075 11068 48076 11108
rect 48116 11068 48117 11108
rect 48075 11059 48117 11068
rect 47404 11024 47444 11033
rect 46924 10564 47060 10604
rect 47211 10604 47253 10613
rect 47211 10564 47212 10604
rect 47252 10564 47253 10604
rect 46924 10268 46964 10564
rect 47211 10555 47253 10564
rect 47020 10436 47060 10445
rect 47404 10436 47444 10984
rect 47691 11024 47733 11033
rect 47691 10984 47692 11024
rect 47732 10984 47733 11024
rect 47691 10975 47733 10984
rect 47060 10396 47444 10436
rect 47020 10387 47060 10396
rect 46924 10228 47156 10268
rect 46923 10100 46965 10109
rect 46923 10060 46924 10100
rect 46964 10060 46965 10100
rect 46923 10051 46965 10060
rect 46924 8177 46964 10051
rect 47020 9428 47060 9437
rect 47020 8672 47060 9388
rect 47116 8849 47156 10228
rect 47692 10109 47732 10975
rect 47788 10193 47828 11059
rect 48076 10772 48116 11059
rect 48076 10361 48116 10732
rect 48075 10352 48117 10361
rect 48075 10312 48076 10352
rect 48116 10312 48117 10352
rect 48075 10303 48117 10312
rect 47787 10184 47829 10193
rect 48172 10184 48212 11143
rect 48268 11033 48308 11118
rect 48267 11024 48309 11033
rect 48267 10984 48268 11024
rect 48308 10984 48309 11024
rect 48267 10975 48309 10984
rect 48364 11024 48404 11395
rect 48556 11192 48596 11201
rect 48459 11108 48501 11117
rect 48459 11068 48460 11108
rect 48500 11068 48501 11108
rect 48459 11059 48501 11068
rect 48364 10975 48404 10984
rect 48460 10974 48500 11059
rect 48363 10856 48405 10865
rect 48363 10816 48364 10856
rect 48404 10816 48405 10856
rect 48363 10807 48405 10816
rect 48267 10772 48309 10781
rect 48267 10732 48268 10772
rect 48308 10732 48309 10772
rect 48267 10723 48309 10732
rect 47787 10144 47788 10184
rect 47828 10144 47829 10184
rect 47787 10135 47829 10144
rect 47884 10144 48172 10184
rect 47691 10100 47733 10109
rect 47691 10060 47692 10100
rect 47732 10060 47733 10100
rect 47691 10051 47733 10060
rect 47788 9512 47828 10135
rect 47788 9463 47828 9472
rect 47307 9260 47349 9269
rect 47307 9220 47308 9260
rect 47348 9220 47349 9260
rect 47307 9211 47349 9220
rect 47115 8840 47157 8849
rect 47115 8800 47116 8840
rect 47156 8800 47157 8840
rect 47115 8791 47157 8800
rect 46923 8168 46965 8177
rect 46923 8128 46924 8168
rect 46964 8128 46965 8168
rect 46923 8119 46965 8128
rect 46924 8000 46964 8009
rect 47020 8000 47060 8632
rect 47115 8672 47157 8681
rect 47115 8632 47116 8672
rect 47156 8632 47157 8672
rect 47115 8623 47157 8632
rect 46964 7960 47060 8000
rect 46924 7589 46964 7960
rect 46923 7580 46965 7589
rect 46923 7540 46924 7580
rect 46964 7540 46965 7580
rect 46923 7531 46965 7540
rect 47020 7160 47060 7169
rect 47116 7160 47156 8623
rect 47308 8000 47348 9211
rect 47884 8672 47924 10144
rect 48172 10135 48212 10144
rect 48172 9680 48212 9689
rect 48268 9680 48308 10723
rect 48364 10722 48404 10807
rect 48556 10781 48596 11152
rect 48844 11192 48884 11647
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 48844 11143 48884 11152
rect 48940 11024 48980 11033
rect 48555 10772 48597 10781
rect 48555 10732 48556 10772
rect 48596 10732 48597 10772
rect 48555 10723 48597 10732
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 48940 10445 48980 10984
rect 49132 10772 49172 10781
rect 49172 10732 49460 10772
rect 49132 10723 49172 10732
rect 48939 10436 48981 10445
rect 48939 10396 48940 10436
rect 48980 10396 48981 10436
rect 48939 10387 48981 10396
rect 49035 10184 49077 10193
rect 49035 10144 49036 10184
rect 49076 10144 49077 10184
rect 49035 10135 49077 10144
rect 49420 10184 49460 10732
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 49420 10135 49460 10144
rect 49036 10050 49076 10135
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 48212 9640 48308 9680
rect 48172 9631 48212 9640
rect 48844 9512 48884 9521
rect 48884 9472 48980 9512
rect 48844 9463 48884 9472
rect 48172 9260 48212 9269
rect 48172 8681 48212 9220
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 48940 8924 48980 9472
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 49036 8924 49076 8933
rect 48940 8884 49036 8924
rect 49036 8875 49076 8884
rect 47884 8623 47924 8632
rect 48171 8672 48213 8681
rect 48171 8632 48172 8672
rect 48212 8632 48213 8672
rect 48171 8623 48213 8632
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 47308 7951 47348 7960
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 47060 7120 47156 7160
rect 47020 7111 47060 7120
rect 46827 6992 46869 7001
rect 46827 6952 46828 6992
rect 46868 6952 46869 6992
rect 46827 6943 46869 6952
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 46732 6439 46772 6448
rect 47115 6488 47157 6497
rect 47115 6448 47116 6488
rect 47156 6448 47157 6488
rect 47115 6439 47157 6448
rect 47116 6354 47156 6439
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 45004 5599 45044 5608
rect 45579 5648 45621 5657
rect 45579 5608 45580 5648
rect 45620 5608 45621 5648
rect 45579 5599 45621 5608
rect 44468 5524 44564 5564
rect 44811 5564 44853 5573
rect 44811 5524 44812 5564
rect 44852 5524 44853 5564
rect 44428 5515 44468 5524
rect 44811 5515 44853 5524
rect 42356 5440 42548 5480
rect 42316 5431 42356 5440
rect 44812 5430 44852 5515
rect 44908 5514 44948 5599
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 41644 4927 41684 4936
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 40780 4339 40820 4348
rect 39627 3968 39669 3977
rect 39627 3928 39628 3968
rect 39668 3928 39669 3968
rect 39627 3919 39669 3928
rect 40491 3968 40533 3977
rect 40491 3928 40492 3968
rect 40532 3928 40533 3968
rect 40491 3919 40533 3928
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 39628 3464 39668 3473
rect 39532 3424 39628 3464
rect 39244 3415 39284 3424
rect 39628 3415 39668 3424
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 38284 2575 38324 2584
rect 38475 2624 38517 2633
rect 38475 2584 38476 2624
rect 38516 2584 38517 2624
rect 38475 2575 38517 2584
rect 37708 2491 37748 2500
rect 37996 2490 38036 2575
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 34060 1903 34100 1912
rect 30124 1818 30164 1903
rect 32812 1818 32852 1903
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 29644 1280 29684 1289
rect 29260 1240 29644 1280
rect 29644 1231 29684 1240
rect 26668 1063 26708 1072
rect 26859 1112 26901 1121
rect 26859 1072 26860 1112
rect 26900 1072 26901 1112
rect 26859 1063 26901 1072
rect 27723 1112 27765 1121
rect 27723 1072 27724 1112
rect 27764 1072 27765 1112
rect 27723 1063 27765 1072
rect 19564 978 19604 1063
rect 26860 978 26900 1063
rect 19372 944 19412 953
rect 19084 904 19372 944
rect 19372 895 19412 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 9676 38368 9716 38408
rect 11884 38368 11924 38408
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 268 37528 308 37568
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 3436 35764 3476 35804
rect 3916 35764 3956 35804
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3340 35176 3380 35216
rect 3244 34924 3284 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 3724 35176 3764 35216
rect 3628 34924 3668 34964
rect 1132 33412 1172 33452
rect 1228 33328 1268 33368
rect 3532 34336 3572 34376
rect 3628 34252 3668 34292
rect 3820 34756 3860 34796
rect 3916 34672 3956 34712
rect 3916 34168 3956 34208
rect 4684 34924 4724 34964
rect 4204 34588 4244 34628
rect 4492 34336 4532 34376
rect 5068 34672 5108 34712
rect 4780 34420 4820 34460
rect 5260 34504 5300 34544
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 4012 33916 4052 33956
rect 3532 33748 3572 33788
rect 3724 33748 3764 33788
rect 4012 33748 4052 33788
rect 2476 33160 2516 33200
rect 1708 33076 1748 33116
rect 1996 32992 2036 33032
rect 2668 32824 2708 32864
rect 2476 32320 2516 32360
rect 2380 32152 2420 32192
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 3244 33076 3284 33116
rect 3820 33664 3860 33704
rect 3628 33580 3668 33620
rect 3820 33412 3860 33452
rect 3724 33076 3764 33116
rect 3052 32908 3092 32948
rect 3532 32908 3572 32948
rect 2956 32824 2996 32864
rect 2860 32740 2900 32780
rect 3244 32824 3284 32864
rect 4108 32908 4148 32948
rect 3724 32320 3764 32360
rect 2860 32152 2900 32192
rect 2764 31564 2804 31604
rect 3532 31900 3572 31940
rect 3916 31900 3956 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 3916 31648 3956 31688
rect 3820 31564 3860 31604
rect 1324 30388 1364 30428
rect 4012 31396 4052 31436
rect 3052 30388 3092 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3724 30220 3764 30260
rect 3820 30136 3860 30176
rect 3724 30052 3764 30092
rect 2668 29800 2708 29840
rect 1324 29212 1364 29252
rect 2572 29128 2612 29168
rect 1132 28960 1172 29000
rect 1708 28960 1748 29000
rect 3724 29716 3764 29756
rect 3532 29128 3572 29168
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 2764 28624 2804 28664
rect 4492 33076 4532 33116
rect 4300 32992 4340 33032
rect 4780 33664 4820 33704
rect 4876 33244 4916 33284
rect 4588 32656 4628 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 4684 32320 4724 32360
rect 4492 31900 4532 31940
rect 4396 31480 4436 31520
rect 4300 31396 4340 31436
rect 4780 31648 4820 31688
rect 5068 33664 5108 33704
rect 5068 33076 5108 33116
rect 4972 32656 5012 32696
rect 4876 31564 4916 31604
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 4588 30640 4628 30680
rect 4972 30808 5012 30848
rect 4972 30640 5012 30680
rect 5260 33832 5300 33872
rect 5164 32824 5204 32864
rect 6316 35680 6356 35720
rect 6604 36604 6644 36644
rect 6988 36520 7028 36560
rect 6700 35848 6740 35888
rect 6892 35848 6932 35888
rect 6796 35680 6836 35720
rect 6412 35596 6452 35636
rect 5452 35176 5492 35216
rect 5452 34756 5492 34796
rect 5644 34504 5684 34544
rect 5452 34000 5492 34040
rect 5548 33916 5588 33956
rect 6316 34420 6356 34460
rect 5644 33664 5684 33704
rect 5836 33664 5876 33704
rect 5644 33328 5684 33368
rect 6220 34336 6260 34376
rect 6124 33832 6164 33872
rect 6028 33580 6068 33620
rect 6124 33412 6164 33452
rect 5932 33160 5972 33200
rect 7084 35596 7124 35636
rect 6604 35092 6644 35132
rect 6892 35092 6932 35132
rect 6796 35008 6836 35048
rect 6508 34672 6548 34712
rect 6796 34588 6836 34628
rect 6508 34252 6548 34292
rect 6316 34168 6356 34208
rect 6508 34084 6548 34124
rect 7468 37276 7508 37316
rect 8332 37276 8372 37316
rect 8044 36604 8084 36644
rect 7564 36520 7604 36560
rect 7372 35008 7412 35048
rect 7276 34924 7316 34964
rect 6988 34504 7028 34544
rect 7468 34924 7508 34964
rect 8140 35932 8180 35972
rect 8332 35848 8372 35888
rect 8140 35680 8180 35720
rect 7756 35092 7796 35132
rect 7660 34756 7700 34796
rect 7372 34420 7412 34460
rect 7084 34336 7124 34376
rect 6988 34000 7028 34040
rect 6220 32908 6260 32948
rect 5356 32740 5396 32780
rect 6124 32404 6164 32444
rect 5740 31984 5780 32024
rect 6316 32656 6356 32696
rect 6604 33412 6644 33452
rect 6508 32824 6548 32864
rect 6316 31564 6356 31604
rect 6700 32992 6740 33032
rect 7276 32992 7316 33032
rect 7564 34336 7604 34376
rect 7468 34168 7508 34208
rect 7468 33664 7508 33704
rect 7756 34168 7796 34208
rect 7372 32236 7412 32276
rect 7180 32152 7220 32192
rect 9100 36436 9140 36476
rect 8908 35764 8948 35804
rect 8524 35680 8564 35720
rect 9772 37696 9812 37736
rect 9580 36604 9620 36644
rect 9196 35932 9236 35972
rect 9388 35848 9428 35888
rect 9676 35932 9716 35972
rect 10732 38032 10772 38072
rect 11404 37948 11444 37988
rect 11596 38032 11636 38072
rect 11500 37780 11540 37820
rect 9868 37612 9908 37652
rect 10540 37612 10580 37652
rect 12844 37948 12884 37988
rect 10060 37192 10100 37232
rect 9868 36772 9908 36812
rect 9964 36436 10004 36476
rect 10444 37192 10484 37232
rect 10828 36772 10868 36812
rect 10636 36604 10676 36644
rect 10156 35932 10196 35972
rect 10156 35764 10196 35804
rect 8428 35176 8468 35216
rect 9388 34504 9428 34544
rect 9868 35176 9908 35216
rect 9580 34420 9620 34460
rect 8044 34252 8084 34292
rect 7948 32740 7988 32780
rect 7948 32152 7988 32192
rect 8140 33748 8180 33788
rect 8428 33748 8468 33788
rect 8140 32656 8180 32696
rect 8236 32236 8276 32276
rect 8140 32152 8180 32192
rect 7948 31984 7988 32024
rect 6508 31480 6548 31520
rect 6892 31480 6932 31520
rect 5452 31396 5492 31436
rect 5932 31228 5972 31268
rect 6124 31144 6164 31184
rect 7660 31144 7700 31184
rect 7564 31060 7604 31100
rect 4396 30136 4436 30176
rect 4204 29884 4244 29924
rect 5356 30640 5396 30680
rect 5548 30640 5588 30680
rect 4876 30220 4916 30260
rect 5068 30220 5108 30260
rect 5356 30220 5396 30260
rect 4684 30136 4724 30176
rect 4588 30052 4628 30092
rect 4588 29800 4628 29840
rect 5260 30052 5300 30092
rect 5164 29884 5204 29924
rect 4012 29716 4052 29756
rect 4300 29716 4340 29756
rect 3916 29212 3956 29252
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 4876 29212 4916 29252
rect 6028 30556 6068 30596
rect 5836 30220 5876 30260
rect 6316 30640 6356 30680
rect 7564 30640 7604 30680
rect 6508 30556 6548 30596
rect 6604 30052 6644 30092
rect 5644 29212 5684 29252
rect 3820 28288 3860 28328
rect 2956 27700 2996 27740
rect 2476 27616 2516 27656
rect 2572 27616 2612 27656
rect 2860 27616 2900 27656
rect 1228 26860 1268 26900
rect 1900 26692 1940 26732
rect 1708 26608 1748 26648
rect 844 26356 884 26396
rect 1036 24760 1076 24800
rect 940 24676 980 24716
rect 2764 27028 2804 27068
rect 3628 27532 3668 27572
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4108 27784 4148 27824
rect 4876 28456 4916 28496
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3916 27364 3956 27404
rect 3820 27028 3860 27068
rect 2284 26440 2324 26480
rect 2572 26440 2612 26480
rect 2956 26440 2996 26480
rect 2188 25852 2228 25892
rect 1996 24760 2036 24800
rect 2092 24592 2132 24632
rect 3148 26440 3188 26480
rect 3628 26776 3668 26816
rect 4780 27532 4820 27572
rect 4684 27364 4724 27404
rect 4492 27280 4532 27320
rect 3820 26692 3860 26732
rect 3532 26608 3572 26648
rect 3436 26524 3476 26564
rect 3628 26440 3668 26480
rect 3340 26356 3380 26396
rect 3052 25852 3092 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 3436 25516 3476 25556
rect 1612 24340 1652 24380
rect 1132 23668 1172 23708
rect 2476 25180 2516 25220
rect 3628 25180 3668 25220
rect 3916 25180 3956 25220
rect 2380 24592 2420 24632
rect 2668 24592 2708 24632
rect 4396 26776 4436 26816
rect 5932 28876 5972 28916
rect 5452 28456 5492 28496
rect 5068 27700 5108 27740
rect 5836 28372 5876 28412
rect 5260 27868 5300 27908
rect 5740 27868 5780 27908
rect 4684 26692 4724 26732
rect 4972 26692 5012 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 4108 26020 4148 26060
rect 4204 25264 4244 25304
rect 4012 25096 4052 25136
rect 4012 24760 4052 24800
rect 4300 25180 4340 25220
rect 4588 25180 4628 25220
rect 4780 25180 4820 25220
rect 4492 25096 4532 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 2572 24508 2612 24548
rect 2860 24340 2900 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 2380 24088 2420 24128
rect 3532 24004 3572 24044
rect 2668 23920 2708 23960
rect 4396 24676 4436 24716
rect 4588 24592 4628 24632
rect 4108 24172 4148 24212
rect 4012 24004 4052 24044
rect 4204 24004 4244 24044
rect 3724 23752 3764 23792
rect 3820 23500 3860 23540
rect 3820 23248 3860 23288
rect 652 22408 692 22448
rect 652 21568 692 21608
rect 268 20896 308 20936
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 1708 22156 1748 22196
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 5164 25012 5204 25052
rect 5164 24760 5204 24800
rect 4780 24424 4820 24464
rect 4780 24004 4820 24044
rect 4684 23668 4724 23708
rect 4108 23080 4148 23120
rect 4012 22240 4052 22280
rect 2092 21400 2132 21440
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 4876 23752 4916 23792
rect 5548 27700 5588 27740
rect 5452 26692 5492 26732
rect 5356 26104 5396 26144
rect 5356 25516 5396 25556
rect 6124 29128 6164 29168
rect 7276 29044 7316 29084
rect 7468 29296 7508 29336
rect 7564 29128 7604 29168
rect 6508 28624 6548 28664
rect 6700 28288 6740 28328
rect 6604 28120 6644 28160
rect 6028 27616 6068 27656
rect 5836 26860 5876 26900
rect 6412 26860 6452 26900
rect 6892 27364 6932 27404
rect 7084 27616 7124 27656
rect 7276 27364 7316 27404
rect 6988 27280 7028 27320
rect 6796 27112 6836 27152
rect 7564 28288 7604 28328
rect 7564 27112 7604 27152
rect 5932 26692 5972 26732
rect 6316 26524 6356 26564
rect 5932 26356 5972 26396
rect 5548 26020 5588 26060
rect 6124 26104 6164 26144
rect 6220 26020 6260 26060
rect 6316 25516 6356 25556
rect 6508 26776 6548 26816
rect 6700 26692 6740 26732
rect 6508 26608 6548 26648
rect 6604 26272 6644 26312
rect 6028 25264 6068 25304
rect 5932 25096 5972 25136
rect 6220 25096 6260 25136
rect 5836 25038 5876 25052
rect 5836 25012 5876 25038
rect 5260 24508 5300 24548
rect 5260 24340 5300 24380
rect 4492 23248 4532 23288
rect 5068 23248 5108 23288
rect 4396 22324 4436 22364
rect 4300 22240 4340 22280
rect 5356 24172 5396 24212
rect 4780 22828 4820 22868
rect 5740 24592 5780 24632
rect 5644 24508 5684 24548
rect 5644 24340 5684 24380
rect 5644 23500 5684 23540
rect 6124 24676 6164 24716
rect 6028 24424 6068 24464
rect 6508 25012 6548 25052
rect 6700 25012 6740 25052
rect 6508 24592 6548 24632
rect 6412 24424 6452 24464
rect 6604 24340 6644 24380
rect 6316 24172 6356 24212
rect 6124 23920 6164 23960
rect 7468 26860 7508 26900
rect 7084 26440 7124 26480
rect 6892 25936 6932 25976
rect 7564 25264 7604 25304
rect 7564 24676 7604 24716
rect 7756 31060 7796 31100
rect 7756 29884 7796 29924
rect 8044 31228 8084 31268
rect 8044 30640 8084 30680
rect 8044 30052 8084 30092
rect 8236 29884 8276 29924
rect 7852 28372 7892 28412
rect 7756 27700 7796 27740
rect 8332 29800 8372 29840
rect 9388 34336 9428 34376
rect 10156 34672 10196 34712
rect 11116 36016 11156 36056
rect 11404 36520 11444 36560
rect 11212 35764 11252 35804
rect 11116 35680 11156 35720
rect 10924 35260 10964 35300
rect 10540 35008 10580 35048
rect 10060 34504 10100 34544
rect 10060 34084 10100 34124
rect 9868 33496 9908 33536
rect 9964 33160 10004 33200
rect 9292 32908 9332 32948
rect 9964 32824 10004 32864
rect 10444 34336 10484 34376
rect 10732 34672 10772 34712
rect 11596 35848 11636 35888
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 13996 37192 14036 37232
rect 15532 36856 15572 36896
rect 14956 36688 14996 36728
rect 15340 36688 15380 36728
rect 11788 36520 11828 36560
rect 11500 35260 11540 35300
rect 11212 35176 11252 35216
rect 11020 34252 11060 34292
rect 10732 34000 10772 34040
rect 13996 36520 14036 36560
rect 14860 36520 14900 36560
rect 12844 35932 12884 35972
rect 11884 35176 11924 35216
rect 12364 35176 12404 35216
rect 11980 34084 12020 34124
rect 12364 34084 12404 34124
rect 11884 34000 11924 34040
rect 11788 33664 11828 33704
rect 11692 33496 11732 33536
rect 10348 33160 10388 33200
rect 10636 32992 10676 33032
rect 10348 32908 10388 32948
rect 11692 32908 11732 32948
rect 8812 32740 8852 32780
rect 8716 32656 8756 32696
rect 8812 32572 8852 32612
rect 9580 32152 9620 32192
rect 9388 31984 9428 32024
rect 9484 31480 9524 31520
rect 10348 31984 10388 32024
rect 10060 31900 10100 31940
rect 9964 31564 10004 31604
rect 9772 31480 9812 31520
rect 10444 31900 10484 31940
rect 10924 32824 10964 32864
rect 11020 32740 11060 32780
rect 11500 32656 11540 32696
rect 10828 31480 10868 31520
rect 11308 31564 11348 31604
rect 11212 31480 11252 31520
rect 11020 31144 11060 31184
rect 10732 30640 10772 30680
rect 9964 30472 10004 30512
rect 8716 30052 8756 30092
rect 8524 29800 8564 29840
rect 8812 29800 8852 29840
rect 8620 29716 8660 29756
rect 9676 29716 9716 29756
rect 11212 30472 11252 30512
rect 11788 32824 11828 32864
rect 12652 33664 12692 33704
rect 12268 32992 12308 33032
rect 12172 32908 12212 32948
rect 12076 32740 12116 32780
rect 11980 32656 12020 32696
rect 11596 31564 11636 31604
rect 12556 32824 12596 32864
rect 12364 32572 12404 32612
rect 12364 32236 12404 32276
rect 12268 31900 12308 31940
rect 12364 31564 12404 31604
rect 12748 32152 12788 32192
rect 12748 31732 12788 31772
rect 12556 31480 12596 31520
rect 12460 31396 12500 31436
rect 13228 35008 13268 35048
rect 13132 33832 13172 33872
rect 13036 33664 13076 33704
rect 12940 33160 12980 33200
rect 13036 32740 13076 32780
rect 12940 32152 12980 32192
rect 13132 32404 13172 32444
rect 13612 35176 13652 35216
rect 13708 33832 13748 33872
rect 13612 32824 13652 32864
rect 14380 35680 14420 35720
rect 14956 35680 14996 35720
rect 13996 34000 14036 34040
rect 14956 35008 14996 35048
rect 14092 33832 14132 33872
rect 14572 34084 14612 34124
rect 14572 33076 14612 33116
rect 14380 32824 14420 32864
rect 13804 32404 13844 32444
rect 13708 32320 13748 32360
rect 13132 32068 13172 32108
rect 12940 31900 12980 31940
rect 12076 31228 12116 31268
rect 12652 31060 12692 31100
rect 12844 31312 12884 31352
rect 12844 31144 12884 31184
rect 12748 30892 12788 30932
rect 10828 30052 10868 30092
rect 10828 29884 10868 29924
rect 12844 30808 12884 30848
rect 12844 30556 12884 30596
rect 12652 30220 12692 30260
rect 12172 29884 12212 29924
rect 11788 29296 11828 29336
rect 11692 28960 11732 29000
rect 10348 28876 10388 28916
rect 11116 28876 11156 28916
rect 11500 28876 11540 28916
rect 8428 28288 8468 28328
rect 8140 28120 8180 28160
rect 8140 27616 8180 27656
rect 8428 27616 8468 27656
rect 7948 27448 7988 27488
rect 7852 27280 7892 27320
rect 7948 27112 7988 27152
rect 7852 26776 7892 26816
rect 8524 27364 8564 27404
rect 8428 27028 8468 27068
rect 8524 26860 8564 26900
rect 8332 26608 8372 26648
rect 7948 26356 7988 26396
rect 7756 26272 7796 26312
rect 7852 26104 7892 26144
rect 9676 28120 9716 28160
rect 10060 27868 10100 27908
rect 9292 27448 9332 27488
rect 10540 27700 10580 27740
rect 10924 27700 10964 27740
rect 9964 27280 10004 27320
rect 8716 26356 8756 26396
rect 9484 27112 9524 27152
rect 9772 27112 9812 27152
rect 8908 26860 8948 26900
rect 7756 25936 7796 25976
rect 9292 26776 9332 26816
rect 9868 26860 9908 26900
rect 10540 27112 10580 27152
rect 10252 26944 10292 26984
rect 9676 26692 9716 26732
rect 10060 26608 10100 26648
rect 10252 26776 10292 26816
rect 10444 26440 10484 26480
rect 10060 26104 10100 26144
rect 8908 25768 8948 25808
rect 7948 24844 7988 24884
rect 7276 24424 7316 24464
rect 7948 24508 7988 24548
rect 7852 24256 7892 24296
rect 8140 24424 8180 24464
rect 8044 23920 8084 23960
rect 5836 23080 5876 23120
rect 5260 22744 5300 22784
rect 4972 22660 5012 22700
rect 5548 22660 5588 22700
rect 5452 22324 5492 22364
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4492 21736 4532 21776
rect 4876 22156 4916 22196
rect 4876 21652 4916 21692
rect 4492 20728 4532 20768
rect 5644 22324 5684 22364
rect 5164 21904 5204 21944
rect 5068 21736 5108 21776
rect 5548 21904 5588 21944
rect 5260 21568 5300 21608
rect 5068 21400 5108 21440
rect 4972 21232 5012 21272
rect 4780 21148 4820 21188
rect 4876 20728 4916 20768
rect 6028 22828 6068 22868
rect 6124 22744 6164 22784
rect 6508 22828 6548 22868
rect 7852 22744 7892 22784
rect 7372 22660 7412 22700
rect 7564 22324 7604 22364
rect 6124 22240 6164 22280
rect 5932 21568 5972 21608
rect 6604 21652 6644 21692
rect 6508 21568 6548 21608
rect 6604 21484 6644 21524
rect 5836 21400 5876 21440
rect 6220 21400 6260 21440
rect 5644 21148 5684 21188
rect 6220 20812 6260 20852
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 5164 20728 5204 20768
rect 4972 20308 5012 20348
rect 4108 20224 4148 20264
rect 3532 20056 3572 20096
rect 2956 19804 2996 19844
rect 844 18796 884 18836
rect 2284 19048 2324 19088
rect 1900 18712 1940 18752
rect 1996 18544 2036 18584
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 1036 17032 1076 17072
rect 652 16528 692 16568
rect 748 15688 788 15728
rect 1228 16360 1268 16400
rect 1228 16108 1268 16148
rect 1132 15940 1172 15980
rect 1132 15520 1172 15560
rect 1036 14848 1076 14888
rect 940 14680 980 14720
rect 1708 17032 1748 17072
rect 1420 16024 1460 16064
rect 1612 16192 1652 16232
rect 2092 16360 2132 16400
rect 2188 16276 2228 16316
rect 2572 18880 2612 18920
rect 2860 18712 2900 18752
rect 2764 18544 2804 18584
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 5260 20560 5300 20600
rect 5164 20224 5204 20264
rect 4876 20056 4916 20096
rect 4012 19972 4052 20012
rect 3244 18964 3284 19004
rect 3148 18880 3188 18920
rect 3820 19216 3860 19256
rect 3820 19048 3860 19088
rect 4876 19804 4916 19844
rect 4012 18964 4052 19004
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3532 18712 3572 18752
rect 4108 18712 4148 18752
rect 2764 18208 2804 18248
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3628 17788 3668 17828
rect 2572 17032 2612 17072
rect 3628 17032 3668 17072
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 2476 15940 2516 15980
rect 2476 15604 2516 15644
rect 1708 15520 1748 15560
rect 2380 15520 2420 15560
rect 2380 15268 2420 15308
rect 3340 16024 3380 16064
rect 3916 15940 3956 15980
rect 5068 18712 5108 18752
rect 5068 18460 5108 18500
rect 4780 17788 4820 17828
rect 4972 17788 5012 17828
rect 4396 17704 4436 17744
rect 4588 17620 4628 17660
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4204 16192 4244 16232
rect 4108 15772 4148 15812
rect 4012 15688 4052 15728
rect 3628 15520 3668 15560
rect 1612 15184 1652 15224
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 3532 14932 3572 14972
rect 4972 17620 5012 17660
rect 4876 17032 4916 17072
rect 4876 16192 4916 16232
rect 5740 20728 5780 20768
rect 5644 20560 5684 20600
rect 5548 20140 5588 20180
rect 5644 20056 5684 20096
rect 6028 19888 6068 19928
rect 5932 19300 5972 19340
rect 5548 19216 5588 19256
rect 5356 18712 5396 18752
rect 5260 18460 5300 18500
rect 5260 18292 5300 18332
rect 5356 17536 5396 17576
rect 5068 16360 5108 16400
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4780 15856 4820 15896
rect 5068 15856 5108 15896
rect 5644 18544 5684 18584
rect 5836 18628 5876 18668
rect 6508 20056 6548 20096
rect 7468 22240 7508 22280
rect 7276 22156 7316 22196
rect 9964 25600 10004 25640
rect 9292 25348 9332 25388
rect 9100 25264 9140 25304
rect 9388 25264 9428 25304
rect 9292 24928 9332 24968
rect 9004 24676 9044 24716
rect 8716 24424 8756 24464
rect 8716 23920 8756 23960
rect 11596 27700 11636 27740
rect 11692 27616 11732 27656
rect 11212 27448 11252 27488
rect 11116 27364 11156 27404
rect 11404 26440 11444 26480
rect 11212 26104 11252 26144
rect 11692 26776 11732 26816
rect 11884 26776 11924 26816
rect 11788 26692 11828 26732
rect 11500 26020 11540 26060
rect 10540 25684 10580 25724
rect 9868 25096 9908 25136
rect 10060 24928 10100 24968
rect 9004 23248 9044 23288
rect 8812 23080 8852 23120
rect 9580 23920 9620 23960
rect 9292 22996 9332 23036
rect 9004 22912 9044 22952
rect 9580 22828 9620 22868
rect 6796 20308 6836 20348
rect 6604 19972 6644 20012
rect 6604 19384 6644 19424
rect 6220 19300 6260 19340
rect 6220 19048 6260 19088
rect 9964 24592 10004 24632
rect 10444 25264 10484 25304
rect 12460 28204 12500 28244
rect 12076 27616 12116 27656
rect 12076 26104 12116 26144
rect 12076 25684 12116 25724
rect 10732 25600 10772 25640
rect 11980 25600 12020 25640
rect 10636 25264 10676 25304
rect 11020 25432 11060 25472
rect 11884 25432 11924 25472
rect 10828 25264 10868 25304
rect 11884 25264 11924 25304
rect 12172 25264 12212 25304
rect 10636 25096 10676 25136
rect 10252 24928 10292 24968
rect 10348 24676 10388 24716
rect 10060 23752 10100 23792
rect 9868 23248 9908 23288
rect 10828 25012 10868 25052
rect 11308 24928 11348 24968
rect 11692 24676 11732 24716
rect 12556 27868 12596 27908
rect 12748 27700 12788 27740
rect 12460 26608 12500 26648
rect 13132 31648 13172 31688
rect 13324 31480 13364 31520
rect 12940 30136 12980 30176
rect 13228 31312 13268 31352
rect 13516 31396 13556 31436
rect 13612 31228 13652 31268
rect 13804 32152 13844 32192
rect 13996 31564 14036 31604
rect 13516 31060 13556 31100
rect 13132 30640 13172 30680
rect 13612 30976 13652 31016
rect 14284 32488 14324 32528
rect 14476 32152 14516 32192
rect 15628 36688 15668 36728
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 16396 36856 16436 36896
rect 16492 36772 16532 36812
rect 17548 36772 17588 36812
rect 16684 36688 16724 36728
rect 16012 36520 16052 36560
rect 15820 35680 15860 35720
rect 15340 35176 15380 35216
rect 16204 35176 16244 35216
rect 16588 35176 16628 35216
rect 16492 35008 16532 35048
rect 15532 33076 15572 33116
rect 14956 32824 14996 32864
rect 14860 32488 14900 32528
rect 14764 32320 14804 32360
rect 14668 32152 14708 32192
rect 14284 32068 14324 32108
rect 14188 31396 14228 31436
rect 14764 31396 14804 31436
rect 14284 31312 14324 31352
rect 14668 31312 14708 31352
rect 15148 32656 15188 32696
rect 14956 31816 14996 31856
rect 15148 31564 15188 31604
rect 14764 31228 14804 31268
rect 13996 30976 14036 31016
rect 13900 30808 13940 30848
rect 13804 30388 13844 30428
rect 13420 30220 13460 30260
rect 13804 30136 13844 30176
rect 13708 29128 13748 29168
rect 12940 28204 12980 28244
rect 13036 27616 13076 27656
rect 13612 28876 13652 28916
rect 13324 27448 13364 27488
rect 13132 26692 13172 26732
rect 13036 26608 13076 26648
rect 13132 26524 13172 26564
rect 13036 26104 13076 26144
rect 12748 25768 12788 25808
rect 12652 25348 12692 25388
rect 12556 25264 12596 25304
rect 12940 25600 12980 25640
rect 12460 24844 12500 24884
rect 11980 24592 12020 24632
rect 12364 24592 12404 24632
rect 12652 24508 12692 24548
rect 11308 24424 11348 24464
rect 11884 23752 11924 23792
rect 11212 23668 11252 23708
rect 11692 23668 11732 23708
rect 10156 23080 10196 23120
rect 9868 22996 9908 23036
rect 10060 22828 10100 22868
rect 8236 22156 8276 22196
rect 8140 21484 8180 21524
rect 7756 20812 7796 20852
rect 8524 21484 8564 21524
rect 8908 20812 8948 20852
rect 9004 20644 9044 20684
rect 6892 20056 6932 20096
rect 7372 20056 7412 20096
rect 6220 18796 6260 18836
rect 5932 18544 5972 18584
rect 5932 18292 5972 18332
rect 5836 18124 5876 18164
rect 5740 17788 5780 17828
rect 6124 17788 6164 17828
rect 6028 17704 6068 17744
rect 5740 17620 5780 17660
rect 5644 17536 5684 17576
rect 7180 18880 7220 18920
rect 6412 18544 6452 18584
rect 6604 18544 6644 18584
rect 6508 18460 6548 18500
rect 6412 18376 6452 18416
rect 6796 18376 6836 18416
rect 6700 17872 6740 17912
rect 6604 17704 6644 17744
rect 6796 17704 6836 17744
rect 7372 18880 7412 18920
rect 8044 19216 8084 19256
rect 7468 18628 7508 18668
rect 7372 18460 7412 18500
rect 6988 17704 7028 17744
rect 6988 17536 7028 17576
rect 6316 16948 6356 16988
rect 5363 16024 5396 16064
rect 5396 16024 5403 16064
rect 5452 15772 5492 15812
rect 4972 15688 5012 15728
rect 4300 15604 4340 15644
rect 3820 15184 3860 15224
rect 4012 15100 4052 15140
rect 2764 14680 2804 14720
rect 3628 14680 3668 14720
rect 4012 14260 4052 14300
rect 4204 15268 4244 15308
rect 5356 15688 5396 15728
rect 4876 15436 4916 15476
rect 4780 15100 4820 15140
rect 1324 14092 1364 14132
rect 652 14008 692 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 652 13168 692 13208
rect 2956 13000 2996 13040
rect 4108 14176 4148 14216
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4492 14176 4532 14216
rect 4684 14176 4724 14216
rect 4204 13924 4244 13964
rect 3820 13840 3860 13880
rect 5452 15520 5492 15560
rect 5260 15436 5300 15476
rect 5164 15352 5204 15392
rect 5164 15184 5204 15224
rect 5452 15016 5492 15056
rect 5356 14932 5396 14972
rect 5260 14848 5300 14888
rect 5932 15856 5972 15896
rect 6220 15856 6260 15896
rect 5644 15688 5684 15728
rect 5644 15100 5684 15140
rect 5644 14932 5684 14972
rect 5068 14008 5108 14048
rect 5356 14344 5396 14384
rect 5548 14512 5588 14552
rect 5452 14008 5492 14048
rect 5740 14008 5780 14048
rect 6028 15772 6068 15812
rect 6412 16360 6452 16400
rect 6412 15940 6452 15980
rect 6604 16948 6644 16988
rect 6988 17116 7028 17156
rect 7180 16948 7220 16988
rect 6796 16864 6836 16904
rect 6700 16696 6740 16736
rect 6508 15856 6548 15896
rect 6604 15688 6644 15728
rect 6220 15436 6260 15476
rect 6124 15184 6164 15224
rect 6316 15268 6356 15308
rect 6412 14932 6452 14972
rect 5260 13924 5300 13964
rect 6124 13840 6164 13880
rect 3628 13168 3668 13208
rect 3532 12580 3572 12620
rect 652 12328 692 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3724 11908 3764 11948
rect 5356 13336 5396 13376
rect 5836 13252 5876 13292
rect 4012 12916 4052 12956
rect 4300 13000 4340 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3916 11908 3956 11948
rect 4012 11824 4052 11864
rect 3820 11656 3860 11696
rect 652 11488 692 11528
rect 3628 11152 3668 11192
rect 2572 10984 2612 11024
rect 1516 10816 1556 10856
rect 652 10648 692 10688
rect 2572 10816 2612 10856
rect 2572 10144 2612 10184
rect 652 9808 692 9848
rect 1612 9472 1652 9512
rect 1036 9220 1076 9260
rect 652 8968 692 9008
rect 1324 8884 1364 8924
rect 652 8128 692 8168
rect 1036 8128 1076 8168
rect 1708 9304 1748 9344
rect 1420 8044 1460 8084
rect 844 7876 884 7916
rect 1132 7792 1172 7832
rect 844 7708 884 7748
rect 652 7288 692 7328
rect 1612 7960 1652 8000
rect 1900 9220 1940 9260
rect 2284 8884 2324 8924
rect 2380 8800 2420 8840
rect 2764 10144 2804 10184
rect 3436 10984 3476 11024
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3532 9976 3572 10016
rect 3532 9472 3572 9512
rect 2860 9388 2900 9428
rect 2668 8800 2708 8840
rect 1708 7876 1748 7916
rect 1996 7876 2036 7916
rect 1804 7708 1844 7748
rect 1228 7288 1268 7328
rect 652 6448 692 6488
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4012 11068 4052 11108
rect 4492 11908 4532 11948
rect 4396 11656 4436 11696
rect 4684 11824 4724 11864
rect 5548 13168 5588 13208
rect 5644 12916 5684 12956
rect 5644 12580 5684 12620
rect 6796 15856 6836 15896
rect 6604 15436 6644 15476
rect 6700 15352 6740 15392
rect 6604 14344 6644 14384
rect 6508 13924 6548 13964
rect 6220 13336 6260 13376
rect 7372 17032 7412 17072
rect 7276 16192 7316 16232
rect 7084 15688 7124 15728
rect 7180 15604 7220 15644
rect 6988 15520 7028 15560
rect 7180 15100 7220 15140
rect 7084 14680 7124 14720
rect 7468 16864 7508 16904
rect 8044 18544 8084 18584
rect 8524 19384 8564 19424
rect 8716 20056 8756 20096
rect 9100 19384 9140 19424
rect 9772 21568 9812 21608
rect 11212 23080 11252 23120
rect 10732 22912 10772 22952
rect 10924 22324 10964 22364
rect 9868 20812 9908 20852
rect 9964 20644 10004 20684
rect 11212 21652 11252 21692
rect 10348 21316 10388 21356
rect 10444 20812 10484 20852
rect 10636 20728 10676 20768
rect 10444 20476 10484 20516
rect 9676 19972 9716 20012
rect 8620 18880 8660 18920
rect 8716 18712 8756 18752
rect 7756 17956 7796 17996
rect 7660 16780 7700 16820
rect 7564 16696 7604 16736
rect 7564 16024 7604 16064
rect 7468 15856 7508 15896
rect 7660 15688 7700 15728
rect 7564 15604 7604 15644
rect 7468 15520 7508 15560
rect 8332 17536 8372 17576
rect 9292 18712 9332 18752
rect 9772 18376 9812 18416
rect 7948 16780 7988 16820
rect 8812 17032 8852 17072
rect 9196 17032 9236 17072
rect 8524 16864 8564 16904
rect 8332 16192 8372 16232
rect 8908 16024 8948 16064
rect 9100 15856 9140 15896
rect 8620 15688 8660 15728
rect 8236 14848 8276 14888
rect 7756 14344 7796 14384
rect 9388 17032 9428 17072
rect 9964 18880 10004 18920
rect 10060 18712 10100 18752
rect 10060 17704 10100 17744
rect 9868 17116 9908 17156
rect 9580 15688 9620 15728
rect 10252 19972 10292 20012
rect 11404 21568 11444 21608
rect 11980 23668 12020 23708
rect 12556 22828 12596 22868
rect 11884 22660 11924 22700
rect 12460 22660 12500 22700
rect 12268 22576 12308 22616
rect 11788 22240 11828 22280
rect 12844 24844 12884 24884
rect 12844 23752 12884 23792
rect 12748 23668 12788 23708
rect 13420 26440 13460 26480
rect 13996 27364 14036 27404
rect 13804 27028 13844 27068
rect 13804 26608 13844 26648
rect 13996 26608 14036 26648
rect 13900 26524 13940 26564
rect 13996 26440 14036 26480
rect 13228 26104 13268 26144
rect 13223 25432 13263 25472
rect 13036 25012 13076 25052
rect 13420 24928 13460 24968
rect 13228 24676 13268 24716
rect 13612 26104 13652 26144
rect 13900 26104 13940 26144
rect 14572 30724 14612 30764
rect 14188 30640 14228 30680
rect 15052 30472 15092 30512
rect 14668 30388 14708 30428
rect 15436 31732 15476 31772
rect 15340 31480 15380 31520
rect 15340 31228 15380 31268
rect 15820 33664 15860 33704
rect 16108 32740 16148 32780
rect 16876 36688 16916 36728
rect 17164 36520 17204 36560
rect 16876 35260 16916 35300
rect 17164 35848 17204 35888
rect 17068 35260 17108 35300
rect 16972 35176 17012 35216
rect 18124 36688 18164 36728
rect 17548 35260 17588 35300
rect 18028 35260 18068 35300
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 18796 36016 18836 36056
rect 19180 36016 19220 36056
rect 18316 35848 18356 35888
rect 17260 35092 17300 35132
rect 16780 35008 16820 35048
rect 16684 34924 16724 34964
rect 16492 33076 16532 33116
rect 16684 33076 16724 33116
rect 16780 32824 16820 32864
rect 16972 34168 17012 34208
rect 16204 32236 16244 32276
rect 16012 32152 16052 32192
rect 16108 31900 16148 31940
rect 15628 31564 15668 31604
rect 16012 31396 16052 31436
rect 15916 31228 15956 31268
rect 16588 32656 16628 32696
rect 16876 32656 16916 32696
rect 17740 34924 17780 34964
rect 17260 34168 17300 34208
rect 17548 34000 17588 34040
rect 17260 32824 17300 32864
rect 17836 34168 17876 34208
rect 17356 32740 17396 32780
rect 16300 32152 16340 32192
rect 16300 31900 16340 31940
rect 16300 31732 16340 31772
rect 16300 31228 16340 31268
rect 15532 30892 15572 30932
rect 15436 30808 15476 30848
rect 15820 30808 15860 30848
rect 15532 30556 15572 30596
rect 15436 30472 15476 30512
rect 14380 29800 14420 29840
rect 14572 29800 14612 29840
rect 15244 29800 15284 29840
rect 15820 30388 15860 30428
rect 15916 30220 15956 30260
rect 15820 29380 15860 29420
rect 14860 29296 14900 29336
rect 14572 29212 14612 29252
rect 14476 29044 14516 29084
rect 14668 28876 14708 28916
rect 14188 28792 14228 28832
rect 14476 27448 14516 27488
rect 14572 27364 14612 27404
rect 15340 28624 15380 28664
rect 15244 28540 15284 28580
rect 14764 27784 14804 27824
rect 14188 26692 14228 26732
rect 15820 28288 15860 28328
rect 15628 27448 15668 27488
rect 14860 27364 14900 27404
rect 14284 26608 14324 26648
rect 14188 26524 14228 26564
rect 14092 26272 14132 26312
rect 13804 25936 13844 25976
rect 13996 25936 14036 25976
rect 13708 25852 13748 25892
rect 13708 25516 13748 25556
rect 13612 25432 13652 25472
rect 13612 25264 13652 25304
rect 13036 22828 13076 22868
rect 12652 22576 12692 22616
rect 12556 22240 12596 22280
rect 12940 22408 12980 22448
rect 11788 21652 11828 21692
rect 13900 25096 13940 25136
rect 13804 24340 13844 24380
rect 14380 26440 14420 26480
rect 14727 26692 14767 26732
rect 14956 26776 14996 26816
rect 15148 26776 15188 26816
rect 15436 26776 15476 26816
rect 16108 28288 16148 28328
rect 16012 27700 16052 27740
rect 15916 27616 15956 27656
rect 15724 27280 15764 27320
rect 14668 26524 14708 26564
rect 14860 26524 14900 26564
rect 14284 25768 14324 25808
rect 14380 25264 14420 25304
rect 14572 26104 14612 26144
rect 15052 26440 15092 26480
rect 14764 26272 14804 26312
rect 14956 26272 14996 26312
rect 14860 26188 14900 26228
rect 14860 25852 14900 25892
rect 15052 25684 15092 25724
rect 15532 26692 15572 26732
rect 15436 26524 15476 26564
rect 15340 26440 15380 26480
rect 15340 26272 15380 26312
rect 15340 26104 15380 26144
rect 15244 26020 15284 26060
rect 15532 25768 15572 25808
rect 15724 26020 15764 26060
rect 16588 31396 16628 31436
rect 17164 31312 17204 31352
rect 16492 30808 16532 30848
rect 16972 30724 17012 30764
rect 16492 30556 16532 30596
rect 16492 29128 16532 29168
rect 16780 29128 16820 29168
rect 16972 29212 17012 29252
rect 16876 28792 16916 28832
rect 17452 32656 17492 32696
rect 17452 32152 17492 32192
rect 17452 31816 17492 31856
rect 18028 33664 18068 33704
rect 18412 35260 18452 35300
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 21196 35680 21236 35720
rect 22348 35680 22388 35720
rect 18988 35260 19028 35300
rect 19660 35176 19700 35216
rect 20044 35176 20084 35216
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 18316 34504 18356 34544
rect 18796 34504 18836 34544
rect 19660 34504 19700 34544
rect 19948 34504 19988 34544
rect 20812 34924 20852 34964
rect 21772 34924 21812 34964
rect 19372 34420 19412 34460
rect 18604 34336 18644 34376
rect 18796 34336 18836 34376
rect 18700 33664 18740 33704
rect 18028 32656 18068 32696
rect 17932 32404 17972 32444
rect 17836 32152 17876 32192
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 18220 33076 18260 33116
rect 18412 32824 18452 32864
rect 19852 34336 19892 34376
rect 20044 34336 20084 34376
rect 20140 34252 20180 34292
rect 19948 34168 19988 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 18796 33076 18836 33116
rect 19852 33076 19892 33116
rect 19660 32992 19700 33032
rect 19276 32908 19316 32948
rect 19372 32824 19412 32864
rect 21676 34504 21716 34544
rect 21196 34336 21236 34376
rect 20524 34168 20564 34208
rect 21388 34252 21428 34292
rect 21580 34168 21620 34208
rect 22156 34252 22196 34292
rect 21772 33832 21812 33872
rect 21580 33748 21620 33788
rect 20236 33664 20276 33704
rect 18412 32404 18452 32444
rect 20524 32992 20564 33032
rect 21292 32992 21332 33032
rect 20236 32740 20276 32780
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 20908 32908 20948 32948
rect 22252 33748 22292 33788
rect 21772 33496 21812 33536
rect 21676 32992 21716 33032
rect 21964 32824 22004 32864
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 23116 35176 23156 35216
rect 24076 35176 24116 35216
rect 26188 35008 26228 35048
rect 23788 34000 23828 34040
rect 23692 33916 23732 33956
rect 22636 33664 22676 33704
rect 22252 32740 22292 32780
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 17836 30808 17876 30848
rect 17548 30556 17588 30596
rect 17644 29632 17684 29672
rect 17644 29380 17684 29420
rect 17452 28540 17492 28580
rect 16588 27532 16628 27572
rect 16108 26440 16148 26480
rect 16108 26272 16148 26312
rect 16012 26104 16052 26144
rect 16588 26776 16628 26816
rect 16396 26104 16436 26144
rect 16588 26104 16628 26144
rect 20716 31480 20756 31520
rect 21100 31480 21140 31520
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 18892 30724 18932 30764
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 18700 29296 18740 29336
rect 19180 30640 19220 30680
rect 19372 30556 19412 30596
rect 19180 29632 19220 29672
rect 19084 29128 19124 29168
rect 18796 29044 18836 29084
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 17260 27784 17300 27824
rect 17740 27784 17780 27824
rect 17452 27700 17492 27740
rect 17548 27532 17588 27572
rect 17356 27448 17396 27488
rect 17836 27364 17876 27404
rect 18604 28540 18644 28580
rect 18796 28540 18836 28580
rect 19084 28372 19124 28412
rect 18988 28288 19028 28328
rect 18796 27448 18836 27488
rect 18508 27364 18548 27404
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 18124 27028 18164 27068
rect 18700 27028 18740 27068
rect 18604 26944 18644 26984
rect 16780 26776 16820 26816
rect 16972 26776 17012 26816
rect 17164 26776 17204 26816
rect 17836 26776 17876 26816
rect 17164 26356 17204 26396
rect 17068 26272 17108 26312
rect 16780 26020 16820 26060
rect 15148 25432 15188 25472
rect 15052 25348 15092 25388
rect 15532 25348 15572 25388
rect 15724 25348 15764 25388
rect 14476 25180 14516 25220
rect 14380 24340 14420 24380
rect 13900 24004 13940 24044
rect 13996 23920 14036 23960
rect 13900 23752 13940 23792
rect 15244 25180 15284 25220
rect 15244 24592 15284 24632
rect 13516 22744 13556 22784
rect 13708 22744 13748 22784
rect 13516 22576 13556 22616
rect 13708 21568 13748 21608
rect 11500 21484 11540 21524
rect 12076 21400 12116 21440
rect 12652 21400 12692 21440
rect 11308 20728 11348 20768
rect 11596 20476 11636 20516
rect 11212 19804 11252 19844
rect 10252 19132 10292 19172
rect 11020 19216 11060 19256
rect 11404 19720 11444 19760
rect 11116 19132 11156 19172
rect 11500 19216 11540 19256
rect 13132 21316 13172 21356
rect 12460 20056 12500 20096
rect 11692 19972 11732 20012
rect 12268 19888 12308 19928
rect 12748 19888 12788 19928
rect 12556 19720 12596 19760
rect 13132 20056 13172 20096
rect 13228 19972 13268 20012
rect 13708 20056 13748 20096
rect 13420 19804 13460 19844
rect 13324 19048 13364 19088
rect 10636 18880 10676 18920
rect 11404 18880 11444 18920
rect 10828 18376 10868 18416
rect 12076 17872 12116 17912
rect 11404 17788 11444 17828
rect 11788 17788 11828 17828
rect 10636 17704 10676 17744
rect 10348 15688 10388 15728
rect 13612 16360 13652 16400
rect 10924 15436 10964 15476
rect 9868 14848 9908 14888
rect 10060 14680 10100 14720
rect 8908 14260 8948 14300
rect 8620 14176 8660 14216
rect 7852 14008 7892 14048
rect 8044 14008 8084 14048
rect 6892 13252 6932 13292
rect 6700 13168 6740 13208
rect 6412 11908 6452 11948
rect 5836 11740 5876 11780
rect 6220 11740 6260 11780
rect 5740 11656 5780 11696
rect 5548 11572 5588 11612
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 4684 11152 4724 11192
rect 4108 10816 4148 10856
rect 3724 10396 3764 10436
rect 3724 8800 3764 8840
rect 3628 8716 3668 8756
rect 2860 8128 2900 8168
rect 3532 8632 3572 8672
rect 3532 8464 3572 8504
rect 3436 8044 3476 8084
rect 2860 7960 2900 8000
rect 3724 8632 3764 8672
rect 4204 10396 4244 10436
rect 3916 10228 3956 10268
rect 5260 10984 5300 11024
rect 4780 10648 4820 10688
rect 4684 10060 4724 10100
rect 3916 9976 3956 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4204 9472 4244 9512
rect 4876 10228 4916 10268
rect 5548 11152 5588 11192
rect 6604 11656 6644 11696
rect 6028 11488 6068 11528
rect 8044 13168 8084 13208
rect 6700 11488 6740 11528
rect 5932 11068 5972 11108
rect 5452 10816 5492 10856
rect 5356 10648 5396 10688
rect 4972 10144 5012 10184
rect 4876 9976 4916 10016
rect 5356 10144 5396 10184
rect 5260 9472 5300 9512
rect 4300 9388 4340 9428
rect 4588 9388 4628 9428
rect 4012 8884 4052 8924
rect 4108 8800 4148 8840
rect 4876 9304 4916 9344
rect 4972 8716 5012 8756
rect 2476 7792 2516 7832
rect 2860 7708 2900 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2764 7288 2804 7328
rect 3628 7708 3668 7748
rect 3532 6952 3572 6992
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4396 8044 4436 8084
rect 5068 8380 5108 8420
rect 4972 8044 5012 8084
rect 4012 7288 4052 7328
rect 2860 6448 2900 6488
rect 1036 5608 1076 5648
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4876 7960 4916 8000
rect 5932 10648 5972 10688
rect 6316 10648 6356 10688
rect 7084 11908 7124 11948
rect 6988 10396 7028 10436
rect 6316 10144 6356 10184
rect 6892 10144 6932 10184
rect 5836 9976 5876 10016
rect 8140 12496 8180 12536
rect 8044 11824 8084 11864
rect 7372 10984 7412 11024
rect 7180 9640 7220 9680
rect 5740 9304 5780 9344
rect 6988 9472 7028 9512
rect 6124 9388 6164 9428
rect 7276 9304 7316 9344
rect 7468 10396 7508 10436
rect 9772 14176 9812 14216
rect 9004 14092 9044 14132
rect 8812 13840 8852 13880
rect 10924 14680 10964 14720
rect 10444 14176 10484 14216
rect 10156 13840 10196 13880
rect 9292 13168 9332 13208
rect 10060 13168 10100 13208
rect 10252 13000 10292 13040
rect 8908 12916 8948 12956
rect 8044 11572 8084 11612
rect 7948 11488 7988 11528
rect 7852 11152 7892 11192
rect 7756 11068 7796 11108
rect 7564 10312 7604 10352
rect 8236 11404 8276 11444
rect 8620 11656 8660 11696
rect 10156 12832 10196 12872
rect 9004 12496 9044 12536
rect 8908 11824 8948 11864
rect 8812 11740 8852 11780
rect 8428 11572 8468 11612
rect 8332 11236 8372 11276
rect 8716 11236 8756 11276
rect 8140 10984 8180 11024
rect 7660 10228 7700 10268
rect 8428 10816 8468 10856
rect 8428 10396 8468 10436
rect 8620 10396 8660 10436
rect 8236 10144 8276 10184
rect 8524 10312 8564 10352
rect 8716 10144 8756 10184
rect 9676 12496 9716 12536
rect 9868 12328 9908 12368
rect 9772 11908 9812 11948
rect 9676 11740 9716 11780
rect 9388 11656 9428 11696
rect 9484 11488 9524 11528
rect 9196 11320 9236 11360
rect 9388 11320 9428 11360
rect 9100 11152 9140 11192
rect 8908 10984 8948 11024
rect 9292 10984 9332 11024
rect 10156 11740 10196 11780
rect 9964 11656 10004 11696
rect 9964 11404 10004 11444
rect 9580 11236 9620 11276
rect 9388 10732 9428 10772
rect 9292 10648 9332 10688
rect 8908 10396 8948 10436
rect 8812 10060 8852 10100
rect 7660 9556 7700 9596
rect 7372 9136 7412 9176
rect 7564 9136 7604 9176
rect 5932 8800 5972 8840
rect 6604 8632 6644 8672
rect 6796 8380 6836 8420
rect 6028 8296 6068 8336
rect 5356 7960 5396 8000
rect 5836 7960 5876 8000
rect 5260 7876 5300 7916
rect 4204 6952 4244 6992
rect 4588 6952 4628 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 4012 6448 4052 6488
rect 4492 6448 4532 6488
rect 4204 6280 4244 6320
rect 4780 5608 4820 5648
rect 4204 5440 4244 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 4972 6280 5012 6320
rect 3724 5020 3764 5060
rect 2956 4936 2996 4976
rect 4684 5104 4724 5144
rect 5164 6364 5204 6404
rect 5068 5440 5108 5480
rect 5164 5188 5204 5228
rect 5164 5020 5204 5060
rect 6028 7876 6068 7916
rect 5548 6784 5588 6824
rect 6028 6952 6068 6992
rect 7084 6448 7124 6488
rect 6028 6280 6068 6320
rect 6604 6280 6644 6320
rect 5452 5608 5492 5648
rect 4204 4852 4244 4892
rect 4684 4852 4724 4892
rect 652 4768 692 4808
rect 5548 4936 5588 4976
rect 6604 4936 6644 4976
rect 4300 4684 4340 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 5932 4684 5972 4724
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 5548 4096 5588 4136
rect 6796 6280 6836 6320
rect 7180 6196 7220 6236
rect 7468 8632 7508 8672
rect 7468 8128 7508 8168
rect 7468 7960 7508 8000
rect 7852 9220 7892 9260
rect 7756 9136 7796 9176
rect 7660 8800 7700 8840
rect 8044 9556 8084 9596
rect 8332 9472 8372 9512
rect 9100 10312 9140 10352
rect 9196 10144 9236 10184
rect 9676 10816 9716 10856
rect 9868 10984 9908 11024
rect 10156 11068 10196 11108
rect 10060 10732 10100 10772
rect 11212 15436 11252 15476
rect 11116 15268 11156 15308
rect 11500 15100 11540 15140
rect 11980 15100 12020 15140
rect 11308 14680 11348 14720
rect 12556 15268 12596 15308
rect 13228 15268 13268 15308
rect 13228 15016 13268 15056
rect 12268 14932 12308 14972
rect 11884 14848 11924 14888
rect 11500 14092 11540 14132
rect 11212 13000 11252 13040
rect 11404 12832 11444 12872
rect 12844 14848 12884 14888
rect 12844 14680 12884 14720
rect 12556 13924 12596 13964
rect 12460 13840 12500 13880
rect 12364 13672 12404 13712
rect 11692 13000 11732 13040
rect 10732 12496 10772 12536
rect 11692 12496 11732 12536
rect 11404 12328 11444 12368
rect 11980 13168 12020 13208
rect 12076 12580 12116 12620
rect 11308 12244 11348 12284
rect 11884 12244 11924 12284
rect 12556 13756 12596 13796
rect 14188 22492 14228 22532
rect 14764 22492 14804 22532
rect 15148 22912 15188 22952
rect 14956 22660 14996 22700
rect 13900 21484 13940 21524
rect 14668 22240 14708 22280
rect 15148 22240 15188 22280
rect 15628 25264 15668 25304
rect 15532 24004 15572 24044
rect 15436 23836 15476 23876
rect 15724 25180 15764 25220
rect 15724 24424 15764 24464
rect 15532 23080 15572 23120
rect 15532 22744 15572 22784
rect 15436 22660 15476 22700
rect 15340 22408 15380 22448
rect 15724 22912 15764 22952
rect 15628 22660 15668 22700
rect 15532 22156 15572 22196
rect 15148 20896 15188 20936
rect 14284 20056 14324 20096
rect 15916 25768 15956 25808
rect 16204 25432 16244 25472
rect 16396 25432 16436 25472
rect 15916 25180 15956 25220
rect 16972 26104 17012 26144
rect 17644 26188 17684 26228
rect 17836 26188 17876 26228
rect 17260 26020 17300 26060
rect 17644 25852 17684 25892
rect 16972 24844 17012 24884
rect 17740 25600 17780 25640
rect 17836 25516 17876 25556
rect 15916 23920 15956 23960
rect 16108 24592 16148 24632
rect 18124 26608 18164 26648
rect 18220 26104 18260 26144
rect 18124 26020 18164 26060
rect 19756 30640 19796 30680
rect 19948 30595 19988 30596
rect 19948 30556 19988 30595
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 19756 29296 19796 29336
rect 19372 28960 19412 29000
rect 19276 27784 19316 27824
rect 19468 28876 19508 28916
rect 19468 28624 19508 28664
rect 20524 29632 20564 29672
rect 20044 29296 20084 29336
rect 19756 28372 19796 28412
rect 19564 28288 19604 28328
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 19468 27784 19508 27824
rect 19084 27532 19124 27572
rect 18988 27364 19028 27404
rect 18796 26608 18836 26648
rect 18316 25852 18356 25892
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 18700 25516 18740 25556
rect 18508 25180 18548 25220
rect 18124 25096 18164 25136
rect 18316 25096 18356 25136
rect 18220 24760 18260 24800
rect 16972 24592 17012 24632
rect 17260 24592 17300 24632
rect 16300 24424 16340 24464
rect 16684 24172 16724 24212
rect 17068 24172 17108 24212
rect 16204 23920 16244 23960
rect 16204 23752 16244 23792
rect 16492 23752 16532 23792
rect 16108 23668 16148 23708
rect 16108 23500 16148 23540
rect 16012 23080 16052 23120
rect 15916 22912 15956 22952
rect 16396 23584 16436 23624
rect 16300 23080 16340 23120
rect 17932 24172 17972 24212
rect 18412 24592 18452 24632
rect 17548 23920 17588 23960
rect 17836 23836 17876 23876
rect 16972 23584 17012 23624
rect 17548 23752 17588 23792
rect 17740 23763 17780 23792
rect 17740 23752 17780 23763
rect 17548 23332 17588 23372
rect 16588 23164 16628 23204
rect 16204 22996 16244 23036
rect 16012 22576 16052 22616
rect 16204 22660 16244 22700
rect 16780 23080 16820 23120
rect 16876 22996 16916 23036
rect 17260 22660 17300 22700
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 18892 26524 18932 26564
rect 19084 26944 19124 26984
rect 20812 29044 20852 29084
rect 20140 28876 20180 28916
rect 21388 30724 21428 30764
rect 22060 31480 22100 31520
rect 22540 31480 22580 31520
rect 21868 30724 21908 30764
rect 21772 29800 21812 29840
rect 22348 31144 22388 31184
rect 23020 33664 23060 33704
rect 23884 33832 23924 33872
rect 23692 33496 23732 33536
rect 23596 32992 23636 33032
rect 23500 32824 23540 32864
rect 24844 34000 24884 34040
rect 24652 33916 24692 33956
rect 24076 33664 24116 33704
rect 24172 33580 24212 33620
rect 24076 33076 24116 33116
rect 23980 32992 24020 33032
rect 22732 31480 22772 31520
rect 23212 31480 23252 31520
rect 22924 31396 22964 31436
rect 22828 30220 22868 30260
rect 23020 31144 23060 31184
rect 23980 32824 24020 32864
rect 24172 32824 24212 32864
rect 25516 33664 25556 33704
rect 25804 33580 25844 33620
rect 25708 33496 25748 33536
rect 24844 33076 24884 33116
rect 24652 32824 24692 32864
rect 24364 32740 24404 32780
rect 25804 33244 25844 33284
rect 25708 32740 25748 32780
rect 26284 33664 26324 33704
rect 26668 35008 26708 35048
rect 27052 34336 27092 34376
rect 26476 33580 26516 33620
rect 26188 33496 26228 33536
rect 25900 32572 25940 32612
rect 25324 32152 25364 32192
rect 23884 31480 23924 31520
rect 23788 31396 23828 31436
rect 22636 29800 22676 29840
rect 22540 29296 22580 29336
rect 22636 29212 22676 29252
rect 21484 29128 21524 29168
rect 22540 29128 22580 29168
rect 23308 29380 23348 29420
rect 23116 29296 23156 29336
rect 23212 29128 23252 29168
rect 23500 29212 23540 29252
rect 20524 28288 20564 28328
rect 21100 28288 21140 28328
rect 19948 27700 19988 27740
rect 19564 27616 19604 27656
rect 20716 27700 20756 27740
rect 19372 26944 19412 26984
rect 20044 27196 20084 27236
rect 19564 26776 19604 26816
rect 20524 27028 20564 27068
rect 20620 26944 20660 26984
rect 20044 26692 20084 26732
rect 19180 26608 19220 26648
rect 19084 26524 19124 26564
rect 18796 23836 18836 23876
rect 18124 22996 18164 23036
rect 17452 22912 17492 22952
rect 17740 22912 17780 22952
rect 17644 22744 17684 22784
rect 17548 22576 17588 22616
rect 18988 23752 19028 23792
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 19372 26104 19412 26144
rect 19276 25264 19316 25304
rect 19180 25180 19220 25220
rect 20140 26188 20180 26228
rect 20428 26608 20468 26648
rect 20332 26104 20372 26144
rect 20236 25768 20276 25808
rect 21100 26272 21140 26312
rect 21100 25852 21140 25892
rect 19084 23584 19124 23624
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 21004 24592 21044 24632
rect 21196 24592 21236 24632
rect 20908 24256 20948 24296
rect 20812 23920 20852 23960
rect 22252 28876 22292 28916
rect 21868 28792 21908 28832
rect 23788 30220 23828 30260
rect 25228 31564 25268 31604
rect 25036 31480 25076 31520
rect 24940 31396 24980 31436
rect 23980 30640 24020 30680
rect 23884 29716 23924 29756
rect 24940 30472 24980 30512
rect 25996 32152 26036 32192
rect 26668 32740 26708 32780
rect 26668 32572 26708 32612
rect 26572 32236 26612 32276
rect 26188 32152 26228 32192
rect 26188 31984 26228 32024
rect 25900 31732 25940 31772
rect 25132 30472 25172 30512
rect 24172 29632 24212 29672
rect 24940 29632 24980 29672
rect 23788 28288 23828 28328
rect 23788 27700 23828 27740
rect 22828 27616 22868 27656
rect 23884 27616 23924 27656
rect 21676 27028 21716 27068
rect 23404 26944 23444 26984
rect 22156 26440 22196 26480
rect 21676 26104 21716 26144
rect 21484 25936 21524 25976
rect 21484 24340 21524 24380
rect 21580 23920 21620 23960
rect 19468 23752 19508 23792
rect 20716 23500 20756 23540
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 21580 23416 21620 23456
rect 19372 23332 19412 23372
rect 20812 23332 20852 23372
rect 18988 23164 19028 23204
rect 18700 22744 18740 22784
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 18220 22324 18260 22364
rect 17836 22240 17876 22280
rect 17548 22072 17588 22112
rect 18220 22156 18260 22196
rect 18700 22072 18740 22112
rect 19660 23080 19700 23120
rect 13804 19804 13844 19844
rect 14284 19804 14324 19844
rect 15820 19804 15860 19844
rect 14764 19216 14804 19256
rect 14380 19048 14420 19088
rect 13996 16360 14036 16400
rect 14188 16192 14228 16232
rect 14476 18040 14516 18080
rect 14764 17620 14804 17660
rect 14668 16192 14708 16232
rect 14764 15016 14804 15056
rect 13804 14932 13844 14972
rect 14092 14848 14132 14888
rect 13804 14092 13844 14132
rect 13228 14008 13268 14048
rect 13132 13840 13172 13880
rect 15244 19048 15284 19088
rect 15340 16360 15380 16400
rect 15052 16276 15092 16316
rect 14956 15268 14996 15308
rect 14860 14932 14900 14972
rect 14284 14680 14324 14720
rect 12748 13672 12788 13712
rect 14764 14008 14804 14048
rect 12940 13336 12980 13376
rect 12844 13168 12884 13208
rect 12460 13000 12500 13040
rect 12268 12244 12308 12284
rect 11116 11740 11156 11780
rect 10828 11656 10868 11696
rect 11404 11572 11444 11612
rect 11308 11152 11348 11192
rect 9772 10396 9812 10436
rect 9676 10312 9716 10352
rect 9772 10228 9812 10268
rect 9676 9976 9716 10016
rect 9292 9304 9332 9344
rect 9388 9136 9428 9176
rect 8332 8800 8372 8840
rect 9004 8800 9044 8840
rect 8044 8716 8084 8756
rect 8140 8128 8180 8168
rect 8908 8632 8948 8672
rect 8620 8380 8660 8420
rect 8524 8128 8564 8168
rect 7852 7960 7892 8000
rect 8044 7708 8084 7748
rect 8428 7708 8468 7748
rect 7948 6952 7988 6992
rect 8332 6952 8372 6992
rect 8716 7540 8756 7580
rect 8812 7372 8852 7412
rect 9868 10144 9908 10184
rect 9964 10060 10004 10100
rect 9772 9640 9812 9680
rect 9484 8800 9524 8840
rect 10636 10396 10676 10436
rect 10540 10144 10580 10184
rect 11308 10312 11348 10352
rect 10732 10144 10772 10184
rect 10252 9556 10292 9596
rect 9868 8632 9908 8672
rect 9676 8380 9716 8420
rect 9388 8128 9428 8168
rect 9004 7624 9044 7664
rect 9100 7540 9140 7580
rect 9292 7708 9332 7748
rect 9196 7204 9236 7244
rect 7468 6364 7508 6404
rect 7372 6280 7412 6320
rect 7468 5776 7508 5816
rect 7372 5608 7412 5648
rect 7468 5524 7508 5564
rect 7180 5440 7220 5480
rect 7372 4936 7412 4976
rect 8332 6616 8372 6656
rect 8428 6448 8468 6488
rect 8332 6364 8372 6404
rect 8236 6280 8276 6320
rect 7660 5608 7700 5648
rect 7948 5608 7988 5648
rect 8140 5608 8180 5648
rect 7756 5524 7796 5564
rect 8428 6280 8468 6320
rect 8716 6952 8756 6992
rect 8812 6532 8852 6572
rect 9004 6532 9044 6572
rect 9100 6448 9140 6488
rect 10060 8800 10100 8840
rect 9772 7960 9812 8000
rect 9580 7372 9620 7412
rect 9388 7288 9428 7328
rect 9388 7120 9428 7160
rect 9676 7120 9716 7160
rect 9772 6952 9812 6992
rect 9484 6868 9524 6908
rect 9580 6700 9620 6740
rect 9484 6448 9524 6488
rect 9196 6280 9236 6320
rect 9292 6196 9332 6236
rect 9004 5776 9044 5816
rect 6604 4096 6644 4136
rect 5356 3760 5396 3800
rect 6700 3928 6740 3968
rect 6796 3760 6836 3800
rect 652 3088 692 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 6604 3424 6644 3464
rect 844 2668 884 2708
rect 7756 4936 7796 4976
rect 8908 5524 8948 5564
rect 8428 5440 8468 5480
rect 9100 5440 9140 5480
rect 8812 5104 8852 5144
rect 7660 4012 7700 4052
rect 7468 3928 7508 3968
rect 7948 3760 7988 3800
rect 7756 3592 7796 3632
rect 7468 2668 7508 2708
rect 7180 2584 7220 2624
rect 7564 2584 7604 2624
rect 8140 3928 8180 3968
rect 8236 3508 8276 3548
rect 8716 4936 8756 4976
rect 9393 5608 9433 5648
rect 9676 6280 9716 6320
rect 9964 7960 10004 8000
rect 10252 8716 10292 8756
rect 10636 8716 10676 8756
rect 10156 8296 10196 8336
rect 10924 9556 10964 9596
rect 11884 11656 11924 11696
rect 11788 11404 11828 11444
rect 12172 11824 12212 11864
rect 12076 11488 12116 11528
rect 11692 10060 11732 10100
rect 12268 11404 12308 11444
rect 12172 11152 12212 11192
rect 12172 10144 12212 10184
rect 12940 12916 12980 12956
rect 12940 12580 12980 12620
rect 13612 12580 13652 12620
rect 13036 11656 13076 11696
rect 13324 11572 13364 11612
rect 13228 11488 13268 11528
rect 13900 10984 13940 11024
rect 11980 9976 12020 10016
rect 10732 8632 10772 8672
rect 11404 8632 11444 8672
rect 10540 7960 10580 8000
rect 10828 8296 10868 8336
rect 11116 8044 11156 8084
rect 11692 8632 11732 8672
rect 11596 8548 11636 8588
rect 11884 8548 11924 8588
rect 11692 8044 11732 8084
rect 12460 9976 12500 10016
rect 14092 13000 14132 13040
rect 14092 11824 14132 11864
rect 15628 15520 15668 15560
rect 15436 15100 15476 15140
rect 15340 14596 15380 14636
rect 16396 19720 16436 19760
rect 16108 19216 16148 19256
rect 15916 19048 15956 19088
rect 18892 21568 18932 21608
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 16972 19888 17012 19928
rect 16300 17620 16340 17660
rect 16108 17452 16148 17492
rect 16012 17200 16052 17240
rect 15916 17032 15956 17072
rect 16780 17032 16820 17072
rect 16012 16108 16052 16148
rect 16588 16192 16628 16232
rect 16972 18712 17012 18752
rect 16972 17536 17012 17576
rect 16972 16276 17012 16316
rect 16396 16108 16436 16148
rect 15820 15520 15860 15560
rect 16204 15520 16244 15560
rect 15724 15016 15764 15056
rect 15724 14680 15764 14720
rect 15820 14596 15860 14636
rect 15244 14092 15284 14132
rect 15820 14092 15860 14132
rect 15724 14008 15764 14048
rect 16300 14680 16340 14720
rect 17548 20056 17588 20096
rect 18316 20056 18356 20096
rect 17452 19972 17492 20012
rect 17356 19888 17396 19928
rect 17164 18964 17204 19004
rect 17452 18880 17492 18920
rect 17260 18796 17300 18836
rect 17356 18712 17396 18752
rect 18796 19972 18836 20012
rect 18988 20560 19028 20600
rect 18892 19888 18932 19928
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 18220 19216 18260 19256
rect 17644 18964 17684 19004
rect 18028 18880 18068 18920
rect 17644 18544 17684 18584
rect 17164 17788 17204 17828
rect 17452 18292 17492 18332
rect 17548 17872 17588 17912
rect 18220 18292 18260 18332
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 19180 19888 19220 19928
rect 19756 22408 19796 22448
rect 20332 22408 20372 22448
rect 21196 22240 21236 22280
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 21292 22072 21332 22112
rect 21964 26020 22004 26060
rect 22252 26020 22292 26060
rect 22060 25852 22100 25892
rect 22156 25600 22196 25640
rect 21772 25432 21812 25472
rect 22924 26272 22964 26312
rect 22636 26020 22676 26060
rect 22540 25936 22580 25976
rect 22348 25432 22388 25472
rect 23596 25516 23636 25556
rect 21868 24844 21908 24884
rect 21964 24424 22004 24464
rect 21772 24340 21812 24380
rect 21676 23080 21716 23120
rect 21484 21736 21524 21776
rect 21484 21400 21524 21440
rect 21676 21400 21716 21440
rect 21292 20980 21332 21020
rect 20524 20728 20564 20768
rect 21676 20812 21716 20852
rect 21388 20728 21428 20768
rect 21580 20742 21620 20768
rect 21580 20728 21620 20742
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 20620 20476 20660 20516
rect 20908 20392 20948 20432
rect 19468 20056 19508 20096
rect 19660 19972 19700 20012
rect 19372 19216 19412 19256
rect 21292 20560 21332 20600
rect 21484 20560 21524 20600
rect 21388 20308 21428 20348
rect 22156 25096 22196 25136
rect 23500 25348 23540 25388
rect 23596 25269 23636 25304
rect 23596 25264 23636 25269
rect 22732 25096 22772 25136
rect 22252 24844 22292 24884
rect 22252 24592 22292 24632
rect 22156 24508 22196 24548
rect 23020 23836 23060 23876
rect 21868 22072 21908 22112
rect 22060 20980 22100 21020
rect 21868 20644 21908 20684
rect 21772 20308 21812 20348
rect 21484 20224 21524 20264
rect 21676 20224 21716 20264
rect 21004 19972 21044 20012
rect 21292 19300 21332 19340
rect 19372 19048 19412 19088
rect 20332 19048 20372 19088
rect 19276 18964 19316 19004
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 19084 18712 19124 18752
rect 19276 18544 19316 18584
rect 19084 18460 19124 18500
rect 18988 18292 19028 18332
rect 18988 17956 19028 17996
rect 17740 17788 17780 17828
rect 17356 17452 17396 17492
rect 17164 17032 17204 17072
rect 17452 17284 17492 17324
rect 18508 17704 18548 17744
rect 18124 17620 18164 17660
rect 18412 17620 18452 17660
rect 18028 17368 18068 17408
rect 17836 17200 17876 17240
rect 17548 16780 17588 16820
rect 18316 17200 18356 17240
rect 18220 17032 18260 17072
rect 18124 16948 18164 16988
rect 18796 17788 18836 17828
rect 18988 17788 19028 17828
rect 18700 17368 18740 17408
rect 19276 18208 19316 18248
rect 21004 19048 21044 19088
rect 21100 18964 21140 19004
rect 20812 18880 20852 18920
rect 20716 18628 20756 18668
rect 20620 18544 20660 18584
rect 19756 18460 19796 18500
rect 20524 18460 20564 18500
rect 19468 18292 19508 18332
rect 19372 17956 19412 17996
rect 19276 17704 19316 17744
rect 20524 17956 20564 17996
rect 19660 17872 19700 17912
rect 21196 18628 21236 18668
rect 20908 18544 20948 18584
rect 20812 18208 20852 18248
rect 20716 18040 20756 18080
rect 19181 17620 19221 17660
rect 19372 17536 19412 17576
rect 19660 17536 19700 17576
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 18700 17200 18740 17240
rect 19084 17200 19124 17240
rect 18796 17116 18836 17156
rect 18892 17032 18932 17072
rect 18604 16780 18644 16820
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 18700 16360 18740 16400
rect 18028 16192 18068 16232
rect 19180 16276 19220 16316
rect 18700 16192 18740 16232
rect 16876 15520 16916 15560
rect 17644 15520 17684 15560
rect 16492 15100 16532 15140
rect 16684 14848 16724 14888
rect 16684 14680 16724 14720
rect 16972 14680 17012 14720
rect 16492 14176 16532 14216
rect 14476 11740 14516 11780
rect 13420 10144 13460 10184
rect 13228 10060 13268 10100
rect 12268 8632 12308 8672
rect 13612 9304 13652 9344
rect 13900 8716 13940 8756
rect 11500 7540 11540 7580
rect 11692 7540 11732 7580
rect 12940 7540 12980 7580
rect 13132 7540 13172 7580
rect 10156 6784 10196 6824
rect 10060 6700 10100 6740
rect 10156 6616 10196 6656
rect 9868 5776 9908 5816
rect 10252 6448 10292 6488
rect 11404 6952 11444 6992
rect 11116 6616 11156 6656
rect 12076 7120 12116 7160
rect 12844 7120 12884 7160
rect 13996 8632 14036 8672
rect 14284 11404 14324 11444
rect 15340 12580 15380 12620
rect 15532 11656 15572 11696
rect 15436 10228 15476 10268
rect 16204 14008 16244 14048
rect 16204 13336 16244 13376
rect 16684 13252 16724 13292
rect 16396 12580 16436 12620
rect 16108 11656 16148 11696
rect 16876 13168 16916 13208
rect 16780 12496 16820 12536
rect 16588 12328 16628 12368
rect 16780 11824 16820 11864
rect 16300 11152 16340 11192
rect 17644 15016 17684 15056
rect 17548 14680 17588 14720
rect 17164 14176 17204 14216
rect 17068 14008 17108 14048
rect 17164 13924 17204 13964
rect 17068 11656 17108 11696
rect 17068 11488 17108 11528
rect 17452 14008 17492 14048
rect 18604 16024 18644 16064
rect 18508 15520 18548 15560
rect 21100 17872 21140 17912
rect 20812 17788 20852 17828
rect 20908 17704 20948 17744
rect 21292 18544 21332 18584
rect 21388 18376 21428 18416
rect 21388 18040 21428 18080
rect 21772 18880 21812 18920
rect 21964 20392 22004 20432
rect 22060 20224 22100 20264
rect 22156 20056 22196 20096
rect 21964 19972 22004 20012
rect 22444 22660 22484 22700
rect 22348 22492 22388 22532
rect 22540 22072 22580 22112
rect 23692 24844 23732 24884
rect 23788 23920 23828 23960
rect 25324 29716 25364 29756
rect 25516 29296 25556 29336
rect 25132 29128 25172 29168
rect 26476 31732 26516 31772
rect 26380 31564 26420 31604
rect 26476 30640 26516 30680
rect 25708 30220 25748 30260
rect 25708 29800 25748 29840
rect 25900 29632 25940 29672
rect 25996 29380 26036 29420
rect 25804 29128 25844 29168
rect 25228 29044 25268 29084
rect 24748 27616 24788 27656
rect 25324 27616 25364 27656
rect 25228 27532 25268 27572
rect 23980 26944 24020 26984
rect 24172 25264 24212 25304
rect 24076 24760 24116 24800
rect 23404 23584 23444 23624
rect 23212 22660 23252 22700
rect 23212 22492 23252 22532
rect 23884 23836 23924 23876
rect 24172 23080 24212 23120
rect 23788 22660 23828 22700
rect 25708 28288 25748 28328
rect 25612 27700 25652 27740
rect 25900 27616 25940 27656
rect 27148 34000 27188 34040
rect 28204 34000 28244 34040
rect 30028 34336 30068 34376
rect 29068 34000 29108 34040
rect 28972 33832 29012 33872
rect 27052 32908 27092 32948
rect 27436 32824 27476 32864
rect 27244 32236 27284 32276
rect 27052 31984 27092 32024
rect 26956 31480 26996 31520
rect 27340 31312 27380 31352
rect 27532 32152 27572 32192
rect 26764 30724 26804 30764
rect 26668 30472 26708 30512
rect 26572 30220 26612 30260
rect 27052 30640 27092 30680
rect 27244 30724 27284 30764
rect 27532 30472 27572 30512
rect 28588 33496 28628 33536
rect 29068 33664 29108 33704
rect 29164 33496 29204 33536
rect 28876 33328 28916 33368
rect 28108 33244 28148 33284
rect 28588 32908 28628 32948
rect 28492 32824 28532 32864
rect 27724 32740 27764 32780
rect 28108 31312 28148 31352
rect 28780 32824 28820 32864
rect 29452 33328 29492 33368
rect 29260 32824 29300 32864
rect 28684 31900 28724 31940
rect 29356 31900 29396 31940
rect 29644 32908 29684 32948
rect 30508 34336 30548 34376
rect 30220 33832 30260 33872
rect 30796 33832 30836 33872
rect 31276 34588 31316 34628
rect 31660 34588 31700 34628
rect 32140 34588 32180 34628
rect 30988 33832 31028 33872
rect 30220 32908 30260 32948
rect 29644 31396 29684 31436
rect 30316 32320 30356 32360
rect 30700 32320 30740 32360
rect 30124 31480 30164 31520
rect 30028 31396 30068 31436
rect 29932 31312 29972 31352
rect 28204 30472 28244 30512
rect 26380 29632 26420 29672
rect 26668 29548 26708 29588
rect 26572 29296 26612 29336
rect 26860 29212 26900 29252
rect 26764 29128 26804 29168
rect 25612 27028 25652 27068
rect 25036 26524 25076 26564
rect 24844 26104 24884 26144
rect 24748 25516 24788 25556
rect 25132 25600 25172 25640
rect 24940 25264 24980 25304
rect 24556 24760 24596 24800
rect 24364 24592 24404 24632
rect 27052 27700 27092 27740
rect 26380 27028 26420 27068
rect 26188 26860 26228 26900
rect 25996 26776 26036 26816
rect 25516 26608 25556 26648
rect 25900 26524 25940 26564
rect 26956 27028 26996 27068
rect 26572 26776 26612 26816
rect 27052 26860 27092 26900
rect 27340 30136 27380 30176
rect 27436 29800 27476 29840
rect 27724 29632 27764 29672
rect 27436 29128 27476 29168
rect 27628 29128 27668 29168
rect 27340 29044 27380 29084
rect 27820 29044 27860 29084
rect 28108 29128 28148 29168
rect 28300 28540 28340 28580
rect 28396 28456 28436 28496
rect 29836 30220 29876 30260
rect 29260 29632 29300 29672
rect 30796 32152 30836 32192
rect 30604 31480 30644 31520
rect 30700 31312 30740 31352
rect 30028 30220 30068 30260
rect 29164 29044 29204 29084
rect 29932 28876 29972 28916
rect 29740 28540 29780 28580
rect 28684 28288 28724 28328
rect 29068 28288 29108 28328
rect 29452 28288 29492 28328
rect 27436 27532 27476 27572
rect 27916 27196 27956 27236
rect 28684 27532 28724 27572
rect 29836 27700 29876 27740
rect 29260 27532 29300 27572
rect 26572 26608 26612 26648
rect 27532 26356 27572 26396
rect 28492 27196 28532 27236
rect 28876 26944 28916 26984
rect 28108 26860 28148 26900
rect 28780 26860 28820 26900
rect 28012 26776 28052 26816
rect 28108 26524 28148 26564
rect 27916 26188 27956 26228
rect 25324 25768 25364 25808
rect 26860 26104 26900 26144
rect 26476 25432 26516 25472
rect 26380 25264 26420 25304
rect 26956 25768 26996 25808
rect 26188 25180 26228 25220
rect 26092 24760 26132 24800
rect 26572 25180 26612 25220
rect 25708 24592 25748 24632
rect 26476 24676 26516 24716
rect 25516 24088 25556 24128
rect 25228 23920 25268 23960
rect 24364 22660 24404 22700
rect 24268 22324 24308 22364
rect 24172 22240 24212 22280
rect 23116 21736 23156 21776
rect 22540 21568 22580 21608
rect 22636 21400 22676 21440
rect 22540 20980 22580 21020
rect 22540 20812 22580 20852
rect 23404 21400 23444 21440
rect 23116 21064 23156 21104
rect 22636 20728 22676 20768
rect 22540 20056 22580 20096
rect 23020 20896 23060 20936
rect 23212 20812 23252 20852
rect 22732 20392 22772 20432
rect 23308 20728 23348 20768
rect 23596 21316 23636 21356
rect 23980 21568 24020 21608
rect 23788 21064 23828 21104
rect 23500 20896 23540 20936
rect 24460 21484 24500 21524
rect 24268 21316 24308 21356
rect 24268 21148 24308 21188
rect 24268 20728 24308 20768
rect 22636 19972 22676 20012
rect 22444 19048 22484 19088
rect 21868 18628 21908 18668
rect 22444 18628 22484 18668
rect 22636 18796 22676 18836
rect 23404 20056 23444 20096
rect 23308 19552 23348 19592
rect 23212 19300 23252 19340
rect 24172 20392 24212 20432
rect 23692 19300 23732 19340
rect 24076 19972 24116 20012
rect 23980 19552 24020 19592
rect 24268 20140 24308 20180
rect 25420 23752 25460 23792
rect 26188 24592 26228 24632
rect 26860 25264 26900 25304
rect 27916 25516 27956 25556
rect 27244 25264 27284 25304
rect 27340 24844 27380 24884
rect 27244 24592 27284 24632
rect 26956 24508 26996 24548
rect 27436 24676 27476 24716
rect 27340 24508 27380 24548
rect 26188 23920 26228 23960
rect 26764 23920 26804 23960
rect 26092 23752 26132 23792
rect 26572 23752 26612 23792
rect 25036 21736 25076 21776
rect 24652 21568 24692 21608
rect 25132 21568 25172 21608
rect 24940 21484 24980 21524
rect 25324 21484 25364 21524
rect 24844 20896 24884 20936
rect 24556 20560 24596 20600
rect 25036 20308 25076 20348
rect 24460 20140 24500 20180
rect 24940 20056 24980 20096
rect 24364 19888 24404 19928
rect 25804 21568 25844 21608
rect 25516 21148 25556 21188
rect 25228 19468 25268 19508
rect 25708 20308 25748 20348
rect 25612 20140 25652 20180
rect 25516 20056 25556 20096
rect 25324 19300 25364 19340
rect 24364 19216 24404 19256
rect 25036 19216 25076 19256
rect 25228 19216 25268 19256
rect 24268 19132 24308 19172
rect 23692 19048 23732 19088
rect 23884 19048 23924 19088
rect 22828 18964 22868 19004
rect 22060 18376 22100 18416
rect 21580 18124 21620 18164
rect 21580 17956 21620 17996
rect 21484 17788 21524 17828
rect 21388 17704 21428 17744
rect 21964 17788 22004 17828
rect 21868 17704 21908 17744
rect 20044 17116 20084 17156
rect 20428 16360 20468 16400
rect 20236 16276 20276 16316
rect 19948 16192 19988 16232
rect 20140 16192 20180 16232
rect 20908 16276 20948 16316
rect 19180 16024 19220 16064
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 18700 15604 18740 15644
rect 18700 15268 18740 15308
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 18604 14932 18644 14972
rect 17644 14176 17684 14216
rect 18508 14680 18548 14720
rect 18700 14680 18740 14720
rect 18892 15436 18932 15476
rect 18988 15268 19028 15308
rect 19276 15520 19316 15560
rect 19468 15352 19508 15392
rect 19756 15268 19796 15308
rect 19276 15100 19316 15140
rect 19756 15100 19796 15140
rect 18988 14848 19028 14888
rect 18892 14680 18932 14720
rect 19180 14848 19220 14888
rect 19372 14680 19412 14720
rect 20140 15688 20180 15728
rect 20140 15520 20180 15560
rect 19948 15184 19988 15224
rect 19852 14764 19892 14804
rect 20140 14764 20180 14804
rect 19084 14596 19124 14636
rect 18796 14428 18836 14468
rect 19276 14428 19316 14468
rect 18412 14176 18452 14216
rect 18988 14176 19028 14216
rect 17932 14008 17972 14048
rect 17356 13168 17396 13208
rect 17644 13252 17684 13292
rect 17548 12580 17588 12620
rect 17452 12244 17492 12284
rect 17740 12580 17780 12620
rect 17740 12160 17780 12200
rect 17740 11908 17780 11948
rect 17644 11656 17684 11696
rect 18124 13924 18164 13964
rect 18700 14092 18740 14132
rect 18604 14008 18644 14048
rect 18508 13840 18548 13880
rect 18700 13840 18740 13880
rect 17932 12832 17972 12872
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18412 13168 18452 13208
rect 18220 12832 18260 12872
rect 18124 12748 18164 12788
rect 18028 12580 18068 12620
rect 17932 12496 17972 12536
rect 18316 12664 18356 12704
rect 18700 13168 18740 13208
rect 19180 14008 19220 14048
rect 19084 13840 19124 13880
rect 18892 13420 18932 13460
rect 19084 13336 19124 13376
rect 19948 14680 19988 14720
rect 19948 14512 19988 14552
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 20044 14260 20084 14300
rect 19660 14176 19700 14216
rect 19948 14176 19988 14216
rect 19372 14008 19412 14048
rect 20044 14092 20084 14132
rect 19948 13840 19988 13880
rect 19468 13420 19508 13460
rect 18604 12748 18644 12788
rect 18220 12412 18260 12452
rect 18508 12412 18548 12452
rect 18028 12244 18068 12284
rect 19756 13252 19796 13292
rect 19948 13336 19988 13376
rect 20140 13336 20180 13376
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 19564 12664 19604 12704
rect 19372 12580 19412 12620
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 20140 13000 20180 13040
rect 20044 12832 20084 12872
rect 20044 12664 20084 12704
rect 19084 12328 19124 12368
rect 18316 11656 18356 11696
rect 17356 11404 17396 11444
rect 17260 11320 17300 11360
rect 17644 11236 17684 11276
rect 16780 10396 16820 10436
rect 15532 9808 15572 9848
rect 15916 9808 15956 9848
rect 14860 9052 14900 9092
rect 15148 9052 15188 9092
rect 14668 8632 14708 8672
rect 15724 9640 15764 9680
rect 16012 9640 16052 9680
rect 15628 9472 15668 9512
rect 16588 9976 16628 10016
rect 16396 9724 16436 9764
rect 16492 9556 16532 9596
rect 16492 9052 16532 9092
rect 16012 8632 16052 8672
rect 16396 8632 16436 8672
rect 15916 8380 15956 8420
rect 15820 8128 15860 8168
rect 14380 7960 14420 8000
rect 11884 6448 11924 6488
rect 12940 6448 12980 6488
rect 10060 6280 10100 6320
rect 9388 5356 9428 5396
rect 9196 5104 9236 5144
rect 9196 4936 9236 4976
rect 8812 4852 8852 4892
rect 9004 4600 9044 4640
rect 8812 3928 8852 3968
rect 8716 3592 8756 3632
rect 9004 3760 9044 3800
rect 9772 5440 9812 5480
rect 9676 5356 9716 5396
rect 9580 5020 9620 5060
rect 9676 4936 9716 4976
rect 9196 3928 9236 3968
rect 9196 3760 9236 3800
rect 9676 3760 9716 3800
rect 8908 3340 8948 3380
rect 9388 3424 9428 3464
rect 8236 2836 8276 2876
rect 9196 2836 9236 2876
rect 9868 4264 9908 4304
rect 11980 5608 12020 5648
rect 10156 4936 10196 4976
rect 10060 4768 10100 4808
rect 10348 5020 10388 5060
rect 10540 4936 10580 4976
rect 10444 4852 10484 4892
rect 10348 4768 10388 4808
rect 11596 4768 11636 4808
rect 11596 4348 11636 4388
rect 10252 4264 10292 4304
rect 10540 4264 10580 4304
rect 11020 4264 11060 4304
rect 11500 4264 11540 4304
rect 10444 4180 10484 4220
rect 10924 4180 10964 4220
rect 9964 3760 10004 3800
rect 10252 3928 10292 3968
rect 10156 3760 10196 3800
rect 10060 3592 10100 3632
rect 9772 3340 9812 3380
rect 11404 4180 11444 4220
rect 12172 5524 12212 5564
rect 11788 4264 11828 4304
rect 11980 4264 12020 4304
rect 11884 4180 11924 4220
rect 11788 4096 11828 4136
rect 12172 4180 12212 4220
rect 10636 3844 10676 3884
rect 11116 3928 11156 3968
rect 11308 3592 11348 3632
rect 10828 3508 10868 3548
rect 12076 3760 12116 3800
rect 12748 3760 12788 3800
rect 12940 5524 12980 5564
rect 13132 5608 13172 5648
rect 14188 5440 14228 5480
rect 13036 5104 13076 5144
rect 13324 4936 13364 4976
rect 14188 4768 14228 4808
rect 13420 4264 13460 4304
rect 13132 4096 13172 4136
rect 13324 4096 13364 4136
rect 13612 4096 13652 4136
rect 14092 3592 14132 3632
rect 14380 7708 14420 7748
rect 14668 6952 14708 6992
rect 15628 6952 15668 6992
rect 14668 6448 14708 6488
rect 16204 7708 16244 7748
rect 16108 6868 16148 6908
rect 15820 5860 15860 5900
rect 15532 5524 15572 5564
rect 16300 6616 16340 6656
rect 16204 5776 16244 5816
rect 16396 6448 16436 6488
rect 16012 5020 16052 5060
rect 15340 4096 15380 4136
rect 15052 4012 15092 4052
rect 15724 3928 15764 3968
rect 14668 3592 14708 3632
rect 16204 5356 16244 5396
rect 16108 4936 16148 4976
rect 16396 5104 16436 5144
rect 16396 4852 16436 4892
rect 16396 4432 16436 4472
rect 16396 4180 16436 4220
rect 16108 4012 16148 4052
rect 16300 3844 16340 3884
rect 15916 3592 15956 3632
rect 16300 3424 16340 3464
rect 16780 9976 16820 10016
rect 16972 10984 17012 11024
rect 17068 9808 17108 9848
rect 16972 9724 17012 9764
rect 17260 9640 17300 9680
rect 17548 10984 17588 11024
rect 17452 10816 17492 10856
rect 17932 11068 17972 11108
rect 17740 10900 17780 10940
rect 17644 10396 17684 10436
rect 17740 10144 17780 10184
rect 18124 11320 18164 11360
rect 18796 11656 18836 11696
rect 18028 10984 18068 11024
rect 18604 11152 18644 11192
rect 18796 10816 18836 10856
rect 18412 10732 18452 10772
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 18220 10396 18260 10436
rect 18700 10396 18740 10436
rect 18604 10312 18644 10352
rect 17356 9556 17396 9596
rect 16780 9472 16820 9512
rect 16684 9220 16724 9260
rect 17068 9472 17108 9512
rect 17260 9220 17300 9260
rect 17548 9472 17588 9512
rect 17740 9472 17780 9512
rect 17644 9304 17684 9344
rect 16972 8464 17012 8504
rect 17356 8632 17396 8672
rect 17260 8380 17300 8420
rect 16588 8212 16628 8252
rect 17068 8212 17108 8252
rect 17836 8800 17876 8840
rect 18028 9304 18068 9344
rect 18508 10060 18548 10100
rect 18316 9472 18356 9512
rect 18220 9304 18260 9344
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 19180 12076 19220 12116
rect 19180 11488 19220 11528
rect 20812 16192 20852 16232
rect 20908 16024 20948 16064
rect 20428 15520 20468 15560
rect 20620 15100 20660 15140
rect 20908 15520 20948 15560
rect 20812 15352 20852 15392
rect 20716 14932 20756 14972
rect 21100 16780 21140 16820
rect 21676 17032 21716 17072
rect 22252 17704 22292 17744
rect 22732 18544 22772 18584
rect 22636 18376 22676 18416
rect 22828 17704 22868 17744
rect 23788 17704 23828 17744
rect 22540 17620 22580 17660
rect 21580 16360 21620 16400
rect 22156 17032 22196 17072
rect 23884 17116 23924 17156
rect 22636 16948 22676 16988
rect 22924 16696 22964 16736
rect 21676 16192 21716 16232
rect 21580 16024 21620 16064
rect 21196 15688 21236 15728
rect 21868 15520 21908 15560
rect 22060 16360 22100 16400
rect 21772 15436 21812 15476
rect 21388 15184 21428 15224
rect 21292 14932 21332 14972
rect 20620 14764 20660 14804
rect 20428 14680 20468 14720
rect 20428 13924 20468 13964
rect 20332 13672 20372 13712
rect 20620 14512 20660 14552
rect 21196 14596 21236 14636
rect 21004 14428 21044 14468
rect 20716 14092 20756 14132
rect 21100 14176 21140 14216
rect 21105 13840 21145 13880
rect 20908 13756 20948 13796
rect 20812 13672 20852 13712
rect 20524 13420 20564 13460
rect 20908 13336 20948 13376
rect 20716 13252 20756 13292
rect 20332 13000 20372 13040
rect 20236 12832 20276 12872
rect 19948 12328 19988 12368
rect 20908 12832 20948 12872
rect 20620 12748 20660 12788
rect 20812 12580 20852 12620
rect 19468 12244 19508 12284
rect 20428 12244 20468 12284
rect 20716 12076 20756 12116
rect 20236 11992 20276 12032
rect 20908 11992 20948 12032
rect 20524 11908 20564 11948
rect 20908 11824 20948 11864
rect 20620 11740 20660 11780
rect 20777 11740 20817 11780
rect 20332 11656 20372 11696
rect 19756 11488 19796 11528
rect 20716 11488 20756 11528
rect 20524 11404 20564 11444
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 20428 11320 20468 11360
rect 19276 11236 19316 11276
rect 19084 11068 19124 11108
rect 19564 11068 19604 11108
rect 19468 10984 19508 11024
rect 19756 10984 19796 11024
rect 20812 11068 20852 11108
rect 21580 14848 21620 14888
rect 21484 14680 21524 14720
rect 21868 14596 21908 14636
rect 21772 14428 21812 14468
rect 21676 14092 21716 14132
rect 21388 14008 21428 14048
rect 21388 13840 21428 13880
rect 21580 13840 21620 13880
rect 21100 13672 21140 13712
rect 22156 15436 22196 15476
rect 22252 15268 22292 15308
rect 22060 14512 22100 14552
rect 21964 14260 22004 14300
rect 21868 13924 21908 13964
rect 21388 13336 21428 13376
rect 21100 12916 21140 12956
rect 21676 12664 21716 12704
rect 21292 12580 21332 12620
rect 21100 12412 21140 12452
rect 21292 12412 21332 12452
rect 21004 11740 21044 11780
rect 21196 11656 21236 11696
rect 21772 12496 21812 12536
rect 21388 12328 21428 12368
rect 21868 12328 21908 12368
rect 22348 14764 22388 14804
rect 22444 14680 22484 14720
rect 22348 14512 22388 14552
rect 22252 14428 22292 14468
rect 22636 14260 22676 14300
rect 22252 13924 22292 13964
rect 22444 13168 22484 13208
rect 22348 12496 22388 12536
rect 22252 12328 22292 12368
rect 22156 12160 22196 12200
rect 22348 12160 22388 12200
rect 21388 11824 21428 11864
rect 21641 11740 21681 11780
rect 22156 11740 22196 11780
rect 21292 11236 21332 11276
rect 19660 10816 19700 10856
rect 18988 10396 19028 10436
rect 19372 10480 19412 10520
rect 19276 10144 19316 10184
rect 19756 10732 19796 10772
rect 20620 10648 20660 10688
rect 20332 10312 20372 10352
rect 20236 10144 20276 10184
rect 18796 9724 18836 9764
rect 19084 9892 19124 9932
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 20332 9808 20372 9848
rect 18892 8800 18932 8840
rect 18316 8632 18356 8672
rect 17836 8212 17876 8252
rect 16588 7456 16628 7496
rect 16876 7204 16916 7244
rect 16876 6952 16916 6992
rect 16780 6448 16820 6488
rect 16684 5776 16724 5816
rect 16780 5608 16820 5648
rect 17260 7960 17300 8000
rect 17644 7456 17684 7496
rect 17548 7120 17588 7160
rect 17356 7036 17396 7076
rect 17164 6868 17204 6908
rect 17452 6784 17492 6824
rect 16982 5692 17022 5732
rect 16972 5356 17012 5396
rect 17260 6112 17300 6152
rect 17356 5944 17396 5984
rect 17452 5860 17492 5900
rect 18508 8044 18548 8084
rect 17932 7036 17972 7076
rect 17836 6700 17876 6740
rect 18796 8464 18836 8504
rect 20140 9136 20180 9176
rect 19084 8632 19124 8672
rect 19756 8632 19796 8672
rect 19852 8464 19892 8504
rect 20044 8380 20084 8420
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 20332 9136 20372 9176
rect 20524 10144 20564 10184
rect 20716 10480 20756 10520
rect 20620 10060 20660 10100
rect 20812 10060 20852 10100
rect 20919 10060 20959 10100
rect 21004 9640 21044 9680
rect 20428 8968 20468 9008
rect 20332 8464 20372 8504
rect 20236 8296 20276 8336
rect 20428 8380 20468 8420
rect 20332 8212 20372 8252
rect 18892 7960 18932 8000
rect 20332 8044 20372 8084
rect 20236 7876 20276 7916
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 18700 7540 18740 7580
rect 18508 7372 18548 7412
rect 18508 7204 18548 7244
rect 18700 7120 18740 7160
rect 18988 7120 19028 7160
rect 18796 6952 18836 6992
rect 17932 6196 17972 6236
rect 17548 5608 17588 5648
rect 16588 4180 16628 4220
rect 16492 4096 16532 4136
rect 17932 5272 17972 5312
rect 18124 6364 18164 6404
rect 18892 6532 18932 6572
rect 17068 5020 17108 5060
rect 17260 5020 17300 5060
rect 17548 4852 17588 4892
rect 17260 4348 17300 4388
rect 17164 4264 17204 4304
rect 17356 4264 17396 4304
rect 16492 3592 16532 3632
rect 17068 3508 17108 3548
rect 15820 3256 15860 3296
rect 15724 3088 15764 3128
rect 14284 2752 14324 2792
rect 11404 2668 11444 2708
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16300 2836 16340 2876
rect 16588 2752 16628 2792
rect 16108 2584 16148 2624
rect 16396 2500 16436 2540
rect 16780 2836 16820 2876
rect 17740 5104 17780 5144
rect 17836 5020 17876 5060
rect 17740 4852 17780 4892
rect 17836 4768 17876 4808
rect 17740 4348 17780 4388
rect 17644 4264 17684 4304
rect 17836 4264 17876 4304
rect 18028 4936 18068 4976
rect 17548 4012 17588 4052
rect 17452 3928 17492 3968
rect 17836 3928 17876 3968
rect 17740 3844 17780 3884
rect 17548 3760 17588 3800
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 18892 5860 18932 5900
rect 19180 6952 19220 6992
rect 19084 6448 19124 6488
rect 19276 6868 19316 6908
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 19468 6616 19508 6656
rect 19756 6616 19796 6656
rect 19852 6364 19892 6404
rect 19564 6112 19604 6152
rect 19756 6112 19796 6152
rect 18988 5776 19028 5816
rect 18508 5440 18548 5480
rect 18604 5188 18644 5228
rect 18892 5440 18932 5480
rect 19180 5860 19220 5900
rect 19276 5776 19316 5816
rect 19084 5356 19124 5396
rect 19948 5944 19988 5984
rect 19852 5776 19892 5816
rect 19660 5608 19700 5648
rect 20044 5776 20084 5816
rect 19372 5272 19412 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 18892 5020 18932 5060
rect 18700 4684 18740 4724
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 18508 4348 18548 4388
rect 18220 4180 18260 4220
rect 18412 4180 18452 4220
rect 18988 4852 19028 4892
rect 19084 4180 19124 4220
rect 18700 4012 18740 4052
rect 18508 3928 18548 3968
rect 18892 3844 18932 3884
rect 18028 3760 18068 3800
rect 17932 3676 17972 3716
rect 18124 3676 18164 3716
rect 17836 3508 17876 3548
rect 18028 3508 18068 3548
rect 17740 3004 17780 3044
rect 17452 2752 17492 2792
rect 16876 2584 16916 2624
rect 16684 2248 16724 2288
rect 17260 2668 17300 2708
rect 17164 2586 17204 2624
rect 17164 2584 17204 2586
rect 17068 2500 17108 2540
rect 17164 2416 17204 2456
rect 16492 2164 16532 2204
rect 16012 2080 16052 2120
rect 16492 1996 16532 2036
rect 16876 1996 16916 2036
rect 17068 1996 17108 2036
rect 17356 2500 17396 2540
rect 17644 2584 17684 2624
rect 17548 2416 17588 2456
rect 17356 2164 17396 2204
rect 17260 1996 17300 2036
rect 16492 1660 16532 1700
rect 16780 1660 16820 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 17548 2248 17588 2288
rect 18028 3004 18068 3044
rect 17932 2836 17972 2876
rect 19276 4936 19316 4976
rect 19372 4768 19412 4808
rect 20140 4852 20180 4892
rect 20236 4432 20276 4472
rect 20428 7960 20468 8000
rect 20428 7792 20468 7832
rect 20812 9472 20852 9512
rect 20812 9304 20852 9344
rect 20716 8884 20756 8924
rect 20620 8548 20660 8588
rect 20620 8380 20660 8420
rect 21004 9052 21044 9092
rect 20908 8800 20948 8840
rect 22636 11572 22676 11612
rect 21484 11404 21524 11444
rect 22348 10900 22388 10940
rect 21580 10312 21620 10352
rect 22156 10312 22196 10352
rect 21388 9388 21428 9428
rect 21292 9052 21332 9092
rect 21484 8632 21524 8672
rect 22060 10228 22100 10268
rect 21868 10144 21908 10184
rect 22252 10144 22292 10184
rect 22636 10396 22676 10436
rect 21964 9640 22004 9680
rect 21964 9304 22004 9344
rect 21964 8884 22004 8924
rect 21868 8716 21908 8756
rect 20908 8464 20948 8504
rect 21100 8464 21140 8504
rect 20620 7876 20660 7916
rect 20812 7876 20852 7916
rect 20524 7624 20564 7664
rect 20428 7372 20468 7412
rect 21196 8128 21236 8168
rect 21100 8044 21140 8084
rect 21004 7792 21044 7832
rect 21580 8464 21620 8504
rect 22060 8296 22100 8336
rect 21676 8128 21716 8168
rect 21484 7960 21524 8000
rect 20524 7120 20564 7160
rect 20620 7036 20660 7076
rect 20524 6448 20564 6488
rect 20812 7120 20852 7160
rect 21004 7036 21044 7076
rect 20812 6112 20852 6152
rect 21388 7036 21428 7076
rect 22540 9472 22580 9512
rect 22732 9640 22772 9680
rect 23020 16192 23060 16232
rect 22924 15016 22964 15056
rect 22924 14512 22964 14552
rect 22924 14092 22964 14132
rect 23884 16192 23924 16232
rect 24268 18796 24308 18836
rect 24172 18544 24212 18584
rect 24172 17704 24212 17744
rect 24460 18796 24500 18836
rect 24844 18796 24884 18836
rect 24652 18544 24692 18584
rect 24460 18376 24500 18416
rect 24364 17704 24404 17744
rect 24844 17872 24884 17912
rect 23692 15268 23732 15308
rect 23116 14764 23156 14804
rect 23020 13168 23060 13208
rect 23308 13168 23348 13208
rect 24748 17200 24788 17240
rect 25708 19468 25748 19508
rect 25996 19888 26036 19928
rect 25996 19300 26036 19340
rect 26572 21568 26612 21608
rect 26188 19972 26228 20012
rect 26572 20056 26612 20096
rect 26860 19804 26900 19844
rect 26476 19300 26516 19340
rect 26188 19216 26228 19256
rect 27340 23668 27380 23708
rect 27052 23080 27092 23120
rect 27052 22660 27092 22700
rect 28588 26608 28628 26648
rect 28492 26272 28532 26312
rect 28492 26104 28532 26144
rect 28684 26440 28724 26480
rect 28972 26860 29012 26900
rect 28876 26524 28916 26564
rect 29068 26524 29108 26564
rect 29644 27364 29684 27404
rect 29548 26776 29588 26816
rect 29836 27028 29876 27068
rect 29356 26608 29396 26648
rect 30220 28372 30260 28412
rect 30028 27616 30068 27656
rect 30412 30388 30452 30428
rect 30412 29548 30452 29588
rect 30412 29044 30452 29084
rect 30700 28960 30740 29000
rect 30892 30388 30932 30428
rect 31084 33664 31124 33704
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 33484 34336 33524 34376
rect 33772 34336 33812 34376
rect 34156 34336 34196 34376
rect 32044 33832 32084 33872
rect 31372 33664 31412 33704
rect 31372 33496 31412 33536
rect 31372 33328 31412 33368
rect 31180 33076 31220 33116
rect 31180 32908 31220 32948
rect 30796 28624 30836 28664
rect 30604 28540 30644 28580
rect 32140 33664 32180 33704
rect 31660 33076 31700 33116
rect 31660 32824 31700 32864
rect 31756 32320 31796 32360
rect 31468 32236 31508 32276
rect 32620 33664 32660 33704
rect 32044 32908 32084 32948
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 33772 33076 33812 33116
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 34924 33328 34964 33368
rect 34348 33076 34388 33116
rect 33676 32992 33716 33032
rect 33292 32908 33332 32948
rect 33196 32824 33236 32864
rect 32140 32656 32180 32696
rect 31756 31900 31796 31940
rect 32236 32320 32276 32360
rect 32236 31480 32276 31520
rect 32044 31396 32084 31436
rect 31084 29884 31124 29924
rect 31468 29884 31508 29924
rect 30988 29296 31028 29336
rect 31084 29128 31124 29168
rect 30220 27532 30260 27572
rect 30124 27028 30164 27068
rect 29260 26272 29300 26312
rect 29548 26272 29588 26312
rect 28204 25348 28244 25388
rect 28108 24844 28148 24884
rect 28204 23752 28244 23792
rect 28108 22744 28148 22784
rect 27436 20728 27476 20768
rect 27148 20476 27188 20516
rect 27820 20140 27860 20180
rect 29356 25936 29396 25976
rect 28972 25600 29012 25640
rect 29260 25348 29300 25388
rect 29644 26188 29684 26228
rect 29836 25852 29876 25892
rect 29836 25180 29876 25220
rect 29740 24340 29780 24380
rect 28876 23836 28916 23876
rect 28972 23332 29012 23372
rect 29164 22912 29204 22952
rect 29164 22744 29204 22784
rect 28588 22660 28628 22700
rect 30124 24340 30164 24380
rect 30508 27616 30548 27656
rect 30796 27616 30836 27656
rect 30508 27364 30548 27404
rect 30988 27028 31028 27068
rect 30892 26860 30932 26900
rect 30700 26776 30740 26816
rect 30604 26104 30644 26144
rect 30796 26440 30836 26480
rect 30604 25852 30644 25892
rect 30412 25516 30452 25556
rect 30316 24844 30356 24884
rect 30412 24760 30452 24800
rect 30412 23752 30452 23792
rect 30220 23332 30260 23372
rect 30412 23080 30452 23120
rect 30316 22912 30356 22952
rect 30316 22660 30356 22700
rect 30220 21568 30260 21608
rect 29836 21400 29876 21440
rect 28684 20728 28724 20768
rect 27532 19468 27572 19508
rect 25996 18712 26036 18752
rect 25708 18376 25748 18416
rect 25516 17956 25556 17996
rect 25132 17872 25172 17912
rect 24652 16696 24692 16736
rect 24268 15520 24308 15560
rect 23980 15016 24020 15056
rect 23596 14680 23636 14720
rect 23500 14008 23540 14048
rect 23788 14512 23828 14552
rect 24076 14680 24116 14720
rect 24172 14512 24212 14552
rect 23980 14428 24020 14468
rect 24844 16024 24884 16064
rect 25324 17200 25364 17240
rect 25612 17200 25652 17240
rect 25804 17956 25844 17996
rect 25612 16696 25652 16736
rect 25228 15520 25268 15560
rect 24940 15016 24980 15056
rect 24748 14764 24788 14804
rect 23692 13336 23732 13376
rect 22924 13084 22964 13124
rect 23596 11656 23636 11696
rect 24268 13084 24308 13124
rect 23500 11236 23540 11276
rect 23404 11152 23444 11192
rect 23020 10816 23060 10856
rect 23980 11656 24020 11696
rect 24172 11236 24212 11276
rect 23884 11152 23924 11192
rect 23692 10816 23732 10856
rect 22924 10228 22964 10268
rect 23404 10144 23444 10184
rect 23697 10228 23737 10268
rect 23308 9976 23348 10016
rect 23596 10144 23636 10184
rect 23308 9640 23348 9680
rect 22828 9136 22868 9176
rect 22732 9052 22772 9092
rect 22828 8884 22868 8924
rect 22444 8800 22484 8840
rect 23116 9220 23156 9260
rect 23020 9136 23060 9176
rect 22732 8632 22772 8672
rect 22348 8548 22388 8588
rect 22348 8380 22388 8420
rect 22540 8380 22580 8420
rect 22444 7960 22484 8000
rect 22919 8464 22959 8504
rect 23212 8800 23252 8840
rect 23404 8632 23444 8672
rect 23308 8548 23348 8588
rect 23020 8380 23060 8420
rect 24076 10984 24116 11024
rect 24652 14680 24692 14720
rect 24460 11488 24500 11528
rect 24364 10984 24404 11024
rect 25132 14848 25172 14888
rect 24940 14680 24980 14720
rect 25516 16024 25556 16064
rect 25708 16024 25748 16064
rect 26380 17956 26420 17996
rect 26572 17200 26612 17240
rect 26380 17032 26420 17072
rect 26572 16948 26612 16988
rect 26572 16696 26612 16736
rect 26092 15772 26132 15812
rect 25324 14512 25364 14552
rect 25804 14428 25844 14468
rect 25516 14092 25556 14132
rect 24652 13084 24692 13124
rect 24844 11908 24884 11948
rect 24748 11152 24788 11192
rect 24556 10984 24596 11024
rect 24556 10396 24596 10436
rect 24076 9976 24116 10016
rect 24364 10144 24404 10184
rect 24268 9976 24308 10016
rect 24172 9892 24212 9932
rect 24844 10984 24884 11024
rect 26188 14680 26228 14720
rect 26092 14512 26132 14552
rect 26092 14260 26132 14300
rect 25900 13924 25940 13964
rect 25612 12664 25652 12704
rect 25036 12076 25076 12116
rect 25036 11404 25076 11444
rect 24748 10396 24788 10436
rect 23692 9472 23732 9512
rect 23596 8800 23636 8840
rect 24172 9472 24212 9512
rect 24076 9388 24116 9428
rect 24172 9220 24212 9260
rect 23788 8884 23828 8924
rect 24364 8884 24404 8924
rect 23692 8632 23732 8672
rect 23884 8632 23924 8672
rect 24364 8716 24404 8756
rect 24076 8632 24116 8672
rect 23116 8296 23156 8336
rect 23596 8296 23636 8336
rect 23020 8212 23060 8252
rect 22156 7624 22196 7664
rect 22060 7540 22100 7580
rect 21676 7288 21716 7328
rect 21484 6364 21524 6404
rect 21388 5776 21428 5816
rect 22348 7204 22388 7244
rect 22252 7120 22292 7160
rect 22732 7792 22772 7832
rect 22732 7540 22772 7580
rect 22636 7456 22676 7496
rect 22540 6868 22580 6908
rect 23212 8128 23252 8168
rect 23308 8044 23348 8084
rect 23788 8296 23828 8336
rect 23500 8128 23540 8168
rect 23692 8044 23732 8084
rect 24268 8632 24308 8672
rect 23884 7960 23924 8000
rect 23020 7540 23060 7580
rect 22924 7372 22964 7412
rect 23596 7624 23636 7664
rect 23212 7288 23252 7328
rect 23404 7288 23444 7328
rect 23116 7204 23156 7244
rect 22828 6952 22868 6992
rect 23308 7204 23348 7244
rect 23596 7120 23636 7160
rect 23788 7120 23828 7160
rect 23980 7792 24020 7832
rect 24172 8128 24212 8168
rect 24364 8548 24404 8588
rect 24364 8212 24404 8252
rect 24268 7624 24308 7664
rect 24172 7288 24212 7328
rect 24081 6952 24121 6992
rect 23692 6868 23732 6908
rect 23212 6784 23252 6824
rect 23116 6616 23156 6656
rect 22828 6532 22868 6572
rect 22732 6448 22772 6488
rect 23116 6448 23156 6488
rect 22636 6364 22676 6404
rect 23500 6532 23540 6572
rect 23788 6616 23828 6656
rect 23212 6364 23252 6404
rect 23404 6364 23444 6404
rect 22828 6280 22868 6320
rect 22060 6196 22100 6236
rect 23020 6196 23060 6236
rect 22444 5692 22484 5732
rect 21580 5524 21620 5564
rect 22348 5524 22388 5564
rect 22732 5776 22772 5816
rect 20908 5188 20948 5228
rect 20332 4264 20372 4304
rect 20044 4180 20084 4220
rect 20332 4096 20372 4136
rect 20236 3928 20276 3968
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 19948 3676 19988 3716
rect 19372 3592 19412 3632
rect 19276 3424 19316 3464
rect 19756 3508 19796 3548
rect 19180 3340 19220 3380
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 17836 2752 17876 2792
rect 18028 2752 18068 2792
rect 18124 2500 18164 2540
rect 17932 2416 17972 2456
rect 18316 2836 18356 2876
rect 18316 2500 18356 2540
rect 19372 2920 19412 2960
rect 18412 2416 18452 2456
rect 19468 2668 19508 2708
rect 19660 2584 19700 2624
rect 19852 2584 19892 2624
rect 20140 3424 20180 3464
rect 20140 3256 20180 3296
rect 20524 4852 20564 4892
rect 20620 4516 20660 4556
rect 21484 5104 21524 5144
rect 21388 4936 21428 4976
rect 20908 4852 20948 4892
rect 20908 4432 20948 4472
rect 20908 4264 20948 4304
rect 20620 3760 20660 3800
rect 20524 3676 20564 3716
rect 18604 2500 18644 2540
rect 18796 1744 18836 1784
rect 17452 1660 17492 1700
rect 17260 1072 17300 1112
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 19372 2416 19412 2456
rect 20140 2584 20180 2624
rect 20428 3424 20468 3464
rect 20620 2668 20660 2708
rect 20428 2584 20468 2624
rect 20236 2416 20276 2456
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 19372 1744 19412 1784
rect 20812 4096 20852 4136
rect 21100 4516 21140 4556
rect 21196 4348 21236 4388
rect 21100 3592 21140 3632
rect 20908 3508 20948 3548
rect 20812 3256 20852 3296
rect 20812 3004 20852 3044
rect 21100 3424 21140 3464
rect 21004 3340 21044 3380
rect 20908 2920 20948 2960
rect 21671 4936 21676 4976
rect 21676 4936 21711 4976
rect 21772 4936 21812 4976
rect 21580 3760 21620 3800
rect 21388 3508 21428 3548
rect 21484 3340 21524 3380
rect 21292 3256 21332 3296
rect 21292 3088 21332 3128
rect 21196 2584 21236 2624
rect 21676 3424 21716 3464
rect 21580 1912 21620 1952
rect 21772 2080 21812 2120
rect 23884 6448 23924 6488
rect 24556 9472 24596 9512
rect 24652 9220 24692 9260
rect 24844 10144 24884 10184
rect 26092 13084 26132 13124
rect 26764 16276 26804 16316
rect 26860 16024 26900 16064
rect 26860 15688 26900 15728
rect 26764 15268 26804 15308
rect 27724 18544 27764 18584
rect 27724 18208 27764 18248
rect 27340 17200 27380 17240
rect 27532 17200 27572 17240
rect 27148 16276 27188 16316
rect 27724 17032 27764 17072
rect 28588 19132 28628 19172
rect 27916 18712 27956 18752
rect 29164 19216 29204 19256
rect 29260 19048 29300 19088
rect 28780 18964 28820 19004
rect 28492 18712 28532 18752
rect 28204 18628 28244 18668
rect 28108 18544 28148 18584
rect 28012 18208 28052 18248
rect 28012 17872 28052 17912
rect 28012 17704 28052 17744
rect 28396 18460 28436 18500
rect 28204 17536 28244 17576
rect 28204 17200 28244 17240
rect 28108 17116 28148 17156
rect 27916 17032 27956 17072
rect 27436 16780 27476 16820
rect 27628 16780 27668 16820
rect 27340 16276 27380 16316
rect 27244 16024 27284 16064
rect 28492 17872 28532 17912
rect 28780 18544 28820 18584
rect 31564 29296 31604 29336
rect 31756 30640 31796 30680
rect 32812 32152 32852 32192
rect 32620 31480 32660 31520
rect 32908 31480 32948 31520
rect 33484 32152 33524 32192
rect 34156 32908 34196 32948
rect 33868 32824 33908 32864
rect 36364 34336 36404 34376
rect 35884 33328 35924 33368
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 33196 31564 33236 31604
rect 33388 31564 33428 31604
rect 33004 30724 33044 30764
rect 31948 30388 31988 30428
rect 32332 30556 32372 30596
rect 32236 29968 32276 30008
rect 32044 29632 32084 29672
rect 31852 29464 31892 29504
rect 33196 30640 33236 30680
rect 32812 30556 32852 30596
rect 32524 30388 32564 30428
rect 32908 30388 32948 30428
rect 33004 29800 33044 29840
rect 32812 29716 32852 29756
rect 32428 29464 32468 29504
rect 32716 29464 32756 29504
rect 31660 29044 31700 29084
rect 32428 28624 32468 28664
rect 31564 28456 31604 28496
rect 32236 28456 32276 28496
rect 31276 28372 31316 28412
rect 32044 28288 32084 28328
rect 31660 28120 31700 28160
rect 31276 27700 31316 27740
rect 31468 27700 31508 27740
rect 31180 27616 31220 27656
rect 31660 27616 31700 27656
rect 32044 27616 32084 27656
rect 31372 27364 31412 27404
rect 31468 26776 31508 26816
rect 31276 26440 31316 26480
rect 31756 26440 31796 26480
rect 31180 26188 31220 26228
rect 31564 25852 31604 25892
rect 31180 25768 31220 25808
rect 34156 32152 34196 32192
rect 34540 32152 34580 32192
rect 35116 32824 35156 32864
rect 36652 34336 36692 34376
rect 36652 33664 36692 33704
rect 35980 32992 36020 33032
rect 36268 32992 36308 33032
rect 35212 32656 35252 32696
rect 35788 32320 35828 32360
rect 35020 32236 35060 32276
rect 35212 32152 35252 32192
rect 35692 32152 35732 32192
rect 36172 32320 36212 32360
rect 36844 32908 36884 32948
rect 36652 32488 36692 32528
rect 36556 32236 36596 32276
rect 34156 31480 34196 31520
rect 34060 30808 34100 30848
rect 33868 30640 33908 30680
rect 34732 31228 34772 31268
rect 36076 31984 36116 32024
rect 35596 31228 35636 31268
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 34540 30808 34580 30848
rect 35020 30808 35060 30848
rect 33772 30556 33812 30596
rect 33676 30472 33716 30512
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 33388 29968 33428 30008
rect 33964 29800 34004 29840
rect 33100 29716 33140 29756
rect 33100 29128 33140 29168
rect 33004 29044 33044 29084
rect 32812 28288 32852 28328
rect 32236 28204 32276 28244
rect 32620 28120 32660 28160
rect 32908 27784 32948 27824
rect 32236 27448 32276 27488
rect 32812 27448 32852 27488
rect 32140 27028 32180 27068
rect 32236 26608 32276 26648
rect 31852 25348 31892 25388
rect 32812 26104 32852 26144
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 33196 28204 33236 28244
rect 34156 30472 34196 30512
rect 34732 30556 34772 30596
rect 34636 30304 34676 30344
rect 36460 32068 36500 32108
rect 36172 31900 36212 31940
rect 36172 31564 36212 31604
rect 35788 30640 35828 30680
rect 35212 30472 35252 30512
rect 35692 29884 35732 29924
rect 35116 29632 35156 29672
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 34444 29296 34484 29336
rect 35116 29128 35156 29168
rect 34060 28372 34100 28412
rect 33772 28288 33812 28328
rect 33964 28204 34004 28244
rect 33868 27448 33908 27488
rect 33100 27364 33140 27404
rect 33292 27364 33332 27404
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 33868 27028 33908 27068
rect 33100 26608 33140 26648
rect 32716 25432 32756 25472
rect 32236 25264 32276 25304
rect 31084 25180 31124 25220
rect 31660 25180 31700 25220
rect 31276 24760 31316 24800
rect 32140 24592 32180 24632
rect 30988 24340 31028 24380
rect 32044 24340 32084 24380
rect 30796 24088 30836 24128
rect 31276 23920 31316 23960
rect 32140 23920 32180 23960
rect 31276 23752 31316 23792
rect 32044 23668 32084 23708
rect 31084 23500 31124 23540
rect 31948 23332 31988 23372
rect 31468 22912 31508 22952
rect 30700 22660 30740 22700
rect 30604 21484 30644 21524
rect 30508 20728 30548 20768
rect 30988 21568 31028 21608
rect 30796 21484 30836 21524
rect 31084 21484 31124 21524
rect 31852 22240 31892 22280
rect 31564 21736 31604 21776
rect 31756 21484 31796 21524
rect 31180 21400 31220 21440
rect 31372 21400 31412 21440
rect 31852 21400 31892 21440
rect 31660 20896 31700 20936
rect 31948 20896 31988 20936
rect 32620 24760 32660 24800
rect 32716 23836 32756 23876
rect 32332 23752 32372 23792
rect 32524 23668 32564 23708
rect 32524 23416 32564 23456
rect 32428 22492 32468 22532
rect 32428 22240 32468 22280
rect 33004 25852 33044 25892
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 33388 25432 33428 25472
rect 32908 24760 32948 24800
rect 32908 23920 32948 23960
rect 33004 23836 33044 23876
rect 32716 23416 32756 23456
rect 32524 21904 32564 21944
rect 32908 22324 32948 22364
rect 32716 22156 32756 22196
rect 32716 21904 32756 21944
rect 32332 21736 32372 21776
rect 32236 21568 32276 21608
rect 32140 21400 32180 21440
rect 32428 21568 32468 21608
rect 32332 21484 32372 21524
rect 32812 21652 32852 21692
rect 32908 21484 32948 21524
rect 33292 24592 33332 24632
rect 34252 27028 34292 27068
rect 34156 26860 34196 26900
rect 33964 26104 34004 26144
rect 34060 26020 34100 26060
rect 35980 31312 36020 31352
rect 36364 30976 36404 31016
rect 36076 30724 36116 30764
rect 36172 30472 36212 30512
rect 35692 29380 35732 29420
rect 36556 30976 36596 31016
rect 36556 30808 36596 30848
rect 36652 30724 36692 30764
rect 36748 30640 36788 30680
rect 36556 30472 36596 30512
rect 36364 29380 36404 29420
rect 35788 29212 35828 29252
rect 35692 29128 35732 29168
rect 36748 29884 36788 29924
rect 36748 29296 36788 29336
rect 35308 28960 35348 29000
rect 36940 32152 36980 32192
rect 37132 32488 37172 32528
rect 37228 32236 37268 32276
rect 37804 34336 37844 34376
rect 37996 34336 38036 34376
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 38764 33664 38804 33704
rect 38668 33412 38708 33452
rect 39628 33412 39668 33452
rect 38188 32656 38228 32696
rect 37036 31900 37076 31940
rect 37228 30808 37268 30848
rect 37036 30304 37076 30344
rect 37132 30136 37172 30176
rect 37036 29800 37076 29840
rect 37420 29884 37460 29924
rect 37324 29800 37364 29840
rect 37228 29716 37268 29756
rect 36940 29632 36980 29672
rect 37324 29296 37364 29336
rect 37420 29212 37460 29252
rect 37516 29128 37556 29168
rect 35692 28372 35732 28412
rect 35980 28372 36020 28412
rect 35404 28288 35444 28328
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 34540 27784 34580 27824
rect 34444 27616 34484 27656
rect 35404 27616 35444 27656
rect 34732 26860 34772 26900
rect 34636 26776 34676 26816
rect 34444 26608 34484 26648
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 34348 26188 34388 26228
rect 34348 25852 34388 25892
rect 34252 25264 34292 25304
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 33484 23836 33524 23876
rect 33196 23752 33236 23792
rect 33100 23248 33140 23288
rect 33676 23752 33716 23792
rect 34060 24172 34100 24212
rect 33676 23500 33716 23540
rect 33484 23248 33524 23288
rect 33868 23416 33908 23456
rect 35308 26776 35348 26816
rect 35980 27700 36020 27740
rect 35596 27028 35636 27068
rect 37036 28876 37076 28916
rect 36556 27448 36596 27488
rect 36844 27448 36884 27488
rect 35116 26440 35156 26480
rect 35500 26440 35540 26480
rect 35404 26188 35444 26228
rect 35212 26020 35252 26060
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 35884 25264 35924 25304
rect 35692 25180 35732 25220
rect 36940 26440 36980 26480
rect 36556 26272 36596 26312
rect 36268 26020 36308 26060
rect 36652 25768 36692 25808
rect 36460 25348 36500 25388
rect 35980 25180 36020 25220
rect 36556 24424 36596 24464
rect 34444 24172 34484 24212
rect 34252 24088 34292 24128
rect 33964 23332 34004 23372
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 34060 22492 34100 22532
rect 34348 23248 34388 23288
rect 34540 23668 34580 23708
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 34540 23248 34580 23288
rect 34156 22408 34196 22448
rect 33196 22324 33236 22364
rect 34060 22240 34100 22280
rect 33772 22156 33812 22196
rect 33100 21652 33140 21692
rect 33100 21484 33140 21524
rect 34156 21568 34196 21608
rect 34444 22324 34484 22364
rect 34924 23164 34964 23204
rect 34732 22912 34772 22952
rect 34828 22492 34868 22532
rect 35404 23248 35444 23288
rect 36364 23668 36404 23708
rect 38188 31984 38228 32024
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 39916 32656 39956 32696
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 39724 32068 39764 32108
rect 38764 31816 38804 31856
rect 39244 31816 39284 31856
rect 38572 31312 38612 31352
rect 38380 30808 38420 30848
rect 38284 30724 38324 30764
rect 39340 31144 39380 31184
rect 38956 30808 38996 30848
rect 39148 30640 39188 30680
rect 38572 30556 38612 30596
rect 38092 30388 38132 30428
rect 39436 30892 39476 30932
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 40588 31144 40628 31184
rect 40780 31144 40820 31184
rect 39628 30556 39668 30596
rect 39820 30388 39860 30428
rect 38956 30304 38996 30344
rect 37900 29128 37940 29168
rect 37708 28288 37748 28328
rect 37324 26524 37364 26564
rect 38092 28960 38132 29000
rect 38380 27700 38420 27740
rect 38764 27532 38804 27572
rect 38188 26776 38228 26816
rect 37996 26608 38036 26648
rect 37420 26272 37460 26312
rect 37228 26020 37268 26060
rect 37804 26188 37844 26228
rect 38860 27448 38900 27488
rect 38476 26692 38516 26732
rect 38380 26440 38420 26480
rect 38284 26188 38324 26228
rect 38476 26188 38516 26228
rect 37900 26020 37940 26060
rect 37228 25852 37268 25892
rect 37132 25516 37172 25556
rect 37612 25348 37652 25388
rect 37036 25180 37076 25220
rect 37708 25096 37748 25136
rect 38188 26104 38228 26144
rect 38188 25852 38228 25892
rect 38092 25768 38132 25808
rect 38092 25264 38132 25304
rect 38476 25768 38516 25808
rect 35692 23164 35732 23204
rect 35212 23080 35252 23120
rect 35020 22408 35060 22448
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 35500 23080 35540 23120
rect 35308 22912 35348 22952
rect 37324 23332 37364 23372
rect 37228 22912 37268 22952
rect 35596 21568 35636 21608
rect 34348 21484 34388 21524
rect 33196 21400 33236 21440
rect 35596 21400 35636 21440
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 29548 19552 29588 19592
rect 30316 19552 30356 19592
rect 29740 19048 29780 19088
rect 29548 18628 29588 18668
rect 28684 18460 28724 18500
rect 28684 18292 28724 18332
rect 28588 17368 28628 17408
rect 28396 17284 28436 17324
rect 29836 18712 29876 18752
rect 30508 19216 30548 19256
rect 29836 18544 29876 18584
rect 30028 18376 30068 18416
rect 28876 17872 28916 17912
rect 28780 17536 28820 17576
rect 28972 17704 29012 17744
rect 29740 17872 29780 17912
rect 28684 17200 28724 17240
rect 28396 17032 28436 17072
rect 28108 16780 28148 16820
rect 27724 16444 27764 16484
rect 28396 16360 28436 16400
rect 27916 16276 27956 16316
rect 27436 16024 27476 16064
rect 27052 15604 27092 15644
rect 27052 14932 27092 14972
rect 26956 14848 26996 14888
rect 26860 14764 26900 14804
rect 26956 14680 26996 14720
rect 26476 13840 26516 13880
rect 26956 14092 26996 14132
rect 27340 15604 27380 15644
rect 28012 16192 28052 16232
rect 27916 16024 27956 16064
rect 27820 15436 27860 15476
rect 27436 15268 27476 15308
rect 27244 15100 27284 15140
rect 27340 14848 27380 14888
rect 27820 14680 27860 14720
rect 27532 14512 27572 14552
rect 27436 14092 27476 14132
rect 27724 14596 27764 14636
rect 27436 13924 27476 13964
rect 27244 13756 27284 13796
rect 26860 12496 26900 12536
rect 26284 12328 26324 12368
rect 26188 12244 26228 12284
rect 26188 11572 26228 11612
rect 25612 10312 25652 10352
rect 27148 12580 27188 12620
rect 26956 11992 26996 12032
rect 27148 11824 27188 11864
rect 26860 11740 26900 11780
rect 26668 11656 26708 11696
rect 26572 11572 26612 11612
rect 26956 10984 26996 11024
rect 27340 12496 27380 12536
rect 27628 14008 27668 14048
rect 27820 13924 27860 13964
rect 28012 14848 28052 14888
rect 27532 13756 27572 13796
rect 27916 13756 27956 13796
rect 27820 13168 27860 13208
rect 28684 17032 28724 17072
rect 28972 17368 29012 17408
rect 28876 17200 28916 17240
rect 29452 17704 29492 17744
rect 30028 17872 30068 17912
rect 29356 17536 29396 17576
rect 29164 17200 29204 17240
rect 29260 17032 29300 17072
rect 29548 17536 29588 17576
rect 29164 16528 29204 16568
rect 29260 16276 29300 16316
rect 29452 16528 29492 16568
rect 30028 17032 30068 17072
rect 29644 16948 29684 16988
rect 29836 16528 29876 16568
rect 29836 16108 29876 16148
rect 28492 15688 28532 15728
rect 28396 15604 28436 15644
rect 28396 15352 28436 15392
rect 28684 15604 28724 15644
rect 28684 15352 28724 15392
rect 29260 15688 29300 15728
rect 29068 15604 29108 15644
rect 29164 15352 29204 15392
rect 28972 15268 29012 15308
rect 29548 15604 29588 15644
rect 28876 15100 28916 15140
rect 29452 15100 29492 15140
rect 28780 14932 28820 14972
rect 28588 14848 28628 14888
rect 28780 14764 28820 14804
rect 28684 14680 28724 14720
rect 28204 14596 28244 14636
rect 28108 14512 28148 14552
rect 28108 13924 28148 13964
rect 28108 13756 28148 13796
rect 27628 12664 27668 12704
rect 28300 14008 28340 14048
rect 29163 14764 29203 14804
rect 28972 14512 29012 14552
rect 29260 14680 29300 14720
rect 29356 14512 29396 14552
rect 28876 14344 28916 14384
rect 27820 12748 27860 12788
rect 27724 12580 27764 12620
rect 27724 12412 27764 12452
rect 27340 11656 27380 11696
rect 27628 11572 27668 11612
rect 27532 11488 27572 11528
rect 27244 10900 27284 10940
rect 25708 10228 25748 10268
rect 26956 10228 26996 10268
rect 25324 10060 25364 10100
rect 25132 9808 25172 9848
rect 25132 9640 25172 9680
rect 24844 9388 24884 9428
rect 25612 10144 25652 10184
rect 25516 9640 25556 9680
rect 25516 9472 25556 9512
rect 25324 9388 25364 9428
rect 25036 9220 25076 9260
rect 24748 8800 24788 8840
rect 24652 8716 24692 8756
rect 24940 8716 24980 8756
rect 24652 8464 24692 8504
rect 24844 8296 24884 8336
rect 24652 8212 24692 8252
rect 24556 8128 24596 8168
rect 24748 7960 24788 8000
rect 24556 7876 24596 7916
rect 24460 7708 24500 7748
rect 24652 7624 24692 7664
rect 24556 7540 24596 7580
rect 24460 7456 24500 7496
rect 24460 7288 24500 7328
rect 24556 7204 24596 7244
rect 24748 7120 24788 7160
rect 25324 9220 25364 9260
rect 25132 8464 25172 8504
rect 24460 6952 24500 6992
rect 24268 6448 24308 6488
rect 23692 6280 23732 6320
rect 23980 6364 24020 6404
rect 24172 6280 24212 6320
rect 23116 5440 23156 5480
rect 23020 5272 23060 5312
rect 23116 4852 23156 4892
rect 23980 5776 24020 5816
rect 23596 5608 23636 5648
rect 24076 5608 24116 5648
rect 24268 6196 24308 6236
rect 25228 8296 25268 8336
rect 25228 7876 25268 7916
rect 25132 7624 25172 7664
rect 25132 7372 25172 7412
rect 28492 13168 28532 13208
rect 28684 13168 28724 13208
rect 28396 12832 28436 12872
rect 29356 13336 29396 13376
rect 29068 13252 29108 13292
rect 28108 12412 28148 12452
rect 28492 12664 28532 12704
rect 28492 12496 28532 12536
rect 28396 12412 28436 12452
rect 28012 11656 28052 11696
rect 28108 10984 28148 11024
rect 27724 10648 27764 10688
rect 27052 10144 27092 10184
rect 27340 10144 27380 10184
rect 28012 10144 28052 10184
rect 26860 10060 26900 10100
rect 26668 9052 26708 9092
rect 25420 8212 25460 8252
rect 25420 7960 25460 8000
rect 25324 7624 25364 7664
rect 25804 8464 25844 8504
rect 26284 8296 26324 8336
rect 25996 8212 26036 8252
rect 25516 7456 25556 7496
rect 26572 8548 26612 8588
rect 26476 8464 26516 8504
rect 26092 7960 26132 8000
rect 26380 7960 26420 8000
rect 26668 8296 26708 8336
rect 26572 8044 26612 8084
rect 26381 7624 26421 7664
rect 26284 7540 26324 7580
rect 25036 7120 25076 7160
rect 25324 7120 25364 7160
rect 26380 7120 26420 7160
rect 24940 6616 24980 6656
rect 24748 6364 24788 6404
rect 24556 6280 24596 6320
rect 24364 5608 24404 5648
rect 24844 5692 24884 5732
rect 23788 5524 23828 5564
rect 26572 7036 26612 7076
rect 26764 7624 26804 7664
rect 26380 5860 26420 5900
rect 26572 6364 26612 6404
rect 23308 5356 23348 5396
rect 23596 5356 23636 5396
rect 23299 5020 23339 5060
rect 23404 5020 23444 5060
rect 23212 4768 23252 4808
rect 22060 4012 22100 4052
rect 22924 4348 22964 4388
rect 22732 4180 22772 4220
rect 22732 3424 22772 3464
rect 23692 5272 23732 5312
rect 23884 5020 23924 5060
rect 24268 4852 24308 4892
rect 23788 4684 23828 4724
rect 23500 4600 23540 4640
rect 23596 4516 23636 4556
rect 24460 5020 24500 5060
rect 24652 5020 24692 5060
rect 24844 5020 24884 5060
rect 26380 5440 26420 5480
rect 26956 9388 26996 9428
rect 27436 9472 27476 9512
rect 27239 8800 27279 8840
rect 27436 8632 27476 8672
rect 27916 9388 27956 9428
rect 27724 8800 27764 8840
rect 28300 11740 28340 11780
rect 28588 12412 28628 12452
rect 28396 11488 28436 11528
rect 28396 10060 28436 10100
rect 28300 9388 28340 9428
rect 28204 9304 28244 9344
rect 28588 9472 28628 9512
rect 28012 8800 28052 8840
rect 27724 8632 27764 8672
rect 27628 8464 27668 8504
rect 27340 8296 27380 8336
rect 27532 8128 27572 8168
rect 27052 7960 27092 8000
rect 27244 7960 27284 8000
rect 27148 7372 27188 7412
rect 27436 7960 27476 8000
rect 28588 8716 28628 8756
rect 28012 8632 28052 8672
rect 28588 8548 28628 8588
rect 28396 8464 28436 8504
rect 27916 8296 27956 8336
rect 27820 7960 27860 8000
rect 27820 7708 27860 7748
rect 27820 7540 27860 7580
rect 27148 7120 27188 7160
rect 27436 7120 27476 7160
rect 27628 7372 27668 7412
rect 27244 6952 27284 6992
rect 27820 6868 27860 6908
rect 27628 6532 27668 6572
rect 27532 6448 27572 6488
rect 28108 8128 28148 8168
rect 28204 7204 28244 7244
rect 28396 6700 28436 6740
rect 28204 6448 28244 6488
rect 28780 12664 28820 12704
rect 28972 12580 29012 12620
rect 28876 12496 28916 12536
rect 29164 13000 29204 13040
rect 30316 18292 30356 18332
rect 31564 18292 31604 18332
rect 30508 17956 30548 17996
rect 31180 17956 31220 17996
rect 30700 17872 30740 17912
rect 30220 16780 30260 16820
rect 30220 16276 30260 16316
rect 30988 17704 31028 17744
rect 31852 18040 31892 18080
rect 32908 19468 32948 19508
rect 32140 19216 32180 19256
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 32812 18964 32852 19004
rect 32332 18712 32372 18752
rect 32428 18544 32468 18584
rect 30988 17032 31028 17072
rect 30700 16864 30740 16904
rect 31084 16612 31124 16652
rect 31372 16948 31412 16988
rect 30508 16360 30548 16400
rect 31180 16360 31220 16400
rect 30892 16276 30932 16316
rect 30316 15856 30356 15896
rect 30220 15772 30260 15812
rect 29740 15352 29780 15392
rect 29740 15184 29780 15224
rect 29644 14680 29684 14720
rect 29932 15352 29972 15392
rect 29836 15016 29876 15056
rect 29932 14848 29972 14888
rect 29836 14764 29876 14804
rect 29932 14176 29972 14216
rect 29740 14092 29780 14132
rect 29836 13924 29876 13964
rect 29548 13000 29588 13040
rect 29452 12916 29492 12956
rect 29068 12496 29108 12536
rect 29068 12328 29108 12368
rect 28780 12160 28820 12200
rect 29356 12412 29396 12452
rect 29260 12328 29300 12368
rect 28876 11824 28916 11864
rect 28972 10984 29012 11024
rect 29164 11488 29204 11528
rect 29164 11236 29204 11276
rect 29068 10816 29108 10856
rect 29452 11488 29492 11528
rect 29740 13000 29780 13040
rect 29836 12328 29876 12368
rect 29740 11404 29780 11444
rect 30124 15688 30164 15728
rect 30316 15520 30356 15560
rect 30220 15352 30260 15392
rect 30508 16192 30548 16232
rect 30796 15604 30836 15644
rect 30700 15520 30740 15560
rect 30700 15352 30740 15392
rect 30412 15100 30452 15140
rect 30316 15016 30356 15056
rect 30028 13840 30068 13880
rect 31564 16360 31604 16400
rect 31372 16276 31412 16316
rect 31084 16192 31124 16232
rect 30988 16108 31028 16148
rect 31276 16108 31316 16148
rect 31564 16024 31604 16064
rect 31468 15856 31508 15896
rect 30892 15184 30932 15224
rect 30796 15016 30836 15056
rect 30508 14596 30548 14636
rect 30412 14008 30452 14048
rect 30892 14932 30932 14972
rect 30892 14680 30932 14720
rect 30796 14428 30836 14468
rect 30700 14008 30740 14048
rect 30508 13840 30548 13880
rect 30220 13672 30260 13712
rect 30124 13420 30164 13460
rect 30305 13168 30345 13208
rect 30604 13168 30644 13208
rect 30028 12916 30068 12956
rect 30796 13588 30836 13628
rect 30796 13252 30836 13292
rect 31372 15688 31412 15728
rect 31276 14932 31316 14972
rect 31756 16192 31796 16232
rect 31660 15688 31700 15728
rect 31084 14848 31124 14888
rect 31756 14932 31796 14972
rect 31084 13756 31124 13796
rect 30220 12916 30260 12956
rect 30796 12916 30836 12956
rect 30700 12580 30740 12620
rect 30796 12496 30836 12536
rect 30508 12076 30548 12116
rect 30700 12076 30740 12116
rect 29260 10312 29300 10352
rect 30124 10984 30164 11024
rect 29452 10228 29492 10268
rect 29644 10144 29684 10184
rect 29260 9892 29300 9932
rect 29068 9388 29108 9428
rect 28876 8548 28916 8588
rect 28972 8464 29012 8504
rect 29740 10060 29780 10100
rect 30412 11656 30452 11696
rect 30796 11992 30836 12032
rect 30796 11404 30836 11444
rect 31084 12748 31124 12788
rect 31468 14512 31508 14552
rect 31756 14344 31796 14384
rect 31756 14008 31796 14048
rect 32908 18712 32948 18752
rect 32812 17788 32852 17828
rect 32524 17704 32564 17744
rect 32428 17620 32468 17660
rect 32236 16948 32276 16988
rect 32140 16780 32180 16820
rect 32140 16276 32180 16316
rect 32044 16108 32084 16148
rect 32140 16024 32180 16064
rect 32524 17032 32564 17072
rect 32620 16780 32660 16820
rect 32428 16612 32468 16652
rect 32332 16444 32372 16484
rect 33100 18544 33140 18584
rect 33772 18544 33812 18584
rect 33676 18292 33716 18332
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 33100 17788 33140 17828
rect 32620 16360 32660 16400
rect 33004 16360 33044 16400
rect 32428 16108 32468 16148
rect 32620 16024 32660 16064
rect 32812 15940 32852 15980
rect 32140 15016 32180 15056
rect 32524 15520 32564 15560
rect 32620 15352 32660 15392
rect 33292 17704 33332 17744
rect 33196 17620 33236 17660
rect 33388 17620 33428 17660
rect 32812 15184 32852 15224
rect 32812 14848 32852 14888
rect 31948 14512 31988 14552
rect 31948 14260 31988 14300
rect 32140 14680 32180 14720
rect 32716 14512 32756 14552
rect 32908 14548 32948 14552
rect 32908 14512 32948 14548
rect 32140 14428 32180 14468
rect 36172 22240 36212 22280
rect 36844 22240 36884 22280
rect 36460 21484 36500 21524
rect 36748 21400 36788 21440
rect 37324 21736 37364 21776
rect 36556 19972 36596 20012
rect 36652 19888 36692 19928
rect 35308 19720 35348 19760
rect 35692 19720 35732 19760
rect 34252 19132 34292 19172
rect 34924 19132 34964 19172
rect 34156 18292 34196 18332
rect 34060 17620 34100 17660
rect 33292 16864 33332 16904
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 35116 19132 35156 19172
rect 34444 17704 34484 17744
rect 34252 16192 34292 16232
rect 33580 16024 33620 16064
rect 33676 15604 33716 15644
rect 34156 15604 34196 15644
rect 33388 15520 33428 15560
rect 33964 15520 34004 15560
rect 33388 15268 33428 15308
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 33868 15100 33908 15140
rect 33868 14932 33908 14972
rect 33100 14848 33140 14888
rect 33196 14764 33236 14804
rect 32908 14344 32948 14384
rect 33009 14344 33049 14384
rect 32236 14092 32276 14132
rect 32044 13924 32084 13964
rect 32524 14008 32564 14048
rect 32716 14008 32756 14048
rect 31660 13504 31700 13544
rect 31756 13168 31796 13208
rect 31564 12664 31604 12704
rect 31372 12496 31412 12536
rect 31276 12412 31316 12452
rect 31660 12496 31700 12536
rect 32332 13840 32372 13880
rect 32236 13756 32276 13796
rect 32524 13672 32564 13712
rect 32044 13252 32084 13292
rect 32236 13168 32276 13208
rect 32332 13084 32372 13124
rect 32428 12916 32468 12956
rect 32140 12748 32180 12788
rect 32428 12664 32468 12704
rect 31852 12160 31892 12200
rect 31564 12076 31604 12116
rect 32044 12076 32084 12116
rect 31564 11908 31604 11948
rect 30988 11740 31028 11780
rect 31372 11740 31412 11780
rect 31084 11656 31124 11696
rect 31084 11404 31124 11444
rect 31660 11824 31700 11864
rect 31852 11824 31892 11864
rect 31468 11572 31508 11612
rect 31564 11404 31604 11444
rect 31564 10984 31604 11024
rect 31756 11152 31796 11192
rect 31372 10312 31412 10352
rect 31756 10312 31796 10352
rect 31660 10228 31700 10268
rect 29836 9640 29876 9680
rect 30220 9556 30260 9596
rect 29644 9388 29684 9428
rect 29356 9304 29396 9344
rect 29932 9304 29972 9344
rect 30412 8968 30452 9008
rect 30316 8884 30356 8924
rect 30700 9556 30740 9596
rect 30892 9388 30932 9428
rect 29164 8716 29204 8756
rect 29164 8464 29204 8504
rect 28876 8128 28916 8168
rect 29068 7540 29108 7580
rect 28780 7204 28820 7244
rect 27436 6280 27476 6320
rect 26284 5356 26324 5396
rect 25036 4684 25076 4724
rect 24940 4516 24980 4556
rect 23596 4264 23636 4304
rect 24076 4264 24116 4304
rect 24844 4264 24884 4304
rect 23308 3760 23348 3800
rect 23500 3676 23540 3716
rect 23980 4096 24020 4136
rect 23788 3928 23828 3968
rect 23788 3592 23828 3632
rect 24172 3676 24212 3716
rect 25420 4600 25460 4640
rect 25420 4348 25460 4388
rect 25324 4264 25364 4304
rect 24364 4012 24404 4052
rect 24268 3592 24308 3632
rect 24076 3508 24116 3548
rect 23692 3424 23732 3464
rect 24268 3424 24308 3464
rect 25612 4096 25652 4136
rect 26092 4768 26132 4808
rect 25900 4180 25940 4220
rect 26284 4768 26324 4808
rect 26476 4936 26516 4976
rect 26380 4180 26420 4220
rect 26092 4096 26132 4136
rect 26188 4012 26228 4052
rect 26476 4012 26516 4052
rect 25516 3592 25556 3632
rect 25420 3508 25460 3548
rect 24460 3340 24500 3380
rect 25324 3340 25364 3380
rect 24172 3256 24212 3296
rect 24364 3256 24404 3296
rect 22636 2752 22676 2792
rect 25132 2920 25172 2960
rect 22444 2080 22484 2120
rect 22540 1996 22580 2036
rect 22444 1912 22484 1952
rect 25420 2752 25460 2792
rect 23020 2416 23060 2456
rect 24076 2416 24116 2456
rect 22924 1996 22964 2036
rect 26380 3928 26420 3968
rect 26860 5608 26900 5648
rect 26668 4852 26708 4892
rect 26668 4096 26708 4136
rect 26860 4936 26900 4976
rect 27244 4936 27284 4976
rect 27148 4768 27188 4808
rect 27340 4768 27380 4808
rect 26764 3760 26804 3800
rect 26572 3508 26612 3548
rect 26764 3424 26804 3464
rect 26572 3172 26612 3212
rect 27244 3508 27284 3548
rect 27148 3088 27188 3128
rect 27244 3004 27284 3044
rect 27628 4432 27668 4472
rect 27628 4096 27668 4136
rect 27532 3928 27572 3968
rect 27436 3844 27476 3884
rect 27628 3844 27668 3884
rect 27532 3760 27572 3800
rect 27436 3508 27476 3548
rect 27436 3172 27476 3212
rect 27628 2836 27668 2876
rect 25324 1240 25364 1280
rect 26860 1912 26900 1952
rect 26284 1240 26324 1280
rect 26668 1240 26708 1280
rect 19564 1072 19604 1112
rect 20716 1072 20756 1112
rect 27916 5608 27956 5648
rect 27820 5440 27860 5480
rect 28588 6448 28628 6488
rect 29548 8632 29588 8672
rect 30700 8800 30740 8840
rect 29740 8548 29780 8588
rect 30065 8548 30105 8588
rect 29836 8128 29876 8168
rect 29452 7960 29492 8000
rect 29836 7960 29876 8000
rect 29356 7372 29396 7412
rect 29260 7204 29300 7244
rect 30028 7960 30068 8000
rect 30124 7624 30164 7664
rect 30316 8632 30356 8672
rect 31084 9220 31124 9260
rect 30604 8716 30644 8756
rect 30988 8716 31028 8756
rect 30508 8464 30548 8504
rect 30988 8128 31028 8168
rect 30604 7960 30644 8000
rect 30412 7876 30452 7916
rect 30028 7540 30068 7580
rect 29740 7204 29780 7244
rect 29548 7120 29588 7160
rect 29452 6784 29492 6824
rect 29356 6700 29396 6740
rect 28972 6448 29012 6488
rect 29164 6448 29204 6488
rect 29836 6868 29876 6908
rect 29548 6364 29588 6404
rect 30220 7540 30260 7580
rect 30124 7456 30164 7496
rect 30028 7288 30068 7328
rect 30508 7456 30548 7496
rect 30412 7288 30452 7328
rect 30412 7120 30452 7160
rect 30316 6868 30356 6908
rect 30220 6784 30260 6824
rect 30124 6700 30164 6740
rect 29740 6364 29780 6404
rect 29644 6280 29684 6320
rect 28108 5104 28148 5144
rect 27916 4600 27956 4640
rect 28300 5020 28340 5060
rect 28492 5608 28532 5648
rect 28396 4852 28436 4892
rect 28204 4684 28244 4724
rect 28108 4432 28148 4472
rect 28972 5608 29012 5648
rect 28780 5440 28820 5480
rect 28972 5440 29012 5480
rect 28780 5188 28820 5228
rect 28876 4936 28916 4976
rect 29260 5440 29300 5480
rect 29164 5104 29204 5144
rect 29740 5440 29780 5480
rect 29548 5272 29588 5312
rect 29260 4936 29300 4976
rect 29452 4936 29492 4976
rect 29356 4852 29396 4892
rect 29068 4768 29108 4808
rect 28972 4684 29012 4724
rect 28780 4600 28820 4640
rect 28684 4348 28724 4388
rect 28108 4096 28148 4136
rect 28012 4012 28052 4052
rect 27916 3760 27956 3800
rect 27820 3424 27860 3464
rect 28108 3424 28148 3464
rect 28396 4096 28436 4136
rect 28588 4096 28628 4136
rect 28588 3844 28628 3884
rect 28492 3676 28532 3716
rect 27820 3172 27860 3212
rect 27916 3088 27956 3128
rect 28012 3004 28052 3044
rect 28396 3424 28436 3464
rect 28300 2836 28340 2876
rect 28108 2584 28148 2624
rect 29068 4096 29108 4136
rect 29068 3844 29108 3884
rect 29164 3760 29204 3800
rect 28972 3592 29012 3632
rect 29452 4600 29492 4640
rect 29836 5188 29876 5228
rect 29835 5020 29875 5060
rect 30028 5020 30068 5060
rect 29740 4936 29780 4976
rect 29932 4936 29972 4976
rect 29644 4852 29684 4892
rect 29356 3844 29396 3884
rect 29260 3676 29300 3716
rect 28684 3508 28724 3548
rect 29356 3424 29396 3464
rect 29548 4180 29588 4220
rect 29740 3928 29780 3968
rect 29644 3844 29684 3884
rect 29836 3424 29876 3464
rect 29260 3340 29300 3380
rect 29932 3340 29972 3380
rect 28972 2584 29012 2624
rect 29740 2752 29780 2792
rect 29356 2584 29396 2624
rect 30220 5608 30260 5648
rect 30700 7288 30740 7328
rect 30796 6868 30836 6908
rect 30796 6700 30836 6740
rect 30892 6616 30932 6656
rect 30892 6448 30932 6488
rect 30604 5944 30644 5984
rect 30508 5440 30548 5480
rect 30412 5104 30452 5144
rect 30508 5020 30548 5060
rect 31084 7456 31124 7496
rect 31564 10144 31604 10184
rect 31564 9976 31604 10016
rect 31756 9724 31796 9764
rect 31276 9556 31316 9596
rect 31276 9304 31316 9344
rect 31372 9220 31412 9260
rect 31372 8800 31412 8840
rect 31660 9388 31700 9428
rect 31564 9052 31604 9092
rect 31564 8884 31604 8924
rect 31468 8632 31508 8672
rect 31660 7960 31700 8000
rect 31180 7372 31220 7412
rect 31276 6700 31316 6740
rect 31372 6532 31412 6572
rect 31660 7540 31700 7580
rect 32140 11656 32180 11696
rect 32524 12244 32564 12284
rect 32332 11824 32372 11864
rect 31948 11572 31988 11612
rect 32236 11572 32276 11612
rect 33004 14008 33044 14048
rect 33292 14512 33332 14552
rect 33676 14596 33716 14636
rect 33484 14512 33524 14552
rect 33676 14260 33716 14300
rect 33388 14176 33428 14216
rect 33580 14092 33620 14132
rect 33004 13756 33044 13796
rect 32908 13588 32948 13628
rect 32812 13168 32852 13208
rect 33388 14008 33428 14048
rect 33484 13924 33524 13964
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 34540 17032 34580 17072
rect 35596 18964 35636 19004
rect 35788 18544 35828 18584
rect 35308 17788 35348 17828
rect 35692 16948 35732 16988
rect 35596 16360 35636 16400
rect 35212 16276 35252 16316
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 34252 15520 34292 15560
rect 34060 15436 34100 15476
rect 34252 15268 34292 15308
rect 34156 15100 34196 15140
rect 34060 14764 34100 14804
rect 34444 15520 34484 15560
rect 34828 15100 34868 15140
rect 34636 14848 34676 14888
rect 34732 14680 34772 14720
rect 34060 14428 34100 14468
rect 33868 14344 33908 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 34156 14260 34196 14300
rect 34060 14092 34100 14132
rect 33772 13924 33812 13964
rect 33196 13672 33236 13712
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 33100 13252 33140 13292
rect 33580 13168 33620 13208
rect 35116 14344 35156 14384
rect 34252 14092 34292 14132
rect 33868 13168 33908 13208
rect 33868 13000 33908 13040
rect 34444 13504 34484 13544
rect 34444 13336 34484 13376
rect 34348 13168 34388 13208
rect 33196 12496 33236 12536
rect 34348 13000 34388 13040
rect 34252 12580 34292 12620
rect 32620 11908 32660 11948
rect 33004 11824 33044 11864
rect 32428 11488 32468 11528
rect 32524 11404 32564 11444
rect 32908 11656 32948 11696
rect 32716 11572 32756 11612
rect 32812 11488 32852 11528
rect 32332 11236 32372 11276
rect 32428 11152 32468 11192
rect 32044 10900 32084 10940
rect 32524 10984 32564 11024
rect 32716 11152 32756 11192
rect 32716 10984 32756 11024
rect 34924 13756 34964 13796
rect 34828 13168 34868 13208
rect 35404 14008 35444 14048
rect 35212 13840 35252 13880
rect 36556 17032 36596 17072
rect 36460 16948 36500 16988
rect 35980 15184 36020 15224
rect 35884 14008 35924 14048
rect 36172 14008 36212 14048
rect 34924 13084 34964 13124
rect 35020 13000 35060 13040
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 34444 12580 34484 12620
rect 35020 12580 35060 12620
rect 35212 13168 35252 13208
rect 35500 13084 35540 13124
rect 35692 13168 35732 13208
rect 36172 13252 36212 13292
rect 35788 13000 35828 13040
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 33292 11740 33332 11780
rect 33196 11236 33236 11276
rect 32236 10564 32276 10604
rect 32140 10480 32180 10520
rect 31948 10312 31988 10352
rect 32524 10312 32564 10352
rect 32428 10144 32468 10184
rect 32908 10648 32948 10688
rect 32812 10480 32852 10520
rect 32812 10228 32852 10268
rect 32140 10060 32180 10100
rect 31948 9892 31988 9932
rect 32051 9472 32091 9512
rect 32044 9304 32084 9344
rect 31948 8800 31988 8840
rect 33196 10984 33236 11024
rect 33388 11572 33428 11612
rect 33676 11488 33716 11528
rect 34156 12160 34196 12200
rect 34252 11824 34292 11864
rect 33868 11488 33908 11528
rect 33868 11236 33908 11276
rect 33772 10816 33812 10856
rect 33100 10564 33140 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 33004 10396 33044 10436
rect 32908 10144 32948 10184
rect 33484 10396 33524 10436
rect 33100 10312 33140 10352
rect 33292 10060 33332 10100
rect 32620 9976 32660 10016
rect 32236 9808 32276 9848
rect 32236 8968 32276 9008
rect 32140 8884 32180 8924
rect 31852 8212 31892 8252
rect 32140 7876 32180 7916
rect 31756 7372 31796 7412
rect 31660 7288 31700 7328
rect 31468 6448 31508 6488
rect 32140 7288 32180 7328
rect 32044 7120 32084 7160
rect 31756 6532 31796 6572
rect 31948 6532 31988 6572
rect 31564 6280 31604 6320
rect 32524 7540 32564 7580
rect 32524 7372 32564 7412
rect 32332 7288 32372 7328
rect 32236 7120 32276 7160
rect 34156 10900 34196 10940
rect 35212 12412 35252 12452
rect 34924 12244 34964 12284
rect 35596 12580 35636 12620
rect 34924 11656 34964 11696
rect 34636 11488 34676 11528
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 35500 11656 35540 11696
rect 35212 11152 35252 11192
rect 34348 10816 34388 10856
rect 34156 10228 34196 10268
rect 34540 10144 34580 10184
rect 35308 11068 35348 11108
rect 34924 10984 34964 11024
rect 35020 10900 35060 10940
rect 36076 13000 36116 13040
rect 35980 11488 36020 11528
rect 35692 11152 35732 11192
rect 35884 11152 35924 11192
rect 36652 16948 36692 16988
rect 36652 16780 36692 16820
rect 36652 16360 36692 16400
rect 36652 15772 36692 15812
rect 38188 23752 38228 23792
rect 38572 24592 38612 24632
rect 38764 26104 38804 26144
rect 41740 30220 41780 30260
rect 42700 30220 42740 30260
rect 40300 29800 40340 29840
rect 40012 29716 40052 29756
rect 39436 28960 39476 29000
rect 40396 29632 40436 29672
rect 40684 29800 40724 29840
rect 41356 29800 41396 29840
rect 40876 29632 40916 29672
rect 41260 29632 41300 29672
rect 40684 29212 40724 29252
rect 39244 28204 39284 28244
rect 39340 27532 39380 27572
rect 39628 27112 39668 27152
rect 39436 27028 39476 27068
rect 39052 26440 39092 26480
rect 39436 26440 39476 26480
rect 39148 26188 39188 26228
rect 39628 26188 39668 26228
rect 38956 26020 38996 26060
rect 38956 25264 38996 25304
rect 39340 26104 39380 26144
rect 39340 25264 39380 25304
rect 38860 24676 38900 24716
rect 38764 24592 38804 24632
rect 38668 24508 38708 24548
rect 37996 21820 38036 21860
rect 38092 21652 38132 21692
rect 38188 21568 38228 21608
rect 39052 24627 39092 24632
rect 39052 24592 39092 24627
rect 39532 24592 39572 24632
rect 40300 27028 40340 27068
rect 40876 28876 40916 28916
rect 40588 28288 40628 28328
rect 40492 27700 40532 27740
rect 40780 27616 40820 27656
rect 40972 27448 41012 27488
rect 41068 26776 41108 26816
rect 42220 29716 42260 29756
rect 42124 29044 42164 29084
rect 41452 28792 41492 28832
rect 41452 28288 41492 28328
rect 41644 28120 41684 28160
rect 41548 27616 41588 27656
rect 41260 26692 41300 26732
rect 40204 26608 40244 26648
rect 40396 26608 40436 26648
rect 40300 25852 40340 25892
rect 40300 25264 40340 25304
rect 40588 26104 40628 26144
rect 41452 26188 41492 26228
rect 41356 26104 41396 26144
rect 40684 25852 40724 25892
rect 40588 25432 40628 25472
rect 40780 25264 40820 25304
rect 40588 25180 40628 25220
rect 40108 24760 40148 24800
rect 40492 24760 40532 24800
rect 40012 24508 40052 24548
rect 39532 24340 39572 24380
rect 39724 24340 39764 24380
rect 39244 23416 39284 23456
rect 40972 24844 41012 24884
rect 40780 24592 40820 24632
rect 41068 24676 41108 24716
rect 40492 24340 40532 24380
rect 41644 26356 41684 26396
rect 42700 29716 42740 29756
rect 42316 29212 42356 29252
rect 42604 29632 42644 29672
rect 42508 28960 42548 29000
rect 42796 29044 42836 29084
rect 42700 28792 42740 28832
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 43372 30388 43412 30428
rect 43084 29044 43124 29084
rect 42988 28792 43028 28832
rect 43276 29800 43316 29840
rect 43276 29296 43316 29336
rect 42988 28372 43028 28412
rect 43180 28288 43220 28328
rect 43756 30136 43796 30176
rect 45772 30388 45812 30428
rect 45292 30220 45332 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 44812 30136 44852 30176
rect 46252 29968 46292 30008
rect 46636 29968 46676 30008
rect 43756 29716 43796 29756
rect 43756 29296 43796 29336
rect 44236 29296 44276 29336
rect 43468 28372 43508 28412
rect 42316 28204 42356 28244
rect 42508 28204 42548 28244
rect 42124 28120 42164 28160
rect 42220 27700 42260 27740
rect 41932 27448 41972 27488
rect 42028 26776 42068 26816
rect 41836 26272 41876 26312
rect 41932 26188 41972 26228
rect 41452 24844 41492 24884
rect 41644 25264 41684 25304
rect 41548 24760 41588 24800
rect 43756 28456 43796 28496
rect 43564 28204 43604 28244
rect 43852 28288 43892 28328
rect 45292 29128 45332 29168
rect 45196 28456 45236 28496
rect 44140 28373 44180 28412
rect 44140 28372 44180 28373
rect 44044 28288 44084 28328
rect 44332 28372 44372 28412
rect 43564 27112 43604 27152
rect 42988 27028 43028 27068
rect 44140 27028 44180 27068
rect 42796 26944 42836 26984
rect 43468 26944 43508 26984
rect 43756 26944 43796 26984
rect 43372 26860 43412 26900
rect 43276 26692 43316 26732
rect 42892 26104 42932 26144
rect 43084 26104 43124 26144
rect 42316 26020 42356 26060
rect 42028 25768 42068 25808
rect 42700 25768 42740 25808
rect 43852 26608 43892 26648
rect 45100 27784 45140 27824
rect 44236 26692 44276 26732
rect 44428 26692 44468 26732
rect 43948 26440 43988 26480
rect 43948 25936 43988 25976
rect 43756 25768 43796 25808
rect 43372 25348 43412 25388
rect 42892 25264 42932 25304
rect 41260 24592 41300 24632
rect 43084 24760 43124 24800
rect 41932 24676 41972 24716
rect 41452 24508 41492 24548
rect 41740 24592 41780 24632
rect 40972 24424 41012 24464
rect 41548 24424 41588 24464
rect 41932 24424 41972 24464
rect 41260 24340 41300 24380
rect 40108 23752 40148 23792
rect 38764 22324 38804 22364
rect 38572 22240 38612 22280
rect 38668 21820 38708 21860
rect 38380 21652 38420 21692
rect 38476 21484 38516 21524
rect 38284 21064 38324 21104
rect 37996 20728 38036 20768
rect 38188 20560 38228 20600
rect 37996 20308 38036 20348
rect 37420 20056 37460 20096
rect 38092 20056 38132 20096
rect 38380 20140 38420 20180
rect 37900 19972 37940 20012
rect 38572 20056 38612 20096
rect 38476 19804 38516 19844
rect 37804 18796 37844 18836
rect 36844 18544 36884 18584
rect 37996 19468 38036 19508
rect 36844 18376 36884 18416
rect 37420 18544 37460 18584
rect 39148 22072 39188 22112
rect 39052 21820 39092 21860
rect 39052 20728 39092 20768
rect 38860 20560 38900 20600
rect 38764 20308 38804 20348
rect 38860 19972 38900 20012
rect 40492 23080 40532 23120
rect 39724 22660 39764 22700
rect 40396 22660 40436 22700
rect 39916 22324 39956 22364
rect 40876 23668 40916 23708
rect 41068 22408 41108 22448
rect 40780 22324 40820 22364
rect 39340 21736 39380 21776
rect 39436 21568 39476 21608
rect 39340 20980 39380 21020
rect 39436 20728 39476 20768
rect 39820 20812 39860 20852
rect 40108 22156 40148 22196
rect 40876 22240 40916 22280
rect 40972 21820 41012 21860
rect 40492 21736 40532 21776
rect 40300 21652 40340 21692
rect 40204 21568 40244 21608
rect 40108 21400 40148 21440
rect 40396 21568 40436 21608
rect 40972 21652 41012 21692
rect 41356 23752 41396 23792
rect 41164 22156 41204 22196
rect 41164 21820 41204 21860
rect 40876 21400 40916 21440
rect 42028 23752 42068 23792
rect 41548 23584 41588 23624
rect 41932 23080 41972 23120
rect 41644 22912 41684 22952
rect 42604 23668 42644 23708
rect 42220 23584 42260 23624
rect 43276 23752 43316 23792
rect 42604 23080 42644 23120
rect 43084 23080 43124 23120
rect 42124 22576 42164 22616
rect 42508 22576 42548 22616
rect 41932 22408 41972 22448
rect 41836 22324 41876 22364
rect 41740 22240 41780 22280
rect 42124 22072 42164 22112
rect 41260 21484 41300 21524
rect 41164 21148 41204 21188
rect 41068 20728 41108 20768
rect 38956 19468 38996 19508
rect 38668 19384 38708 19424
rect 38380 19300 38420 19340
rect 38476 19216 38516 19256
rect 38956 19300 38996 19340
rect 38860 19132 38900 19172
rect 38956 18964 38996 19004
rect 39628 19636 39668 19676
rect 40108 19384 40148 19424
rect 39532 19216 39572 19256
rect 39628 19132 39668 19172
rect 38284 18880 38324 18920
rect 39148 18880 39188 18920
rect 38476 18796 38516 18836
rect 37708 17704 37748 17744
rect 36844 16780 36884 16820
rect 37036 16948 37076 16988
rect 36940 16024 36980 16064
rect 36940 15436 36980 15476
rect 36844 15184 36884 15224
rect 36748 15100 36788 15140
rect 36940 14848 36980 14888
rect 36652 14008 36692 14048
rect 36844 14008 36884 14048
rect 36556 13840 36596 13880
rect 36652 13756 36692 13796
rect 36460 13168 36500 13208
rect 36364 13084 36404 13124
rect 36268 11488 36308 11528
rect 36172 11320 36212 11360
rect 37228 16108 37268 16148
rect 37420 16024 37460 16064
rect 37420 15520 37460 15560
rect 37036 13336 37076 13376
rect 36940 13168 36980 13208
rect 36652 12076 36692 12116
rect 37324 13420 37364 13460
rect 37324 13168 37364 13208
rect 37996 15352 38036 15392
rect 37612 14932 37652 14972
rect 37804 14932 37844 14972
rect 37516 14764 37556 14804
rect 37900 14848 37940 14888
rect 37612 14512 37652 14552
rect 38284 15520 38324 15560
rect 38380 14848 38420 14888
rect 38188 14764 38228 14804
rect 38284 14176 38324 14216
rect 39148 18544 39188 18584
rect 38860 17704 38900 17744
rect 40012 19216 40052 19256
rect 40492 19216 40532 19256
rect 40396 19132 40436 19172
rect 39916 18880 39956 18920
rect 40204 18880 40244 18920
rect 41740 20308 41780 20348
rect 41644 20056 41684 20096
rect 41932 20224 41972 20264
rect 41260 19804 41300 19844
rect 41836 19720 41876 19760
rect 40684 18880 40724 18920
rect 40300 18292 40340 18332
rect 38572 17032 38612 17072
rect 41932 19216 41972 19256
rect 42220 20560 42260 20600
rect 42508 21736 42548 21776
rect 44332 26356 44372 26396
rect 44236 26188 44276 26228
rect 43564 25180 43604 25220
rect 44332 25180 44372 25220
rect 44524 26440 44564 26480
rect 44716 26944 44756 26984
rect 44716 26440 44756 26480
rect 44620 26272 44660 26312
rect 44620 26020 44660 26060
rect 45388 27616 45428 27656
rect 45292 27364 45332 27404
rect 45004 26860 45044 26900
rect 45388 26944 45428 26984
rect 45580 27196 45620 27236
rect 45004 26608 45044 26648
rect 47116 29128 47156 29168
rect 47404 28456 47444 28496
rect 46540 28288 46580 28328
rect 47116 28288 47156 28328
rect 45868 28204 45908 28244
rect 46060 27196 46100 27236
rect 45964 26944 46004 26984
rect 45868 26776 45908 26816
rect 45964 26692 46004 26732
rect 45580 26524 45620 26564
rect 46060 26272 46100 26312
rect 45964 25936 46004 25976
rect 45580 25852 45620 25892
rect 47500 27700 47540 27740
rect 46252 27616 46292 27656
rect 46732 27364 46772 27404
rect 46540 27028 46580 27068
rect 46732 26944 46772 26984
rect 46444 26356 46484 26396
rect 46252 25516 46292 25556
rect 46156 25348 46196 25388
rect 45772 25180 45812 25220
rect 45964 25180 46004 25220
rect 45484 25096 45524 25136
rect 43564 22828 43604 22868
rect 43660 22744 43700 22784
rect 42988 22324 43028 22364
rect 42412 20560 42452 20600
rect 42316 19384 42356 19424
rect 42220 19216 42260 19256
rect 43948 23080 43988 23120
rect 44236 22912 44276 22952
rect 44140 22828 44180 22868
rect 45676 23836 45716 23876
rect 45196 23752 45236 23792
rect 44428 22660 44468 22700
rect 45196 22576 45236 22616
rect 43852 22408 43892 22448
rect 44044 22408 44084 22448
rect 44524 22408 44564 22448
rect 45004 22408 45044 22448
rect 43756 22324 43796 22364
rect 43660 22240 43700 22280
rect 43468 22156 43508 22196
rect 43180 22072 43220 22112
rect 42892 21400 42932 21440
rect 42892 20980 42932 21020
rect 43372 21568 43412 21608
rect 43852 22156 43892 22196
rect 43468 21484 43508 21524
rect 42796 20560 42836 20600
rect 43276 20728 43316 20768
rect 43084 20224 43124 20264
rect 42508 19720 42548 19760
rect 43180 19636 43220 19676
rect 42892 19384 42932 19424
rect 41644 18544 41684 18584
rect 42124 18544 42164 18584
rect 41068 18292 41108 18332
rect 41356 17704 41396 17744
rect 42892 17704 42932 17744
rect 42988 17620 43028 17660
rect 40300 17032 40340 17072
rect 43372 20056 43412 20096
rect 44140 22240 44180 22280
rect 44236 21568 44276 21608
rect 44332 21484 44372 21524
rect 44044 21400 44084 21440
rect 43756 20560 43796 20600
rect 44524 21400 44564 21440
rect 44620 20560 44660 20600
rect 43948 20308 43988 20348
rect 43852 19636 43892 19676
rect 43852 19468 43892 19508
rect 44236 19384 44276 19424
rect 43852 19216 43892 19256
rect 45772 23752 45812 23792
rect 45388 22408 45428 22448
rect 45388 22156 45428 22196
rect 45004 21652 45044 21692
rect 45292 21568 45332 21608
rect 44908 21148 44948 21188
rect 45388 20728 45428 20768
rect 45964 23752 46004 23792
rect 45868 23500 45908 23540
rect 46156 25180 46196 25220
rect 46444 25264 46484 25304
rect 46348 25180 46388 25220
rect 46540 25096 46580 25136
rect 47020 26860 47060 26900
rect 46828 26440 46868 26480
rect 47212 26440 47252 26480
rect 47404 26440 47444 26480
rect 47404 26188 47444 26228
rect 47116 26104 47156 26144
rect 47020 25516 47060 25556
rect 46924 25348 46964 25388
rect 47404 25684 47444 25724
rect 47212 25600 47252 25640
rect 46828 25180 46868 25220
rect 46732 24676 46772 24716
rect 46540 24592 46580 24632
rect 47692 28288 47732 28328
rect 47692 26356 47732 26396
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 47884 29296 47924 29336
rect 48460 29296 48500 29336
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 48268 28456 48308 28496
rect 49228 28456 49268 28496
rect 48940 28372 48980 28412
rect 48748 28288 48788 28328
rect 50284 28288 50324 28328
rect 50572 28288 50612 28328
rect 49036 27784 49076 27824
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 49132 27028 49172 27068
rect 48172 26944 48212 26984
rect 47980 26692 48020 26732
rect 48940 26692 48980 26732
rect 47884 26440 47924 26480
rect 48268 26272 48308 26312
rect 48076 26104 48116 26144
rect 49036 26104 49076 26144
rect 47884 26020 47924 26060
rect 47884 25768 47924 25808
rect 47788 25684 47828 25724
rect 47596 25600 47636 25640
rect 47500 25432 47540 25472
rect 47596 25264 47636 25304
rect 47788 25264 47828 25304
rect 48076 25936 48116 25976
rect 49132 25936 49172 25976
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 50284 27700 50324 27740
rect 49708 26776 49748 26816
rect 49324 26692 49364 26732
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 48268 25600 48308 25640
rect 48844 25516 48884 25556
rect 48268 25432 48308 25472
rect 47212 24592 47252 24632
rect 46540 23836 46580 23876
rect 47308 23836 47348 23876
rect 46156 23584 46196 23624
rect 45676 22660 45716 22700
rect 46060 22660 46100 22700
rect 45772 22576 45812 22616
rect 47212 23668 47252 23708
rect 46540 23500 46580 23540
rect 46348 23248 46388 23288
rect 46252 22324 46292 22364
rect 46348 22240 46388 22280
rect 46828 23248 46868 23288
rect 47020 23332 47060 23372
rect 46924 23080 46964 23120
rect 47116 23248 47156 23288
rect 47020 22240 47060 22280
rect 47500 24424 47540 24464
rect 47692 24424 47732 24464
rect 47788 24340 47828 24380
rect 47596 23584 47636 23624
rect 47404 23332 47444 23372
rect 47308 22912 47348 22952
rect 47212 22660 47252 22700
rect 46540 22156 46580 22196
rect 47596 23080 47636 23120
rect 47500 22744 47540 22784
rect 47500 22576 47540 22616
rect 48748 24676 48788 24716
rect 48364 24340 48404 24380
rect 49420 25516 49460 25556
rect 50092 25852 50132 25892
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 50572 27028 50612 27068
rect 51148 27028 51188 27068
rect 50476 25768 50516 25808
rect 49804 25264 49844 25304
rect 50956 26104 50996 26144
rect 51724 27028 51764 27068
rect 51436 26776 51476 26816
rect 51244 26524 51284 26564
rect 50764 25516 50804 25556
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 51148 25432 51188 25472
rect 49420 25180 49460 25220
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 48172 23920 48212 23960
rect 47884 23836 47924 23876
rect 50476 23836 50516 23876
rect 48172 23080 48212 23120
rect 48364 22912 48404 22952
rect 48076 22744 48116 22784
rect 46252 21736 46292 21776
rect 47212 21736 47252 21776
rect 47404 21736 47444 21776
rect 45580 21652 45620 21692
rect 46348 21652 46388 21692
rect 47020 21568 47060 21608
rect 46540 21400 46580 21440
rect 46348 20728 46388 20768
rect 45484 20056 45524 20096
rect 46348 20056 46388 20096
rect 47596 21652 47636 21692
rect 47692 21568 47732 21608
rect 50188 23584 50228 23624
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 49036 23080 49076 23120
rect 51820 25264 51860 25304
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 51724 23920 51764 23960
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 50476 23080 50516 23120
rect 48940 22744 48980 22784
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 49036 22408 49076 22448
rect 47980 22156 48020 22196
rect 49228 22156 49268 22196
rect 49036 22072 49076 22112
rect 47980 21652 48020 21692
rect 48652 21484 48692 21524
rect 49036 21400 49076 21440
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 51628 22408 51668 22448
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 50284 21484 50324 21524
rect 49900 21400 49940 21440
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 49036 20728 49076 20768
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 47116 20560 47156 20600
rect 47788 20560 47828 20600
rect 45100 19384 45140 19424
rect 44236 19216 44276 19256
rect 44716 18544 44756 18584
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 47788 19888 47828 19928
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 46348 19384 46388 19424
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 46732 18544 46772 18584
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 44620 17620 44660 17660
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 39532 16948 39572 16988
rect 39724 16948 39764 16988
rect 38956 14848 38996 14888
rect 39724 14848 39764 14888
rect 37996 14092 38036 14132
rect 37612 13756 37652 13796
rect 37804 13168 37844 13208
rect 38572 14092 38612 14132
rect 37324 12496 37364 12536
rect 36940 11992 36980 12032
rect 37132 12160 37172 12200
rect 37228 12076 37268 12116
rect 37036 11740 37076 11780
rect 36652 11488 36692 11528
rect 36556 11404 36596 11444
rect 36652 11236 36692 11276
rect 36172 11152 36212 11192
rect 36364 11152 36404 11192
rect 35596 10900 35636 10940
rect 34924 10480 34964 10520
rect 35308 10480 35348 10520
rect 35020 10312 35060 10352
rect 34060 10060 34100 10100
rect 35404 10144 35444 10184
rect 35692 10144 35732 10184
rect 35793 10144 35833 10184
rect 35308 10060 35348 10100
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 33580 9220 33620 9260
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 33580 8800 33620 8840
rect 34060 8800 34100 8840
rect 33772 8716 33812 8756
rect 32812 8296 32852 8336
rect 32524 6784 32564 6824
rect 32332 6532 32372 6572
rect 32043 6280 32083 6320
rect 31660 6196 31700 6236
rect 31084 5944 31124 5984
rect 32044 6028 32084 6068
rect 31948 5944 31988 5984
rect 31180 5776 31220 5816
rect 31564 5776 31604 5816
rect 31852 5776 31892 5816
rect 31084 5608 31124 5648
rect 30316 4852 30356 4892
rect 30988 5020 31028 5060
rect 31084 4936 31124 4976
rect 30892 4768 30932 4808
rect 30988 4180 31028 4220
rect 30796 3676 30836 3716
rect 31948 5608 31988 5648
rect 32140 5524 32180 5564
rect 31564 4936 31604 4976
rect 31468 4852 31508 4892
rect 31852 4516 31892 4556
rect 31660 4096 31700 4136
rect 31468 3928 31508 3968
rect 31276 3844 31316 3884
rect 31084 3760 31124 3800
rect 31180 3676 31220 3716
rect 31372 3676 31412 3716
rect 30988 3424 31028 3464
rect 29932 3004 29972 3044
rect 30124 3004 30164 3044
rect 30316 3004 30356 3044
rect 31276 3424 31316 3464
rect 31660 3844 31700 3884
rect 31372 3340 31412 3380
rect 31564 3424 31604 3464
rect 31468 2752 31508 2792
rect 31180 2584 31220 2624
rect 28876 2500 28916 2540
rect 30124 1912 30164 1952
rect 31756 3760 31796 3800
rect 31948 3760 31988 3800
rect 32044 3424 32084 3464
rect 34732 8968 34772 9008
rect 34348 8884 34388 8924
rect 34252 8716 34292 8756
rect 34060 8380 34100 8420
rect 33868 8212 33908 8252
rect 35116 9472 35156 9512
rect 35020 9304 35060 9344
rect 34924 8716 34964 8756
rect 35020 8632 35060 8672
rect 34444 8464 34484 8504
rect 35212 8632 35252 8672
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 33580 7792 33620 7832
rect 34060 7792 34100 7832
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 32812 6868 32852 6908
rect 32716 6448 32756 6488
rect 32428 6112 32468 6152
rect 32620 6112 32660 6152
rect 32620 5944 32660 5984
rect 32524 5776 32564 5816
rect 32332 5440 32372 5480
rect 33004 6196 33044 6236
rect 32812 6112 32852 6152
rect 32620 5356 32660 5396
rect 32236 5272 32276 5312
rect 32716 5020 32756 5060
rect 32908 6028 32948 6068
rect 33196 7120 33236 7160
rect 34348 7792 34388 7832
rect 34252 7540 34292 7580
rect 34348 7372 34388 7412
rect 34828 8128 34868 8168
rect 35308 8128 35348 8168
rect 34540 7372 34580 7412
rect 34156 7120 34196 7160
rect 34828 7960 34868 8000
rect 34636 7204 34676 7244
rect 33196 6784 33236 6824
rect 34060 6868 34100 6908
rect 34540 7120 34580 7160
rect 36172 10984 36212 11024
rect 36364 10984 36404 11024
rect 36268 10816 36308 10856
rect 36076 10312 36116 10352
rect 35980 10144 36020 10184
rect 35596 9808 35636 9848
rect 35884 9640 35924 9680
rect 35788 9472 35828 9512
rect 35884 9304 35924 9344
rect 35596 8632 35636 8672
rect 35788 9136 35828 9176
rect 37036 11236 37076 11276
rect 36940 11068 36980 11108
rect 36844 10984 36884 11024
rect 36652 10900 36692 10940
rect 37132 11068 37172 11108
rect 37324 11992 37364 12032
rect 37516 12580 37556 12620
rect 38188 12580 38228 12620
rect 37996 12496 38036 12536
rect 37516 12412 37556 12452
rect 38188 12244 38228 12284
rect 37612 12160 37652 12200
rect 36748 10816 36788 10856
rect 37228 10732 37268 10772
rect 36556 10396 36596 10436
rect 36364 10312 36404 10352
rect 36844 10312 36884 10352
rect 36556 10228 36596 10268
rect 36364 10144 36404 10184
rect 36268 9640 36308 9680
rect 36748 10144 36788 10184
rect 37324 10396 37364 10436
rect 37900 11656 37940 11696
rect 37612 11236 37652 11276
rect 37516 10984 37556 11024
rect 37516 10648 37556 10688
rect 37420 10312 37460 10352
rect 37420 10144 37460 10184
rect 37708 10816 37748 10856
rect 37612 10564 37652 10604
rect 37708 10396 37748 10436
rect 36652 9976 36692 10016
rect 35500 8464 35540 8504
rect 37228 9976 37268 10016
rect 35788 8296 35828 8336
rect 35596 8128 35636 8168
rect 35116 7792 35156 7832
rect 35116 7624 35156 7664
rect 35020 7204 35060 7244
rect 35404 7204 35444 7244
rect 35308 7120 35348 7160
rect 35116 7036 35156 7076
rect 34156 6784 34196 6824
rect 34348 6784 34388 6824
rect 33196 6280 33236 6320
rect 33868 6280 33908 6320
rect 33100 6112 33140 6152
rect 33004 5608 33044 5648
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 33484 5776 33524 5816
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 34636 6616 34676 6656
rect 35020 6616 35060 6656
rect 34732 6532 34772 6572
rect 34540 5944 34580 5984
rect 35020 6448 35060 6488
rect 35308 6952 35348 6992
rect 34828 5944 34868 5984
rect 32812 4768 32852 4808
rect 33676 4768 33716 4808
rect 32908 4684 32948 4724
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 33868 4348 33908 4388
rect 32716 4180 32756 4220
rect 32908 4096 32948 4136
rect 32140 3004 32180 3044
rect 32044 2920 32084 2960
rect 33580 3592 33620 3632
rect 34924 5608 34964 5648
rect 35020 5440 35060 5480
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 35308 6280 35348 6320
rect 35404 6196 35444 6236
rect 35212 5608 35252 5648
rect 34252 4936 34292 4976
rect 34252 4348 34292 4388
rect 34924 5020 34964 5060
rect 35116 5020 35156 5060
rect 34540 4432 34580 4472
rect 35404 5776 35444 5816
rect 36076 8380 36116 8420
rect 36556 8380 36596 8420
rect 35884 8128 35924 8168
rect 35692 7540 35732 7580
rect 35980 7960 36020 8000
rect 35884 7876 35924 7916
rect 35884 7624 35924 7664
rect 35788 7288 35828 7328
rect 36212 8128 36252 8168
rect 36364 8128 36404 8168
rect 36364 7876 36404 7916
rect 36460 7792 36500 7832
rect 36556 7708 36596 7748
rect 35980 7036 36020 7076
rect 35980 6784 36020 6824
rect 35596 6532 35636 6572
rect 35788 6532 35828 6572
rect 35884 6448 35924 6488
rect 35788 6280 35828 6320
rect 35692 5944 35732 5984
rect 35404 5608 35444 5648
rect 35500 5524 35540 5564
rect 34060 3592 34100 3632
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 33292 2836 33332 2876
rect 32812 2584 32852 2624
rect 33100 2584 33140 2624
rect 32236 2500 32276 2540
rect 32812 1912 32852 1952
rect 34444 3928 34484 3968
rect 34924 3928 34964 3968
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 35308 3928 35348 3968
rect 36076 6616 36116 6656
rect 36076 6280 36116 6320
rect 35980 5608 36020 5648
rect 36268 6952 36308 6992
rect 36364 5776 36404 5816
rect 36172 5440 36212 5480
rect 36364 4936 36404 4976
rect 36940 7960 36980 8000
rect 37708 10228 37748 10268
rect 37996 11068 38036 11108
rect 37804 9388 37844 9428
rect 37036 7876 37076 7916
rect 36940 7792 36980 7832
rect 37324 7372 37364 7412
rect 36844 7120 36884 7160
rect 37420 7288 37460 7328
rect 36748 6868 36788 6908
rect 36748 6616 36788 6656
rect 36652 5524 36692 5564
rect 35884 4096 35924 4136
rect 36268 3928 36308 3968
rect 36172 3424 36212 3464
rect 34540 2584 34580 2624
rect 36652 4096 36692 4136
rect 36652 3424 36692 3464
rect 36460 2584 36500 2624
rect 37996 9304 38036 9344
rect 37900 8800 37940 8840
rect 38380 10984 38420 11024
rect 38860 14008 38900 14048
rect 38668 13924 38708 13964
rect 38668 12580 38708 12620
rect 39724 14344 39764 14384
rect 39628 14008 39668 14048
rect 39052 13756 39092 13796
rect 38956 12664 38996 12704
rect 38860 12580 38900 12620
rect 38764 12496 38804 12536
rect 39244 12496 39284 12536
rect 41644 15520 41684 15560
rect 42604 15520 42644 15560
rect 43948 15520 43988 15560
rect 40972 14848 41012 14888
rect 41260 14764 41300 14804
rect 40492 14680 40532 14720
rect 40684 14512 40724 14552
rect 40876 14548 40916 14552
rect 40876 14512 40916 14548
rect 41068 14176 41108 14216
rect 40972 13924 41012 13964
rect 39436 12328 39476 12368
rect 38956 12244 38996 12284
rect 39244 12244 39284 12284
rect 40684 12580 40724 12620
rect 40396 12412 40436 12452
rect 38764 11656 38804 11696
rect 38572 11068 38612 11108
rect 38188 10732 38228 10772
rect 38188 10480 38228 10520
rect 38956 11152 38996 11192
rect 38764 10648 38804 10688
rect 38188 10144 38228 10184
rect 38668 10060 38708 10100
rect 38572 9388 38612 9428
rect 39148 10396 39188 10436
rect 39052 10060 39092 10100
rect 39436 11656 39476 11696
rect 39532 11152 39572 11192
rect 40300 11656 40340 11696
rect 39724 11572 39764 11612
rect 39628 10144 39668 10184
rect 38668 9304 38708 9344
rect 39244 9388 39284 9428
rect 37611 7204 37651 7244
rect 37900 7960 37940 8000
rect 37804 7540 37844 7580
rect 38092 7540 38132 7580
rect 37996 7372 38036 7412
rect 37900 7204 37940 7244
rect 37612 6952 37652 6992
rect 37324 6532 37364 6572
rect 37516 6532 37556 6572
rect 36844 6448 36884 6488
rect 36940 6196 36980 6236
rect 37612 6448 37652 6488
rect 38092 7204 38132 7244
rect 38284 8464 38324 8504
rect 38284 7960 38324 8000
rect 38956 8800 38996 8840
rect 38956 8296 38996 8336
rect 38764 8212 38804 8252
rect 38572 7540 38612 7580
rect 38188 7120 38228 7160
rect 37900 6700 37940 6740
rect 37804 6364 37844 6404
rect 37132 5608 37172 5648
rect 37228 4264 37268 4304
rect 37612 5608 37652 5648
rect 37420 5020 37460 5060
rect 37900 6196 37940 6236
rect 38380 5776 38420 5816
rect 40012 11152 40052 11192
rect 40204 10984 40244 11024
rect 39820 10648 39860 10688
rect 41356 14008 41396 14048
rect 41452 12916 41492 12956
rect 41452 12496 41492 12536
rect 40492 11572 40532 11612
rect 40684 11488 40724 11528
rect 40684 10984 40724 11024
rect 41068 9892 41108 9932
rect 41164 8800 41204 8840
rect 40012 8632 40052 8672
rect 39436 8128 39476 8168
rect 38764 7288 38804 7328
rect 38668 7204 38708 7244
rect 38572 6700 38612 6740
rect 38572 6448 38612 6488
rect 39436 7120 39476 7160
rect 38476 5692 38516 5732
rect 38668 5608 38708 5648
rect 37804 5104 37844 5144
rect 37612 3760 37652 3800
rect 37420 2836 37460 2876
rect 37804 4012 37844 4052
rect 37900 3844 37940 3884
rect 38188 5356 38228 5396
rect 38284 5104 38324 5144
rect 38380 4936 38420 4976
rect 38380 3928 38420 3968
rect 38284 3844 38324 3884
rect 38092 3760 38132 3800
rect 37996 2836 38036 2876
rect 37996 2584 38036 2624
rect 38668 5020 38708 5060
rect 39628 8044 39668 8084
rect 40204 8464 40244 8504
rect 40876 8296 40916 8336
rect 41068 8296 41108 8336
rect 41068 8128 41108 8168
rect 40204 7960 40244 8000
rect 41356 9976 41396 10016
rect 41548 12328 41588 12368
rect 41548 11488 41588 11528
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 42124 14764 42164 14804
rect 42988 14680 43028 14720
rect 41836 14176 41876 14216
rect 41740 13924 41780 13964
rect 41932 14008 41972 14048
rect 42028 13840 42068 13880
rect 41740 13000 41780 13040
rect 42028 13168 42068 13208
rect 42508 13840 42548 13880
rect 42796 13840 42836 13880
rect 42412 13336 42452 13376
rect 42124 13000 42164 13040
rect 41836 12580 41876 12620
rect 41932 12412 41972 12452
rect 41836 12328 41876 12368
rect 41740 11572 41780 11612
rect 41644 11068 41684 11108
rect 41644 10312 41684 10352
rect 42508 13168 42548 13208
rect 42508 12664 42548 12704
rect 42124 12328 42164 12368
rect 42028 12076 42068 12116
rect 42700 12496 42740 12536
rect 42604 12328 42644 12368
rect 42508 12244 42548 12284
rect 42700 12244 42740 12284
rect 42412 11992 42452 12032
rect 42028 11908 42068 11948
rect 42220 11908 42260 11948
rect 42700 11992 42740 12032
rect 42508 11740 42548 11780
rect 42124 11656 42164 11696
rect 42220 11404 42260 11444
rect 42124 11236 42164 11276
rect 42508 11320 42548 11360
rect 41356 9388 41396 9428
rect 41740 9892 41780 9932
rect 41740 9640 41780 9680
rect 41548 8800 41588 8840
rect 41452 8716 41492 8756
rect 41356 8632 41396 8672
rect 41452 8044 41492 8084
rect 41260 7960 41300 8000
rect 41740 8464 41780 8504
rect 41644 7288 41684 7328
rect 40588 7204 40628 7244
rect 42220 10312 42260 10352
rect 42316 10228 42356 10268
rect 41932 7960 41972 8000
rect 42412 9472 42452 9512
rect 42604 10144 42644 10184
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 44428 14848 44468 14888
rect 44620 14764 44660 14804
rect 44236 14344 44276 14384
rect 43276 14008 43316 14048
rect 43180 13336 43220 13376
rect 43084 12580 43124 12620
rect 42988 12496 43028 12536
rect 42892 12328 42932 12368
rect 42892 12076 42932 12116
rect 42796 11320 42836 11360
rect 44140 14008 44180 14048
rect 43468 12580 43508 12620
rect 43468 12412 43508 12452
rect 43084 12076 43124 12116
rect 43852 13168 43892 13208
rect 44236 12580 44276 12620
rect 43564 12328 43604 12368
rect 43948 12076 43988 12116
rect 42892 10732 42932 10772
rect 42892 10396 42932 10436
rect 43180 10312 43220 10352
rect 43660 10984 43700 11024
rect 44428 13168 44468 13208
rect 43660 10732 43700 10772
rect 43564 10144 43604 10184
rect 43084 10060 43124 10100
rect 42988 9640 43028 9680
rect 42700 9304 42740 9344
rect 42508 8380 42548 8420
rect 41260 7036 41300 7076
rect 40972 6952 41012 6992
rect 39916 6028 39956 6068
rect 39532 5860 39572 5900
rect 38860 5524 38900 5564
rect 39820 5356 39860 5396
rect 39628 5020 39668 5060
rect 38764 4936 38804 4976
rect 39244 4936 39284 4976
rect 40684 6448 40724 6488
rect 40780 5692 40820 5732
rect 40876 5608 40916 5648
rect 41260 6448 41300 6488
rect 41644 6448 41684 6488
rect 41644 5860 41684 5900
rect 40492 5440 40532 5480
rect 40780 5356 40820 5396
rect 38764 4096 38804 4136
rect 39244 4096 39284 4136
rect 41932 7120 41972 7160
rect 42028 6364 42068 6404
rect 42220 6364 42260 6404
rect 42220 6028 42260 6068
rect 41836 5608 41876 5648
rect 42796 8800 42836 8840
rect 42700 8212 42740 8252
rect 42796 7960 42836 8000
rect 42988 9472 43028 9512
rect 43372 10012 43412 10016
rect 43372 9976 43412 10012
rect 43276 9388 43316 9428
rect 43180 9304 43220 9344
rect 42988 7792 43028 7832
rect 42700 7288 42740 7328
rect 42604 5608 42644 5648
rect 42892 7288 42932 7328
rect 43468 8716 43508 8756
rect 43372 8632 43412 8672
rect 43468 8464 43508 8504
rect 43468 7792 43508 7832
rect 44716 11908 44756 11948
rect 44812 11740 44852 11780
rect 45292 12496 45332 12536
rect 45100 12244 45140 12284
rect 45100 11320 45140 11360
rect 45676 13840 45716 13880
rect 45676 12496 45716 12536
rect 45772 11824 45812 11864
rect 46444 11824 46484 11864
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 46732 12496 46772 12536
rect 46636 11740 46676 11780
rect 46540 11656 46580 11696
rect 46444 11404 46484 11444
rect 45388 11152 45428 11192
rect 45964 11152 46004 11192
rect 46636 11152 46676 11192
rect 45004 10984 45044 11024
rect 45772 10816 45812 10856
rect 44428 10732 44468 10772
rect 44908 10732 44948 10772
rect 44140 10144 44180 10184
rect 44428 10144 44468 10184
rect 44044 9472 44084 9512
rect 44716 10060 44756 10100
rect 44428 9472 44468 9512
rect 45676 10312 45716 10352
rect 44620 9388 44660 9428
rect 45484 10060 45524 10100
rect 46156 10984 46196 11024
rect 46348 10564 46388 10604
rect 46636 10228 46676 10268
rect 45868 9220 45908 9260
rect 44236 8800 44276 8840
rect 43180 7036 43220 7076
rect 43468 6952 43508 6992
rect 43276 5608 43316 5648
rect 43948 8296 43988 8336
rect 45484 8632 45524 8672
rect 44812 8548 44852 8588
rect 45196 8548 45236 8588
rect 44044 7540 44084 7580
rect 43756 7120 43796 7160
rect 45772 8380 45812 8420
rect 46444 8800 46484 8840
rect 44524 6448 44564 6488
rect 44716 6448 44756 6488
rect 45292 6448 45332 6488
rect 44716 6280 44756 6320
rect 44236 6028 44276 6068
rect 43948 5608 43988 5648
rect 43660 5524 43700 5564
rect 45004 6028 45044 6068
rect 44908 5608 44948 5648
rect 46636 8128 46676 8168
rect 46732 7540 46772 7580
rect 46252 6532 46292 6572
rect 47116 11656 47156 11696
rect 47596 12496 47636 12536
rect 47308 11068 47348 11108
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 48652 12244 48692 12284
rect 49324 12160 49364 12200
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 47980 11404 48020 11444
rect 48844 11656 48884 11696
rect 48364 11404 48404 11444
rect 48172 11152 48212 11192
rect 47788 11068 47828 11108
rect 48076 11068 48116 11108
rect 47212 10564 47252 10604
rect 47692 10984 47732 11024
rect 46924 10060 46964 10100
rect 48076 10312 48116 10352
rect 48268 10984 48308 11024
rect 48460 11068 48500 11108
rect 48364 10816 48404 10856
rect 48268 10732 48308 10772
rect 47788 10144 47828 10184
rect 47692 10060 47732 10100
rect 47308 9220 47348 9260
rect 47116 8800 47156 8840
rect 46924 8128 46964 8168
rect 47116 8632 47156 8672
rect 46924 7540 46964 7580
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 48556 10732 48596 10772
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 48940 10396 48980 10436
rect 49036 10144 49076 10184
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 48172 8632 48212 8672
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 46828 6952 46868 6992
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 47116 6448 47156 6488
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 45580 5608 45620 5648
rect 44812 5524 44852 5564
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 39628 3928 39668 3968
rect 40492 3928 40532 3968
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 38476 2584 38516 2624
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 26860 1072 26900 1112
rect 27724 1072 27764 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 9667 38368 9676 38408
rect 9716 38368 11884 38408
rect 11924 38368 11933 38408
rect 10723 38032 10732 38072
rect 10772 38032 11596 38072
rect 11636 38032 11645 38072
rect 11395 37948 11404 37988
rect 11444 37948 12844 37988
rect 12884 37948 12893 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 11320 37780 11500 37820
rect 11540 37780 11549 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 11320 37736 11360 37780
rect 9763 37696 9772 37736
rect 9812 37696 11360 37736
rect 9859 37612 9868 37652
rect 9908 37612 10540 37652
rect 10580 37612 10589 37652
rect 0 37568 80 37588
rect 0 37528 268 37568
rect 308 37528 317 37568
rect 0 37508 80 37528
rect 7459 37276 7468 37316
rect 7508 37276 8332 37316
rect 8372 37276 8381 37316
rect 10051 37192 10060 37232
rect 10100 37192 10444 37232
rect 10484 37192 13996 37232
rect 14036 37192 14045 37232
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 15523 36856 15532 36896
rect 15572 36856 16396 36896
rect 16436 36856 16445 36896
rect 9859 36772 9868 36812
rect 9908 36772 10828 36812
rect 10868 36772 10877 36812
rect 16483 36772 16492 36812
rect 16532 36772 17548 36812
rect 17588 36772 17597 36812
rect 0 36729 80 36748
rect 0 36728 125 36729
rect 0 36688 76 36728
rect 116 36688 125 36728
rect 14947 36688 14956 36728
rect 14996 36688 15340 36728
rect 15380 36688 15389 36728
rect 15619 36688 15628 36728
rect 15668 36688 16684 36728
rect 16724 36688 16733 36728
rect 16867 36688 16876 36728
rect 16916 36688 18124 36728
rect 18164 36688 18173 36728
rect 0 36687 125 36688
rect 0 36668 80 36687
rect 6595 36604 6604 36644
rect 6644 36604 8044 36644
rect 8084 36604 8093 36644
rect 9571 36604 9580 36644
rect 9620 36604 10636 36644
rect 10676 36604 10685 36644
rect 6979 36520 6988 36560
rect 7028 36520 7564 36560
rect 7604 36520 7613 36560
rect 11395 36520 11404 36560
rect 11444 36520 11788 36560
rect 11828 36520 11837 36560
rect 13987 36520 13996 36560
rect 14036 36520 14860 36560
rect 14900 36520 14909 36560
rect 16003 36520 16012 36560
rect 16052 36520 17164 36560
rect 17204 36520 17213 36560
rect 9091 36436 9100 36476
rect 9140 36436 9964 36476
rect 10004 36436 10013 36476
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 11107 36016 11116 36056
rect 11156 36016 11360 36056
rect 18787 36016 18796 36056
rect 18836 36016 19180 36056
rect 19220 36016 19229 36056
rect 11320 35972 11360 36016
rect 6700 35932 8140 35972
rect 8180 35932 9196 35972
rect 9236 35932 9676 35972
rect 9716 35932 10156 35972
rect 10196 35932 10205 35972
rect 11320 35932 12844 35972
rect 12884 35932 12893 35972
rect 0 35828 80 35908
rect 6700 35888 6740 35932
rect 6691 35848 6700 35888
rect 6740 35848 6749 35888
rect 6883 35848 6892 35888
rect 6932 35848 6941 35888
rect 8323 35848 8332 35888
rect 8372 35848 9388 35888
rect 9428 35848 9437 35888
rect 11587 35848 11596 35888
rect 11636 35848 11645 35888
rect 17155 35848 17164 35888
rect 17204 35848 18316 35888
rect 18356 35848 18365 35888
rect 6892 35804 6932 35848
rect 11596 35804 11636 35848
rect 3427 35764 3436 35804
rect 3476 35764 3916 35804
rect 3956 35764 3965 35804
rect 6892 35764 8908 35804
rect 8948 35764 8957 35804
rect 10147 35764 10156 35804
rect 10196 35764 11212 35804
rect 11252 35764 11636 35804
rect 6307 35680 6316 35720
rect 6356 35680 6796 35720
rect 6836 35680 6845 35720
rect 8131 35680 8140 35720
rect 8180 35680 8524 35720
rect 8564 35680 8573 35720
rect 11107 35680 11116 35720
rect 11156 35680 14380 35720
rect 14420 35680 14956 35720
rect 14996 35680 15820 35720
rect 15860 35680 15869 35720
rect 21187 35680 21196 35720
rect 21236 35680 22348 35720
rect 22388 35680 22397 35720
rect 6403 35596 6412 35636
rect 6452 35596 7084 35636
rect 7124 35596 7133 35636
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 10915 35260 10924 35300
rect 10964 35260 11500 35300
rect 11540 35260 11549 35300
rect 16867 35260 16876 35300
rect 16916 35260 17068 35300
rect 17108 35260 17117 35300
rect 17539 35260 17548 35300
rect 17588 35260 18028 35300
rect 18068 35260 18077 35300
rect 18403 35260 18412 35300
rect 18452 35260 18988 35300
rect 19028 35260 19037 35300
rect 3331 35176 3340 35216
rect 3380 35176 3724 35216
rect 3764 35176 3773 35216
rect 5443 35176 5452 35216
rect 5492 35176 8428 35216
rect 8468 35176 8477 35216
rect 9859 35176 9868 35216
rect 9908 35176 11212 35216
rect 11252 35176 11261 35216
rect 11875 35176 11884 35216
rect 11924 35176 12364 35216
rect 12404 35176 13612 35216
rect 13652 35176 15340 35216
rect 15380 35176 15389 35216
rect 16195 35176 16204 35216
rect 16244 35176 16588 35216
rect 16628 35176 16637 35216
rect 16963 35176 16972 35216
rect 17012 35176 19660 35216
rect 19700 35176 20044 35216
rect 20084 35176 20093 35216
rect 23107 35176 23116 35216
rect 23156 35176 24076 35216
rect 24116 35176 24125 35216
rect 6595 35092 6604 35132
rect 6644 35092 6892 35132
rect 6932 35092 7756 35132
rect 7796 35092 7805 35132
rect 0 34988 80 35068
rect 6787 35048 6845 35049
rect 9868 35048 9908 35176
rect 10540 35048 10580 35176
rect 16588 35132 16628 35176
rect 16588 35092 17260 35132
rect 17300 35092 17309 35132
rect 6702 35008 6796 35048
rect 6836 35008 6845 35048
rect 7363 35008 7372 35048
rect 7412 35008 9908 35048
rect 10531 35008 10540 35048
rect 10580 35008 10589 35048
rect 13219 35008 13228 35048
rect 13268 35008 14956 35048
rect 14996 35008 15005 35048
rect 16483 35008 16492 35048
rect 16532 35008 16780 35048
rect 16820 35008 16829 35048
rect 26179 35008 26188 35048
rect 26228 35008 26668 35048
rect 26708 35008 26717 35048
rect 6787 35007 6845 35008
rect 3235 34924 3244 34964
rect 3284 34924 3628 34964
rect 3668 34924 3677 34964
rect 4675 34924 4684 34964
rect 4724 34924 7276 34964
rect 7316 34924 7468 34964
rect 7508 34924 7517 34964
rect 16675 34924 16684 34964
rect 16724 34924 17740 34964
rect 17780 34924 20812 34964
rect 20852 34924 21772 34964
rect 21812 34924 21821 34964
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 3811 34756 3820 34796
rect 3860 34756 5452 34796
rect 5492 34756 7660 34796
rect 7700 34756 7709 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 3907 34672 3916 34712
rect 3956 34672 5068 34712
rect 5108 34672 6508 34712
rect 6548 34672 6557 34712
rect 10147 34672 10156 34712
rect 10196 34672 10732 34712
rect 10772 34672 10781 34712
rect 4195 34588 4204 34628
rect 4244 34588 6796 34628
rect 6836 34588 6845 34628
rect 31267 34588 31276 34628
rect 31316 34588 31660 34628
rect 31700 34588 32140 34628
rect 32180 34588 32189 34628
rect 5251 34504 5260 34544
rect 5300 34504 5644 34544
rect 5684 34504 6988 34544
rect 7028 34504 7037 34544
rect 9379 34504 9388 34544
rect 9428 34504 10060 34544
rect 10100 34504 10109 34544
rect 18307 34504 18316 34544
rect 18356 34504 18365 34544
rect 18787 34504 18796 34544
rect 18836 34504 19660 34544
rect 19700 34504 19709 34544
rect 19939 34504 19948 34544
rect 19988 34504 21676 34544
rect 21716 34504 21725 34544
rect 18316 34460 18356 34504
rect 4771 34420 4780 34460
rect 4820 34420 6316 34460
rect 6356 34420 7372 34460
rect 7412 34420 7421 34460
rect 7564 34420 9580 34460
rect 9620 34420 9629 34460
rect 18316 34420 19372 34460
rect 19412 34420 19421 34460
rect 7564 34376 7604 34420
rect 3523 34336 3532 34376
rect 3572 34336 4492 34376
rect 4532 34336 4541 34376
rect 6211 34336 6220 34376
rect 6260 34336 7084 34376
rect 7124 34336 7133 34376
rect 7555 34336 7564 34376
rect 7604 34336 7613 34376
rect 9379 34336 9388 34376
rect 9428 34336 10444 34376
rect 10484 34336 10493 34376
rect 18595 34336 18604 34376
rect 18644 34336 18653 34376
rect 18787 34336 18796 34376
rect 18836 34336 19852 34376
rect 19892 34336 19901 34376
rect 20035 34336 20044 34376
rect 20084 34336 21196 34376
rect 21236 34336 21245 34376
rect 27043 34336 27052 34376
rect 27092 34336 30028 34376
rect 30068 34336 30508 34376
rect 30548 34336 33484 34376
rect 33524 34336 33772 34376
rect 33812 34336 33821 34376
rect 34147 34336 34156 34376
rect 34196 34336 36364 34376
rect 36404 34336 36413 34376
rect 36643 34336 36652 34376
rect 36692 34336 37804 34376
rect 37844 34336 37996 34376
rect 38036 34336 38045 34376
rect 18604 34292 18644 34336
rect 3619 34252 3628 34292
rect 3668 34252 6356 34292
rect 6499 34252 6508 34292
rect 6548 34252 8044 34292
rect 8084 34252 11020 34292
rect 11060 34252 11069 34292
rect 18604 34252 20140 34292
rect 20180 34252 21332 34292
rect 21379 34252 21388 34292
rect 21428 34252 22156 34292
rect 22196 34252 22205 34292
rect 0 34148 80 34228
rect 6316 34208 6356 34252
rect 21292 34208 21332 34252
rect 3907 34168 3916 34208
rect 3956 34168 3965 34208
rect 6307 34168 6316 34208
rect 6356 34168 6365 34208
rect 7459 34168 7468 34208
rect 7508 34168 7756 34208
rect 7796 34168 7805 34208
rect 16963 34168 16972 34208
rect 17012 34168 17260 34208
rect 17300 34168 17836 34208
rect 17876 34168 17885 34208
rect 19939 34168 19948 34208
rect 19988 34168 20524 34208
rect 20564 34168 20573 34208
rect 21292 34168 21580 34208
rect 21620 34168 21629 34208
rect 3916 34124 3956 34168
rect 6787 34124 6845 34125
rect 3916 34084 5492 34124
rect 6499 34084 6508 34124
rect 6548 34084 6796 34124
rect 6836 34084 6845 34124
rect 10051 34084 10060 34124
rect 10100 34084 11980 34124
rect 12020 34084 12029 34124
rect 12355 34084 12364 34124
rect 12404 34084 14572 34124
rect 14612 34084 14621 34124
rect 5452 34040 5492 34084
rect 6787 34083 6845 34084
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 5443 34000 5452 34040
rect 5492 34000 6988 34040
rect 7028 34000 7037 34040
rect 10723 34000 10732 34040
rect 10772 34000 11884 34040
rect 11924 34000 11933 34040
rect 13987 34000 13996 34040
rect 14036 34000 17548 34040
rect 17588 34000 17597 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 23779 34000 23788 34040
rect 23828 34000 24844 34040
rect 24884 34000 24893 34040
rect 27139 34000 27148 34040
rect 27188 34000 28204 34040
rect 28244 34000 29068 34040
rect 29108 34000 29117 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 4003 33916 4012 33956
rect 4052 33916 5548 33956
rect 5588 33916 5597 33956
rect 23683 33916 23692 33956
rect 23732 33916 24652 33956
rect 24692 33916 24701 33956
rect 5251 33832 5260 33872
rect 5300 33832 6124 33872
rect 6164 33832 6173 33872
rect 13123 33832 13132 33872
rect 13172 33832 13708 33872
rect 13748 33832 14092 33872
rect 14132 33832 14141 33872
rect 21763 33832 21772 33872
rect 21812 33832 23884 33872
rect 23924 33832 23933 33872
rect 28963 33832 28972 33872
rect 29012 33832 30220 33872
rect 30260 33832 30269 33872
rect 30787 33832 30796 33872
rect 30836 33832 30988 33872
rect 31028 33832 32044 33872
rect 32084 33832 32093 33872
rect 3523 33748 3532 33788
rect 3572 33748 3724 33788
rect 3764 33748 4012 33788
rect 4052 33748 5108 33788
rect 8131 33748 8140 33788
rect 8180 33748 8428 33788
rect 8468 33748 8477 33788
rect 21571 33748 21580 33788
rect 21620 33748 22252 33788
rect 22292 33748 22301 33788
rect 5068 33704 5108 33748
rect 3811 33664 3820 33704
rect 3860 33664 4780 33704
rect 4820 33664 4829 33704
rect 5059 33664 5068 33704
rect 5108 33664 5644 33704
rect 5684 33664 5836 33704
rect 5876 33664 5885 33704
rect 7459 33664 7468 33704
rect 7508 33664 7517 33704
rect 11779 33664 11788 33704
rect 11828 33664 12652 33704
rect 12692 33664 13036 33704
rect 13076 33664 15820 33704
rect 15860 33664 15869 33704
rect 18019 33664 18028 33704
rect 18068 33664 18700 33704
rect 18740 33664 18749 33704
rect 20227 33664 20236 33704
rect 20276 33664 22636 33704
rect 22676 33664 22685 33704
rect 23011 33664 23020 33704
rect 23060 33664 24076 33704
rect 24116 33664 24125 33704
rect 25507 33664 25516 33704
rect 25556 33664 26284 33704
rect 26324 33664 26333 33704
rect 29059 33664 29068 33704
rect 29108 33664 31084 33704
rect 31124 33664 31133 33704
rect 31363 33664 31372 33704
rect 31412 33664 32140 33704
rect 32180 33664 32620 33704
rect 32660 33664 32669 33704
rect 36643 33664 36652 33704
rect 36692 33664 38764 33704
rect 38804 33664 38813 33704
rect 7468 33620 7508 33664
rect 3619 33580 3628 33620
rect 3668 33580 6028 33620
rect 6068 33580 7508 33620
rect 24163 33580 24172 33620
rect 24212 33580 25804 33620
rect 25844 33580 26476 33620
rect 26516 33580 26525 33620
rect 9859 33496 9868 33536
rect 9908 33496 11692 33536
rect 11732 33496 11741 33536
rect 21763 33496 21772 33536
rect 21812 33496 23692 33536
rect 23732 33496 23741 33536
rect 25699 33496 25708 33536
rect 25748 33496 26188 33536
rect 26228 33496 26237 33536
rect 28579 33496 28588 33536
rect 28628 33496 29164 33536
rect 29204 33496 29213 33536
rect 29452 33496 31372 33536
rect 31412 33496 31421 33536
rect 1123 33412 1132 33452
rect 1172 33412 3820 33452
rect 3860 33412 3869 33452
rect 6115 33412 6124 33452
rect 6164 33412 6604 33452
rect 6644 33412 6653 33452
rect 0 33308 80 33388
rect 29452 33368 29492 33496
rect 38659 33412 38668 33452
rect 38708 33412 39628 33452
rect 39668 33412 39677 33452
rect 1219 33328 1228 33368
rect 1268 33328 5644 33368
rect 5684 33328 5693 33368
rect 28867 33328 28876 33368
rect 28916 33328 29452 33368
rect 29492 33328 29501 33368
rect 31363 33328 31372 33368
rect 31412 33328 34924 33368
rect 34964 33328 35884 33368
rect 35924 33328 35933 33368
rect 4867 33284 4925 33285
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 4782 33244 4876 33284
rect 4916 33244 4925 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 25795 33244 25804 33284
rect 25844 33244 28108 33284
rect 28148 33244 28157 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 4867 33243 4925 33244
rect 2467 33160 2476 33200
rect 2516 33160 5932 33200
rect 5972 33160 5981 33200
rect 9955 33160 9964 33200
rect 10004 33160 10348 33200
rect 10388 33160 12940 33200
rect 12980 33160 12989 33200
rect 1699 33076 1708 33116
rect 1748 33076 3244 33116
rect 3284 33076 3293 33116
rect 3715 33076 3724 33116
rect 3764 33076 4492 33116
rect 4532 33076 5068 33116
rect 5108 33076 5117 33116
rect 14563 33076 14572 33116
rect 14612 33076 15532 33116
rect 15572 33076 16492 33116
rect 16532 33076 16684 33116
rect 16724 33076 18220 33116
rect 18260 33076 18269 33116
rect 18787 33076 18796 33116
rect 18836 33076 19852 33116
rect 19892 33076 19901 33116
rect 24067 33076 24076 33116
rect 24116 33076 24844 33116
rect 24884 33076 24893 33116
rect 31171 33076 31180 33116
rect 31220 33076 31229 33116
rect 31651 33076 31660 33116
rect 31700 33076 33772 33116
rect 33812 33076 34348 33116
rect 34388 33076 34397 33116
rect 21283 33032 21341 33033
rect 31180 33032 31220 33076
rect 1987 32992 1996 33032
rect 2036 32992 4300 33032
rect 4340 32992 4349 33032
rect 6691 32992 6700 33032
rect 6740 32992 7276 33032
rect 7316 32992 7325 33032
rect 10627 32992 10636 33032
rect 10676 32992 12268 33032
rect 12308 32992 12317 33032
rect 19651 32992 19660 33032
rect 19700 32992 20524 33032
rect 20564 32992 20573 33032
rect 21198 32992 21292 33032
rect 21332 32992 21341 33032
rect 21667 32992 21676 33032
rect 21716 32992 23596 33032
rect 23636 32992 23980 33032
rect 24020 32992 24029 33032
rect 31180 32992 32780 33032
rect 33667 32992 33676 33032
rect 33716 32992 35980 33032
rect 36020 32992 36268 33032
rect 36308 32992 36317 33032
rect 21283 32991 21341 32992
rect 32740 32948 32780 32992
rect 3043 32908 3052 32948
rect 3092 32908 3532 32948
rect 3572 32908 3581 32948
rect 4099 32908 4108 32948
rect 4148 32908 6220 32948
rect 6260 32908 6269 32948
rect 9283 32908 9292 32948
rect 9332 32908 10348 32948
rect 10388 32908 10397 32948
rect 10924 32908 11692 32948
rect 11732 32908 12172 32948
rect 12212 32908 12221 32948
rect 19267 32908 19276 32948
rect 19316 32908 20908 32948
rect 20948 32908 20957 32948
rect 27043 32908 27052 32948
rect 27092 32908 28588 32948
rect 28628 32908 29644 32948
rect 29684 32908 29693 32948
rect 30211 32908 30220 32948
rect 30260 32908 31180 32948
rect 31220 32908 32044 32948
rect 32084 32908 32093 32948
rect 32740 32908 33292 32948
rect 33332 32908 33341 32948
rect 34147 32908 34156 32948
rect 34196 32908 36844 32948
rect 36884 32908 36893 32948
rect 10924 32864 10964 32908
rect 2659 32824 2668 32864
rect 2708 32824 2956 32864
rect 2996 32824 3005 32864
rect 3235 32824 3244 32864
rect 3284 32824 5164 32864
rect 5204 32824 5213 32864
rect 6499 32824 6508 32864
rect 6548 32824 9964 32864
rect 10004 32824 10013 32864
rect 10915 32824 10924 32864
rect 10964 32824 10973 32864
rect 11320 32824 11788 32864
rect 11828 32824 11837 32864
rect 12547 32824 12556 32864
rect 12596 32824 13612 32864
rect 13652 32824 13661 32864
rect 14371 32824 14380 32864
rect 14420 32824 14956 32864
rect 14996 32824 15005 32864
rect 16771 32824 16780 32864
rect 16820 32824 17260 32864
rect 17300 32824 17309 32864
rect 18403 32824 18412 32864
rect 18452 32824 19372 32864
rect 19412 32824 19421 32864
rect 21955 32824 21964 32864
rect 22004 32824 23500 32864
rect 23540 32824 23549 32864
rect 23971 32824 23980 32864
rect 24020 32824 24172 32864
rect 24212 32824 24221 32864
rect 24643 32824 24652 32864
rect 24692 32824 27436 32864
rect 27476 32824 28492 32864
rect 28532 32824 28541 32864
rect 28771 32824 28780 32864
rect 28820 32824 29260 32864
rect 29300 32824 29309 32864
rect 31651 32824 31660 32864
rect 31700 32824 33196 32864
rect 33236 32824 33245 32864
rect 33859 32824 33868 32864
rect 33908 32824 35116 32864
rect 35156 32824 35165 32864
rect 11320 32780 11360 32824
rect 19372 32780 19412 32824
rect 2851 32740 2860 32780
rect 2900 32740 5356 32780
rect 5396 32740 5405 32780
rect 7939 32740 7948 32780
rect 7988 32740 8812 32780
rect 8852 32740 8861 32780
rect 11011 32740 11020 32780
rect 11060 32740 11360 32780
rect 12067 32740 12076 32780
rect 12116 32740 13036 32780
rect 13076 32740 13085 32780
rect 16099 32740 16108 32780
rect 16148 32740 17356 32780
rect 17396 32740 17405 32780
rect 19372 32740 20236 32780
rect 20276 32740 20285 32780
rect 22243 32740 22252 32780
rect 22292 32740 24364 32780
rect 24404 32740 25708 32780
rect 25748 32740 25757 32780
rect 26659 32740 26668 32780
rect 26708 32740 27724 32780
rect 27764 32740 27773 32780
rect 4579 32656 4588 32696
rect 4628 32656 4972 32696
rect 5012 32656 6316 32696
rect 6356 32656 6365 32696
rect 8131 32656 8140 32696
rect 8180 32656 8716 32696
rect 8756 32656 8765 32696
rect 11491 32656 11500 32696
rect 11540 32656 11980 32696
rect 12020 32656 12029 32696
rect 15139 32656 15148 32696
rect 15188 32656 16588 32696
rect 16628 32656 16637 32696
rect 16867 32656 16876 32696
rect 16916 32656 17452 32696
rect 17492 32656 18028 32696
rect 18068 32656 18077 32696
rect 32131 32656 32140 32696
rect 32180 32656 35212 32696
rect 35252 32656 35261 32696
rect 38179 32656 38188 32696
rect 38228 32656 39916 32696
rect 39956 32656 39965 32696
rect 8803 32572 8812 32612
rect 8852 32572 12364 32612
rect 12404 32572 12413 32612
rect 25891 32572 25900 32612
rect 25940 32572 26668 32612
rect 26708 32572 26717 32612
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 14275 32488 14284 32528
rect 14324 32488 14860 32528
rect 14900 32488 14909 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 36643 32488 36652 32528
rect 36692 32488 37132 32528
rect 37172 32488 37181 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 13603 32444 13661 32445
rect 6115 32404 6124 32444
rect 6164 32404 13132 32444
rect 13172 32404 13181 32444
rect 13603 32404 13612 32444
rect 13652 32404 13804 32444
rect 13844 32404 17932 32444
rect 17972 32404 18412 32444
rect 18452 32404 18461 32444
rect 13603 32403 13661 32404
rect 4867 32360 4925 32361
rect 2467 32320 2476 32360
rect 2516 32320 3724 32360
rect 3764 32320 3773 32360
rect 4675 32320 4684 32360
rect 4724 32320 4876 32360
rect 4916 32320 4925 32360
rect 13699 32320 13708 32360
rect 13748 32320 14764 32360
rect 14804 32320 14813 32360
rect 30307 32320 30316 32360
rect 30356 32320 30700 32360
rect 30740 32320 31756 32360
rect 31796 32320 32236 32360
rect 32276 32320 32285 32360
rect 35779 32320 35788 32360
rect 35828 32320 36172 32360
rect 36212 32320 36221 32360
rect 4867 32319 4925 32320
rect 7363 32236 7372 32276
rect 7412 32236 8236 32276
rect 8276 32236 8285 32276
rect 12355 32236 12364 32276
rect 12404 32236 16204 32276
rect 16244 32236 16253 32276
rect 25996 32236 26572 32276
rect 26612 32236 27244 32276
rect 27284 32236 27293 32276
rect 31459 32236 31468 32276
rect 31508 32236 35020 32276
rect 35060 32236 35069 32276
rect 36547 32236 36556 32276
rect 36596 32236 37228 32276
rect 37268 32236 37277 32276
rect 25996 32192 26036 32236
rect 2371 32152 2380 32192
rect 2420 32152 2860 32192
rect 2900 32152 2909 32192
rect 7171 32152 7180 32192
rect 7220 32152 7948 32192
rect 7988 32152 7997 32192
rect 8131 32152 8140 32192
rect 8180 32152 9580 32192
rect 9620 32152 9629 32192
rect 12739 32152 12748 32192
rect 12788 32152 12940 32192
rect 12980 32152 12989 32192
rect 13795 32152 13804 32192
rect 13844 32152 14476 32192
rect 14516 32152 14525 32192
rect 14659 32152 14668 32192
rect 14708 32152 16012 32192
rect 16052 32152 16300 32192
rect 16340 32152 16349 32192
rect 17443 32152 17452 32192
rect 17492 32152 17836 32192
rect 17876 32152 17885 32192
rect 25315 32152 25324 32192
rect 25364 32152 25996 32192
rect 26036 32152 26045 32192
rect 26179 32152 26188 32192
rect 26228 32152 27532 32192
rect 27572 32152 27581 32192
rect 30787 32152 30796 32192
rect 30836 32152 32812 32192
rect 32852 32152 32861 32192
rect 33475 32152 33484 32192
rect 33524 32152 34156 32192
rect 34196 32152 34540 32192
rect 34580 32152 34589 32192
rect 35203 32152 35212 32192
rect 35252 32152 35692 32192
rect 35732 32152 36940 32192
rect 36980 32152 36989 32192
rect 13123 32068 13132 32108
rect 13172 32068 14284 32108
rect 14324 32068 14333 32108
rect 36451 32068 36460 32108
rect 36500 32068 39724 32108
rect 39764 32068 39773 32108
rect 5731 31984 5740 32024
rect 5780 31984 7948 32024
rect 7988 31984 7997 32024
rect 9379 31984 9388 32024
rect 9428 31984 10348 32024
rect 10388 31984 10397 32024
rect 26179 31984 26188 32024
rect 26228 31984 27052 32024
rect 27092 31984 27101 32024
rect 36067 31984 36076 32024
rect 36116 31984 38188 32024
rect 38228 31984 38237 32024
rect 31747 31940 31805 31941
rect 3523 31900 3532 31940
rect 3572 31900 3916 31940
rect 3956 31900 4492 31940
rect 4532 31900 4541 31940
rect 10051 31900 10060 31940
rect 10100 31900 10444 31940
rect 10484 31900 10493 31940
rect 12259 31900 12268 31940
rect 12308 31900 12940 31940
rect 12980 31900 12989 31940
rect 16099 31900 16108 31940
rect 16148 31900 16300 31940
rect 16340 31900 16349 31940
rect 28675 31900 28684 31940
rect 28724 31900 29356 31940
rect 29396 31900 29405 31940
rect 31662 31900 31756 31940
rect 31796 31900 31805 31940
rect 36163 31900 36172 31940
rect 36212 31900 37036 31940
rect 37076 31900 37085 31940
rect 31747 31899 31805 31900
rect 14947 31816 14956 31856
rect 14996 31816 17452 31856
rect 17492 31816 17501 31856
rect 38755 31816 38764 31856
rect 38804 31816 39244 31856
rect 39284 31816 39293 31856
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 12739 31732 12748 31772
rect 12788 31732 15436 31772
rect 15476 31732 16300 31772
rect 16340 31732 16349 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 25891 31732 25900 31772
rect 25940 31732 26476 31772
rect 26516 31732 26525 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31628 80 31708
rect 3907 31648 3916 31688
rect 3956 31648 4780 31688
rect 4820 31648 4829 31688
rect 13123 31648 13132 31688
rect 13172 31648 13181 31688
rect 13132 31604 13172 31648
rect 13987 31604 14045 31605
rect 2755 31564 2764 31604
rect 2804 31564 3820 31604
rect 3860 31564 3869 31604
rect 4867 31564 4876 31604
rect 4916 31564 6316 31604
rect 6356 31564 6365 31604
rect 9955 31564 9964 31604
rect 10004 31564 11308 31604
rect 11348 31564 11357 31604
rect 11587 31564 11596 31604
rect 11636 31564 12364 31604
rect 12404 31564 13172 31604
rect 13902 31564 13996 31604
rect 14036 31564 14045 31604
rect 15139 31564 15148 31604
rect 15188 31564 15628 31604
rect 15668 31564 15677 31604
rect 25219 31564 25228 31604
rect 25268 31564 26380 31604
rect 26420 31564 26429 31604
rect 33187 31564 33196 31604
rect 33236 31564 33388 31604
rect 33428 31564 36172 31604
rect 36212 31564 36221 31604
rect 13987 31563 14045 31564
rect 4387 31480 4396 31520
rect 4436 31480 6508 31520
rect 6548 31480 6557 31520
rect 6883 31480 6892 31520
rect 6932 31480 9484 31520
rect 9524 31480 9533 31520
rect 9763 31480 9772 31520
rect 9812 31480 10828 31520
rect 10868 31480 10877 31520
rect 11203 31480 11212 31520
rect 11252 31480 12556 31520
rect 12596 31480 12605 31520
rect 13315 31480 13324 31520
rect 13364 31480 15340 31520
rect 15380 31480 15389 31520
rect 20707 31480 20716 31520
rect 20756 31480 21100 31520
rect 21140 31480 22060 31520
rect 22100 31480 22540 31520
rect 22580 31480 22732 31520
rect 22772 31480 22781 31520
rect 23203 31480 23212 31520
rect 23252 31480 23884 31520
rect 23924 31480 23933 31520
rect 25027 31480 25036 31520
rect 25076 31480 26956 31520
rect 26996 31480 27005 31520
rect 30115 31480 30124 31520
rect 30164 31480 30173 31520
rect 30595 31480 30604 31520
rect 30644 31480 32236 31520
rect 32276 31480 32285 31520
rect 32611 31480 32620 31520
rect 32660 31480 32908 31520
rect 32948 31480 34156 31520
rect 34196 31480 34205 31520
rect 30124 31436 30164 31480
rect 4003 31396 4012 31436
rect 4052 31396 4300 31436
rect 4340 31396 5452 31436
rect 5492 31396 5501 31436
rect 12451 31396 12460 31436
rect 12500 31396 13516 31436
rect 13556 31396 13565 31436
rect 14179 31396 14188 31436
rect 14228 31396 14420 31436
rect 14755 31396 14764 31436
rect 14804 31396 16012 31436
rect 16052 31396 16588 31436
rect 16628 31396 16637 31436
rect 22915 31396 22924 31436
rect 22964 31396 23788 31436
rect 23828 31396 24940 31436
rect 24980 31396 24989 31436
rect 29635 31396 29644 31436
rect 29684 31396 30028 31436
rect 30068 31396 30077 31436
rect 30124 31396 32044 31436
rect 32084 31396 32093 31436
rect 12835 31352 12893 31353
rect 12750 31312 12844 31352
rect 12884 31312 12893 31352
rect 13219 31312 13228 31352
rect 13268 31312 14284 31352
rect 14324 31312 14333 31352
rect 12835 31311 12893 31312
rect 14380 31268 14420 31396
rect 14659 31312 14668 31352
rect 14708 31312 17164 31352
rect 17204 31312 17213 31352
rect 27331 31312 27340 31352
rect 27380 31312 28108 31352
rect 28148 31312 28157 31352
rect 29923 31312 29932 31352
rect 29972 31312 30700 31352
rect 30740 31312 30749 31352
rect 35971 31312 35980 31352
rect 36020 31312 38572 31352
rect 38612 31312 38621 31352
rect 5923 31228 5932 31268
rect 5972 31228 8044 31268
rect 8084 31228 8093 31268
rect 12067 31228 12076 31268
rect 12116 31228 13612 31268
rect 13652 31228 14764 31268
rect 14804 31228 15340 31268
rect 15380 31228 15389 31268
rect 15907 31228 15916 31268
rect 15956 31228 16300 31268
rect 16340 31228 16349 31268
rect 34723 31228 34732 31268
rect 34772 31228 35596 31268
rect 35636 31228 35645 31268
rect 6115 31144 6124 31184
rect 6164 31144 7660 31184
rect 7700 31144 7709 31184
rect 11011 31144 11020 31184
rect 11060 31144 12844 31184
rect 12884 31144 12893 31184
rect 22339 31144 22348 31184
rect 22388 31144 23020 31184
rect 23060 31144 23069 31184
rect 39331 31144 39340 31184
rect 39380 31144 40588 31184
rect 40628 31144 40780 31184
rect 40820 31144 40829 31184
rect 7555 31060 7564 31100
rect 7604 31060 7756 31100
rect 7796 31060 12652 31100
rect 12692 31060 13516 31100
rect 13556 31060 13565 31100
rect 13603 31016 13661 31017
rect 13987 31016 14045 31017
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 13518 30976 13612 31016
rect 13652 30976 13661 31016
rect 13902 30976 13996 31016
rect 14036 30976 14045 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 36355 30976 36364 31016
rect 36404 30976 36556 31016
rect 36596 30976 36605 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 13603 30975 13661 30976
rect 13987 30975 14045 30976
rect 12739 30892 12748 30932
rect 12788 30892 15532 30932
rect 15572 30892 15581 30932
rect 37228 30892 39436 30932
rect 39476 30892 39485 30932
rect 0 30788 80 30868
rect 37228 30848 37268 30892
rect 4588 30808 4972 30848
rect 5012 30808 5021 30848
rect 12835 30808 12844 30848
rect 12884 30808 13900 30848
rect 13940 30808 13949 30848
rect 15427 30808 15436 30848
rect 15476 30808 15820 30848
rect 15860 30808 16492 30848
rect 16532 30808 17836 30848
rect 17876 30808 17885 30848
rect 34051 30808 34060 30848
rect 34100 30808 34540 30848
rect 34580 30808 35020 30848
rect 35060 30808 36556 30848
rect 36596 30808 37228 30848
rect 37268 30808 37277 30848
rect 38371 30808 38380 30848
rect 38420 30808 38956 30848
rect 38996 30808 39005 30848
rect 4588 30680 4628 30808
rect 11320 30724 14572 30764
rect 14612 30724 14621 30764
rect 16963 30724 16972 30764
rect 17012 30724 18892 30764
rect 18932 30724 18941 30764
rect 21379 30724 21388 30764
rect 21428 30724 21868 30764
rect 21908 30724 21917 30764
rect 26755 30724 26764 30764
rect 26804 30724 27244 30764
rect 27284 30724 27293 30764
rect 32995 30724 33004 30764
rect 33044 30724 36076 30764
rect 36116 30724 36125 30764
rect 36643 30724 36652 30764
rect 36692 30724 38284 30764
rect 38324 30724 38333 30764
rect 11320 30680 11360 30724
rect 4579 30640 4588 30680
rect 4628 30640 4637 30680
rect 4963 30640 4972 30680
rect 5012 30640 5356 30680
rect 5396 30640 5405 30680
rect 5539 30640 5548 30680
rect 5588 30640 6316 30680
rect 6356 30640 6365 30680
rect 7555 30640 7564 30680
rect 7604 30640 8044 30680
rect 8084 30640 8093 30680
rect 10723 30640 10732 30680
rect 10772 30640 11360 30680
rect 13123 30640 13132 30680
rect 13172 30640 14188 30680
rect 14228 30640 14237 30680
rect 19171 30640 19180 30680
rect 19220 30640 19756 30680
rect 19796 30640 23980 30680
rect 24020 30640 24029 30680
rect 26467 30640 26476 30680
rect 26516 30640 27052 30680
rect 27092 30640 27101 30680
rect 31747 30640 31756 30680
rect 31796 30640 33196 30680
rect 33236 30640 33245 30680
rect 33859 30640 33868 30680
rect 33908 30640 35788 30680
rect 35828 30640 35837 30680
rect 36739 30640 36748 30680
rect 36788 30640 39148 30680
rect 39188 30640 39197 30680
rect 12835 30596 12893 30597
rect 6019 30556 6028 30596
rect 6068 30556 6508 30596
rect 6548 30556 6557 30596
rect 12750 30556 12844 30596
rect 12884 30556 12893 30596
rect 15523 30556 15532 30596
rect 15572 30556 16492 30596
rect 16532 30556 17548 30596
rect 17588 30556 17597 30596
rect 19363 30556 19372 30596
rect 19412 30556 19948 30596
rect 19988 30556 19997 30596
rect 32323 30556 32332 30596
rect 32372 30556 32812 30596
rect 32852 30556 33772 30596
rect 33812 30556 34732 30596
rect 34772 30556 34781 30596
rect 38563 30556 38572 30596
rect 38612 30556 39628 30596
rect 39668 30556 39677 30596
rect 12835 30555 12893 30556
rect 9955 30472 9964 30512
rect 10004 30472 11212 30512
rect 11252 30472 11261 30512
rect 15043 30472 15052 30512
rect 15092 30472 15436 30512
rect 15476 30472 15485 30512
rect 24931 30472 24940 30512
rect 24980 30472 25132 30512
rect 25172 30472 26668 30512
rect 26708 30472 27532 30512
rect 27572 30472 28204 30512
rect 28244 30472 28253 30512
rect 33667 30472 33676 30512
rect 33716 30472 34156 30512
rect 34196 30472 35212 30512
rect 35252 30472 35261 30512
rect 36163 30472 36172 30512
rect 36212 30472 36556 30512
rect 36596 30472 36605 30512
rect 13891 30428 13949 30429
rect 1315 30388 1324 30428
rect 1364 30388 3052 30428
rect 3092 30388 3101 30428
rect 13795 30388 13804 30428
rect 13844 30388 13900 30428
rect 13940 30388 13949 30428
rect 14659 30388 14668 30428
rect 14708 30388 15820 30428
rect 15860 30388 15869 30428
rect 30403 30388 30412 30428
rect 30452 30388 30892 30428
rect 30932 30388 30941 30428
rect 31939 30388 31948 30428
rect 31988 30388 32524 30428
rect 32564 30388 32908 30428
rect 32948 30388 32957 30428
rect 38083 30388 38092 30428
rect 38132 30388 39820 30428
rect 39860 30388 39869 30428
rect 43363 30388 43372 30428
rect 43412 30388 45772 30428
rect 45812 30388 45821 30428
rect 13891 30387 13949 30388
rect 30892 30344 30932 30388
rect 30892 30304 34636 30344
rect 34676 30304 34685 30344
rect 37027 30304 37036 30344
rect 37076 30304 38956 30344
rect 38996 30304 39005 30344
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 3715 30220 3724 30260
rect 3764 30220 4876 30260
rect 4916 30220 4925 30260
rect 5059 30220 5068 30260
rect 5108 30220 5356 30260
rect 5396 30220 5836 30260
rect 5876 30220 5885 30260
rect 12643 30220 12652 30260
rect 12692 30220 13420 30260
rect 13460 30220 15916 30260
rect 15956 30220 15965 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 22819 30220 22828 30260
rect 22868 30220 23788 30260
rect 23828 30220 25708 30260
rect 25748 30220 25757 30260
rect 26563 30220 26572 30260
rect 26612 30220 29836 30260
rect 29876 30220 30028 30260
rect 30068 30220 30077 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 41731 30220 41740 30260
rect 41780 30220 42700 30260
rect 42740 30220 45292 30260
rect 45332 30220 45341 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 5068 30176 5108 30220
rect 27340 30176 27380 30220
rect 3811 30136 3820 30176
rect 3860 30136 4396 30176
rect 4436 30136 4684 30176
rect 4724 30136 5108 30176
rect 12931 30136 12940 30176
rect 12980 30136 13804 30176
rect 13844 30136 13853 30176
rect 27331 30136 27340 30176
rect 27380 30136 27389 30176
rect 37123 30136 37132 30176
rect 37172 30136 37181 30176
rect 43747 30136 43756 30176
rect 43796 30136 44812 30176
rect 44852 30136 44861 30176
rect 3715 30052 3724 30092
rect 3764 30052 4588 30092
rect 4628 30052 5260 30092
rect 5300 30052 5309 30092
rect 6595 30052 6604 30092
rect 6644 30052 8044 30092
rect 8084 30052 8716 30092
rect 8756 30052 10828 30092
rect 10868 30052 11360 30092
rect 0 29948 80 30028
rect 11320 29924 11360 30052
rect 32227 29968 32236 30008
rect 32276 29968 33388 30008
rect 33428 29968 33437 30008
rect 37132 29924 37172 30136
rect 46243 29968 46252 30008
rect 46292 29968 46636 30008
rect 46676 29968 46685 30008
rect 4195 29884 4204 29924
rect 4244 29884 5164 29924
rect 5204 29884 7756 29924
rect 7796 29884 8236 29924
rect 8276 29884 10828 29924
rect 10868 29884 10877 29924
rect 11320 29884 12172 29924
rect 12212 29884 12221 29924
rect 31075 29884 31084 29924
rect 31124 29884 31468 29924
rect 31508 29884 35692 29924
rect 35732 29884 35741 29924
rect 36739 29884 36748 29924
rect 36788 29884 37420 29924
rect 37460 29884 37469 29924
rect 2659 29800 2668 29840
rect 2708 29800 4588 29840
rect 4628 29800 4637 29840
rect 8323 29800 8332 29840
rect 8372 29800 8524 29840
rect 8564 29800 8573 29840
rect 8803 29800 8812 29840
rect 8852 29800 14380 29840
rect 14420 29800 14429 29840
rect 14563 29800 14572 29840
rect 14612 29800 15244 29840
rect 15284 29800 15293 29840
rect 21763 29800 21772 29840
rect 21812 29800 22636 29840
rect 22676 29800 22685 29840
rect 25699 29800 25708 29840
rect 25748 29800 27436 29840
rect 27476 29800 27485 29840
rect 32995 29800 33004 29840
rect 33044 29800 33964 29840
rect 34004 29800 34013 29840
rect 37027 29800 37036 29840
rect 37076 29800 37324 29840
rect 37364 29800 37373 29840
rect 40291 29800 40300 29840
rect 40340 29800 40684 29840
rect 40724 29800 40733 29840
rect 41347 29800 41356 29840
rect 41396 29800 43276 29840
rect 43316 29800 43325 29840
rect 3715 29716 3724 29756
rect 3764 29716 4012 29756
rect 4052 29716 4300 29756
rect 4340 29716 4349 29756
rect 8611 29716 8620 29756
rect 8660 29716 9676 29756
rect 9716 29716 9725 29756
rect 23875 29716 23884 29756
rect 23924 29716 25324 29756
rect 25364 29716 25373 29756
rect 32803 29716 32812 29756
rect 32852 29716 33100 29756
rect 33140 29716 33149 29756
rect 37219 29716 37228 29756
rect 37268 29716 40012 29756
rect 40052 29716 40061 29756
rect 42211 29716 42220 29756
rect 42260 29716 42700 29756
rect 42740 29716 43756 29756
rect 43796 29716 43805 29756
rect 17635 29632 17644 29672
rect 17684 29632 19180 29672
rect 19220 29632 20524 29672
rect 20564 29632 20573 29672
rect 24163 29632 24172 29672
rect 24212 29632 24940 29672
rect 24980 29632 25900 29672
rect 25940 29632 25949 29672
rect 26371 29632 26380 29672
rect 26420 29632 27724 29672
rect 27764 29632 27773 29672
rect 29251 29632 29260 29672
rect 29300 29632 32044 29672
rect 32084 29632 32093 29672
rect 35107 29632 35116 29672
rect 35156 29632 36940 29672
rect 36980 29632 36989 29672
rect 40387 29632 40396 29672
rect 40436 29632 40876 29672
rect 40916 29632 40925 29672
rect 41251 29632 41260 29672
rect 41300 29632 42604 29672
rect 42644 29632 42653 29672
rect 26659 29548 26668 29588
rect 26708 29548 30412 29588
rect 30452 29548 30461 29588
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 31843 29464 31852 29504
rect 31892 29464 32428 29504
rect 32468 29464 32716 29504
rect 32756 29464 32765 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 15811 29380 15820 29420
rect 15860 29380 17644 29420
rect 17684 29380 17693 29420
rect 23299 29380 23308 29420
rect 23348 29380 25996 29420
rect 26036 29380 29000 29420
rect 35683 29380 35692 29420
rect 35732 29380 36364 29420
rect 36404 29380 37364 29420
rect 7459 29296 7468 29336
rect 7508 29296 11788 29336
rect 11828 29296 11837 29336
rect 14851 29296 14860 29336
rect 14900 29296 18700 29336
rect 18740 29296 18749 29336
rect 19747 29296 19756 29336
rect 19796 29296 20044 29336
rect 20084 29296 20093 29336
rect 22531 29296 22540 29336
rect 22580 29296 23116 29336
rect 23156 29296 23165 29336
rect 25507 29296 25516 29336
rect 25556 29296 26572 29336
rect 26612 29296 26621 29336
rect 1315 29212 1324 29252
rect 1364 29212 3916 29252
rect 3956 29212 3965 29252
rect 4867 29212 4876 29252
rect 4916 29212 5644 29252
rect 5684 29212 5693 29252
rect 14563 29212 14572 29252
rect 14612 29212 16972 29252
rect 17012 29212 17021 29252
rect 22627 29212 22636 29252
rect 22676 29212 23500 29252
rect 23540 29212 23549 29252
rect 25132 29212 26860 29252
rect 26900 29212 26909 29252
rect 0 29108 80 29188
rect 25132 29168 25172 29212
rect 2563 29128 2572 29168
rect 2612 29128 3532 29168
rect 3572 29128 6124 29168
rect 6164 29128 6173 29168
rect 7555 29128 7564 29168
rect 7604 29128 13708 29168
rect 13748 29128 13757 29168
rect 16483 29128 16492 29168
rect 16532 29128 16541 29168
rect 16771 29128 16780 29168
rect 16820 29128 19084 29168
rect 19124 29128 19133 29168
rect 21475 29128 21484 29168
rect 21524 29128 22540 29168
rect 22580 29128 23212 29168
rect 23252 29128 23261 29168
rect 25123 29128 25132 29168
rect 25172 29128 25181 29168
rect 25795 29128 25804 29168
rect 25844 29128 26764 29168
rect 26804 29128 27436 29168
rect 27476 29128 27485 29168
rect 27619 29128 27628 29168
rect 27668 29128 28108 29168
rect 28148 29128 28157 29168
rect 16492 29084 16532 29128
rect 23212 29084 23252 29128
rect 28960 29084 29000 29380
rect 37324 29336 37364 29380
rect 30979 29296 30988 29336
rect 31028 29296 31564 29336
rect 31604 29296 34444 29336
rect 34484 29296 34493 29336
rect 35692 29296 36748 29336
rect 36788 29296 36797 29336
rect 37315 29296 37324 29336
rect 37364 29296 37373 29336
rect 43267 29296 43276 29336
rect 43316 29296 43756 29336
rect 43796 29296 43805 29336
rect 44227 29296 44236 29336
rect 44276 29296 47884 29336
rect 47924 29296 48460 29336
rect 48500 29296 48509 29336
rect 35692 29252 35732 29296
rect 32740 29212 35732 29252
rect 35779 29212 35788 29252
rect 35828 29212 37420 29252
rect 37460 29212 37469 29252
rect 40675 29212 40684 29252
rect 40724 29212 42316 29252
rect 42356 29212 42365 29252
rect 32740 29168 32780 29212
rect 31075 29128 31084 29168
rect 31124 29128 32780 29168
rect 33091 29128 33100 29168
rect 33140 29128 35116 29168
rect 35156 29128 35692 29168
rect 35732 29128 35741 29168
rect 37507 29128 37516 29168
rect 37556 29128 37900 29168
rect 37940 29128 37949 29168
rect 45283 29128 45292 29168
rect 45332 29128 47116 29168
rect 47156 29128 47165 29168
rect 5644 29044 7276 29084
rect 7316 29044 7325 29084
rect 11692 29044 14476 29084
rect 14516 29044 14525 29084
rect 16492 29044 18796 29084
rect 18836 29044 18845 29084
rect 19372 29044 20812 29084
rect 20852 29044 20861 29084
rect 23212 29044 25228 29084
rect 25268 29044 25277 29084
rect 27331 29044 27340 29084
rect 27380 29044 27820 29084
rect 27860 29044 27869 29084
rect 28960 29044 29164 29084
rect 29204 29044 29213 29084
rect 30403 29044 30412 29084
rect 30452 29044 31660 29084
rect 31700 29044 33004 29084
rect 33044 29044 33053 29084
rect 42115 29044 42124 29084
rect 42164 29044 42796 29084
rect 42836 29044 43084 29084
rect 43124 29044 43133 29084
rect 1123 28960 1132 29000
rect 1172 28960 1708 29000
rect 1748 28960 1757 29000
rect 5644 28916 5684 29044
rect 11692 29000 11732 29044
rect 19372 29000 19412 29044
rect 11652 28960 11692 29000
rect 11732 28960 11741 29000
rect 19332 28960 19372 29000
rect 19412 28960 19421 29000
rect 30691 28960 30700 29000
rect 30740 28960 30749 29000
rect 35299 28960 35308 29000
rect 35348 28960 35357 29000
rect 38083 28960 38092 29000
rect 38132 28960 38141 29000
rect 39427 28960 39436 29000
rect 39476 28960 39485 29000
rect 42499 28960 42508 29000
rect 42548 28960 42557 29000
rect 30700 28916 30740 28960
rect 5644 28876 5932 28916
rect 5972 28876 5981 28916
rect 10339 28876 10348 28916
rect 10388 28876 11116 28916
rect 11156 28876 11500 28916
rect 11540 28876 11549 28916
rect 13603 28876 13612 28916
rect 13652 28876 14668 28916
rect 14708 28876 14717 28916
rect 19459 28876 19468 28916
rect 19508 28876 20140 28916
rect 20180 28876 22252 28916
rect 22292 28876 22301 28916
rect 29923 28876 29932 28916
rect 29972 28876 30740 28916
rect 35308 28916 35348 28960
rect 38092 28916 38132 28960
rect 39436 28916 39476 28960
rect 42508 28916 42548 28960
rect 35308 28876 37036 28916
rect 37076 28876 37085 28916
rect 38092 28876 39476 28916
rect 40867 28876 40876 28916
rect 40916 28876 42548 28916
rect 14179 28792 14188 28832
rect 14228 28792 16876 28832
rect 16916 28792 21868 28832
rect 21908 28792 21917 28832
rect 41443 28792 41452 28832
rect 41492 28792 42700 28832
rect 42740 28792 42988 28832
rect 43028 28792 43037 28832
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 2755 28624 2764 28664
rect 2804 28624 6508 28664
rect 6548 28624 6557 28664
rect 15331 28624 15340 28664
rect 15380 28624 19468 28664
rect 19508 28624 19517 28664
rect 30787 28624 30796 28664
rect 30836 28624 32428 28664
rect 32468 28624 32477 28664
rect 15235 28540 15244 28580
rect 15284 28540 17452 28580
rect 17492 28540 17501 28580
rect 18595 28540 18604 28580
rect 18644 28540 18796 28580
rect 18836 28540 18845 28580
rect 28291 28540 28300 28580
rect 28340 28540 29740 28580
rect 29780 28540 30604 28580
rect 30644 28540 30653 28580
rect 4867 28456 4876 28496
rect 4916 28456 5452 28496
rect 5492 28456 5501 28496
rect 28387 28456 28396 28496
rect 28436 28456 31564 28496
rect 31604 28456 32236 28496
rect 32276 28456 32285 28496
rect 37780 28456 43756 28496
rect 43796 28456 45196 28496
rect 45236 28456 47404 28496
rect 47444 28456 47453 28496
rect 48259 28456 48268 28496
rect 48308 28456 49228 28496
rect 49268 28456 49277 28496
rect 37780 28412 37820 28456
rect 47404 28412 47444 28456
rect 5827 28372 5836 28412
rect 5876 28372 7852 28412
rect 7892 28372 7901 28412
rect 19075 28372 19084 28412
rect 19124 28372 19756 28412
rect 19796 28372 19805 28412
rect 30211 28372 30220 28412
rect 30260 28372 31276 28412
rect 31316 28372 31325 28412
rect 34051 28372 34060 28412
rect 34100 28372 35692 28412
rect 35732 28372 35741 28412
rect 35971 28372 35980 28412
rect 36020 28372 37820 28412
rect 42979 28372 42988 28412
rect 43028 28372 43468 28412
rect 43508 28372 44140 28412
rect 44180 28372 44332 28412
rect 44372 28372 44381 28412
rect 47404 28372 48940 28412
rect 48980 28372 48989 28412
rect 0 28268 80 28348
rect 3811 28288 3820 28328
rect 3860 28288 6700 28328
rect 6740 28288 6749 28328
rect 7555 28288 7564 28328
rect 7604 28288 8428 28328
rect 8468 28288 15820 28328
rect 15860 28288 16108 28328
rect 16148 28288 16157 28328
rect 18979 28288 18988 28328
rect 19028 28288 19564 28328
rect 19604 28288 19613 28328
rect 20515 28288 20524 28328
rect 20564 28288 21100 28328
rect 21140 28288 21149 28328
rect 23779 28288 23788 28328
rect 23828 28288 25708 28328
rect 25748 28288 28684 28328
rect 28724 28288 29068 28328
rect 29108 28288 29452 28328
rect 29492 28288 29501 28328
rect 32035 28288 32044 28328
rect 32084 28288 32812 28328
rect 32852 28288 33772 28328
rect 33812 28288 33821 28328
rect 35395 28288 35404 28328
rect 35444 28288 37708 28328
rect 37748 28288 37757 28328
rect 40579 28288 40588 28328
rect 40628 28288 41452 28328
rect 41492 28288 41501 28328
rect 43171 28288 43180 28328
rect 43220 28288 43852 28328
rect 43892 28288 43901 28328
rect 44035 28288 44044 28328
rect 44084 28288 46540 28328
rect 46580 28288 47116 28328
rect 47156 28288 47165 28328
rect 47683 28288 47692 28328
rect 47732 28288 48748 28328
rect 48788 28288 48797 28328
rect 50275 28288 50284 28328
rect 50324 28288 50572 28328
rect 50612 28288 50621 28328
rect 12451 28204 12460 28244
rect 12500 28204 12940 28244
rect 12980 28204 12989 28244
rect 32227 28204 32236 28244
rect 32276 28204 33196 28244
rect 33236 28204 33964 28244
rect 34004 28204 34013 28244
rect 39235 28204 39244 28244
rect 39284 28204 42316 28244
rect 42356 28204 42508 28244
rect 42548 28204 42557 28244
rect 43555 28204 43564 28244
rect 43604 28204 45868 28244
rect 45908 28204 45917 28244
rect 6595 28120 6604 28160
rect 6644 28120 8140 28160
rect 8180 28120 9676 28160
rect 9716 28120 9725 28160
rect 31651 28120 31660 28160
rect 31700 28120 32620 28160
rect 32660 28120 32669 28160
rect 41635 28120 41644 28160
rect 41684 28120 42124 28160
rect 42164 28120 42173 28160
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 5251 27868 5260 27908
rect 5300 27868 5740 27908
rect 5780 27868 5789 27908
rect 10051 27868 10060 27908
rect 10100 27868 12556 27908
rect 12596 27868 12605 27908
rect 4099 27784 4108 27824
rect 4148 27784 4157 27824
rect 14755 27784 14764 27824
rect 14804 27784 14813 27824
rect 17251 27784 17260 27824
rect 17300 27784 17740 27824
rect 17780 27784 19276 27824
rect 19316 27784 19468 27824
rect 19508 27784 19517 27824
rect 32899 27784 32908 27824
rect 32948 27784 34540 27824
rect 34580 27784 34589 27824
rect 45091 27784 45100 27824
rect 45140 27784 49036 27824
rect 49076 27784 49085 27824
rect 4108 27740 4148 27784
rect 14764 27740 14804 27784
rect 2947 27700 2956 27740
rect 2996 27700 5068 27740
rect 5108 27700 5117 27740
rect 5539 27700 5548 27740
rect 5588 27700 7756 27740
rect 7796 27700 7805 27740
rect 10531 27700 10540 27740
rect 10580 27700 10924 27740
rect 10964 27700 11596 27740
rect 11636 27700 11645 27740
rect 12739 27700 12748 27740
rect 12788 27700 14804 27740
rect 16003 27700 16012 27740
rect 16052 27700 17452 27740
rect 17492 27700 17501 27740
rect 19939 27700 19948 27740
rect 19988 27700 20716 27740
rect 20756 27700 20765 27740
rect 23779 27700 23788 27740
rect 23828 27700 25612 27740
rect 25652 27700 27052 27740
rect 27092 27700 27101 27740
rect 29827 27700 29836 27740
rect 29876 27700 31276 27740
rect 31316 27700 31468 27740
rect 31508 27700 31517 27740
rect 35971 27700 35980 27740
rect 36020 27700 38380 27740
rect 38420 27700 38429 27740
rect 40483 27700 40492 27740
rect 40532 27700 42220 27740
rect 42260 27700 42269 27740
rect 47491 27700 47500 27740
rect 47540 27700 50284 27740
rect 50324 27700 50333 27740
rect 2467 27616 2476 27656
rect 2516 27616 2572 27656
rect 2612 27616 2860 27656
rect 2900 27616 2909 27656
rect 6019 27616 6028 27656
rect 6068 27616 6077 27656
rect 7075 27616 7084 27656
rect 7124 27616 8140 27656
rect 8180 27616 8189 27656
rect 8419 27616 8428 27656
rect 8468 27616 11692 27656
rect 11732 27616 12076 27656
rect 12116 27616 12125 27656
rect 13027 27616 13036 27656
rect 13076 27616 15916 27656
rect 15956 27616 19564 27656
rect 19604 27616 19613 27656
rect 22819 27616 22828 27656
rect 22868 27616 23884 27656
rect 23924 27616 23933 27656
rect 24739 27616 24748 27656
rect 24788 27616 25324 27656
rect 25364 27616 25900 27656
rect 25940 27616 25949 27656
rect 30019 27616 30028 27656
rect 30068 27616 30508 27656
rect 30548 27616 30557 27656
rect 30787 27616 30796 27656
rect 30836 27616 31180 27656
rect 31220 27616 31660 27656
rect 31700 27616 32044 27656
rect 32084 27616 32093 27656
rect 34435 27616 34444 27656
rect 34484 27616 35404 27656
rect 35444 27616 35453 27656
rect 40771 27616 40780 27656
rect 40820 27616 41548 27656
rect 41588 27616 41597 27656
rect 45379 27616 45388 27656
rect 45428 27616 46252 27656
rect 46292 27616 46301 27656
rect 6028 27572 6068 27616
rect 30796 27572 30836 27616
rect 3619 27532 3628 27572
rect 3668 27532 4780 27572
rect 4820 27532 6068 27572
rect 16579 27532 16588 27572
rect 16628 27532 17548 27572
rect 17588 27532 19084 27572
rect 19124 27532 19133 27572
rect 25219 27532 25228 27572
rect 25268 27532 27436 27572
rect 27476 27532 27485 27572
rect 28675 27532 28684 27572
rect 28724 27532 29260 27572
rect 29300 27532 29309 27572
rect 30211 27532 30220 27572
rect 30260 27532 30836 27572
rect 38755 27532 38764 27572
rect 38804 27532 39340 27572
rect 39380 27532 39389 27572
rect 0 27428 80 27508
rect 11395 27488 11453 27489
rect 7939 27448 7948 27488
rect 7988 27448 9292 27488
rect 9332 27448 9341 27488
rect 11203 27448 11212 27488
rect 11252 27448 11404 27488
rect 11444 27448 13324 27488
rect 13364 27448 13373 27488
rect 14467 27448 14476 27488
rect 14516 27448 15628 27488
rect 15668 27448 15677 27488
rect 17347 27448 17356 27488
rect 17396 27448 18796 27488
rect 18836 27448 18845 27488
rect 32227 27448 32236 27488
rect 32276 27448 32812 27488
rect 32852 27448 32861 27488
rect 33859 27448 33868 27488
rect 33908 27448 36556 27488
rect 36596 27448 36844 27488
rect 36884 27448 36893 27488
rect 38851 27448 38860 27488
rect 38900 27448 40972 27488
rect 41012 27448 41932 27488
rect 41972 27448 41981 27488
rect 11395 27447 11453 27448
rect 3907 27364 3916 27404
rect 3956 27364 4684 27404
rect 4724 27364 4733 27404
rect 6883 27364 6892 27404
rect 6932 27364 7276 27404
rect 7316 27364 8524 27404
rect 8564 27364 11116 27404
rect 11156 27364 11165 27404
rect 13987 27364 13996 27404
rect 14036 27364 14572 27404
rect 14612 27364 14621 27404
rect 14851 27364 14860 27404
rect 14900 27364 17836 27404
rect 17876 27364 17885 27404
rect 18499 27364 18508 27404
rect 18548 27364 18988 27404
rect 19028 27364 19037 27404
rect 29635 27364 29644 27404
rect 29684 27364 30508 27404
rect 30548 27364 30557 27404
rect 31363 27364 31372 27404
rect 31412 27364 33100 27404
rect 33140 27364 33292 27404
rect 33332 27364 33341 27404
rect 45283 27364 45292 27404
rect 45332 27364 46732 27404
rect 46772 27364 46781 27404
rect 18508 27320 18548 27364
rect 4483 27280 4492 27320
rect 4532 27280 6988 27320
rect 7028 27280 7852 27320
rect 7892 27280 9964 27320
rect 10004 27280 10013 27320
rect 15715 27280 15724 27320
rect 15764 27280 18548 27320
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 20035 27196 20044 27236
rect 20084 27196 27916 27236
rect 27956 27196 28492 27236
rect 28532 27196 28541 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 45571 27196 45580 27236
rect 45620 27196 46060 27236
rect 46100 27196 46109 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 6787 27112 6796 27152
rect 6836 27112 7564 27152
rect 7604 27112 7948 27152
rect 7988 27112 9484 27152
rect 9524 27112 9772 27152
rect 9812 27112 10540 27152
rect 10580 27112 10589 27152
rect 39619 27112 39628 27152
rect 39668 27112 43564 27152
rect 43604 27112 46100 27152
rect 30787 27068 30845 27069
rect 2755 27028 2764 27068
rect 2804 27028 3820 27068
rect 3860 27028 3869 27068
rect 8419 27028 8428 27068
rect 8468 27028 13804 27068
rect 13844 27028 13853 27068
rect 18115 27028 18124 27068
rect 18164 27028 18700 27068
rect 18740 27028 20524 27068
rect 20564 27028 21676 27068
rect 21716 27028 21725 27068
rect 25603 27028 25612 27068
rect 25652 27028 26380 27068
rect 26420 27028 26956 27068
rect 26996 27028 29836 27068
rect 29876 27028 30124 27068
rect 30164 27028 30173 27068
rect 30787 27028 30796 27068
rect 30836 27028 30988 27068
rect 31028 27028 31037 27068
rect 32131 27028 32140 27068
rect 32180 27028 33868 27068
rect 33908 27028 34252 27068
rect 34292 27028 35596 27068
rect 35636 27028 35645 27068
rect 39427 27028 39436 27068
rect 39476 27028 40300 27068
rect 40340 27028 40349 27068
rect 42979 27028 42988 27068
rect 43028 27028 44140 27068
rect 44180 27028 44189 27068
rect 30787 27027 30845 27028
rect 46060 26984 46100 27112
rect 46531 27028 46540 27068
rect 46580 27028 49132 27068
rect 49172 27028 50572 27068
rect 50612 27028 50621 27068
rect 51139 27028 51148 27068
rect 51188 27028 51724 27068
rect 51764 27028 51773 27068
rect 10243 26944 10252 26984
rect 10292 26944 10332 26984
rect 18595 26944 18604 26984
rect 18644 26944 19084 26984
rect 19124 26944 19133 26984
rect 19363 26944 19372 26984
rect 19412 26944 20620 26984
rect 20660 26944 20669 26984
rect 23395 26944 23404 26984
rect 23444 26944 23980 26984
rect 24020 26944 24029 26984
rect 28867 26944 28876 26984
rect 28916 26944 29108 26984
rect 42787 26944 42796 26984
rect 42836 26944 43468 26984
rect 43508 26944 43756 26984
rect 43796 26944 44716 26984
rect 44756 26944 45388 26984
rect 45428 26944 45964 26984
rect 46004 26944 46013 26984
rect 46060 26944 46732 26984
rect 46772 26944 48172 26984
rect 48212 26944 48221 26984
rect 10252 26900 10292 26944
rect 29068 26900 29108 26944
rect 1219 26860 1228 26900
rect 1268 26860 5836 26900
rect 5876 26860 5885 26900
rect 6403 26860 6412 26900
rect 6452 26860 7468 26900
rect 7508 26860 8524 26900
rect 8564 26860 8908 26900
rect 8948 26860 8957 26900
rect 9859 26860 9868 26900
rect 9908 26860 11360 26900
rect 26179 26860 26188 26900
rect 26228 26860 27052 26900
rect 27092 26860 27101 26900
rect 28099 26860 28108 26900
rect 28148 26860 28157 26900
rect 28771 26860 28780 26900
rect 28820 26860 28972 26900
rect 29012 26860 29021 26900
rect 29068 26860 30892 26900
rect 30932 26860 30941 26900
rect 34147 26860 34156 26900
rect 34196 26860 34732 26900
rect 34772 26860 34781 26900
rect 43363 26860 43372 26900
rect 43412 26860 45004 26900
rect 45044 26860 47020 26900
rect 47060 26860 47069 26900
rect 11320 26816 11360 26860
rect 17155 26816 17213 26817
rect 28108 26816 28148 26860
rect 3619 26776 3628 26816
rect 3668 26776 4396 26816
rect 4436 26776 4445 26816
rect 6499 26776 6508 26816
rect 6548 26776 7852 26816
rect 7892 26776 7901 26816
rect 9283 26776 9292 26816
rect 9332 26776 10252 26816
rect 10292 26776 10301 26816
rect 11320 26776 11692 26816
rect 11732 26776 11741 26816
rect 11875 26776 11884 26816
rect 11924 26776 14956 26816
rect 14996 26776 15005 26816
rect 15139 26776 15148 26816
rect 15188 26776 15436 26816
rect 15476 26776 16588 26816
rect 16628 26776 16637 26816
rect 16771 26776 16780 26816
rect 16820 26776 16972 26816
rect 17012 26776 17021 26816
rect 17070 26776 17164 26816
rect 17204 26776 17213 26816
rect 17827 26776 17836 26816
rect 17876 26776 19564 26816
rect 19604 26776 19613 26816
rect 25987 26776 25996 26816
rect 26036 26776 26572 26816
rect 26612 26776 26621 26816
rect 28003 26776 28012 26816
rect 28052 26776 28061 26816
rect 28108 26776 29548 26816
rect 29588 26776 29597 26816
rect 30691 26776 30700 26816
rect 30740 26776 31468 26816
rect 31508 26776 31517 26816
rect 34627 26776 34636 26816
rect 34676 26776 35308 26816
rect 35348 26776 35357 26816
rect 38179 26776 38188 26816
rect 38228 26776 41068 26816
rect 41108 26776 41117 26816
rect 42019 26776 42028 26816
rect 42068 26776 45868 26816
rect 45908 26776 45917 26816
rect 49699 26776 49708 26816
rect 49748 26776 51436 26816
rect 51476 26776 51485 26816
rect 13123 26732 13181 26733
rect 16972 26732 17012 26776
rect 17155 26775 17213 26776
rect 28012 26732 28052 26776
rect 1891 26692 1900 26732
rect 1940 26692 3820 26732
rect 3860 26692 3869 26732
rect 4675 26692 4684 26732
rect 4724 26692 4972 26732
rect 5012 26692 5452 26732
rect 5492 26692 5932 26732
rect 5972 26692 6700 26732
rect 6740 26692 6749 26732
rect 9667 26692 9676 26732
rect 9716 26692 11788 26732
rect 11828 26692 11837 26732
rect 13038 26692 13132 26732
rect 13172 26692 13181 26732
rect 14179 26692 14188 26732
rect 14228 26692 14237 26732
rect 14718 26692 14727 26732
rect 14767 26692 15532 26732
rect 15572 26692 15581 26732
rect 16972 26692 20044 26732
rect 20084 26692 20093 26732
rect 28012 26692 38476 26732
rect 38516 26692 38525 26732
rect 41251 26692 41260 26732
rect 41300 26692 43276 26732
rect 43316 26692 44236 26732
rect 44276 26692 44428 26732
rect 44468 26692 44477 26732
rect 45955 26692 45964 26732
rect 46004 26692 47980 26732
rect 48020 26692 48029 26732
rect 48931 26692 48940 26732
rect 48980 26692 49324 26732
rect 49364 26692 49373 26732
rect 0 26588 80 26668
rect 1699 26608 1708 26648
rect 1748 26608 3532 26648
rect 3572 26608 3581 26648
rect 4684 26564 4724 26692
rect 13123 26691 13181 26692
rect 13795 26648 13853 26649
rect 14188 26648 14228 26692
rect 14755 26648 14813 26649
rect 6499 26608 6508 26648
rect 6548 26608 8332 26648
rect 8372 26608 8381 26648
rect 10051 26608 10060 26648
rect 10100 26608 12460 26648
rect 12500 26608 12509 26648
rect 13027 26608 13036 26648
rect 13076 26608 13268 26648
rect 13710 26608 13804 26648
rect 13844 26608 13853 26648
rect 13987 26608 13996 26648
rect 14036 26608 14228 26648
rect 14275 26608 14284 26648
rect 14324 26608 14764 26648
rect 14804 26608 14813 26648
rect 18115 26608 18124 26648
rect 18164 26608 18796 26648
rect 18836 26608 18845 26648
rect 19171 26608 19180 26648
rect 19220 26608 20428 26648
rect 20468 26608 20477 26648
rect 25507 26608 25516 26648
rect 25556 26608 26572 26648
rect 26612 26608 26621 26648
rect 28579 26608 28588 26648
rect 28628 26608 29356 26648
rect 29396 26608 29405 26648
rect 32227 26608 32236 26648
rect 32276 26608 33100 26648
rect 33140 26608 34444 26648
rect 34484 26608 34493 26648
rect 37987 26608 37996 26648
rect 38036 26608 40204 26648
rect 40244 26608 40396 26648
rect 40436 26608 40445 26648
rect 43843 26608 43852 26648
rect 43892 26608 45004 26648
rect 45044 26608 45053 26648
rect 13228 26564 13268 26608
rect 13795 26607 13853 26608
rect 14755 26607 14813 26608
rect 3427 26524 3436 26564
rect 3476 26524 4724 26564
rect 6307 26524 6316 26564
rect 6356 26524 13132 26564
rect 13172 26524 13181 26564
rect 13228 26524 13900 26564
rect 13940 26524 14188 26564
rect 14228 26524 14668 26564
rect 14708 26524 14860 26564
rect 14900 26524 15436 26564
rect 15476 26524 15485 26564
rect 18883 26524 18892 26564
rect 18932 26524 19084 26564
rect 19124 26524 19133 26564
rect 25027 26524 25036 26564
rect 25076 26524 25900 26564
rect 25940 26524 25949 26564
rect 28099 26524 28108 26564
rect 28148 26524 28876 26564
rect 28916 26524 28925 26564
rect 29059 26524 29068 26564
rect 29108 26524 37324 26564
rect 37364 26524 37373 26564
rect 45571 26524 45580 26564
rect 45620 26524 51244 26564
rect 51284 26524 51293 26564
rect 30787 26480 30845 26481
rect 31267 26480 31325 26481
rect 31747 26480 31805 26481
rect 2275 26440 2284 26480
rect 2324 26440 2572 26480
rect 2612 26440 2956 26480
rect 2996 26440 3005 26480
rect 3139 26440 3148 26480
rect 3188 26440 3628 26480
rect 3668 26440 3677 26480
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 7075 26440 7084 26480
rect 7124 26440 7988 26480
rect 10435 26440 10444 26480
rect 10484 26440 11404 26480
rect 11444 26440 11453 26480
rect 13411 26440 13420 26480
rect 13460 26440 13996 26480
rect 14036 26440 14045 26480
rect 14371 26440 14380 26480
rect 14420 26440 15052 26480
rect 15092 26440 15101 26480
rect 15331 26440 15340 26480
rect 15380 26440 16108 26480
rect 16148 26440 16157 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 22147 26440 22156 26480
rect 22196 26440 28684 26480
rect 28724 26440 28733 26480
rect 30702 26440 30796 26480
rect 30836 26440 30845 26480
rect 31182 26440 31276 26480
rect 31316 26440 31325 26480
rect 31662 26440 31756 26480
rect 31796 26440 31805 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 35107 26440 35116 26480
rect 35156 26440 35500 26480
rect 35540 26440 35549 26480
rect 36931 26440 36940 26480
rect 36980 26440 38380 26480
rect 38420 26440 38429 26480
rect 39043 26440 39052 26480
rect 39092 26440 39436 26480
rect 39476 26440 39485 26480
rect 43939 26440 43948 26480
rect 43988 26440 44524 26480
rect 44564 26440 44573 26480
rect 44707 26440 44716 26480
rect 44756 26440 46828 26480
rect 46868 26440 47212 26480
rect 47252 26440 47261 26480
rect 47395 26440 47404 26480
rect 47444 26440 47884 26480
rect 47924 26440 47933 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 7948 26396 7988 26440
rect 30787 26439 30845 26440
rect 31267 26439 31325 26440
rect 31747 26439 31805 26440
rect 835 26356 844 26396
rect 884 26356 3340 26396
rect 3380 26356 5932 26396
rect 5972 26356 5981 26396
rect 7939 26356 7948 26396
rect 7988 26356 7997 26396
rect 8707 26356 8716 26396
rect 8756 26356 17164 26396
rect 17204 26356 17213 26396
rect 27523 26356 27532 26396
rect 27572 26356 41644 26396
rect 41684 26356 41693 26396
rect 44323 26356 44332 26396
rect 44372 26356 46444 26396
rect 46484 26356 47692 26396
rect 47732 26356 47741 26396
rect 14755 26312 14813 26313
rect 6595 26272 6604 26312
rect 6644 26272 7756 26312
rect 7796 26272 7805 26312
rect 14083 26272 14092 26312
rect 14132 26272 14612 26312
rect 13891 26144 13949 26145
rect 14572 26144 14612 26272
rect 14755 26272 14764 26312
rect 14804 26272 14898 26312
rect 14947 26272 14956 26312
rect 14996 26272 15340 26312
rect 15380 26272 15389 26312
rect 16099 26272 16108 26312
rect 16148 26272 17068 26312
rect 17108 26272 17117 26312
rect 21091 26272 21100 26312
rect 21140 26272 22924 26312
rect 22964 26272 22973 26312
rect 28483 26272 28492 26312
rect 28532 26272 28541 26312
rect 29251 26272 29260 26312
rect 29300 26272 29548 26312
rect 29588 26272 36556 26312
rect 36596 26272 36605 26312
rect 37411 26272 37420 26312
rect 37460 26272 41836 26312
rect 41876 26272 41885 26312
rect 41932 26272 44620 26312
rect 44660 26272 44669 26312
rect 46051 26272 46060 26312
rect 46100 26272 48268 26312
rect 48308 26272 48317 26312
rect 14755 26271 14813 26272
rect 17635 26228 17693 26229
rect 28492 26228 28532 26272
rect 41932 26228 41972 26272
rect 14851 26188 14860 26228
rect 14900 26188 16436 26228
rect 17550 26188 17644 26228
rect 17684 26188 17693 26228
rect 17827 26188 17836 26228
rect 17876 26188 20140 26228
rect 20180 26188 20189 26228
rect 27907 26188 27916 26228
rect 27956 26188 29644 26228
rect 29684 26188 31180 26228
rect 31220 26188 31229 26228
rect 34339 26188 34348 26228
rect 34388 26188 35404 26228
rect 35444 26188 35453 26228
rect 37795 26188 37804 26228
rect 37844 26188 38284 26228
rect 38324 26188 38333 26228
rect 38467 26188 38476 26228
rect 38516 26188 39148 26228
rect 39188 26188 39628 26228
rect 39668 26188 39677 26228
rect 40588 26188 41452 26228
rect 41492 26188 41501 26228
rect 41923 26188 41932 26228
rect 41972 26188 41981 26228
rect 44227 26188 44236 26228
rect 44276 26188 47404 26228
rect 47444 26188 47453 26228
rect 16396 26144 16436 26188
rect 17635 26187 17693 26188
rect 28483 26144 28541 26145
rect 30595 26144 30653 26145
rect 40588 26144 40628 26188
rect 5347 26104 5356 26144
rect 5396 26104 6124 26144
rect 6164 26104 6173 26144
rect 7843 26104 7852 26144
rect 7892 26104 10060 26144
rect 10100 26104 10109 26144
rect 11203 26104 11212 26144
rect 11252 26104 12076 26144
rect 12116 26104 12125 26144
rect 13027 26104 13036 26144
rect 13076 26104 13228 26144
rect 13268 26104 13612 26144
rect 13652 26104 13661 26144
rect 13806 26104 13900 26144
rect 13940 26104 13949 26144
rect 14563 26104 14572 26144
rect 14612 26104 14621 26144
rect 15331 26104 15340 26144
rect 15380 26104 16012 26144
rect 16052 26104 16061 26144
rect 16387 26104 16396 26144
rect 16436 26104 16588 26144
rect 16628 26104 16972 26144
rect 17012 26104 17021 26144
rect 18211 26104 18220 26144
rect 18260 26104 19372 26144
rect 19412 26104 20332 26144
rect 20372 26104 20381 26144
rect 21667 26104 21676 26144
rect 21716 26104 24844 26144
rect 24884 26104 26860 26144
rect 26900 26104 26909 26144
rect 28398 26104 28492 26144
rect 28532 26104 28541 26144
rect 30510 26104 30604 26144
rect 30644 26104 30653 26144
rect 32803 26104 32812 26144
rect 32852 26104 33964 26144
rect 34004 26104 38188 26144
rect 38228 26104 38237 26144
rect 38755 26104 38764 26144
rect 38804 26104 39340 26144
rect 39380 26104 40588 26144
rect 40628 26104 40637 26144
rect 41347 26104 41356 26144
rect 41396 26104 42892 26144
rect 42932 26104 43084 26144
rect 43124 26104 43133 26144
rect 47107 26104 47116 26144
rect 47156 26104 48076 26144
rect 48116 26104 48125 26144
rect 49027 26104 49036 26144
rect 49076 26104 50956 26144
rect 50996 26104 51005 26144
rect 13891 26103 13949 26104
rect 28483 26103 28541 26104
rect 30595 26103 30653 26104
rect 49036 26060 49076 26104
rect 4099 26020 4108 26060
rect 4148 26020 5548 26060
rect 5588 26020 6220 26060
rect 6260 26020 6269 26060
rect 11491 26020 11500 26060
rect 11540 26020 15244 26060
rect 15284 26020 15293 26060
rect 15715 26020 15724 26060
rect 15764 26020 15773 26060
rect 16771 26020 16780 26060
rect 16820 26020 17260 26060
rect 17300 26020 18124 26060
rect 18164 26020 18173 26060
rect 20140 26020 21964 26060
rect 22004 26020 22252 26060
rect 22292 26020 22636 26060
rect 22676 26020 22685 26060
rect 34051 26020 34060 26060
rect 34100 26020 35212 26060
rect 35252 26020 35261 26060
rect 36259 26020 36268 26060
rect 36308 26020 37228 26060
rect 37268 26020 37277 26060
rect 37891 26020 37900 26060
rect 37940 26020 38956 26060
rect 38996 26020 39005 26060
rect 42307 26020 42316 26060
rect 42356 26020 44620 26060
rect 44660 26020 46004 26060
rect 47875 26020 47884 26060
rect 47924 26020 49076 26060
rect 15724 25976 15764 26020
rect 20140 25976 20180 26020
rect 45964 25976 46004 26020
rect 6883 25936 6892 25976
rect 6932 25936 7756 25976
rect 7796 25936 7805 25976
rect 13795 25936 13804 25976
rect 13844 25936 13996 25976
rect 14036 25936 20180 25976
rect 21475 25936 21484 25976
rect 21524 25936 22540 25976
rect 22580 25936 22589 25976
rect 29347 25936 29356 25976
rect 29396 25936 43948 25976
rect 43988 25936 43997 25976
rect 45955 25936 45964 25976
rect 46004 25936 46013 25976
rect 48067 25936 48076 25976
rect 48116 25936 49132 25976
rect 49172 25936 49181 25976
rect 2179 25852 2188 25892
rect 2228 25852 3052 25892
rect 3092 25852 3101 25892
rect 13699 25852 13708 25892
rect 13748 25852 14860 25892
rect 14900 25852 14909 25892
rect 17635 25852 17644 25892
rect 17684 25852 18316 25892
rect 18356 25852 18365 25892
rect 21091 25852 21100 25892
rect 21140 25852 22060 25892
rect 22100 25852 22109 25892
rect 29827 25852 29836 25892
rect 29876 25852 30604 25892
rect 30644 25852 31564 25892
rect 31604 25852 31613 25892
rect 32995 25852 33004 25892
rect 33044 25852 34348 25892
rect 34388 25852 34397 25892
rect 37219 25852 37228 25892
rect 37268 25852 38188 25892
rect 38228 25852 38237 25892
rect 40291 25852 40300 25892
rect 40340 25852 40684 25892
rect 40724 25852 40733 25892
rect 45571 25852 45580 25892
rect 45620 25852 50092 25892
rect 50132 25852 50141 25892
rect 0 25748 80 25828
rect 8899 25768 8908 25808
rect 8948 25768 12748 25808
rect 12788 25768 12797 25808
rect 14275 25768 14284 25808
rect 14324 25768 15532 25808
rect 15572 25768 15916 25808
rect 15956 25768 20236 25808
rect 20276 25768 25324 25808
rect 25364 25768 26956 25808
rect 26996 25768 27005 25808
rect 31171 25768 31180 25808
rect 31220 25768 36652 25808
rect 36692 25768 36701 25808
rect 38083 25768 38092 25808
rect 38132 25768 38476 25808
rect 38516 25768 38525 25808
rect 42019 25768 42028 25808
rect 42068 25768 42700 25808
rect 42740 25768 43756 25808
rect 43796 25768 43805 25808
rect 47875 25768 47884 25808
rect 47924 25768 50476 25808
rect 50516 25768 50525 25808
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 10531 25684 10540 25724
rect 10580 25684 12076 25724
rect 12116 25684 12125 25724
rect 15043 25684 15052 25724
rect 15092 25684 17876 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 47395 25684 47404 25724
rect 47444 25684 47788 25724
rect 47828 25684 47837 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 17836 25640 17876 25684
rect 9955 25600 9964 25640
rect 10004 25600 10732 25640
rect 10772 25600 11980 25640
rect 12020 25600 12940 25640
rect 12980 25600 12989 25640
rect 13516 25600 17740 25640
rect 17780 25600 17789 25640
rect 17836 25600 22156 25640
rect 22196 25600 22205 25640
rect 25123 25600 25132 25640
rect 25172 25600 28972 25640
rect 29012 25600 29021 25640
rect 47203 25600 47212 25640
rect 47252 25600 47596 25640
rect 47636 25600 48268 25640
rect 48308 25600 48317 25640
rect 13516 25556 13556 25600
rect 13699 25556 13757 25557
rect 3427 25516 3436 25556
rect 3476 25516 5356 25556
rect 5396 25516 5405 25556
rect 6307 25516 6316 25556
rect 6356 25516 13556 25556
rect 13614 25516 13708 25556
rect 13748 25516 13757 25556
rect 17827 25516 17836 25556
rect 17876 25516 18700 25556
rect 18740 25516 18749 25556
rect 23587 25516 23596 25556
rect 23636 25516 24748 25556
rect 24788 25516 24797 25556
rect 27907 25516 27916 25556
rect 27956 25516 30412 25556
rect 30452 25516 30461 25556
rect 37123 25516 37132 25556
rect 37172 25516 46252 25556
rect 46292 25516 46301 25556
rect 47011 25516 47020 25556
rect 47060 25516 48844 25556
rect 48884 25516 48893 25556
rect 49411 25516 49420 25556
rect 49460 25516 50764 25556
rect 50804 25516 50813 25556
rect 13699 25515 13757 25516
rect 26467 25472 26525 25473
rect 11011 25432 11020 25472
rect 11060 25432 11884 25472
rect 11924 25432 11933 25472
rect 13214 25432 13223 25472
rect 13263 25432 13612 25472
rect 13652 25432 13661 25472
rect 15139 25432 15148 25472
rect 15188 25432 16204 25472
rect 16244 25432 16253 25472
rect 16387 25432 16396 25472
rect 16436 25432 21772 25472
rect 21812 25432 21821 25472
rect 22339 25432 22348 25472
rect 22388 25432 23636 25472
rect 26382 25432 26476 25472
rect 26516 25432 26525 25472
rect 23596 25388 23636 25432
rect 26467 25431 26525 25432
rect 26572 25432 32660 25472
rect 32707 25432 32716 25472
rect 32756 25432 33388 25472
rect 33428 25432 33437 25472
rect 40579 25432 40588 25472
rect 40628 25432 47500 25472
rect 47540 25432 47549 25472
rect 48259 25432 48268 25472
rect 48308 25432 51148 25472
rect 51188 25432 51197 25472
rect 26572 25388 26612 25432
rect 32620 25388 32660 25432
rect 9283 25348 9292 25388
rect 9332 25348 12212 25388
rect 12643 25348 12652 25388
rect 12692 25348 12980 25388
rect 15043 25348 15052 25388
rect 15092 25348 15532 25388
rect 15572 25348 15581 25388
rect 15715 25348 15724 25388
rect 15764 25348 23500 25388
rect 23540 25348 23549 25388
rect 23596 25348 26612 25388
rect 28195 25348 28204 25388
rect 28244 25348 29260 25388
rect 29300 25348 31852 25388
rect 31892 25348 31901 25388
rect 32620 25348 36460 25388
rect 36500 25348 36509 25388
rect 37603 25348 37612 25388
rect 37652 25348 43372 25388
rect 43412 25348 43421 25388
rect 46147 25348 46156 25388
rect 46196 25348 46924 25388
rect 46964 25348 46973 25388
rect 12172 25304 12212 25348
rect 4195 25264 4204 25304
rect 4244 25264 6028 25304
rect 6068 25264 6077 25304
rect 7555 25264 7564 25304
rect 7604 25264 9100 25304
rect 9140 25264 9149 25304
rect 9379 25264 9388 25304
rect 9428 25264 10444 25304
rect 10484 25264 10493 25304
rect 10540 25264 10636 25304
rect 10676 25264 10685 25304
rect 10819 25264 10828 25304
rect 10868 25264 11884 25304
rect 11924 25264 11933 25304
rect 12163 25264 12172 25304
rect 12212 25264 12221 25304
rect 12268 25264 12556 25304
rect 12596 25264 12605 25304
rect 2467 25180 2476 25220
rect 2516 25180 3628 25220
rect 3668 25180 3677 25220
rect 3907 25180 3916 25220
rect 3956 25180 4300 25220
rect 4340 25180 4349 25220
rect 4396 25180 4588 25220
rect 4628 25180 4780 25220
rect 4820 25180 4829 25220
rect 4396 25136 4436 25180
rect 4003 25096 4012 25136
rect 4052 25096 4436 25136
rect 4483 25096 4492 25136
rect 4532 25096 5932 25136
rect 5972 25096 5981 25136
rect 6211 25096 6220 25136
rect 6260 25096 9868 25136
rect 9908 25096 9917 25136
rect 10540 25052 10580 25264
rect 12268 25220 12308 25264
rect 10636 25180 12308 25220
rect 12940 25220 12980 25348
rect 13603 25264 13612 25304
rect 13652 25264 14380 25304
rect 14420 25264 14429 25304
rect 15619 25264 15628 25304
rect 15668 25264 19276 25304
rect 19316 25264 19325 25304
rect 23587 25264 23596 25304
rect 23636 25264 24172 25304
rect 24212 25264 24221 25304
rect 24931 25264 24940 25304
rect 24980 25264 26380 25304
rect 26420 25264 26429 25304
rect 26851 25264 26860 25304
rect 26900 25264 27244 25304
rect 27284 25264 27293 25304
rect 32227 25264 32236 25304
rect 32276 25264 34252 25304
rect 34292 25264 34301 25304
rect 35875 25264 35884 25304
rect 35924 25264 38092 25304
rect 38132 25264 38141 25304
rect 38947 25264 38956 25304
rect 38996 25264 39340 25304
rect 39380 25264 39389 25304
rect 40291 25264 40300 25304
rect 40340 25264 40780 25304
rect 40820 25264 40829 25304
rect 41635 25264 41644 25304
rect 41684 25264 42892 25304
rect 42932 25264 42941 25304
rect 46435 25264 46444 25304
rect 46484 25264 47596 25304
rect 47636 25264 47788 25304
rect 47828 25264 47837 25304
rect 49795 25264 49804 25304
rect 49844 25264 51820 25304
rect 51860 25264 51869 25304
rect 45763 25220 45821 25221
rect 12940 25180 14476 25220
rect 14516 25180 14525 25220
rect 15235 25180 15244 25220
rect 15284 25180 15724 25220
rect 15764 25180 15916 25220
rect 15956 25180 15965 25220
rect 18499 25180 18508 25220
rect 18548 25180 19180 25220
rect 19220 25180 19229 25220
rect 26179 25180 26188 25220
rect 26228 25180 26572 25220
rect 26612 25180 26621 25220
rect 29827 25180 29836 25220
rect 29876 25180 31084 25220
rect 31124 25180 31660 25220
rect 31700 25180 35692 25220
rect 35732 25180 35980 25220
rect 36020 25180 36029 25220
rect 37027 25180 37036 25220
rect 37076 25180 40588 25220
rect 40628 25180 40637 25220
rect 43555 25180 43564 25220
rect 43604 25180 44332 25220
rect 44372 25180 44381 25220
rect 45678 25180 45772 25220
rect 45812 25180 45821 25220
rect 45955 25180 45964 25220
rect 46004 25180 46156 25220
rect 46196 25180 46348 25220
rect 46388 25180 46397 25220
rect 46819 25180 46828 25220
rect 46868 25180 49420 25220
rect 49460 25180 49469 25220
rect 10636 25136 10676 25180
rect 35980 25136 36020 25180
rect 45763 25179 45821 25180
rect 10627 25096 10636 25136
rect 10676 25096 10685 25136
rect 10828 25096 13900 25136
rect 13940 25096 13949 25136
rect 18115 25096 18124 25136
rect 18164 25096 18316 25136
rect 18356 25096 22156 25136
rect 22196 25096 22732 25136
rect 22772 25096 22781 25136
rect 35980 25096 37708 25136
rect 37748 25096 37757 25136
rect 45475 25096 45484 25136
rect 45524 25096 46540 25136
rect 46580 25096 46589 25136
rect 10828 25052 10868 25096
rect 5155 25012 5164 25052
rect 5204 25012 5836 25052
rect 5876 25012 5885 25052
rect 6499 25012 6508 25052
rect 6548 25012 6700 25052
rect 6740 25012 6749 25052
rect 10540 25012 10828 25052
rect 10868 25012 10877 25052
rect 11116 25012 13036 25052
rect 13076 25012 13085 25052
rect 0 24908 80 24988
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 9283 24928 9292 24968
rect 9332 24928 10060 24968
rect 10100 24928 10252 24968
rect 10292 24928 10301 24968
rect 11116 24884 11156 25012
rect 11299 24928 11308 24968
rect 11348 24928 13420 24968
rect 13460 24928 13469 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 7939 24844 7948 24884
rect 7988 24844 11156 24884
rect 12451 24844 12460 24884
rect 12500 24844 12844 24884
rect 12884 24844 12893 24884
rect 16963 24844 16972 24884
rect 17012 24844 20180 24884
rect 21859 24844 21868 24884
rect 21908 24844 22252 24884
rect 22292 24844 22301 24884
rect 23683 24844 23692 24884
rect 23732 24844 26324 24884
rect 27331 24844 27340 24884
rect 27380 24844 28108 24884
rect 28148 24844 30316 24884
rect 30356 24844 30365 24884
rect 40963 24844 40972 24884
rect 41012 24844 41452 24884
rect 41492 24844 41501 24884
rect 20140 24800 20180 24844
rect 26284 24800 26324 24844
rect 1027 24760 1036 24800
rect 1076 24760 1996 24800
rect 2036 24760 2045 24800
rect 4003 24760 4012 24800
rect 4052 24760 5164 24800
rect 5204 24760 5213 24800
rect 6028 24760 18220 24800
rect 18260 24760 18269 24800
rect 20140 24760 24076 24800
rect 24116 24760 24125 24800
rect 24547 24760 24556 24800
rect 24596 24760 26092 24800
rect 26132 24760 26141 24800
rect 26284 24760 30412 24800
rect 30452 24760 30461 24800
rect 31267 24760 31276 24800
rect 31316 24760 32620 24800
rect 32660 24760 32908 24800
rect 32948 24760 32957 24800
rect 40099 24760 40108 24800
rect 40148 24760 40492 24800
rect 40532 24760 40541 24800
rect 41539 24760 41548 24800
rect 41588 24760 43084 24800
rect 43124 24760 43133 24800
rect 931 24676 940 24716
rect 980 24676 4396 24716
rect 4436 24676 4445 24716
rect 6028 24632 6068 24760
rect 6115 24676 6124 24716
rect 6164 24676 7564 24716
rect 7604 24676 7613 24716
rect 8995 24676 9004 24716
rect 9044 24676 10348 24716
rect 10388 24676 10397 24716
rect 11683 24676 11692 24716
rect 11732 24676 13228 24716
rect 13268 24676 13277 24716
rect 26467 24676 26476 24716
rect 26516 24676 27436 24716
rect 27476 24676 27485 24716
rect 28960 24676 38860 24716
rect 38900 24676 38909 24716
rect 41059 24676 41068 24716
rect 41108 24676 41932 24716
rect 41972 24676 41981 24716
rect 46723 24676 46732 24716
rect 46772 24676 48748 24716
rect 48788 24676 48797 24716
rect 9004 24632 9044 24676
rect 28960 24632 29000 24676
rect 2083 24592 2092 24632
rect 2132 24592 2380 24632
rect 2420 24592 2429 24632
rect 2659 24592 2668 24632
rect 2708 24592 4588 24632
rect 4628 24592 4637 24632
rect 5731 24592 5740 24632
rect 5780 24592 6068 24632
rect 6499 24592 6508 24632
rect 6548 24592 9044 24632
rect 9955 24592 9964 24632
rect 10004 24592 10013 24632
rect 11971 24592 11980 24632
rect 12020 24592 12364 24632
rect 12404 24592 15244 24632
rect 15284 24592 15293 24632
rect 16099 24592 16108 24632
rect 16148 24592 16972 24632
rect 17012 24592 17260 24632
rect 17300 24592 17309 24632
rect 18403 24592 18412 24632
rect 18452 24592 21004 24632
rect 21044 24592 21053 24632
rect 21187 24592 21196 24632
rect 21236 24592 22252 24632
rect 22292 24592 22301 24632
rect 24355 24592 24364 24632
rect 24404 24592 25708 24632
rect 25748 24592 26188 24632
rect 26228 24592 26237 24632
rect 27235 24592 27244 24632
rect 27284 24592 29000 24632
rect 32131 24592 32140 24632
rect 32180 24592 33292 24632
rect 33332 24592 33341 24632
rect 38563 24592 38572 24632
rect 38612 24592 38764 24632
rect 38804 24592 39052 24632
rect 39092 24592 39101 24632
rect 39523 24592 39532 24632
rect 39572 24592 40780 24632
rect 40820 24592 40829 24632
rect 41251 24592 41260 24632
rect 41300 24592 41740 24632
rect 41780 24592 41789 24632
rect 46531 24592 46540 24632
rect 46580 24592 47212 24632
rect 47252 24592 47261 24632
rect 9964 24548 10004 24592
rect 11395 24548 11453 24549
rect 40780 24548 40820 24592
rect 2563 24508 2572 24548
rect 2612 24508 5260 24548
rect 5300 24508 5309 24548
rect 5635 24508 5644 24548
rect 5684 24508 7948 24548
rect 7988 24508 7997 24548
rect 9964 24508 11404 24548
rect 11444 24508 12652 24548
rect 12692 24508 12701 24548
rect 22147 24508 22156 24548
rect 22196 24508 26956 24548
rect 26996 24508 27340 24548
rect 27380 24508 27389 24548
rect 38659 24508 38668 24548
rect 38708 24508 40012 24548
rect 40052 24508 40061 24548
rect 40780 24508 41452 24548
rect 41492 24508 41501 24548
rect 11395 24507 11453 24508
rect 4771 24424 4780 24464
rect 4820 24424 6028 24464
rect 6068 24424 6412 24464
rect 6452 24424 6461 24464
rect 7267 24424 7276 24464
rect 7316 24424 8140 24464
rect 8180 24424 8189 24464
rect 8707 24424 8716 24464
rect 8756 24424 11308 24464
rect 11348 24424 11357 24464
rect 15715 24424 15724 24464
rect 15764 24424 16300 24464
rect 16340 24424 16349 24464
rect 21955 24424 21964 24464
rect 22004 24424 36556 24464
rect 36596 24424 36605 24464
rect 40963 24424 40972 24464
rect 41012 24424 41548 24464
rect 41588 24424 41932 24464
rect 41972 24424 41981 24464
rect 47491 24424 47500 24464
rect 47540 24424 47692 24464
rect 47732 24424 47741 24464
rect 41260 24380 41300 24424
rect 1603 24340 1612 24380
rect 1652 24340 2860 24380
rect 2900 24340 2909 24380
rect 5251 24340 5260 24380
rect 5300 24340 5644 24380
rect 5684 24340 6604 24380
rect 6644 24340 6653 24380
rect 13795 24340 13804 24380
rect 13844 24340 14380 24380
rect 14420 24340 14429 24380
rect 21475 24340 21484 24380
rect 21524 24340 21772 24380
rect 21812 24340 21821 24380
rect 29731 24340 29740 24380
rect 29780 24340 30124 24380
rect 30164 24340 30173 24380
rect 30979 24340 30988 24380
rect 31028 24340 32044 24380
rect 32084 24340 32093 24380
rect 39523 24340 39532 24380
rect 39572 24340 39724 24380
rect 39764 24340 40492 24380
rect 40532 24340 40541 24380
rect 41251 24340 41260 24380
rect 41300 24340 41340 24380
rect 47779 24340 47788 24380
rect 47828 24340 48364 24380
rect 48404 24340 48413 24380
rect 7843 24256 7852 24296
rect 7892 24256 20908 24296
rect 20948 24256 20957 24296
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 4099 24172 4108 24212
rect 4148 24172 5356 24212
rect 5396 24172 6316 24212
rect 6356 24172 6365 24212
rect 16675 24172 16684 24212
rect 16724 24172 17068 24212
rect 17108 24172 17932 24212
rect 17972 24172 17981 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 34051 24172 34060 24212
rect 34100 24172 34444 24212
rect 34484 24172 34493 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 0 24068 80 24148
rect 2371 24088 2380 24128
rect 2420 24088 4244 24128
rect 25507 24088 25516 24128
rect 25556 24088 30796 24128
rect 30836 24088 30845 24128
rect 33580 24088 34252 24128
rect 34292 24088 34301 24128
rect 4204 24044 4244 24088
rect 3523 24004 3532 24044
rect 3572 24004 4012 24044
rect 4052 24004 4061 24044
rect 4195 24004 4204 24044
rect 4244 24004 4780 24044
rect 4820 24004 4829 24044
rect 13891 24004 13900 24044
rect 13940 24004 13949 24044
rect 15523 24004 15532 24044
rect 15572 24004 17780 24044
rect 2659 23920 2668 23960
rect 2708 23920 6124 23960
rect 6164 23920 8044 23960
rect 8084 23920 8093 23960
rect 8707 23920 8716 23960
rect 8756 23920 9580 23960
rect 9620 23920 9629 23960
rect 13900 23876 13940 24004
rect 13987 23920 13996 23960
rect 14036 23920 15916 23960
rect 15956 23920 15965 23960
rect 16195 23920 16204 23960
rect 16244 23920 17548 23960
rect 17588 23920 17597 23960
rect 13900 23836 15436 23876
rect 15476 23836 15485 23876
rect 17740 23792 17780 24004
rect 20803 23920 20812 23960
rect 20852 23920 21580 23960
rect 21620 23920 21629 23960
rect 23779 23920 23788 23960
rect 23828 23920 25228 23960
rect 25268 23920 25277 23960
rect 26179 23920 26188 23960
rect 26228 23920 26764 23960
rect 26804 23920 26813 23960
rect 31267 23920 31276 23960
rect 31316 23920 32140 23960
rect 32180 23920 32189 23960
rect 32899 23920 32908 23960
rect 32948 23920 33524 23960
rect 33484 23876 33524 23920
rect 17827 23836 17836 23876
rect 17876 23836 18796 23876
rect 18836 23836 18845 23876
rect 23011 23836 23020 23876
rect 23060 23836 23884 23876
rect 23924 23836 28876 23876
rect 28916 23836 28925 23876
rect 32707 23836 32716 23876
rect 32756 23836 33004 23876
rect 33044 23836 33053 23876
rect 33475 23836 33484 23876
rect 33524 23836 33533 23876
rect 33580 23792 33620 24088
rect 48132 23920 48172 23960
rect 48212 23920 48221 23960
rect 51684 23920 51724 23960
rect 51764 23920 51773 23960
rect 48172 23876 48212 23920
rect 51724 23876 51764 23920
rect 45667 23836 45676 23876
rect 45716 23836 46540 23876
rect 46580 23836 46589 23876
rect 47299 23836 47308 23876
rect 47348 23836 47884 23876
rect 47924 23836 47933 23876
rect 48172 23836 50476 23876
rect 50516 23836 51764 23876
rect 3715 23752 3724 23792
rect 3764 23752 4876 23792
rect 4916 23752 4925 23792
rect 10051 23752 10060 23792
rect 10100 23752 11884 23792
rect 11924 23752 11933 23792
rect 12835 23752 12844 23792
rect 12884 23752 13900 23792
rect 13940 23752 16204 23792
rect 16244 23752 16253 23792
rect 16483 23752 16492 23792
rect 16532 23752 17548 23792
rect 17588 23752 17597 23792
rect 17731 23752 17740 23792
rect 17780 23752 17789 23792
rect 18979 23752 18988 23792
rect 19028 23752 19468 23792
rect 19508 23752 19517 23792
rect 25411 23752 25420 23792
rect 25460 23752 26092 23792
rect 26132 23752 26572 23792
rect 26612 23752 26621 23792
rect 28195 23752 28204 23792
rect 28244 23752 30412 23792
rect 30452 23752 30461 23792
rect 31267 23752 31276 23792
rect 31316 23752 32332 23792
rect 32372 23752 32381 23792
rect 33187 23752 33196 23792
rect 33236 23752 33620 23792
rect 33667 23752 33676 23792
rect 33716 23752 38188 23792
rect 38228 23752 38237 23792
rect 40099 23752 40108 23792
rect 40148 23752 41356 23792
rect 41396 23752 41405 23792
rect 42019 23752 42028 23792
rect 42068 23752 43276 23792
rect 43316 23752 43325 23792
rect 45187 23752 45196 23792
rect 45236 23752 45772 23792
rect 45812 23752 45821 23792
rect 45955 23752 45964 23792
rect 46004 23752 46640 23792
rect 13123 23708 13181 23709
rect 17740 23708 17780 23752
rect 46600 23708 46640 23752
rect 1123 23668 1132 23708
rect 1172 23668 4684 23708
rect 4724 23668 4733 23708
rect 11203 23668 11212 23708
rect 11252 23668 11692 23708
rect 11732 23668 11980 23708
rect 12020 23668 12029 23708
rect 12739 23668 12748 23708
rect 12788 23668 13132 23708
rect 13172 23668 16108 23708
rect 16148 23668 16157 23708
rect 17740 23668 27340 23708
rect 27380 23668 27389 23708
rect 32035 23668 32044 23708
rect 32084 23668 32524 23708
rect 32564 23668 33716 23708
rect 34531 23668 34540 23708
rect 34580 23668 36364 23708
rect 36404 23668 36413 23708
rect 40867 23668 40876 23708
rect 40916 23668 42604 23708
rect 42644 23668 42653 23708
rect 46600 23668 47212 23708
rect 47252 23668 47261 23708
rect 13123 23667 13181 23668
rect 16387 23584 16396 23624
rect 16436 23584 16972 23624
rect 17012 23584 19084 23624
rect 19124 23584 23404 23624
rect 23444 23584 23453 23624
rect 33676 23540 33716 23668
rect 41539 23584 41548 23624
rect 41588 23584 42220 23624
rect 42260 23584 42269 23624
rect 46147 23584 46156 23624
rect 46196 23584 47596 23624
rect 47636 23584 50188 23624
rect 50228 23584 50237 23624
rect 3811 23500 3820 23540
rect 3860 23500 5644 23540
rect 5684 23500 5693 23540
rect 16099 23500 16108 23540
rect 16148 23500 20716 23540
rect 20756 23500 20765 23540
rect 31075 23500 31084 23540
rect 31124 23500 32852 23540
rect 33667 23500 33676 23540
rect 33716 23500 33725 23540
rect 45859 23500 45868 23540
rect 45908 23500 46540 23540
rect 46580 23500 46589 23540
rect 32812 23456 32852 23500
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 21571 23416 21580 23456
rect 21620 23416 32524 23456
rect 32564 23416 32716 23456
rect 32756 23416 32765 23456
rect 32812 23416 33868 23456
rect 33908 23416 33917 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 37780 23416 39244 23456
rect 39284 23416 39293 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 37780 23372 37820 23416
rect 17539 23332 17548 23372
rect 17588 23332 19372 23372
rect 19412 23332 20812 23372
rect 20852 23332 20861 23372
rect 28963 23332 28972 23372
rect 29012 23332 30220 23372
rect 30260 23332 31948 23372
rect 31988 23332 31997 23372
rect 33955 23332 33964 23372
rect 34004 23332 37324 23372
rect 37364 23332 37820 23372
rect 47011 23332 47020 23372
rect 47060 23332 47404 23372
rect 47444 23332 47453 23372
rect 0 23228 80 23308
rect 3811 23248 3820 23288
rect 3860 23248 4492 23288
rect 4532 23248 5068 23288
rect 5108 23248 5117 23288
rect 8995 23248 9004 23288
rect 9044 23248 9868 23288
rect 9908 23248 9917 23288
rect 33091 23248 33100 23288
rect 33140 23248 33484 23288
rect 33524 23248 34348 23288
rect 34388 23248 34397 23288
rect 34531 23248 34540 23288
rect 34580 23248 35404 23288
rect 35444 23248 35453 23288
rect 46339 23248 46348 23288
rect 46388 23248 46828 23288
rect 46868 23248 47116 23288
rect 47156 23248 47165 23288
rect 16579 23164 16588 23204
rect 16628 23164 18988 23204
rect 19028 23164 19037 23204
rect 34915 23164 34924 23204
rect 34964 23164 35692 23204
rect 35732 23164 35741 23204
rect 4099 23080 4108 23120
rect 4148 23080 5836 23120
rect 5876 23080 5885 23120
rect 8803 23080 8812 23120
rect 8852 23080 10156 23120
rect 10196 23080 11212 23120
rect 11252 23080 11261 23120
rect 15523 23080 15532 23120
rect 15572 23080 16012 23120
rect 16052 23080 16061 23120
rect 16291 23080 16300 23120
rect 16340 23080 16780 23120
rect 16820 23080 16829 23120
rect 19651 23080 19660 23120
rect 19700 23080 21676 23120
rect 21716 23080 21725 23120
rect 24163 23080 24172 23120
rect 24212 23080 27052 23120
rect 27092 23080 27101 23120
rect 30403 23080 30412 23120
rect 30452 23080 35212 23120
rect 35252 23080 35500 23120
rect 35540 23080 35549 23120
rect 40483 23080 40492 23120
rect 40532 23080 41932 23120
rect 41972 23080 42604 23120
rect 42644 23080 43084 23120
rect 43124 23080 43133 23120
rect 43939 23080 43948 23120
rect 43988 23080 46924 23120
rect 46964 23080 46973 23120
rect 47587 23080 47596 23120
rect 47636 23080 48172 23120
rect 48212 23080 48221 23120
rect 49027 23080 49036 23120
rect 49076 23080 50476 23120
rect 50516 23080 50525 23120
rect 9283 22996 9292 23036
rect 9332 22996 9868 23036
rect 9908 22996 9917 23036
rect 16195 22996 16204 23036
rect 16244 22996 16876 23036
rect 16916 22996 18124 23036
rect 18164 22996 18173 23036
rect 17740 22952 17780 22996
rect 8995 22912 9004 22952
rect 9044 22912 10732 22952
rect 10772 22912 10781 22952
rect 15139 22912 15148 22952
rect 15188 22912 15724 22952
rect 15764 22912 15916 22952
rect 15956 22912 17452 22952
rect 17492 22912 17501 22952
rect 17731 22912 17740 22952
rect 17780 22912 17820 22952
rect 29155 22912 29164 22952
rect 29204 22912 30316 22952
rect 30356 22912 31468 22952
rect 31508 22912 31517 22952
rect 34723 22912 34732 22952
rect 34772 22912 35308 22952
rect 35348 22912 35357 22952
rect 37219 22912 37228 22952
rect 37268 22912 41644 22952
rect 41684 22912 41693 22952
rect 44227 22912 44236 22952
rect 44276 22912 47308 22952
rect 47348 22912 48364 22952
rect 48404 22912 48413 22952
rect 4867 22868 4925 22869
rect 4771 22828 4780 22868
rect 4820 22828 4876 22868
rect 4916 22828 4925 22868
rect 6019 22828 6028 22868
rect 6068 22828 6508 22868
rect 6548 22828 6557 22868
rect 9571 22828 9580 22868
rect 9620 22828 10060 22868
rect 10100 22828 10109 22868
rect 12547 22828 12556 22868
rect 12596 22828 13036 22868
rect 13076 22828 13085 22868
rect 43555 22828 43564 22868
rect 43604 22828 44140 22868
rect 44180 22828 44189 22868
rect 4867 22827 4925 22828
rect 5251 22744 5260 22784
rect 5300 22744 6124 22784
rect 6164 22744 7852 22784
rect 7892 22744 13516 22784
rect 13556 22744 13565 22784
rect 13699 22744 13708 22784
rect 13748 22744 15532 22784
rect 15572 22744 15581 22784
rect 17635 22744 17644 22784
rect 17684 22744 18700 22784
rect 18740 22744 18749 22784
rect 28099 22744 28108 22784
rect 28148 22744 29164 22784
rect 29204 22744 29213 22784
rect 43651 22744 43660 22784
rect 43700 22744 47444 22784
rect 47491 22744 47500 22784
rect 47540 22744 48076 22784
rect 48116 22744 48125 22784
rect 48364 22744 48940 22784
rect 48980 22744 48989 22784
rect 4771 22700 4829 22701
rect 47404 22700 47444 22744
rect 48364 22700 48404 22744
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 4771 22660 4780 22700
rect 4820 22660 4972 22700
rect 5012 22660 5021 22700
rect 5539 22660 5548 22700
rect 5588 22660 7372 22700
rect 7412 22660 7421 22700
rect 11875 22660 11884 22700
rect 11924 22660 12460 22700
rect 12500 22660 12509 22700
rect 14947 22660 14956 22700
rect 14996 22660 15436 22700
rect 15476 22660 15485 22700
rect 15619 22660 15628 22700
rect 15668 22660 16204 22700
rect 16244 22660 17260 22700
rect 17300 22660 17309 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 22435 22660 22444 22700
rect 22484 22660 23212 22700
rect 23252 22660 23261 22700
rect 23779 22660 23788 22700
rect 23828 22660 24364 22700
rect 24404 22660 24413 22700
rect 27043 22660 27052 22700
rect 27092 22660 28588 22700
rect 28628 22660 30316 22700
rect 30356 22660 30700 22700
rect 30740 22660 30749 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 39715 22660 39724 22700
rect 39764 22660 40396 22700
rect 40436 22660 40445 22700
rect 44419 22660 44428 22700
rect 44468 22660 45676 22700
rect 45716 22660 45725 22700
rect 45772 22660 46060 22700
rect 46100 22660 47212 22700
rect 47252 22660 47261 22700
rect 47404 22660 48404 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 4771 22659 4829 22660
rect 45772 22616 45812 22660
rect 47500 22616 47540 22660
rect 12259 22576 12268 22616
rect 12308 22576 12652 22616
rect 12692 22576 13516 22616
rect 13556 22576 13565 22616
rect 16003 22576 16012 22616
rect 16052 22576 17548 22616
rect 17588 22576 17597 22616
rect 42115 22576 42124 22616
rect 42164 22576 42508 22616
rect 42548 22576 45196 22616
rect 45236 22576 45245 22616
rect 45763 22576 45772 22616
rect 45812 22576 45821 22616
rect 47491 22576 47500 22616
rect 47540 22576 47549 22616
rect 14179 22492 14188 22532
rect 14228 22492 14764 22532
rect 14804 22492 14813 22532
rect 22339 22492 22348 22532
rect 22388 22492 23212 22532
rect 23252 22492 23261 22532
rect 32419 22492 32428 22532
rect 32468 22492 34060 22532
rect 34100 22492 34828 22532
rect 34868 22492 34877 22532
rect 0 22448 80 22468
rect 0 22408 652 22448
rect 692 22408 701 22448
rect 12931 22408 12940 22448
rect 12980 22408 15340 22448
rect 15380 22408 15389 22448
rect 19747 22408 19756 22448
rect 19796 22408 20332 22448
rect 20372 22408 20381 22448
rect 34147 22408 34156 22448
rect 34196 22408 35020 22448
rect 35060 22408 35069 22448
rect 41059 22408 41068 22448
rect 41108 22408 41932 22448
rect 41972 22408 43852 22448
rect 43892 22408 43901 22448
rect 44035 22408 44044 22448
rect 44084 22408 44524 22448
rect 44564 22408 44573 22448
rect 44995 22408 45004 22448
rect 45044 22408 45388 22448
rect 45428 22408 45437 22448
rect 49027 22408 49036 22448
rect 49076 22408 51628 22448
rect 51668 22408 51677 22448
rect 0 22388 80 22408
rect 44524 22364 44564 22408
rect 4387 22324 4396 22364
rect 4436 22324 5452 22364
rect 5492 22324 5644 22364
rect 5684 22324 5693 22364
rect 7555 22324 7564 22364
rect 7604 22324 10924 22364
rect 10964 22324 10973 22364
rect 18211 22324 18220 22364
rect 18260 22324 24268 22364
rect 24308 22324 24317 22364
rect 32899 22324 32908 22364
rect 32948 22324 33196 22364
rect 33236 22324 34444 22364
rect 34484 22324 34493 22364
rect 38755 22324 38764 22364
rect 38804 22324 39916 22364
rect 39956 22324 40780 22364
rect 40820 22324 41836 22364
rect 41876 22324 42988 22364
rect 43028 22324 43756 22364
rect 43796 22324 43805 22364
rect 44524 22324 46252 22364
rect 46292 22324 46301 22364
rect 4003 22240 4012 22280
rect 4052 22240 4300 22280
rect 4340 22240 4349 22280
rect 6115 22240 6124 22280
rect 6164 22240 7468 22280
rect 7508 22240 7517 22280
rect 11779 22240 11788 22280
rect 11828 22240 12556 22280
rect 12596 22240 12605 22280
rect 14659 22240 14668 22280
rect 14708 22240 15148 22280
rect 15188 22240 15197 22280
rect 17827 22240 17836 22280
rect 17876 22240 21196 22280
rect 21236 22240 24172 22280
rect 24212 22240 24221 22280
rect 31843 22240 31852 22280
rect 31892 22240 32428 22280
rect 32468 22240 32477 22280
rect 34051 22240 34060 22280
rect 34100 22240 36172 22280
rect 36212 22240 36844 22280
rect 36884 22240 38572 22280
rect 38612 22240 38621 22280
rect 40867 22240 40876 22280
rect 40916 22240 41740 22280
rect 41780 22240 41789 22280
rect 43651 22240 43660 22280
rect 43700 22240 44140 22280
rect 44180 22240 44189 22280
rect 46339 22240 46348 22280
rect 46388 22240 47020 22280
rect 47060 22240 47069 22280
rect 1699 22156 1708 22196
rect 1748 22156 4876 22196
rect 4916 22156 4925 22196
rect 7267 22156 7276 22196
rect 7316 22156 8236 22196
rect 8276 22156 8285 22196
rect 15523 22156 15532 22196
rect 15572 22156 18220 22196
rect 18260 22156 18269 22196
rect 32707 22156 32716 22196
rect 32756 22156 33772 22196
rect 33812 22156 33821 22196
rect 40099 22156 40108 22196
rect 40148 22156 41164 22196
rect 41204 22156 41213 22196
rect 43459 22156 43468 22196
rect 43508 22156 43852 22196
rect 43892 22156 43901 22196
rect 45379 22156 45388 22196
rect 45428 22156 46540 22196
rect 46580 22156 46589 22196
rect 47971 22156 47980 22196
rect 48020 22156 49228 22196
rect 49268 22156 49277 22196
rect 17539 22072 17548 22112
rect 17588 22072 18700 22112
rect 18740 22072 21292 22112
rect 21332 22072 21341 22112
rect 21859 22072 21868 22112
rect 21908 22072 22540 22112
rect 22580 22072 22589 22112
rect 39139 22072 39148 22112
rect 39188 22072 42124 22112
rect 42164 22072 42173 22112
rect 43171 22072 43180 22112
rect 43220 22072 49036 22112
rect 49076 22072 49085 22112
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 5155 21904 5164 21944
rect 5204 21904 5548 21944
rect 5588 21904 5597 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 32515 21904 32524 21944
rect 32564 21904 32716 21944
rect 32756 21904 32765 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 37987 21820 37996 21860
rect 38036 21820 38668 21860
rect 38708 21820 39052 21860
rect 39092 21820 40532 21860
rect 40963 21820 40972 21860
rect 41012 21820 41164 21860
rect 41204 21820 41213 21860
rect 4771 21776 4829 21777
rect 5059 21776 5117 21777
rect 21475 21776 21533 21777
rect 23107 21776 23165 21777
rect 40492 21776 40532 21820
rect 4483 21736 4492 21776
rect 4532 21736 4780 21776
rect 4820 21736 4829 21776
rect 4974 21736 5068 21776
rect 5108 21736 5117 21776
rect 21390 21736 21484 21776
rect 21524 21736 21533 21776
rect 23022 21736 23116 21776
rect 23156 21736 23165 21776
rect 25027 21736 25036 21776
rect 25076 21736 31564 21776
rect 31604 21736 32332 21776
rect 32372 21736 32381 21776
rect 37315 21736 37324 21776
rect 37364 21736 39340 21776
rect 39380 21736 39389 21776
rect 40483 21736 40492 21776
rect 40532 21736 42508 21776
rect 42548 21736 42557 21776
rect 46243 21736 46252 21776
rect 46292 21736 47212 21776
rect 47252 21736 47404 21776
rect 47444 21736 47453 21776
rect 4771 21735 4829 21736
rect 5059 21735 5117 21736
rect 21475 21735 21533 21736
rect 23107 21735 23165 21736
rect 6019 21692 6077 21693
rect 4867 21652 4876 21692
rect 4916 21652 6028 21692
rect 6068 21652 6604 21692
rect 6644 21652 6653 21692
rect 9772 21652 11212 21692
rect 11252 21652 11788 21692
rect 11828 21652 11837 21692
rect 22540 21652 26612 21692
rect 32803 21652 32812 21692
rect 32852 21652 33100 21692
rect 33140 21652 33149 21692
rect 38083 21652 38092 21692
rect 38132 21652 38380 21692
rect 38420 21652 38429 21692
rect 39436 21652 40300 21692
rect 40340 21652 40972 21692
rect 41012 21652 41021 21692
rect 44995 21652 45004 21692
rect 45044 21652 45580 21692
rect 45620 21652 46348 21692
rect 46388 21652 46397 21692
rect 47587 21652 47596 21692
rect 47636 21652 47980 21692
rect 48020 21652 48029 21692
rect 6019 21651 6077 21652
rect 0 21608 80 21628
rect 9772 21608 9812 21652
rect 22540 21608 22580 21652
rect 26572 21608 26612 21652
rect 39436 21608 39476 21652
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 5251 21568 5260 21608
rect 5300 21568 5309 21608
rect 5923 21568 5932 21608
rect 5972 21568 6508 21608
rect 6548 21568 6557 21608
rect 9763 21568 9772 21608
rect 9812 21568 9821 21608
rect 11395 21568 11404 21608
rect 11444 21568 13708 21608
rect 13748 21568 13757 21608
rect 18883 21568 18892 21608
rect 18932 21568 22540 21608
rect 22580 21568 22589 21608
rect 23971 21568 23980 21608
rect 24020 21568 24652 21608
rect 24692 21568 24701 21608
rect 25123 21568 25132 21608
rect 25172 21568 25804 21608
rect 25844 21568 25853 21608
rect 26563 21568 26572 21608
rect 26612 21568 30220 21608
rect 30260 21568 30269 21608
rect 30979 21568 30988 21608
rect 31028 21568 32236 21608
rect 32276 21568 32285 21608
rect 32419 21568 32428 21608
rect 32468 21568 34156 21608
rect 34196 21568 34205 21608
rect 35587 21568 35596 21608
rect 35636 21568 35645 21608
rect 38179 21568 38188 21608
rect 38228 21568 39436 21608
rect 39476 21568 39485 21608
rect 40195 21568 40204 21608
rect 40244 21568 40396 21608
rect 40436 21568 43372 21608
rect 43412 21568 43421 21608
rect 44227 21568 44236 21608
rect 44276 21568 45292 21608
rect 45332 21568 45341 21608
rect 47011 21568 47020 21608
rect 47060 21568 47692 21608
rect 47732 21568 47741 21608
rect 0 21548 80 21568
rect 5260 21440 5300 21568
rect 6595 21484 6604 21524
rect 6644 21484 8140 21524
rect 8180 21484 8524 21524
rect 8564 21484 8573 21524
rect 11491 21484 11500 21524
rect 11540 21484 13900 21524
rect 13940 21484 13949 21524
rect 23980 21440 24020 21568
rect 35596 21524 35636 21568
rect 24451 21484 24460 21524
rect 24500 21484 24940 21524
rect 24980 21484 25324 21524
rect 25364 21484 30604 21524
rect 30644 21484 30796 21524
rect 30836 21484 30845 21524
rect 31075 21484 31084 21524
rect 31124 21484 31756 21524
rect 31796 21484 32332 21524
rect 32372 21484 32908 21524
rect 32948 21484 33100 21524
rect 33140 21484 34348 21524
rect 34388 21484 35636 21524
rect 36451 21484 36460 21524
rect 36500 21484 38476 21524
rect 38516 21484 38525 21524
rect 41251 21484 41260 21524
rect 41300 21484 43468 21524
rect 43508 21484 44332 21524
rect 44372 21484 44381 21524
rect 48643 21484 48652 21524
rect 48692 21484 50284 21524
rect 50324 21484 50333 21524
rect 2083 21400 2092 21440
rect 2132 21400 5068 21440
rect 5108 21400 5117 21440
rect 5260 21400 5836 21440
rect 5876 21400 6220 21440
rect 6260 21400 6269 21440
rect 12067 21400 12076 21440
rect 12116 21400 12652 21440
rect 12692 21400 12701 21440
rect 21475 21400 21484 21440
rect 21524 21400 21676 21440
rect 21716 21400 21725 21440
rect 22627 21400 22636 21440
rect 22676 21400 23404 21440
rect 23444 21400 24020 21440
rect 29827 21400 29836 21440
rect 29876 21400 31180 21440
rect 31220 21400 31229 21440
rect 31363 21400 31372 21440
rect 31412 21400 31852 21440
rect 31892 21400 31901 21440
rect 32131 21400 32140 21440
rect 32180 21400 33196 21440
rect 33236 21400 33245 21440
rect 35587 21400 35596 21440
rect 35636 21400 36748 21440
rect 36788 21400 36797 21440
rect 40099 21400 40108 21440
rect 40148 21400 40876 21440
rect 40916 21400 40925 21440
rect 42883 21400 42892 21440
rect 42932 21400 44044 21440
rect 44084 21400 44093 21440
rect 44515 21400 44524 21440
rect 44564 21400 46540 21440
rect 46580 21400 46589 21440
rect 49027 21400 49036 21440
rect 49076 21400 49900 21440
rect 49940 21400 49949 21440
rect 10339 21316 10348 21356
rect 10388 21316 13132 21356
rect 13172 21316 13181 21356
rect 23587 21316 23596 21356
rect 23636 21316 24268 21356
rect 24308 21316 24317 21356
rect 5059 21272 5117 21273
rect 4963 21232 4972 21272
rect 5012 21232 5068 21272
rect 5108 21232 5117 21272
rect 5059 21231 5117 21232
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 4771 21148 4780 21188
rect 4820 21148 5644 21188
rect 5684 21148 5693 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 24259 21148 24268 21188
rect 24308 21148 25516 21188
rect 25556 21148 25565 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 41155 21148 41164 21188
rect 41204 21148 44908 21188
rect 44948 21148 44957 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 23107 21064 23116 21104
rect 23156 21064 23788 21104
rect 23828 21064 23837 21104
rect 37780 21064 38284 21104
rect 38324 21064 38333 21104
rect 21283 20980 21292 21020
rect 21332 20980 22060 21020
rect 22100 20980 22540 21020
rect 22580 20980 22589 21020
rect 37780 20936 37820 21064
rect 39331 20980 39340 21020
rect 39380 20980 42892 21020
rect 42932 20980 42941 21020
rect 259 20896 268 20936
rect 308 20896 15148 20936
rect 15188 20896 15197 20936
rect 21676 20896 23020 20936
rect 23060 20896 23500 20936
rect 23540 20896 23549 20936
rect 24835 20896 24844 20936
rect 24884 20896 24893 20936
rect 31651 20896 31660 20936
rect 31700 20896 31948 20936
rect 31988 20896 37820 20936
rect 21676 20852 21716 20896
rect 24844 20852 24884 20896
rect 6211 20812 6220 20852
rect 6260 20812 7756 20852
rect 7796 20812 8908 20852
rect 8948 20812 9868 20852
rect 9908 20812 10444 20852
rect 10484 20812 10493 20852
rect 21667 20812 21676 20852
rect 21716 20812 21725 20852
rect 22531 20812 22540 20852
rect 22580 20812 23212 20852
rect 23252 20812 24884 20852
rect 39052 20812 39820 20852
rect 39860 20812 39869 20852
rect 0 20768 80 20788
rect 4867 20768 4925 20769
rect 39052 20768 39092 20812
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 4483 20728 4492 20768
rect 4532 20728 4876 20768
rect 4916 20728 4925 20768
rect 5155 20728 5164 20768
rect 5204 20728 5740 20768
rect 5780 20728 5789 20768
rect 10627 20728 10636 20768
rect 10676 20728 11308 20768
rect 11348 20728 11357 20768
rect 20515 20728 20524 20768
rect 20564 20728 21388 20768
rect 21428 20728 21437 20768
rect 21571 20728 21580 20768
rect 21620 20728 22636 20768
rect 22676 20728 22685 20768
rect 23299 20728 23308 20768
rect 23348 20728 24268 20768
rect 24308 20728 24317 20768
rect 27427 20728 27436 20768
rect 27476 20728 28684 20768
rect 28724 20728 30508 20768
rect 30548 20728 30557 20768
rect 37987 20728 37996 20768
rect 38036 20728 39052 20768
rect 39092 20728 39101 20768
rect 39427 20728 39436 20768
rect 39476 20728 41068 20768
rect 41108 20728 41117 20768
rect 43267 20728 43276 20768
rect 43316 20728 45388 20768
rect 45428 20728 45437 20768
rect 46339 20728 46348 20768
rect 46388 20728 49036 20768
rect 49076 20728 49085 20768
rect 0 20708 80 20728
rect 4867 20727 4925 20728
rect 8995 20644 9004 20684
rect 9044 20644 9964 20684
rect 10004 20644 10013 20684
rect 21859 20644 21868 20684
rect 21908 20644 21917 20684
rect 21868 20600 21908 20644
rect 5251 20560 5260 20600
rect 5300 20560 5644 20600
rect 5684 20560 5693 20600
rect 18979 20560 18988 20600
rect 19028 20560 21292 20600
rect 21332 20560 21341 20600
rect 21475 20560 21484 20600
rect 21524 20560 21908 20600
rect 24547 20560 24556 20600
rect 24596 20560 38188 20600
rect 38228 20560 38237 20600
rect 38851 20560 38860 20600
rect 38900 20560 42220 20600
rect 42260 20560 42412 20600
rect 42452 20560 42796 20600
rect 42836 20560 42845 20600
rect 43747 20560 43756 20600
rect 43796 20560 44620 20600
rect 44660 20560 44669 20600
rect 47107 20560 47116 20600
rect 47156 20560 47788 20600
rect 47828 20560 47837 20600
rect 10435 20476 10444 20516
rect 10484 20476 11596 20516
rect 11636 20476 11645 20516
rect 20611 20476 20620 20516
rect 20660 20476 27148 20516
rect 27188 20476 27197 20516
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 20899 20392 20908 20432
rect 20948 20392 21964 20432
rect 22004 20392 22013 20432
rect 22723 20392 22732 20432
rect 22772 20392 24172 20432
rect 24212 20392 24221 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 4963 20308 4972 20348
rect 5012 20308 6796 20348
rect 6836 20308 6845 20348
rect 21379 20308 21388 20348
rect 21428 20308 21772 20348
rect 21812 20308 21821 20348
rect 25027 20308 25036 20348
rect 25076 20308 25708 20348
rect 25748 20308 25757 20348
rect 37987 20308 37996 20348
rect 38036 20308 38764 20348
rect 38804 20308 38813 20348
rect 41731 20308 41740 20348
rect 41780 20308 43948 20348
rect 43988 20308 43997 20348
rect 21475 20264 21533 20265
rect 4099 20224 4108 20264
rect 4148 20224 5164 20264
rect 5204 20224 5213 20264
rect 21390 20224 21484 20264
rect 21524 20224 21533 20264
rect 21667 20224 21676 20264
rect 21716 20224 22060 20264
rect 22100 20224 22109 20264
rect 24268 20224 27860 20264
rect 21475 20223 21533 20224
rect 24268 20180 24308 20224
rect 25612 20180 25652 20224
rect 27820 20180 27860 20224
rect 37780 20224 38420 20264
rect 41923 20224 41932 20264
rect 41972 20224 43084 20264
rect 43124 20224 43133 20264
rect 37780 20180 37820 20224
rect 38380 20180 38420 20224
rect 5539 20140 5548 20180
rect 5588 20140 5597 20180
rect 24259 20140 24268 20180
rect 24308 20140 24317 20180
rect 24420 20140 24460 20180
rect 24500 20140 24509 20180
rect 25603 20140 25612 20180
rect 25652 20140 25661 20180
rect 27811 20140 27820 20180
rect 27860 20140 27869 20180
rect 37612 20140 37820 20180
rect 38371 20140 38380 20180
rect 38420 20140 38429 20180
rect 3523 20056 3532 20096
rect 3572 20056 4876 20096
rect 4916 20056 4925 20096
rect 5548 20012 5588 20140
rect 23107 20096 23165 20097
rect 24460 20096 24500 20140
rect 26563 20096 26621 20097
rect 37612 20096 37652 20140
rect 5635 20056 5644 20096
rect 5684 20056 6508 20096
rect 6548 20056 6557 20096
rect 6883 20056 6892 20096
rect 6932 20056 7372 20096
rect 7412 20056 8716 20096
rect 8756 20056 8765 20096
rect 12451 20056 12460 20096
rect 12500 20056 13132 20096
rect 13172 20056 13181 20096
rect 13699 20056 13708 20096
rect 13748 20056 14284 20096
rect 14324 20056 14333 20096
rect 17539 20056 17548 20096
rect 17588 20056 18316 20096
rect 18356 20056 18365 20096
rect 19459 20056 19468 20096
rect 19508 20056 22156 20096
rect 22196 20056 22205 20096
rect 22531 20056 22540 20096
rect 22580 20056 23116 20096
rect 23156 20056 23165 20096
rect 23395 20056 23404 20096
rect 23444 20056 24500 20096
rect 24931 20056 24940 20096
rect 24980 20056 25516 20096
rect 25556 20056 25565 20096
rect 26478 20056 26572 20096
rect 26612 20056 26621 20096
rect 37411 20056 37420 20096
rect 37460 20056 37652 20096
rect 37780 20056 38092 20096
rect 38132 20056 38572 20096
rect 38612 20056 38621 20096
rect 41635 20056 41644 20096
rect 41684 20056 43372 20096
rect 43412 20056 45484 20096
rect 45524 20056 46348 20096
rect 46388 20056 46397 20096
rect 23107 20055 23165 20056
rect 26563 20055 26621 20056
rect 23116 20012 23156 20055
rect 37780 20012 37820 20056
rect 4003 19972 4012 20012
rect 4052 19972 5588 20012
rect 6595 19972 6604 20012
rect 6644 19972 9676 20012
rect 9716 19972 10252 20012
rect 10292 19972 10301 20012
rect 11683 19972 11692 20012
rect 11732 19972 13228 20012
rect 13268 19972 13277 20012
rect 17443 19972 17452 20012
rect 17492 19972 17501 20012
rect 18787 19972 18796 20012
rect 18836 19972 19660 20012
rect 19700 19972 19709 20012
rect 19756 19972 21004 20012
rect 21044 19972 21053 20012
rect 21955 19972 21964 20012
rect 22004 19972 22636 20012
rect 22676 19972 22685 20012
rect 23116 19972 24076 20012
rect 24116 19972 26188 20012
rect 26228 19972 26237 20012
rect 36547 19972 36556 20012
rect 36596 19972 37820 20012
rect 37891 19972 37900 20012
rect 37940 19972 38860 20012
rect 38900 19972 38909 20012
rect 39148 19972 41600 20012
rect 0 19928 80 19948
rect 6019 19928 6077 19929
rect 17452 19928 17492 19972
rect 19756 19928 19796 19972
rect 39148 19928 39188 19972
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 5934 19888 6028 19928
rect 6068 19888 6077 19928
rect 12259 19888 12268 19928
rect 12308 19888 12748 19928
rect 12788 19888 12797 19928
rect 16963 19888 16972 19928
rect 17012 19888 17356 19928
rect 17396 19888 17405 19928
rect 17452 19888 18892 19928
rect 18932 19888 18941 19928
rect 19171 19888 19180 19928
rect 19220 19888 19796 19928
rect 24355 19888 24364 19928
rect 24404 19888 25996 19928
rect 26036 19888 26045 19928
rect 36643 19888 36652 19928
rect 36692 19888 39188 19928
rect 41560 19928 41600 19972
rect 41560 19888 47788 19928
rect 47828 19888 47837 19928
rect 0 19868 80 19888
rect 6019 19887 6077 19888
rect 2947 19804 2956 19844
rect 2996 19804 4876 19844
rect 4916 19804 4925 19844
rect 11203 19804 11212 19844
rect 11252 19804 13420 19844
rect 13460 19804 13804 19844
rect 13844 19804 14284 19844
rect 14324 19804 14333 19844
rect 15811 19804 15820 19844
rect 15860 19804 26860 19844
rect 26900 19804 26909 19844
rect 38467 19804 38476 19844
rect 38516 19804 41260 19844
rect 41300 19804 41600 19844
rect 41560 19760 41600 19804
rect 11395 19720 11404 19760
rect 11444 19720 12556 19760
rect 12596 19720 12605 19760
rect 16387 19720 16396 19760
rect 16436 19720 35308 19760
rect 35348 19720 35692 19760
rect 35732 19720 35741 19760
rect 41560 19720 41836 19760
rect 41876 19720 42508 19760
rect 42548 19720 42557 19760
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 39619 19636 39628 19676
rect 39668 19636 43180 19676
rect 43220 19636 43852 19676
rect 43892 19636 43901 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 23299 19552 23308 19592
rect 23348 19552 23980 19592
rect 24020 19552 24029 19592
rect 29539 19552 29548 19592
rect 29588 19552 30316 19592
rect 30356 19552 30365 19592
rect 25219 19468 25228 19508
rect 25268 19468 25708 19508
rect 25748 19468 25757 19508
rect 27523 19468 27532 19508
rect 27572 19468 32908 19508
rect 32948 19468 37996 19508
rect 38036 19468 38045 19508
rect 38947 19468 38956 19508
rect 38996 19468 43852 19508
rect 43892 19468 43901 19508
rect 6595 19384 6604 19424
rect 6644 19384 6653 19424
rect 8515 19384 8524 19424
rect 8564 19384 9100 19424
rect 9140 19384 9149 19424
rect 38659 19384 38668 19424
rect 38708 19384 40108 19424
rect 40148 19384 40157 19424
rect 41560 19384 42316 19424
rect 42356 19384 42365 19424
rect 42883 19384 42892 19424
rect 42932 19384 44236 19424
rect 44276 19384 44285 19424
rect 45091 19384 45100 19424
rect 45140 19384 46348 19424
rect 46388 19384 46397 19424
rect 6604 19340 6644 19384
rect 5923 19300 5932 19340
rect 5972 19300 6220 19340
rect 6260 19300 6644 19340
rect 21283 19300 21292 19340
rect 21332 19300 23212 19340
rect 23252 19300 23261 19340
rect 23683 19300 23692 19340
rect 23732 19300 25324 19340
rect 25364 19300 25373 19340
rect 25987 19300 25996 19340
rect 26036 19300 26476 19340
rect 26516 19300 26525 19340
rect 38371 19300 38380 19340
rect 38420 19300 38956 19340
rect 38996 19300 39005 19340
rect 25996 19256 26036 19300
rect 41560 19256 41600 19384
rect 3811 19216 3820 19256
rect 3860 19216 5548 19256
rect 5588 19216 5597 19256
rect 6220 19216 8044 19256
rect 8084 19216 8093 19256
rect 11011 19216 11020 19256
rect 11060 19216 11500 19256
rect 11540 19216 11549 19256
rect 14755 19216 14764 19256
rect 14804 19216 16108 19256
rect 16148 19216 16157 19256
rect 18211 19216 18220 19256
rect 18260 19216 19372 19256
rect 19412 19216 19421 19256
rect 24355 19216 24364 19256
rect 24404 19216 25036 19256
rect 25076 19216 25228 19256
rect 25268 19216 26036 19256
rect 26179 19216 26188 19256
rect 26228 19216 29164 19256
rect 29204 19216 29213 19256
rect 30499 19216 30508 19256
rect 30548 19216 32140 19256
rect 32180 19216 32189 19256
rect 38467 19216 38476 19256
rect 38516 19216 39532 19256
rect 39572 19216 39581 19256
rect 40003 19216 40012 19256
rect 40052 19216 40492 19256
rect 40532 19216 41600 19256
rect 41923 19216 41932 19256
rect 41972 19216 42220 19256
rect 42260 19216 42269 19256
rect 43843 19216 43852 19256
rect 43892 19216 44236 19256
rect 44276 19216 44285 19256
rect 0 19088 80 19108
rect 6220 19088 6260 19216
rect 10243 19132 10252 19172
rect 10292 19132 11116 19172
rect 11156 19132 11165 19172
rect 23920 19132 24268 19172
rect 24308 19132 24317 19172
rect 28579 19132 28588 19172
rect 28628 19132 34252 19172
rect 34292 19132 34924 19172
rect 34964 19132 35116 19172
rect 35156 19132 35165 19172
rect 38851 19132 38860 19172
rect 38900 19132 39628 19172
rect 39668 19132 40396 19172
rect 40436 19132 40445 19172
rect 23920 19088 23960 19132
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 2275 19048 2284 19088
rect 2324 19048 3820 19088
rect 3860 19048 3869 19088
rect 6211 19048 6220 19088
rect 6260 19048 6269 19088
rect 13315 19048 13324 19088
rect 13364 19048 14380 19088
rect 14420 19048 15244 19088
rect 15284 19048 15916 19088
rect 15956 19048 15965 19088
rect 19363 19048 19372 19088
rect 19412 19048 20332 19088
rect 20372 19048 20381 19088
rect 20995 19048 21004 19088
rect 21044 19048 22444 19088
rect 22484 19048 23692 19088
rect 23732 19048 23741 19088
rect 23875 19048 23884 19088
rect 23924 19048 23960 19088
rect 29251 19048 29260 19088
rect 29300 19048 29740 19088
rect 29780 19048 29789 19088
rect 0 19028 80 19048
rect 3235 18964 3244 19004
rect 3284 18964 4012 19004
rect 4052 18964 4061 19004
rect 17155 18964 17164 19004
rect 17204 18964 17644 19004
rect 17684 18964 17693 19004
rect 19267 18964 19276 19004
rect 19316 18964 21100 19004
rect 21140 18964 22828 19004
rect 22868 18964 22877 19004
rect 28771 18964 28780 19004
rect 28820 18964 32812 19004
rect 32852 18964 35596 19004
rect 35636 18964 35645 19004
rect 38947 18964 38956 19004
rect 38996 18964 39956 19004
rect 6403 18920 6461 18921
rect 39916 18920 39956 18964
rect 2563 18880 2572 18920
rect 2612 18880 3148 18920
rect 3188 18880 3197 18920
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 6403 18880 6412 18920
rect 6452 18880 7180 18920
rect 7220 18880 7229 18920
rect 7363 18880 7372 18920
rect 7412 18880 8620 18920
rect 8660 18880 9964 18920
rect 10004 18880 10013 18920
rect 10627 18880 10636 18920
rect 10676 18880 11404 18920
rect 11444 18880 11453 18920
rect 17443 18880 17452 18920
rect 17492 18880 18028 18920
rect 18068 18880 18077 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 20803 18880 20812 18920
rect 20852 18880 21772 18920
rect 21812 18880 21821 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 38275 18880 38284 18920
rect 38324 18880 39148 18920
rect 39188 18880 39197 18920
rect 39907 18880 39916 18920
rect 39956 18880 40204 18920
rect 40244 18880 40684 18920
rect 40724 18880 40733 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 6403 18879 6461 18880
rect 835 18796 844 18836
rect 884 18796 6220 18836
rect 6260 18796 6269 18836
rect 17251 18796 17260 18836
rect 17300 18796 19124 18836
rect 22627 18796 22636 18836
rect 22676 18796 24268 18836
rect 24308 18796 24460 18836
rect 24500 18796 24844 18836
rect 24884 18796 24893 18836
rect 37795 18796 37804 18836
rect 37844 18796 38476 18836
rect 38516 18796 38525 18836
rect 19084 18752 19124 18796
rect 1891 18712 1900 18752
rect 1940 18712 2860 18752
rect 2900 18712 2909 18752
rect 3523 18712 3532 18752
rect 3572 18712 4108 18752
rect 4148 18712 5068 18752
rect 5108 18712 5356 18752
rect 5396 18712 5405 18752
rect 8707 18712 8716 18752
rect 8756 18712 9292 18752
rect 9332 18712 10060 18752
rect 10100 18712 10109 18752
rect 16963 18712 16972 18752
rect 17012 18712 17356 18752
rect 17396 18712 17405 18752
rect 19075 18712 19084 18752
rect 19124 18712 19133 18752
rect 25987 18712 25996 18752
rect 26036 18712 27916 18752
rect 27956 18712 28492 18752
rect 28532 18712 28541 18752
rect 29827 18712 29836 18752
rect 29876 18712 29885 18752
rect 32323 18712 32332 18752
rect 32372 18712 32908 18752
rect 32948 18712 32957 18752
rect 29836 18668 29876 18712
rect 5827 18628 5836 18668
rect 5876 18628 7468 18668
rect 7508 18628 7517 18668
rect 20707 18628 20716 18668
rect 20756 18628 21196 18668
rect 21236 18628 21868 18668
rect 21908 18628 22444 18668
rect 22484 18628 22493 18668
rect 28195 18628 28204 18668
rect 28244 18628 29548 18668
rect 29588 18628 29876 18668
rect 6403 18584 6461 18585
rect 20611 18584 20669 18585
rect 1987 18544 1996 18584
rect 2036 18544 2764 18584
rect 2804 18544 2813 18584
rect 5635 18544 5644 18584
rect 5684 18544 5932 18584
rect 5972 18544 6412 18584
rect 6452 18544 6461 18584
rect 6595 18544 6604 18584
rect 6644 18544 8044 18584
rect 8084 18544 8093 18584
rect 17635 18544 17644 18584
rect 17684 18544 19276 18584
rect 19316 18544 19325 18584
rect 20526 18544 20620 18584
rect 20660 18544 20669 18584
rect 20899 18544 20908 18584
rect 20948 18544 21292 18584
rect 21332 18544 22732 18584
rect 22772 18544 22781 18584
rect 24163 18544 24172 18584
rect 24212 18544 24652 18584
rect 24692 18544 24701 18584
rect 27715 18544 27724 18584
rect 27764 18544 28108 18584
rect 28148 18544 28780 18584
rect 28820 18544 29836 18584
rect 29876 18544 29885 18584
rect 32419 18544 32428 18584
rect 32468 18544 33100 18584
rect 33140 18544 33149 18584
rect 33763 18544 33772 18584
rect 33812 18544 35788 18584
rect 35828 18544 36844 18584
rect 36884 18544 37420 18584
rect 37460 18544 37469 18584
rect 39139 18544 39148 18584
rect 39188 18544 41644 18584
rect 41684 18544 42124 18584
rect 42164 18544 42173 18584
rect 44707 18544 44716 18584
rect 44756 18544 46732 18584
rect 46772 18544 46781 18584
rect 6403 18543 6461 18544
rect 20611 18543 20669 18544
rect 5059 18460 5068 18500
rect 5108 18460 5260 18500
rect 5300 18460 5309 18500
rect 6499 18460 6508 18500
rect 6548 18460 7372 18500
rect 7412 18460 7421 18500
rect 19075 18460 19084 18500
rect 19124 18460 19756 18500
rect 19796 18460 20524 18500
rect 20564 18460 20573 18500
rect 28387 18460 28396 18500
rect 28436 18460 28684 18500
rect 28724 18460 28733 18500
rect 6403 18376 6412 18416
rect 6452 18376 6796 18416
rect 6836 18376 6845 18416
rect 9763 18376 9772 18416
rect 9812 18376 10828 18416
rect 10868 18376 10877 18416
rect 21379 18376 21388 18416
rect 21428 18376 22060 18416
rect 22100 18376 22636 18416
rect 22676 18376 22685 18416
rect 24451 18376 24460 18416
rect 24500 18376 25708 18416
rect 25748 18376 25757 18416
rect 28960 18376 30028 18416
rect 30068 18376 36844 18416
rect 36884 18376 36893 18416
rect 19363 18332 19421 18333
rect 28960 18332 29000 18376
rect 5251 18292 5260 18332
rect 5300 18292 5932 18332
rect 5972 18292 5981 18332
rect 17443 18292 17452 18332
rect 17492 18292 18220 18332
rect 18260 18292 18269 18332
rect 18979 18292 18988 18332
rect 19028 18292 19372 18332
rect 19412 18292 19468 18332
rect 19508 18292 19517 18332
rect 28675 18292 28684 18332
rect 28724 18292 29000 18332
rect 30307 18292 30316 18332
rect 30356 18292 31564 18332
rect 31604 18292 31613 18332
rect 33667 18292 33676 18332
rect 33716 18292 34156 18332
rect 34196 18292 34205 18332
rect 40291 18292 40300 18332
rect 40340 18292 41068 18332
rect 41108 18292 41117 18332
rect 19363 18291 19421 18292
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 2755 18208 2764 18248
rect 2804 18208 5204 18248
rect 19267 18208 19276 18248
rect 19316 18208 20812 18248
rect 20852 18208 20861 18248
rect 27715 18208 27724 18248
rect 27764 18208 28012 18248
rect 28052 18208 28061 18248
rect 0 18188 80 18208
rect 5164 18165 5204 18208
rect 5155 18164 5213 18165
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 5155 18124 5164 18164
rect 5204 18124 5836 18164
rect 5876 18124 5885 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 20620 18124 21580 18164
rect 21620 18124 21629 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 5155 18123 5213 18124
rect 20620 18080 20660 18124
rect 14467 18040 14476 18080
rect 14516 18040 20660 18080
rect 20707 18040 20716 18080
rect 20756 18040 21388 18080
rect 21428 18040 21437 18080
rect 28960 18040 31852 18080
rect 31892 18040 31901 18080
rect 28960 17996 29000 18040
rect 6604 17956 7756 17996
rect 7796 17956 7805 17996
rect 18979 17956 18988 17996
rect 19028 17956 19372 17996
rect 19412 17956 19421 17996
rect 20515 17956 20524 17996
rect 20564 17956 21580 17996
rect 21620 17956 25516 17996
rect 25556 17956 25804 17996
rect 25844 17956 25853 17996
rect 26371 17956 26380 17996
rect 26420 17956 29000 17996
rect 29932 17956 30508 17996
rect 30548 17956 31180 17996
rect 31220 17956 31229 17996
rect 3619 17788 3628 17828
rect 3668 17788 4780 17828
rect 4820 17788 4829 17828
rect 4963 17788 4972 17828
rect 5012 17788 5740 17828
rect 5780 17788 6124 17828
rect 6164 17788 6173 17828
rect 6604 17744 6644 17956
rect 20323 17912 20381 17913
rect 6691 17872 6700 17912
rect 6740 17872 12076 17912
rect 12116 17872 12125 17912
rect 17539 17872 17548 17912
rect 17588 17872 19660 17912
rect 19700 17872 19709 17912
rect 20323 17872 20332 17912
rect 20372 17872 21100 17912
rect 21140 17872 21149 17912
rect 24835 17872 24844 17912
rect 24884 17872 25132 17912
rect 25172 17872 25181 17912
rect 28003 17872 28012 17912
rect 28052 17872 28492 17912
rect 28532 17872 28876 17912
rect 28916 17872 29740 17912
rect 29780 17872 29789 17912
rect 20323 17871 20381 17872
rect 28867 17828 28925 17829
rect 29932 17828 29972 17956
rect 30019 17872 30028 17912
rect 30068 17872 30700 17912
rect 30740 17872 30749 17912
rect 6796 17788 11404 17828
rect 11444 17788 11788 17828
rect 11828 17788 11837 17828
rect 17155 17788 17164 17828
rect 17204 17788 17740 17828
rect 17780 17788 17789 17828
rect 18316 17788 18796 17828
rect 18836 17788 18845 17828
rect 18979 17788 18988 17828
rect 19028 17788 20812 17828
rect 20852 17788 20861 17828
rect 20908 17788 21484 17828
rect 21524 17788 21964 17828
rect 22004 17788 24212 17828
rect 6796 17744 6836 17788
rect 4387 17704 4396 17744
rect 4436 17704 6028 17744
rect 6068 17704 6077 17744
rect 6595 17704 6604 17744
rect 6644 17704 6653 17744
rect 6787 17704 6796 17744
rect 6836 17704 6845 17744
rect 6979 17704 6988 17744
rect 7028 17704 7037 17744
rect 10051 17704 10060 17744
rect 10100 17704 10636 17744
rect 10676 17704 10685 17744
rect 6988 17660 7028 17704
rect 18316 17660 18356 17788
rect 20908 17744 20948 17788
rect 24172 17744 24212 17788
rect 28867 17788 28876 17828
rect 28916 17788 29972 17828
rect 32803 17788 32812 17828
rect 32852 17788 33100 17828
rect 33140 17788 33149 17828
rect 35299 17788 35308 17828
rect 35348 17788 43028 17828
rect 28867 17787 28925 17788
rect 18499 17704 18508 17744
rect 18548 17704 19276 17744
rect 19316 17704 19325 17744
rect 20899 17704 20908 17744
rect 20948 17704 20957 17744
rect 21379 17704 21388 17744
rect 21428 17704 21868 17744
rect 21908 17704 21917 17744
rect 22243 17704 22252 17744
rect 22292 17704 22828 17744
rect 22868 17704 22877 17744
rect 23779 17704 23788 17744
rect 23828 17704 23960 17744
rect 24163 17704 24172 17744
rect 24212 17704 24364 17744
rect 24404 17704 24413 17744
rect 28003 17704 28012 17744
rect 28052 17704 28972 17744
rect 29012 17704 29452 17744
rect 29492 17704 29501 17744
rect 30979 17704 30988 17744
rect 31028 17704 31037 17744
rect 32515 17704 32524 17744
rect 32564 17704 33292 17744
rect 33332 17704 34444 17744
rect 34484 17704 34493 17744
rect 37699 17704 37708 17744
rect 37748 17704 38860 17744
rect 38900 17704 38909 17744
rect 41347 17704 41356 17744
rect 41396 17704 42892 17744
rect 42932 17704 42941 17744
rect 21868 17660 21908 17704
rect 23920 17660 23960 17704
rect 28867 17660 28925 17661
rect 30988 17660 31028 17704
rect 42988 17660 43028 17788
rect 4579 17620 4588 17660
rect 4628 17620 4972 17660
rect 5012 17620 5021 17660
rect 5731 17620 5740 17660
rect 5780 17620 7028 17660
rect 14755 17620 14764 17660
rect 14804 17620 16300 17660
rect 16340 17620 16349 17660
rect 18115 17620 18124 17660
rect 18164 17620 18356 17660
rect 18403 17620 18412 17660
rect 18452 17620 19181 17660
rect 19221 17620 19230 17660
rect 21868 17620 22540 17660
rect 22580 17620 22589 17660
rect 23920 17620 28876 17660
rect 28916 17620 28925 17660
rect 28867 17619 28925 17620
rect 28972 17620 31028 17660
rect 32419 17620 32428 17660
rect 32468 17620 33196 17660
rect 33236 17620 33245 17660
rect 33379 17620 33388 17660
rect 33428 17620 34060 17660
rect 34100 17620 34109 17660
rect 42979 17620 42988 17660
rect 43028 17620 44620 17660
rect 44660 17620 44669 17660
rect 5347 17536 5356 17576
rect 5396 17536 5644 17576
rect 5684 17536 5693 17576
rect 6979 17536 6988 17576
rect 7028 17536 8332 17576
rect 8372 17536 8381 17576
rect 16963 17536 16972 17576
rect 17012 17536 19372 17576
rect 19412 17536 19421 17576
rect 19651 17536 19660 17576
rect 19700 17536 19709 17576
rect 28195 17536 28204 17576
rect 28244 17536 28780 17576
rect 28820 17536 28829 17576
rect 19660 17492 19700 17536
rect 16099 17452 16108 17492
rect 16148 17452 17356 17492
rect 17396 17452 19700 17492
rect 0 17408 80 17428
rect 28003 17408 28061 17409
rect 28972 17408 29012 17620
rect 29347 17536 29356 17576
rect 29396 17536 29548 17576
rect 29588 17536 29597 17576
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 18019 17368 18028 17408
rect 18068 17368 18700 17408
rect 18740 17368 18749 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 28003 17368 28012 17408
rect 28052 17368 28588 17408
rect 28628 17368 28637 17408
rect 28963 17368 28972 17408
rect 29012 17368 29021 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 28003 17367 28061 17368
rect 19363 17324 19421 17325
rect 17443 17284 17452 17324
rect 17492 17284 19372 17324
rect 19412 17284 19421 17324
rect 19363 17283 19421 17284
rect 28108 17284 28396 17324
rect 28436 17284 28445 17324
rect 16003 17200 16012 17240
rect 16052 17200 17836 17240
rect 17876 17200 17885 17240
rect 18307 17200 18316 17240
rect 18356 17200 18700 17240
rect 18740 17200 19084 17240
rect 19124 17200 19133 17240
rect 24739 17200 24748 17240
rect 24788 17200 25324 17240
rect 25364 17200 25612 17240
rect 25652 17200 25661 17240
rect 26563 17200 26572 17240
rect 26612 17200 27340 17240
rect 27380 17200 27532 17240
rect 27572 17200 27581 17240
rect 28108 17156 28148 17284
rect 28195 17200 28204 17240
rect 28244 17200 28684 17240
rect 28724 17200 28733 17240
rect 28867 17200 28876 17240
rect 28916 17200 29164 17240
rect 29204 17200 29213 17240
rect 6979 17116 6988 17156
rect 7028 17116 9868 17156
rect 9908 17116 9917 17156
rect 18787 17116 18796 17156
rect 18836 17116 20044 17156
rect 20084 17116 23884 17156
rect 23924 17116 23933 17156
rect 28099 17116 28108 17156
rect 28148 17116 28157 17156
rect 1027 17032 1036 17072
rect 1076 17032 1708 17072
rect 1748 17032 1757 17072
rect 2563 17032 2572 17072
rect 2612 17032 3628 17072
rect 3668 17032 3677 17072
rect 4867 17032 4876 17072
rect 4916 17032 7372 17072
rect 7412 17032 8812 17072
rect 8852 17032 8861 17072
rect 9187 17032 9196 17072
rect 9236 17032 9388 17072
rect 9428 17032 9437 17072
rect 15907 17032 15916 17072
rect 15956 17032 16780 17072
rect 16820 17032 17164 17072
rect 17204 17032 17213 17072
rect 18211 17032 18220 17072
rect 18260 17032 18892 17072
rect 18932 17032 18941 17072
rect 21667 17032 21676 17072
rect 21716 17032 22156 17072
rect 22196 17032 22676 17072
rect 18115 16988 18173 16989
rect 22636 16988 22676 17032
rect 23920 17032 26380 17072
rect 26420 17032 26429 17072
rect 27715 17032 27724 17072
rect 27764 17032 27916 17072
rect 27956 17032 27965 17072
rect 28387 17032 28396 17072
rect 28436 17032 28684 17072
rect 28724 17032 28733 17072
rect 29251 17032 29260 17072
rect 29300 17032 30028 17072
rect 30068 17032 30077 17072
rect 30979 17032 30988 17072
rect 31028 17032 32524 17072
rect 32564 17032 32573 17072
rect 34531 17032 34540 17072
rect 34580 17032 36556 17072
rect 36596 17032 38572 17072
rect 38612 17032 40300 17072
rect 40340 17032 40349 17072
rect 23920 16988 23960 17032
rect 6307 16948 6316 16988
rect 6356 16948 6604 16988
rect 6644 16948 6653 16988
rect 7171 16948 7180 16988
rect 7220 16948 7229 16988
rect 18030 16948 18124 16988
rect 18164 16948 18173 16988
rect 22627 16948 22636 16988
rect 22676 16948 23960 16988
rect 26563 16948 26572 16988
rect 26612 16948 29644 16988
rect 29684 16948 29693 16988
rect 30604 16948 31372 16988
rect 31412 16948 32236 16988
rect 32276 16948 32285 16988
rect 35683 16948 35692 16988
rect 35732 16948 36460 16988
rect 36500 16948 36652 16988
rect 36692 16948 36701 16988
rect 37027 16948 37036 16988
rect 37076 16948 39532 16988
rect 39572 16948 39724 16988
rect 39764 16948 39773 16988
rect 7180 16904 7220 16948
rect 18115 16947 18173 16948
rect 30604 16904 30644 16948
rect 6787 16864 6796 16904
rect 6836 16864 7220 16904
rect 7459 16864 7468 16904
rect 7508 16864 8524 16904
rect 8564 16864 8573 16904
rect 23920 16864 30644 16904
rect 30691 16864 30700 16904
rect 30740 16864 33292 16904
rect 33332 16864 33341 16904
rect 23920 16820 23960 16864
rect 7651 16780 7660 16820
rect 7700 16780 7948 16820
rect 7988 16780 7997 16820
rect 17539 16780 17548 16820
rect 17588 16780 18604 16820
rect 18644 16780 18653 16820
rect 21091 16780 21100 16820
rect 21140 16780 23960 16820
rect 24556 16780 27436 16820
rect 27476 16780 27628 16820
rect 27668 16780 27677 16820
rect 28099 16780 28108 16820
rect 28148 16780 30220 16820
rect 30260 16780 30269 16820
rect 32131 16780 32140 16820
rect 32180 16780 32620 16820
rect 32660 16780 32669 16820
rect 36643 16780 36652 16820
rect 36692 16780 36844 16820
rect 36884 16780 36893 16820
rect 24556 16736 24596 16780
rect 6691 16696 6700 16736
rect 6740 16696 7564 16736
rect 7604 16696 7613 16736
rect 22915 16696 22924 16736
rect 22964 16696 24596 16736
rect 24643 16696 24652 16736
rect 24692 16696 25612 16736
rect 25652 16696 26572 16736
rect 26612 16696 26621 16736
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 31075 16612 31084 16652
rect 31124 16612 32428 16652
rect 32468 16612 32477 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 31651 16568 31709 16569
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 29155 16528 29164 16568
rect 29204 16528 29452 16568
rect 29492 16528 29501 16568
rect 29827 16528 29836 16568
rect 29876 16528 31660 16568
rect 31700 16528 31709 16568
rect 0 16508 80 16528
rect 31651 16527 31709 16528
rect 27715 16444 27724 16484
rect 27764 16444 32332 16484
rect 32372 16444 32381 16484
rect 1219 16360 1228 16400
rect 1268 16360 2092 16400
rect 2132 16360 2141 16400
rect 2188 16360 5068 16400
rect 5108 16360 5117 16400
rect 6403 16360 6412 16400
rect 6452 16360 6461 16400
rect 13603 16360 13612 16400
rect 13652 16360 13996 16400
rect 14036 16360 14045 16400
rect 15331 16360 15340 16400
rect 15380 16360 18700 16400
rect 18740 16360 18749 16400
rect 20419 16360 20428 16400
rect 20468 16360 21580 16400
rect 21620 16360 22060 16400
rect 22100 16360 22109 16400
rect 28387 16360 28396 16400
rect 28436 16360 30508 16400
rect 30548 16360 30557 16400
rect 31171 16360 31180 16400
rect 31220 16360 31564 16400
rect 31604 16360 31613 16400
rect 31660 16360 32564 16400
rect 32611 16360 32620 16400
rect 32660 16360 33004 16400
rect 33044 16360 33053 16400
rect 35587 16360 35596 16400
rect 35636 16360 36652 16400
rect 36692 16360 36701 16400
rect 2188 16316 2228 16360
rect 2179 16276 2188 16316
rect 2228 16276 2237 16316
rect 1603 16192 1612 16232
rect 1652 16192 4204 16232
rect 4244 16192 4253 16232
rect 4867 16192 4876 16232
rect 4916 16192 4925 16232
rect 4876 16148 4916 16192
rect 1219 16108 1228 16148
rect 1268 16108 4916 16148
rect 6412 16064 6452 16360
rect 28867 16316 28925 16317
rect 31660 16316 31700 16360
rect 32131 16316 32189 16317
rect 15043 16276 15052 16316
rect 15092 16276 16972 16316
rect 17012 16276 18836 16316
rect 19171 16276 19180 16316
rect 19220 16276 20236 16316
rect 20276 16276 20908 16316
rect 20948 16276 23060 16316
rect 26755 16276 26764 16316
rect 26804 16276 27148 16316
rect 27188 16276 27197 16316
rect 27331 16276 27340 16316
rect 27380 16276 27916 16316
rect 27956 16276 27965 16316
rect 28867 16276 28876 16316
rect 28916 16276 29260 16316
rect 29300 16276 29309 16316
rect 30211 16276 30220 16316
rect 30260 16276 30892 16316
rect 30932 16276 31372 16316
rect 31412 16276 31700 16316
rect 32046 16276 32140 16316
rect 32180 16276 32189 16316
rect 32524 16316 32564 16360
rect 34147 16316 34205 16317
rect 32524 16276 34156 16316
rect 34196 16276 35212 16316
rect 35252 16276 35261 16316
rect 18796 16232 18836 16276
rect 19939 16232 19997 16233
rect 23020 16232 23060 16276
rect 28867 16275 28925 16276
rect 32131 16275 32189 16276
rect 34147 16275 34205 16276
rect 7267 16192 7276 16232
rect 7316 16192 8332 16232
rect 8372 16192 8381 16232
rect 14179 16192 14188 16232
rect 14228 16192 14668 16232
rect 14708 16192 14717 16232
rect 16579 16192 16588 16232
rect 16628 16192 18028 16232
rect 18068 16192 18700 16232
rect 18740 16192 18749 16232
rect 18796 16192 19948 16232
rect 19988 16192 19997 16232
rect 20131 16192 20140 16232
rect 20180 16192 20812 16232
rect 20852 16192 21676 16232
rect 21716 16192 21725 16232
rect 23011 16192 23020 16232
rect 23060 16192 23884 16232
rect 23924 16192 23933 16232
rect 28003 16192 28012 16232
rect 28052 16192 30508 16232
rect 30548 16192 31084 16232
rect 31124 16192 31133 16232
rect 31747 16192 31756 16232
rect 31796 16192 34252 16232
rect 34292 16192 34301 16232
rect 19939 16191 19997 16192
rect 16003 16108 16012 16148
rect 16052 16108 16396 16148
rect 16436 16108 16445 16148
rect 29827 16108 29836 16148
rect 29876 16108 30988 16148
rect 31028 16108 31276 16148
rect 31316 16108 31325 16148
rect 31948 16108 32044 16148
rect 32084 16108 32093 16148
rect 32419 16108 32428 16148
rect 32468 16108 37228 16148
rect 37268 16108 37277 16148
rect 31948 16065 31988 16108
rect 31939 16064 31997 16065
rect 1411 16024 1420 16064
rect 1460 16024 3340 16064
rect 3380 16024 3389 16064
rect 5354 16024 5363 16064
rect 5403 16024 6836 16064
rect 7555 16024 7564 16064
rect 7604 16024 8908 16064
rect 8948 16024 8957 16064
rect 18595 16024 18604 16064
rect 18644 16024 19180 16064
rect 19220 16024 19229 16064
rect 20899 16024 20908 16064
rect 20948 16024 21580 16064
rect 21620 16024 21629 16064
rect 24835 16024 24844 16064
rect 24884 16024 25516 16064
rect 25556 16024 25565 16064
rect 25699 16024 25708 16064
rect 25748 16024 26860 16064
rect 26900 16024 26909 16064
rect 27235 16024 27244 16064
rect 27284 16024 27293 16064
rect 27427 16024 27436 16064
rect 27476 16024 27916 16064
rect 27956 16024 27965 16064
rect 31555 16024 31564 16064
rect 31604 16024 31948 16064
rect 31988 16024 31997 16064
rect 32131 16024 32140 16064
rect 32180 16024 32620 16064
rect 32660 16024 33580 16064
rect 33620 16024 33629 16064
rect 36931 16024 36940 16064
rect 36980 16024 37420 16064
rect 37460 16024 37469 16064
rect 1123 15940 1132 15980
rect 1172 15940 2476 15980
rect 2516 15940 2525 15980
rect 3907 15940 3916 15980
rect 3956 15940 6412 15980
rect 6452 15940 6461 15980
rect 4771 15896 4829 15897
rect 6796 15896 6836 16024
rect 27244 15896 27284 16024
rect 31939 16023 31997 16024
rect 28960 15940 32812 15980
rect 32852 15940 32861 15980
rect 28960 15896 29000 15940
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 4771 15856 4780 15896
rect 4820 15856 4914 15896
rect 5059 15856 5068 15896
rect 5108 15856 5932 15896
rect 5972 15856 5981 15896
rect 6211 15856 6220 15896
rect 6260 15856 6508 15896
rect 6548 15856 6557 15896
rect 6787 15856 6796 15896
rect 6836 15856 7468 15896
rect 7508 15856 9100 15896
rect 9140 15856 9149 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 27244 15856 29000 15896
rect 30307 15856 30316 15896
rect 30356 15856 31468 15896
rect 31508 15856 31517 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 4771 15855 4829 15856
rect 5068 15812 5108 15856
rect 4099 15772 4108 15812
rect 4148 15772 5108 15812
rect 5260 15772 5452 15812
rect 5492 15772 6028 15812
rect 6068 15772 6077 15812
rect 26083 15772 26092 15812
rect 26132 15772 29000 15812
rect 30211 15772 30220 15812
rect 30260 15772 36652 15812
rect 36692 15772 36701 15812
rect 0 15728 80 15748
rect 0 15688 748 15728
rect 788 15688 797 15728
rect 4003 15688 4012 15728
rect 4052 15688 4972 15728
rect 5012 15688 5021 15728
rect 0 15668 80 15688
rect 5260 15644 5300 15772
rect 5347 15688 5356 15728
rect 5396 15688 5644 15728
rect 5684 15688 5693 15728
rect 6595 15688 6604 15728
rect 6644 15688 7084 15728
rect 7124 15688 7133 15728
rect 7651 15688 7660 15728
rect 7700 15688 8620 15728
rect 8660 15688 8669 15728
rect 9571 15688 9580 15728
rect 9620 15688 10348 15728
rect 10388 15688 10397 15728
rect 20131 15688 20140 15728
rect 20180 15688 21196 15728
rect 21236 15688 21245 15728
rect 26851 15688 26860 15728
rect 26900 15688 28492 15728
rect 28532 15688 28541 15728
rect 28960 15644 29000 15772
rect 29251 15688 29260 15728
rect 29300 15688 30124 15728
rect 30164 15688 30173 15728
rect 31363 15688 31372 15728
rect 31412 15688 31660 15728
rect 31700 15688 31709 15728
rect 2467 15604 2476 15644
rect 2516 15604 4300 15644
rect 4340 15604 5300 15644
rect 7171 15604 7180 15644
rect 7220 15604 7564 15644
rect 7604 15604 7613 15644
rect 18691 15604 18700 15644
rect 18740 15604 20180 15644
rect 27043 15604 27052 15644
rect 27092 15604 27340 15644
rect 27380 15604 27389 15644
rect 28387 15604 28396 15644
rect 28436 15604 28684 15644
rect 28724 15604 28733 15644
rect 28960 15604 29068 15644
rect 29108 15604 29548 15644
rect 29588 15604 30796 15644
rect 30836 15604 33676 15644
rect 33716 15604 34156 15644
rect 34196 15604 37460 15644
rect 20140 15560 20180 15604
rect 34339 15560 34397 15561
rect 37420 15560 37460 15604
rect 1123 15520 1132 15560
rect 1172 15520 1708 15560
rect 1748 15520 1757 15560
rect 2371 15520 2380 15560
rect 2420 15520 3628 15560
rect 3668 15520 3677 15560
rect 5443 15520 5452 15560
rect 5492 15520 6988 15560
rect 7028 15520 7468 15560
rect 7508 15520 7517 15560
rect 15619 15520 15628 15560
rect 15668 15520 15820 15560
rect 15860 15520 15869 15560
rect 16195 15520 16204 15560
rect 16244 15520 16876 15560
rect 16916 15520 17644 15560
rect 17684 15520 17693 15560
rect 18499 15520 18508 15560
rect 18548 15520 19276 15560
rect 19316 15520 19325 15560
rect 20131 15520 20140 15560
rect 20180 15520 20189 15560
rect 20419 15520 20428 15560
rect 20468 15520 20477 15560
rect 20899 15520 20908 15560
rect 20948 15520 21868 15560
rect 21908 15520 21917 15560
rect 24259 15520 24268 15560
rect 24308 15520 25228 15560
rect 25268 15520 30316 15560
rect 30356 15520 30365 15560
rect 30691 15520 30700 15560
rect 30740 15520 32524 15560
rect 32564 15520 32573 15560
rect 33379 15520 33388 15560
rect 33428 15520 33964 15560
rect 34004 15520 34013 15560
rect 34243 15520 34252 15560
rect 34292 15520 34348 15560
rect 34388 15520 34444 15560
rect 34484 15520 34512 15560
rect 37411 15520 37420 15560
rect 37460 15520 38284 15560
rect 38324 15520 38333 15560
rect 41635 15520 41644 15560
rect 41684 15520 42604 15560
rect 42644 15520 43948 15560
rect 43988 15520 43997 15560
rect 4867 15436 4876 15476
rect 4916 15436 5260 15476
rect 5300 15436 5309 15476
rect 6211 15436 6220 15476
rect 6260 15436 6604 15476
rect 6644 15436 6653 15476
rect 10915 15436 10924 15476
rect 10964 15436 11212 15476
rect 11252 15436 11261 15476
rect 5155 15392 5213 15393
rect 5070 15352 5164 15392
rect 5204 15352 5213 15392
rect 5155 15351 5213 15352
rect 6403 15392 6461 15393
rect 17644 15392 17684 15520
rect 19075 15476 19133 15477
rect 20428 15476 20468 15520
rect 18883 15436 18892 15476
rect 18932 15436 19084 15476
rect 19124 15436 20468 15476
rect 21763 15436 21772 15476
rect 21812 15436 22156 15476
rect 22196 15436 22205 15476
rect 27811 15436 27820 15476
rect 27860 15436 29876 15476
rect 19075 15435 19133 15436
rect 29731 15392 29789 15393
rect 6403 15352 6412 15392
rect 6452 15352 6700 15392
rect 6740 15352 6749 15392
rect 17644 15352 19412 15392
rect 19459 15352 19468 15392
rect 19508 15352 20812 15392
rect 20852 15352 20861 15392
rect 27148 15352 28396 15392
rect 28436 15352 28445 15392
rect 28675 15352 28684 15392
rect 28724 15352 29164 15392
rect 29204 15352 29213 15392
rect 29646 15352 29740 15392
rect 29780 15352 29789 15392
rect 6403 15351 6461 15352
rect 19372 15309 19412 15352
rect 19363 15308 19421 15309
rect 2371 15268 2380 15308
rect 2420 15268 4204 15308
rect 4244 15268 4253 15308
rect 6307 15268 6316 15308
rect 6356 15268 6365 15308
rect 11107 15268 11116 15308
rect 11156 15268 12556 15308
rect 12596 15268 12605 15308
rect 13219 15268 13228 15308
rect 13268 15268 14956 15308
rect 14996 15268 15005 15308
rect 18691 15268 18700 15308
rect 18740 15268 18988 15308
rect 19028 15268 19037 15308
rect 19278 15268 19372 15308
rect 19412 15268 19756 15308
rect 19796 15268 21524 15308
rect 22243 15268 22252 15308
rect 22292 15268 22301 15308
rect 23683 15268 23692 15308
rect 23732 15268 26764 15308
rect 26804 15268 26813 15308
rect 6316 15224 6356 15268
rect 19363 15267 19421 15268
rect 20131 15224 20189 15225
rect 1603 15184 1612 15224
rect 1652 15184 3764 15224
rect 3811 15184 3820 15224
rect 3860 15184 5164 15224
rect 5204 15184 6124 15224
rect 6164 15184 6356 15224
rect 18892 15184 19948 15224
rect 19988 15184 20140 15224
rect 20180 15184 20189 15224
rect 3724 15140 3764 15184
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 3724 15100 4012 15140
rect 4052 15100 4061 15140
rect 4771 15100 4780 15140
rect 4820 15100 5644 15140
rect 5684 15100 5693 15140
rect 6412 15100 7180 15140
rect 7220 15100 7229 15140
rect 11491 15100 11500 15140
rect 11540 15100 11980 15140
rect 12020 15100 12029 15140
rect 15427 15100 15436 15140
rect 15476 15100 16492 15140
rect 16532 15100 16541 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 5443 15016 5452 15056
rect 5492 15016 5501 15056
rect 5452 14972 5492 15016
rect 6412 14972 6452 15100
rect 18892 15056 18932 15184
rect 20131 15183 20189 15184
rect 20620 15184 21388 15224
rect 21428 15184 21437 15224
rect 20620 15140 20660 15184
rect 19267 15100 19276 15140
rect 19316 15100 19756 15140
rect 19796 15100 19805 15140
rect 20580 15100 20620 15140
rect 20660 15100 20669 15140
rect 13219 15016 13228 15056
rect 13268 15016 14764 15056
rect 14804 15016 15724 15056
rect 15764 15016 15773 15056
rect 17635 15016 17644 15056
rect 17684 15016 18932 15056
rect 20035 15056 20093 15057
rect 21484 15056 21524 15268
rect 22252 15224 22292 15268
rect 27148 15224 27188 15352
rect 29731 15351 29789 15352
rect 29836 15308 29876 15436
rect 30316 15392 30356 15520
rect 34339 15519 34397 15520
rect 32524 15436 34060 15476
rect 34100 15436 36940 15476
rect 36980 15436 36989 15476
rect 29923 15352 29932 15392
rect 29972 15352 30220 15392
rect 30260 15352 30269 15392
rect 30316 15352 30700 15392
rect 30740 15352 30749 15392
rect 32524 15308 32564 15436
rect 32611 15352 32620 15392
rect 32660 15352 37996 15392
rect 38036 15352 38045 15392
rect 27427 15268 27436 15308
rect 27476 15268 28972 15308
rect 29012 15268 29021 15308
rect 29836 15268 32564 15308
rect 33379 15268 33388 15308
rect 33428 15268 34252 15308
rect 34292 15268 34301 15308
rect 22252 15184 27188 15224
rect 27244 15184 29012 15224
rect 29731 15184 29740 15224
rect 29780 15184 30892 15224
rect 30932 15184 30941 15224
rect 32803 15184 32812 15224
rect 32852 15184 33812 15224
rect 35971 15184 35980 15224
rect 36020 15184 36844 15224
rect 36884 15184 36893 15224
rect 27244 15140 27284 15184
rect 28867 15140 28925 15141
rect 27204 15100 27244 15140
rect 27284 15100 27293 15140
rect 28782 15100 28876 15140
rect 28916 15100 28925 15140
rect 28867 15099 28925 15100
rect 28972 15056 29012 15184
rect 29443 15100 29452 15140
rect 29492 15100 30412 15140
rect 30452 15100 30461 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 33772 15056 33812 15184
rect 33859 15100 33868 15140
rect 33908 15100 34156 15140
rect 34196 15100 34205 15140
rect 34819 15100 34828 15140
rect 34868 15100 36748 15140
rect 36788 15100 36797 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 20035 15016 20044 15056
rect 20084 15016 21428 15056
rect 21484 15016 22924 15056
rect 22964 15016 22973 15056
rect 23971 15016 23980 15056
rect 24020 15016 24940 15056
rect 24980 15016 24989 15056
rect 28972 15016 29836 15056
rect 29876 15016 30316 15056
rect 30356 15016 30365 15056
rect 30787 15016 30796 15056
rect 30836 15016 32140 15056
rect 32180 15016 32189 15056
rect 33772 15016 33908 15056
rect 20035 15015 20093 15016
rect 21388 14972 21428 15016
rect 33868 14972 33908 15016
rect 3523 14932 3532 14972
rect 3572 14932 5356 14972
rect 5396 14932 5405 14972
rect 5452 14932 5644 14972
rect 5684 14932 5693 14972
rect 6403 14932 6412 14972
rect 6452 14932 6461 14972
rect 12259 14932 12268 14972
rect 12308 14932 13804 14972
rect 13844 14932 14860 14972
rect 14900 14932 14909 14972
rect 18595 14932 18604 14972
rect 18644 14932 20716 14972
rect 20756 14932 21292 14972
rect 21332 14932 21341 14972
rect 21388 14932 27052 14972
rect 27092 14932 27101 14972
rect 28771 14932 28780 14972
rect 28820 14932 28829 14972
rect 30883 14932 30892 14972
rect 30932 14932 31276 14972
rect 31316 14932 31756 14972
rect 31796 14932 31805 14972
rect 33859 14932 33868 14972
rect 33908 14932 33917 14972
rect 37603 14932 37612 14972
rect 37652 14932 37804 14972
rect 37844 14932 37853 14972
rect 0 14888 80 14908
rect 28780 14888 28820 14932
rect 32899 14888 32957 14889
rect 0 14848 1036 14888
rect 1076 14848 1085 14888
rect 5251 14848 5260 14888
rect 5300 14848 8236 14888
rect 8276 14848 8285 14888
rect 9859 14848 9868 14888
rect 9908 14848 11884 14888
rect 11924 14848 11933 14888
rect 12835 14848 12844 14888
rect 12884 14848 14092 14888
rect 14132 14848 14141 14888
rect 16675 14848 16684 14888
rect 16724 14848 18988 14888
rect 19028 14848 19037 14888
rect 19171 14848 19180 14888
rect 19220 14848 21580 14888
rect 21620 14848 25132 14888
rect 25172 14848 25181 14888
rect 26764 14848 26956 14888
rect 26996 14848 27340 14888
rect 27380 14848 27389 14888
rect 28003 14848 28012 14888
rect 28052 14848 28588 14888
rect 28628 14848 28637 14888
rect 28780 14848 29876 14888
rect 29923 14848 29932 14888
rect 29972 14848 31084 14888
rect 31124 14848 31133 14888
rect 32803 14848 32812 14888
rect 32852 14848 32908 14888
rect 32948 14848 32957 14888
rect 33091 14848 33100 14888
rect 33140 14848 34636 14888
rect 34676 14848 34685 14888
rect 36931 14848 36940 14888
rect 36980 14848 37900 14888
rect 37940 14848 37949 14888
rect 38371 14848 38380 14888
rect 38420 14848 38956 14888
rect 38996 14848 39005 14888
rect 39715 14848 39724 14888
rect 39764 14848 40972 14888
rect 41012 14848 41021 14888
rect 44419 14848 44428 14888
rect 44468 14848 44477 14888
rect 0 14828 80 14848
rect 23971 14804 24029 14805
rect 19660 14764 19852 14804
rect 19892 14764 19901 14804
rect 20131 14764 20140 14804
rect 20180 14764 20620 14804
rect 20660 14764 20669 14804
rect 22339 14764 22348 14804
rect 22388 14764 23116 14804
rect 23156 14764 23165 14804
rect 23971 14764 23980 14804
rect 24020 14764 24748 14804
rect 24788 14764 24797 14804
rect 12835 14720 12893 14721
rect 931 14680 940 14720
rect 980 14680 2764 14720
rect 2804 14680 2813 14720
rect 3619 14680 3628 14720
rect 3668 14680 7084 14720
rect 7124 14680 7133 14720
rect 10051 14680 10060 14720
rect 10100 14680 10924 14720
rect 10964 14680 11308 14720
rect 11348 14680 11357 14720
rect 12750 14680 12844 14720
rect 12884 14680 12893 14720
rect 14275 14680 14284 14720
rect 14324 14680 15724 14720
rect 15764 14680 15773 14720
rect 16291 14680 16300 14720
rect 16340 14680 16684 14720
rect 16724 14680 16972 14720
rect 17012 14680 17021 14720
rect 17539 14680 17548 14720
rect 17588 14680 18508 14720
rect 18548 14680 18700 14720
rect 18740 14680 18749 14720
rect 18883 14680 18892 14720
rect 18932 14680 19372 14720
rect 19412 14680 19421 14720
rect 12835 14679 12893 14680
rect 19660 14636 19700 14764
rect 23971 14763 24029 14764
rect 19939 14680 19948 14720
rect 19988 14680 19997 14720
rect 20419 14680 20428 14720
rect 20468 14680 21484 14720
rect 21524 14680 21533 14720
rect 22435 14680 22444 14720
rect 22484 14680 22493 14720
rect 23587 14680 23596 14720
rect 23636 14680 24076 14720
rect 24116 14680 24125 14720
rect 24643 14680 24652 14720
rect 24692 14680 24940 14720
rect 24980 14680 26188 14720
rect 26228 14680 26237 14720
rect 19948 14636 19988 14680
rect 22444 14636 22484 14680
rect 15331 14596 15340 14636
rect 15380 14596 15820 14636
rect 15860 14596 15869 14636
rect 19075 14596 19084 14636
rect 19124 14596 19700 14636
rect 19852 14596 19988 14636
rect 21187 14596 21196 14636
rect 21236 14596 21868 14636
rect 21908 14596 22484 14636
rect 22531 14636 22589 14637
rect 26764 14636 26804 14848
rect 29836 14804 29876 14848
rect 32899 14847 32957 14848
rect 33100 14804 33140 14848
rect 44428 14804 44468 14848
rect 26851 14764 26860 14804
rect 26900 14764 28780 14804
rect 28820 14764 29163 14804
rect 29203 14764 29212 14804
rect 29827 14764 29836 14804
rect 29876 14764 29885 14804
rect 30892 14764 33140 14804
rect 33187 14764 33196 14804
rect 33236 14764 34060 14804
rect 34100 14764 34109 14804
rect 37507 14764 37516 14804
rect 37556 14764 38188 14804
rect 38228 14764 41260 14804
rect 41300 14764 42124 14804
rect 42164 14764 44620 14804
rect 44660 14764 44669 14804
rect 30892 14720 30932 14764
rect 26947 14680 26956 14720
rect 26996 14680 27820 14720
rect 27860 14680 27869 14720
rect 28675 14680 28684 14720
rect 28724 14680 29260 14720
rect 29300 14680 29309 14720
rect 29635 14680 29644 14720
rect 29684 14680 30892 14720
rect 30932 14680 30941 14720
rect 32131 14680 32140 14720
rect 32180 14680 34732 14720
rect 34772 14680 34781 14720
rect 40483 14680 40492 14720
rect 40532 14680 42988 14720
rect 43028 14680 43037 14720
rect 22531 14596 22540 14636
rect 22580 14596 26804 14636
rect 27715 14596 27724 14636
rect 27764 14596 28204 14636
rect 28244 14596 28253 14636
rect 30499 14596 30508 14636
rect 30548 14596 33676 14636
rect 33716 14596 33725 14636
rect 5155 14552 5213 14553
rect 5155 14512 5164 14552
rect 5204 14512 5548 14552
rect 5588 14512 5597 14552
rect 5155 14511 5213 14512
rect 19852 14468 19892 14596
rect 22531 14595 22589 14596
rect 23971 14552 24029 14553
rect 40867 14552 40925 14553
rect 19939 14512 19948 14552
rect 19988 14512 20620 14552
rect 20660 14512 20669 14552
rect 22051 14512 22060 14552
rect 22100 14512 22348 14552
rect 22388 14512 22397 14552
rect 22915 14512 22924 14552
rect 22964 14512 23788 14552
rect 23828 14512 23980 14552
rect 24020 14512 24029 14552
rect 24163 14512 24172 14552
rect 24212 14512 25324 14552
rect 25364 14512 26092 14552
rect 26132 14512 27532 14552
rect 27572 14512 28108 14552
rect 28148 14512 28157 14552
rect 28963 14512 28972 14552
rect 29012 14512 29356 14552
rect 29396 14512 29405 14552
rect 31459 14512 31468 14552
rect 31508 14512 31948 14552
rect 31988 14512 32716 14552
rect 32756 14512 32765 14552
rect 32899 14512 32908 14552
rect 32948 14512 33292 14552
rect 33332 14512 33341 14552
rect 33475 14512 33484 14552
rect 33524 14512 37612 14552
rect 37652 14512 37661 14552
rect 40675 14512 40684 14552
rect 40724 14512 40876 14552
rect 40916 14512 40925 14552
rect 23971 14511 24029 14512
rect 40867 14511 40925 14512
rect 18787 14428 18796 14468
rect 18836 14428 19276 14468
rect 19316 14428 19325 14468
rect 19852 14428 19988 14468
rect 20995 14428 21004 14468
rect 21044 14428 21772 14468
rect 21812 14428 22252 14468
rect 22292 14428 22301 14468
rect 23920 14428 23980 14468
rect 24020 14428 25804 14468
rect 25844 14428 25853 14468
rect 25900 14428 30796 14468
rect 30836 14428 30845 14468
rect 32131 14428 32140 14468
rect 32180 14428 34060 14468
rect 34100 14428 34109 14468
rect 19948 14384 19988 14428
rect 23920 14384 23960 14428
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 5347 14344 5356 14384
rect 5396 14344 6604 14384
rect 6644 14344 7756 14384
rect 7796 14344 7805 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 19948 14344 23960 14384
rect 4003 14260 4012 14300
rect 4052 14260 8908 14300
rect 8948 14260 8957 14300
rect 4771 14216 4829 14217
rect 19363 14216 19421 14217
rect 19948 14216 19988 14344
rect 20035 14260 20044 14300
rect 20084 14260 21964 14300
rect 22004 14260 22636 14300
rect 22676 14260 22685 14300
rect 21091 14216 21149 14217
rect 25900 14216 25940 14428
rect 28867 14384 28925 14385
rect 35011 14384 35069 14385
rect 28782 14344 28876 14384
rect 28916 14344 28925 14384
rect 31747 14344 31756 14384
rect 31796 14344 32908 14384
rect 32948 14344 32957 14384
rect 33000 14344 33009 14384
rect 33049 14344 33868 14384
rect 33908 14344 33917 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 35011 14344 35020 14384
rect 35060 14344 35116 14384
rect 35156 14344 39724 14384
rect 39764 14344 39773 14384
rect 44227 14344 44236 14384
rect 44276 14344 44285 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 28867 14343 28925 14344
rect 35011 14343 35069 14344
rect 26083 14260 26092 14300
rect 26132 14260 29000 14300
rect 31939 14260 31948 14300
rect 31988 14260 33676 14300
rect 33716 14260 34156 14300
rect 34196 14260 38324 14300
rect 4099 14176 4108 14216
rect 4148 14176 4492 14216
rect 4532 14176 4541 14216
rect 4675 14176 4684 14216
rect 4724 14176 4780 14216
rect 4820 14176 4829 14216
rect 8611 14176 8620 14216
rect 8660 14176 9772 14216
rect 9812 14176 10444 14216
rect 10484 14176 10493 14216
rect 16483 14176 16492 14216
rect 16532 14176 17164 14216
rect 17204 14176 17644 14216
rect 17684 14176 17693 14216
rect 18403 14176 18412 14216
rect 18452 14176 18988 14216
rect 19028 14176 19037 14216
rect 19363 14176 19372 14216
rect 19412 14176 19660 14216
rect 19700 14176 19709 14216
rect 19939 14176 19948 14216
rect 19988 14176 19997 14216
rect 21006 14176 21100 14216
rect 21140 14176 21149 14216
rect 4771 14175 4829 14176
rect 19363 14175 19421 14176
rect 21091 14175 21149 14176
rect 23920 14176 25940 14216
rect 28960 14216 29000 14260
rect 38284 14216 38324 14260
rect 28960 14176 29932 14216
rect 29972 14176 31316 14216
rect 20035 14132 20093 14133
rect 1315 14092 1324 14132
rect 1364 14092 2540 14132
rect 0 14048 80 14068
rect 2500 14048 2540 14092
rect 5740 14092 9004 14132
rect 9044 14092 9053 14132
rect 11491 14092 11500 14132
rect 11540 14092 13804 14132
rect 13844 14092 13853 14132
rect 15235 14092 15244 14132
rect 15284 14092 15820 14132
rect 15860 14092 15869 14132
rect 18691 14092 18700 14132
rect 18740 14092 20044 14132
rect 20084 14092 20093 14132
rect 20707 14092 20716 14132
rect 20756 14092 21676 14132
rect 21716 14092 22924 14132
rect 22964 14092 22973 14132
rect 5740 14048 5780 14092
rect 20035 14091 20093 14092
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 2500 14008 5068 14048
rect 5108 14008 5452 14048
rect 5492 14008 5501 14048
rect 5731 14008 5740 14048
rect 5780 14008 5789 14048
rect 7843 14008 7852 14048
rect 7892 14008 8044 14048
rect 8084 14008 13228 14048
rect 13268 14008 13277 14048
rect 14755 14008 14764 14048
rect 14804 14008 15724 14048
rect 15764 14008 15773 14048
rect 16195 14008 16204 14048
rect 16244 14008 17068 14048
rect 17108 14008 17452 14048
rect 17492 14008 17501 14048
rect 17923 14008 17932 14048
rect 17972 14008 18604 14048
rect 18644 14008 18653 14048
rect 19171 14008 19180 14048
rect 19220 14008 19372 14048
rect 19412 14008 21388 14048
rect 21428 14008 23500 14048
rect 23540 14008 23549 14048
rect 0 13988 80 14008
rect 4204 13964 4244 14008
rect 22531 13964 22589 13965
rect 4195 13924 4204 13964
rect 4244 13924 4253 13964
rect 5251 13924 5260 13964
rect 5300 13924 6508 13964
rect 6548 13924 6557 13964
rect 12460 13924 12556 13964
rect 12596 13924 12605 13964
rect 17155 13924 17164 13964
rect 17204 13924 18124 13964
rect 18164 13924 19796 13964
rect 20419 13924 20428 13964
rect 20468 13924 21868 13964
rect 21908 13924 21917 13964
rect 22243 13924 22252 13964
rect 22292 13924 22540 13964
rect 22580 13924 22589 13964
rect 12460 13880 12500 13924
rect 19756 13880 19796 13924
rect 22531 13923 22589 13924
rect 23920 13880 23960 14176
rect 25507 14132 25565 14133
rect 25422 14092 25516 14132
rect 25556 14092 26956 14132
rect 26996 14092 27005 14132
rect 27427 14092 27436 14132
rect 27476 14092 29740 14132
rect 29780 14092 29789 14132
rect 25507 14091 25565 14092
rect 27619 14008 27628 14048
rect 27668 14008 28300 14048
rect 28340 14008 28349 14048
rect 30403 14008 30412 14048
rect 30452 14008 30700 14048
rect 30740 14008 30749 14048
rect 31276 13964 31316 14176
rect 31756 14176 33388 14216
rect 33428 14176 33437 14216
rect 38275 14176 38284 14216
rect 38324 14176 41068 14216
rect 41108 14176 41836 14216
rect 41876 14176 41885 14216
rect 31756 14049 31796 14176
rect 44236 14132 44276 14344
rect 32227 14092 32236 14132
rect 32276 14092 33580 14132
rect 33620 14092 33629 14132
rect 34051 14092 34060 14132
rect 34100 14092 34252 14132
rect 34292 14092 36884 14132
rect 37987 14092 37996 14132
rect 38036 14092 38572 14132
rect 38612 14092 44276 14132
rect 31747 14048 31805 14049
rect 32707 14048 32765 14049
rect 36844 14048 36884 14092
rect 31662 14008 31756 14048
rect 31796 14008 31805 14048
rect 31747 14007 31805 14008
rect 31852 14008 32524 14048
rect 32564 14008 32573 14048
rect 32707 14008 32716 14048
rect 32756 14008 32850 14048
rect 32995 14008 33004 14048
rect 33044 14008 33388 14048
rect 33428 14008 35404 14048
rect 35444 14008 35884 14048
rect 35924 14008 35933 14048
rect 36163 14008 36172 14048
rect 36212 14008 36652 14048
rect 36692 14008 36701 14048
rect 36835 14008 36844 14048
rect 36884 14008 38804 14048
rect 38851 14008 38860 14048
rect 38900 14008 39628 14048
rect 39668 14008 39677 14048
rect 41347 14008 41356 14048
rect 41396 14008 41932 14048
rect 41972 14008 41981 14048
rect 43267 14008 43276 14048
rect 43316 14008 44140 14048
rect 44180 14008 44189 14048
rect 31852 13964 31892 14008
rect 32707 14007 32765 14008
rect 35884 13964 35924 14008
rect 38764 13964 38804 14008
rect 25891 13924 25900 13964
rect 25940 13924 27436 13964
rect 27476 13924 27820 13964
rect 27860 13924 27869 13964
rect 28099 13924 28108 13964
rect 28148 13924 29836 13964
rect 29876 13924 29885 13964
rect 31276 13924 31892 13964
rect 32035 13924 32044 13964
rect 32084 13924 33484 13964
rect 33524 13924 33533 13964
rect 33763 13924 33772 13964
rect 33812 13924 33821 13964
rect 35884 13924 38668 13964
rect 38708 13924 38717 13964
rect 38764 13924 40972 13964
rect 41012 13924 41740 13964
rect 41780 13924 42836 13964
rect 26476 13880 26516 13924
rect 30019 13880 30077 13881
rect 30691 13880 30749 13881
rect 33772 13880 33812 13924
rect 42796 13880 42836 13924
rect 3811 13840 3820 13880
rect 3860 13840 6124 13880
rect 6164 13840 6173 13880
rect 8803 13840 8812 13880
rect 8852 13840 10156 13880
rect 10196 13840 10205 13880
rect 12451 13840 12460 13880
rect 12500 13840 12509 13880
rect 12556 13840 13132 13880
rect 13172 13840 13181 13880
rect 18499 13840 18508 13880
rect 18548 13840 18700 13880
rect 18740 13840 19084 13880
rect 19124 13840 19133 13880
rect 19756 13840 19892 13880
rect 19939 13840 19948 13880
rect 19988 13840 21105 13880
rect 21145 13840 21388 13880
rect 21428 13840 21437 13880
rect 21571 13840 21580 13880
rect 21620 13840 23960 13880
rect 26467 13840 26476 13880
rect 26516 13840 26525 13880
rect 29934 13840 30028 13880
rect 30068 13840 30077 13880
rect 30499 13840 30508 13880
rect 30548 13840 30700 13880
rect 30740 13840 30749 13880
rect 32323 13840 32332 13880
rect 32372 13840 33812 13880
rect 35203 13840 35212 13880
rect 35252 13840 36556 13880
rect 36596 13840 36605 13880
rect 42019 13840 42028 13880
rect 42068 13840 42508 13880
rect 42548 13840 42557 13880
rect 42787 13840 42796 13880
rect 42836 13840 45676 13880
rect 45716 13840 45725 13880
rect 12556 13796 12596 13840
rect 19852 13796 19892 13840
rect 30019 13839 30077 13840
rect 30691 13839 30749 13840
rect 12547 13756 12556 13796
rect 12596 13756 12605 13796
rect 19852 13756 20908 13796
rect 20948 13756 20957 13796
rect 27235 13756 27244 13796
rect 27284 13756 27532 13796
rect 27572 13756 27581 13796
rect 27907 13756 27916 13796
rect 27956 13756 28108 13796
rect 28148 13756 28157 13796
rect 31075 13756 31084 13796
rect 31124 13756 32236 13796
rect 32276 13756 32285 13796
rect 32995 13756 33004 13796
rect 33044 13756 34924 13796
rect 34964 13756 36652 13796
rect 36692 13756 36701 13796
rect 37603 13756 37612 13796
rect 37652 13756 39052 13796
rect 39092 13756 39101 13796
rect 30595 13712 30653 13713
rect 12355 13672 12364 13712
rect 12404 13672 12748 13712
rect 12788 13672 12797 13712
rect 20323 13672 20332 13712
rect 20372 13672 20812 13712
rect 20852 13672 21100 13712
rect 21140 13672 21149 13712
rect 30211 13672 30220 13712
rect 30260 13672 30604 13712
rect 30644 13672 30653 13712
rect 32515 13672 32524 13712
rect 32564 13672 33196 13712
rect 33236 13672 33245 13712
rect 30595 13671 30653 13672
rect 32899 13628 32957 13629
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 30787 13588 30796 13628
rect 30836 13588 31796 13628
rect 32814 13588 32908 13628
rect 32948 13588 32957 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 31651 13544 31709 13545
rect 31566 13504 31660 13544
rect 31700 13504 31709 13544
rect 31756 13544 31796 13588
rect 32899 13587 32957 13588
rect 31756 13504 34444 13544
rect 34484 13504 34493 13544
rect 31651 13503 31709 13504
rect 18883 13420 18892 13460
rect 18932 13420 19468 13460
rect 19508 13420 19517 13460
rect 20515 13420 20524 13460
rect 20564 13420 20756 13460
rect 30115 13420 30124 13460
rect 30164 13420 37324 13460
rect 37364 13420 37373 13460
rect 5347 13336 5356 13376
rect 5396 13336 6220 13376
rect 6260 13336 6269 13376
rect 12931 13336 12940 13376
rect 12980 13336 16204 13376
rect 16244 13336 16253 13376
rect 19075 13336 19084 13376
rect 19124 13336 19948 13376
rect 19988 13336 19997 13376
rect 20044 13336 20140 13376
rect 20180 13336 20189 13376
rect 5827 13252 5836 13292
rect 5876 13252 6892 13292
rect 6932 13252 6941 13292
rect 16675 13252 16684 13292
rect 16724 13252 17644 13292
rect 17684 13252 19756 13292
rect 19796 13252 19805 13292
rect 0 13208 80 13228
rect 18691 13208 18749 13209
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 3619 13168 3628 13208
rect 3668 13168 5548 13208
rect 5588 13168 5597 13208
rect 6691 13168 6700 13208
rect 6740 13168 8044 13208
rect 8084 13168 8093 13208
rect 9283 13168 9292 13208
rect 9332 13168 10060 13208
rect 10100 13168 10109 13208
rect 11971 13168 11980 13208
rect 12020 13168 12844 13208
rect 12884 13168 12893 13208
rect 16867 13168 16876 13208
rect 16916 13168 17356 13208
rect 17396 13168 18412 13208
rect 18452 13168 18461 13208
rect 18606 13168 18700 13208
rect 18740 13168 18749 13208
rect 0 13148 80 13168
rect 2947 13000 2956 13040
rect 2996 13000 4300 13040
rect 4340 13000 4349 13040
rect 5644 13000 10252 13040
rect 10292 13000 11212 13040
rect 11252 13000 11261 13040
rect 11683 13000 11692 13040
rect 11732 13000 12460 13040
rect 12500 13000 14092 13040
rect 14132 13000 14141 13040
rect 5644 12956 5684 13000
rect 18412 12956 18452 13168
rect 18691 13167 18749 13168
rect 20044 12956 20084 13336
rect 20716 13292 20756 13420
rect 20899 13336 20908 13376
rect 20948 13336 21388 13376
rect 21428 13336 21437 13376
rect 23683 13336 23692 13376
rect 23732 13336 23741 13376
rect 29347 13336 29356 13376
rect 29396 13336 33620 13376
rect 34435 13336 34444 13376
rect 34484 13336 37036 13376
rect 37076 13336 37085 13376
rect 42403 13336 42412 13376
rect 42452 13336 43180 13376
rect 43220 13336 43229 13376
rect 23692 13292 23732 13336
rect 20707 13252 20716 13292
rect 20756 13252 29068 13292
rect 29108 13252 29117 13292
rect 30787 13252 30796 13292
rect 30836 13252 30845 13292
rect 32035 13252 32044 13292
rect 32084 13252 33100 13292
rect 33140 13252 33149 13292
rect 23971 13208 24029 13209
rect 30595 13208 30653 13209
rect 22435 13168 22444 13208
rect 22484 13168 23020 13208
rect 23060 13168 23069 13208
rect 23299 13168 23308 13208
rect 23348 13168 23980 13208
rect 24020 13168 24029 13208
rect 27811 13168 27820 13208
rect 27860 13168 28492 13208
rect 28532 13168 28541 13208
rect 28675 13168 28684 13208
rect 28724 13168 30305 13208
rect 30345 13168 30354 13208
rect 30510 13168 30604 13208
rect 30644 13168 30653 13208
rect 23971 13167 24029 13168
rect 30595 13167 30653 13168
rect 30796 13124 30836 13252
rect 33580 13208 33620 13336
rect 34828 13252 36172 13292
rect 36212 13252 36221 13292
rect 34828 13208 34868 13252
rect 31747 13168 31756 13208
rect 31796 13168 32236 13208
rect 32276 13168 32285 13208
rect 32803 13168 32812 13208
rect 32852 13168 32861 13208
rect 33571 13168 33580 13208
rect 33620 13168 33868 13208
rect 33908 13168 33917 13208
rect 34339 13168 34348 13208
rect 34388 13168 34828 13208
rect 34868 13168 34877 13208
rect 35203 13168 35212 13208
rect 35252 13168 35692 13208
rect 35732 13168 35741 13208
rect 36451 13168 36460 13208
rect 36500 13168 36940 13208
rect 36980 13168 36989 13208
rect 37315 13168 37324 13208
rect 37364 13168 37804 13208
rect 37844 13168 37853 13208
rect 42019 13168 42028 13208
rect 42068 13168 42508 13208
rect 42548 13168 42557 13208
rect 43843 13168 43852 13208
rect 43892 13168 44428 13208
rect 44468 13168 44477 13208
rect 22915 13084 22924 13124
rect 22964 13084 24268 13124
rect 24308 13084 24652 13124
rect 24692 13084 24701 13124
rect 26083 13084 26092 13124
rect 26132 13084 30836 13124
rect 31843 13124 31901 13125
rect 32812 13124 32852 13168
rect 31843 13084 31852 13124
rect 31892 13084 32332 13124
rect 32372 13084 32852 13124
rect 33868 13124 33908 13168
rect 33868 13084 34924 13124
rect 34964 13084 34973 13124
rect 35491 13084 35500 13124
rect 35540 13084 36364 13124
rect 36404 13084 36413 13124
rect 31843 13083 31901 13084
rect 29731 13040 29789 13041
rect 34924 13040 34964 13084
rect 20131 13000 20140 13040
rect 20180 13000 20332 13040
rect 20372 13000 20381 13040
rect 29155 13000 29164 13040
rect 29204 13000 29548 13040
rect 29588 13000 29597 13040
rect 29731 13000 29740 13040
rect 29780 13000 29874 13040
rect 33859 13000 33868 13040
rect 33908 13000 34348 13040
rect 34388 13000 34397 13040
rect 34924 13000 35020 13040
rect 35060 13000 35069 13040
rect 35779 13000 35788 13040
rect 35828 13000 36076 13040
rect 36116 13000 36125 13040
rect 41731 13000 41740 13040
rect 41780 13000 42124 13040
rect 42164 13000 42173 13040
rect 29731 12999 29789 13000
rect 4003 12916 4012 12956
rect 4052 12916 5644 12956
rect 5684 12916 5693 12956
rect 8899 12916 8908 12956
rect 8948 12916 12940 12956
rect 12980 12916 12989 12956
rect 18412 12916 21100 12956
rect 21140 12916 21149 12956
rect 29443 12916 29452 12956
rect 29492 12916 30028 12956
rect 30068 12916 30077 12956
rect 30211 12916 30220 12956
rect 30260 12916 30796 12956
rect 30836 12916 30845 12956
rect 32419 12916 32428 12956
rect 32468 12916 41452 12956
rect 41492 12916 41501 12956
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 10147 12832 10156 12872
rect 10196 12832 11404 12872
rect 11444 12832 11453 12872
rect 17923 12832 17932 12872
rect 17972 12832 18220 12872
rect 18260 12832 18269 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 20035 12832 20044 12872
rect 20084 12832 20124 12872
rect 20227 12832 20236 12872
rect 20276 12832 20908 12872
rect 20948 12832 20957 12872
rect 27820 12832 28396 12872
rect 28436 12832 28445 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 20044 12788 20084 12832
rect 27619 12788 27677 12789
rect 27820 12788 27860 12832
rect 18115 12748 18124 12788
rect 18164 12748 18604 12788
rect 18644 12748 18653 12788
rect 19564 12748 20620 12788
rect 20660 12748 20669 12788
rect 26440 12748 27628 12788
rect 27668 12748 27764 12788
rect 27811 12748 27820 12788
rect 27860 12748 27869 12788
rect 28396 12748 31084 12788
rect 31124 12748 31133 12788
rect 31468 12748 32140 12788
rect 32180 12748 32564 12788
rect 19564 12704 19604 12748
rect 26440 12704 26480 12748
rect 27619 12747 27677 12748
rect 27724 12704 27764 12748
rect 28396 12704 28436 12748
rect 17932 12664 18316 12704
rect 18356 12664 19564 12704
rect 19604 12664 19613 12704
rect 20035 12664 20044 12704
rect 20084 12664 21676 12704
rect 21716 12664 21725 12704
rect 25603 12664 25612 12704
rect 25652 12664 26480 12704
rect 27619 12664 27628 12704
rect 27668 12664 27677 12704
rect 27724 12664 28436 12704
rect 28483 12664 28492 12704
rect 28532 12664 28780 12704
rect 28820 12664 28829 12704
rect 17932 12620 17972 12664
rect 3523 12580 3532 12620
rect 3572 12580 5644 12620
rect 5684 12580 5693 12620
rect 12067 12580 12076 12620
rect 12116 12580 12940 12620
rect 12980 12580 12989 12620
rect 13603 12580 13612 12620
rect 13652 12580 15340 12620
rect 15380 12580 15389 12620
rect 16387 12580 16396 12620
rect 16436 12580 17548 12620
rect 17588 12580 17740 12620
rect 17780 12580 17789 12620
rect 17836 12580 17972 12620
rect 18019 12620 18077 12621
rect 20227 12620 20285 12621
rect 23971 12620 24029 12621
rect 18019 12580 18028 12620
rect 18068 12580 18162 12620
rect 19363 12580 19372 12620
rect 19412 12580 20236 12620
rect 20276 12580 20285 12620
rect 20803 12580 20812 12620
rect 20852 12580 21292 12620
rect 21332 12580 21341 12620
rect 23971 12580 23980 12620
rect 24020 12580 27148 12620
rect 27188 12580 27197 12620
rect 17836 12536 17876 12580
rect 18019 12579 18077 12580
rect 20227 12579 20285 12580
rect 23971 12579 24029 12580
rect 18691 12536 18749 12537
rect 21763 12536 21821 12537
rect 27628 12536 27668 12664
rect 31468 12620 31508 12748
rect 31555 12664 31564 12704
rect 31604 12664 32428 12704
rect 32468 12664 32477 12704
rect 27715 12580 27724 12620
rect 27764 12580 28972 12620
rect 29012 12580 29021 12620
rect 30691 12580 30700 12620
rect 30740 12580 31508 12620
rect 32524 12620 32564 12748
rect 38764 12664 38956 12704
rect 38996 12664 39005 12704
rect 42499 12664 42508 12704
rect 42548 12664 42557 12704
rect 38764 12620 38804 12664
rect 42508 12620 42548 12664
rect 32524 12580 34252 12620
rect 34292 12580 34301 12620
rect 34435 12580 34444 12620
rect 34484 12580 34964 12620
rect 35011 12580 35020 12620
rect 35060 12580 35596 12620
rect 35636 12580 35645 12620
rect 37507 12580 37516 12620
rect 37556 12580 38188 12620
rect 38228 12580 38668 12620
rect 38708 12580 38804 12620
rect 38851 12580 38860 12620
rect 38900 12580 40684 12620
rect 40724 12580 40733 12620
rect 41827 12580 41836 12620
rect 41876 12580 43084 12620
rect 43124 12580 43133 12620
rect 43459 12580 43468 12620
rect 43508 12580 44236 12620
rect 44276 12580 44285 12620
rect 29539 12536 29597 12537
rect 8131 12496 8140 12536
rect 8180 12496 9004 12536
rect 9044 12496 9053 12536
rect 9667 12496 9676 12536
rect 9716 12496 10732 12536
rect 10772 12496 10781 12536
rect 11320 12496 11692 12536
rect 11732 12496 11741 12536
rect 16771 12496 16780 12536
rect 16820 12496 17876 12536
rect 17923 12496 17932 12536
rect 17972 12496 18700 12536
rect 18740 12496 18749 12536
rect 21678 12496 21772 12536
rect 21812 12496 22348 12536
rect 22388 12496 22397 12536
rect 26851 12496 26860 12536
rect 26900 12496 27340 12536
rect 27380 12496 27389 12536
rect 27628 12496 28492 12536
rect 28532 12496 28876 12536
rect 28916 12496 28925 12536
rect 29059 12496 29068 12536
rect 29108 12496 29548 12536
rect 29588 12496 29597 12536
rect 30787 12496 30796 12536
rect 30836 12496 31372 12536
rect 31412 12496 31421 12536
rect 31651 12496 31660 12536
rect 31700 12496 33196 12536
rect 33236 12496 33245 12536
rect 11320 12452 11360 12496
rect 18691 12495 18749 12496
rect 21763 12495 21821 12496
rect 29539 12495 29597 12496
rect 31660 12452 31700 12496
rect 9868 12412 11360 12452
rect 18211 12412 18220 12452
rect 18260 12412 18269 12452
rect 18499 12412 18508 12452
rect 18548 12412 19988 12452
rect 21091 12412 21100 12452
rect 21140 12412 21292 12452
rect 21332 12412 21341 12452
rect 27715 12412 27724 12452
rect 27764 12412 28108 12452
rect 28148 12412 28396 12452
rect 28436 12412 28445 12452
rect 28579 12412 28588 12452
rect 28628 12412 29356 12452
rect 29396 12412 29405 12452
rect 31267 12412 31276 12452
rect 31316 12412 31700 12452
rect 34924 12452 34964 12580
rect 37315 12496 37324 12536
rect 37364 12496 37996 12536
rect 38036 12496 38045 12536
rect 38755 12496 38764 12536
rect 38804 12496 39244 12536
rect 39284 12496 39293 12536
rect 41443 12496 41452 12536
rect 41492 12496 42700 12536
rect 42740 12496 42749 12536
rect 42979 12496 42988 12536
rect 43028 12496 45292 12536
rect 45332 12496 45676 12536
rect 45716 12496 45725 12536
rect 46723 12496 46732 12536
rect 46772 12496 47596 12536
rect 47636 12496 47645 12536
rect 34924 12412 35212 12452
rect 35252 12412 35261 12452
rect 37507 12412 37516 12452
rect 37556 12412 37565 12452
rect 37780 12412 40396 12452
rect 40436 12412 41932 12452
rect 41972 12412 43468 12452
rect 43508 12412 43517 12452
rect 0 12368 80 12388
rect 9868 12368 9908 12412
rect 11395 12368 11453 12369
rect 18220 12368 18260 12412
rect 19075 12368 19133 12369
rect 19948 12368 19988 12412
rect 37516 12368 37556 12412
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 9859 12328 9868 12368
rect 9908 12328 9917 12368
rect 11395 12328 11404 12368
rect 11444 12328 11538 12368
rect 16579 12328 16588 12368
rect 16628 12328 18260 12368
rect 18990 12328 19084 12368
rect 19124 12328 19133 12368
rect 19939 12328 19948 12368
rect 19988 12328 19997 12368
rect 20140 12328 21388 12368
rect 21428 12328 21437 12368
rect 21859 12328 21868 12368
rect 21908 12328 22252 12368
rect 22292 12328 26284 12368
rect 26324 12328 26333 12368
rect 29059 12328 29068 12368
rect 29108 12328 29260 12368
rect 29300 12328 29309 12368
rect 29827 12328 29836 12368
rect 29876 12328 37556 12368
rect 0 12308 80 12328
rect 11395 12327 11453 12328
rect 18220 12284 18260 12328
rect 19075 12327 19133 12328
rect 20140 12284 20180 12328
rect 23011 12284 23069 12285
rect 26179 12284 26237 12285
rect 37780 12284 37820 12412
rect 39427 12328 39436 12368
rect 39476 12328 41548 12368
rect 41588 12328 41836 12368
rect 41876 12328 41885 12368
rect 42115 12328 42124 12368
rect 42164 12328 42604 12368
rect 42644 12328 42653 12368
rect 42883 12328 42892 12368
rect 42932 12328 43564 12368
rect 43604 12328 43613 12368
rect 11299 12244 11308 12284
rect 11348 12244 11884 12284
rect 11924 12244 12268 12284
rect 12308 12244 12317 12284
rect 17443 12244 17452 12284
rect 17492 12244 18028 12284
rect 18068 12244 18077 12284
rect 18220 12244 19468 12284
rect 19508 12244 20180 12284
rect 20419 12244 20428 12284
rect 20468 12244 23020 12284
rect 23060 12244 23069 12284
rect 26094 12244 26188 12284
rect 26228 12244 26237 12284
rect 32515 12244 32524 12284
rect 32564 12244 34924 12284
rect 34964 12244 37820 12284
rect 38179 12244 38188 12284
rect 38228 12244 38956 12284
rect 38996 12244 39005 12284
rect 39235 12244 39244 12284
rect 39284 12244 42508 12284
rect 42548 12244 42557 12284
rect 42691 12244 42700 12284
rect 42740 12244 45100 12284
rect 45140 12244 45149 12284
rect 48643 12244 48652 12284
rect 48692 12244 48701 12284
rect 23011 12243 23069 12244
rect 26179 12243 26237 12244
rect 18019 12200 18077 12201
rect 31843 12200 31901 12201
rect 34147 12200 34205 12201
rect 48652 12200 48692 12244
rect 17731 12160 17740 12200
rect 17780 12160 18028 12200
rect 18068 12160 22156 12200
rect 22196 12160 22205 12200
rect 22339 12160 22348 12200
rect 22388 12160 28780 12200
rect 28820 12160 28829 12200
rect 31758 12160 31852 12200
rect 31892 12160 31901 12200
rect 34062 12160 34156 12200
rect 34196 12160 34205 12200
rect 37123 12160 37132 12200
rect 37172 12160 37612 12200
rect 37652 12160 37661 12200
rect 41560 12160 49324 12200
rect 49364 12160 49373 12200
rect 18019 12159 18077 12160
rect 31843 12159 31901 12160
rect 34147 12159 34205 12160
rect 30691 12116 30749 12117
rect 41560 12116 41600 12160
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 19171 12076 19180 12116
rect 19220 12076 20716 12116
rect 20756 12076 20765 12116
rect 25027 12076 25036 12116
rect 25076 12076 30508 12116
rect 30548 12076 30557 12116
rect 30691 12076 30700 12116
rect 30740 12076 30834 12116
rect 31555 12076 31564 12116
rect 31604 12076 32044 12116
rect 32084 12076 32093 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 36643 12076 36652 12116
rect 36692 12076 37228 12116
rect 37268 12076 41600 12116
rect 42019 12076 42028 12116
rect 42068 12076 42892 12116
rect 42932 12076 42941 12116
rect 43075 12076 43084 12116
rect 43124 12076 43948 12116
rect 43988 12076 43997 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 30691 12075 30749 12076
rect 20227 12032 20285 12033
rect 20142 11992 20236 12032
rect 20276 11992 20285 12032
rect 20227 11991 20285 11992
rect 20524 11992 20908 12032
rect 20948 11992 20957 12032
rect 26947 11992 26956 12032
rect 26996 11992 30796 12032
rect 30836 11992 30845 12032
rect 36931 11992 36940 12032
rect 36980 11992 37324 12032
rect 37364 11992 37373 12032
rect 42403 11992 42412 12032
rect 42452 11992 42700 12032
rect 42740 11992 42749 12032
rect 20524 11948 20564 11992
rect 31459 11948 31517 11949
rect 3715 11908 3724 11948
rect 3764 11908 3916 11948
rect 3956 11908 4492 11948
rect 4532 11908 6412 11948
rect 6452 11908 6461 11948
rect 7075 11908 7084 11948
rect 7124 11908 9772 11948
rect 9812 11908 9821 11948
rect 17731 11908 17740 11948
rect 17780 11908 20524 11948
rect 20564 11908 20573 11948
rect 24835 11908 24844 11948
rect 24884 11908 31468 11948
rect 31508 11908 31564 11948
rect 31604 11908 31632 11948
rect 32611 11908 32620 11948
rect 32660 11908 42028 11948
rect 42068 11908 42077 11948
rect 42211 11908 42220 11948
rect 42260 11908 44716 11948
rect 44756 11908 44765 11948
rect 31459 11907 31517 11908
rect 4003 11824 4012 11864
rect 4052 11824 4684 11864
rect 4724 11824 4733 11864
rect 8035 11824 8044 11864
rect 8084 11824 8908 11864
rect 8948 11824 8957 11864
rect 12163 11824 12172 11864
rect 12212 11824 14092 11864
rect 14132 11824 14141 11864
rect 16771 11824 16780 11864
rect 16820 11824 20908 11864
rect 20948 11824 21388 11864
rect 21428 11824 21437 11864
rect 27139 11824 27148 11864
rect 27188 11824 28876 11864
rect 28916 11824 28925 11864
rect 31651 11824 31660 11864
rect 31700 11824 31852 11864
rect 31892 11824 32332 11864
rect 32372 11824 32381 11864
rect 32995 11824 33004 11864
rect 33044 11824 34252 11864
rect 34292 11824 45772 11864
rect 45812 11824 46444 11864
rect 46484 11824 46493 11864
rect 14467 11780 14525 11781
rect 33004 11780 33044 11824
rect 4396 11740 5836 11780
rect 5876 11740 6220 11780
rect 6260 11740 6269 11780
rect 8803 11740 8812 11780
rect 8852 11740 9676 11780
rect 9716 11740 9725 11780
rect 10147 11740 10156 11780
rect 10196 11740 11116 11780
rect 11156 11740 11165 11780
rect 14382 11740 14476 11780
rect 14516 11740 14525 11780
rect 4396 11696 4436 11740
rect 14467 11739 14525 11740
rect 20236 11740 20620 11780
rect 20660 11740 20669 11780
rect 20768 11740 20777 11780
rect 20817 11740 21004 11780
rect 21044 11740 21053 11780
rect 21632 11740 21641 11780
rect 21681 11740 22156 11780
rect 22196 11740 22205 11780
rect 26851 11740 26860 11780
rect 26900 11740 28300 11780
rect 28340 11740 28349 11780
rect 30979 11740 30988 11780
rect 31028 11740 31372 11780
rect 31412 11740 33044 11780
rect 33283 11740 33292 11780
rect 33332 11740 37036 11780
rect 37076 11740 37085 11780
rect 42499 11740 42508 11780
rect 42548 11740 44812 11780
rect 44852 11740 46636 11780
rect 46676 11740 46685 11780
rect 11875 11696 11933 11697
rect 20236 11696 20276 11740
rect 26563 11696 26621 11697
rect 28003 11696 28061 11697
rect 3811 11656 3820 11696
rect 3860 11656 4396 11696
rect 4436 11656 4445 11696
rect 5731 11656 5740 11696
rect 5780 11656 6604 11696
rect 6644 11656 6653 11696
rect 8611 11656 8620 11696
rect 8660 11656 9388 11696
rect 9428 11656 9437 11696
rect 9955 11656 9964 11696
rect 10004 11656 10828 11696
rect 10868 11656 10877 11696
rect 11790 11656 11884 11696
rect 11924 11656 11933 11696
rect 13027 11656 13036 11696
rect 13076 11656 15532 11696
rect 15572 11656 15581 11696
rect 16099 11656 16108 11696
rect 16148 11656 17068 11696
rect 17108 11656 17117 11696
rect 17635 11656 17644 11696
rect 17684 11656 18316 11696
rect 18356 11656 18365 11696
rect 18787 11656 18796 11696
rect 18836 11656 20276 11696
rect 20323 11656 20332 11696
rect 20372 11656 21196 11696
rect 21236 11656 21245 11696
rect 23587 11656 23596 11696
rect 23636 11656 23980 11696
rect 24020 11656 24029 11696
rect 26563 11656 26572 11696
rect 26612 11656 26668 11696
rect 26708 11656 27340 11696
rect 27380 11656 27389 11696
rect 27918 11656 28012 11696
rect 28052 11656 28061 11696
rect 30403 11656 30412 11696
rect 30452 11656 31084 11696
rect 31124 11656 31133 11696
rect 32131 11656 32140 11696
rect 32180 11656 32908 11696
rect 32948 11656 32957 11696
rect 34915 11656 34924 11696
rect 34964 11656 35500 11696
rect 35540 11656 35549 11696
rect 37891 11656 37900 11696
rect 37940 11656 38764 11696
rect 38804 11656 39436 11696
rect 39476 11656 39485 11696
rect 40291 11656 40300 11696
rect 40340 11656 42124 11696
rect 42164 11656 42173 11696
rect 46531 11656 46540 11696
rect 46580 11656 47116 11696
rect 47156 11656 48844 11696
rect 48884 11656 48893 11696
rect 11875 11655 11933 11656
rect 17068 11612 17108 11656
rect 26563 11655 26621 11656
rect 28003 11655 28061 11656
rect 28012 11612 28052 11655
rect 32323 11612 32381 11613
rect 5539 11572 5548 11612
rect 5588 11572 8044 11612
rect 8084 11572 8428 11612
rect 8468 11572 8477 11612
rect 11395 11572 11404 11612
rect 11444 11572 13324 11612
rect 13364 11572 13373 11612
rect 17068 11572 22636 11612
rect 22676 11572 22685 11612
rect 26179 11572 26188 11612
rect 26228 11572 26572 11612
rect 26612 11572 27628 11612
rect 27668 11572 27677 11612
rect 28012 11572 31468 11612
rect 31508 11572 31948 11612
rect 31988 11572 31997 11612
rect 32227 11572 32236 11612
rect 32276 11572 32332 11612
rect 32372 11572 32381 11612
rect 32707 11572 32716 11612
rect 32756 11572 33388 11612
rect 33428 11572 33437 11612
rect 39715 11572 39724 11612
rect 39764 11572 40492 11612
rect 40532 11572 41740 11612
rect 41780 11572 41789 11612
rect 32323 11571 32381 11572
rect 0 11528 80 11548
rect 24451 11528 24509 11529
rect 33187 11528 33245 11529
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 6019 11488 6028 11528
rect 6068 11488 6700 11528
rect 6740 11488 6749 11528
rect 7939 11488 7948 11528
rect 7988 11488 9484 11528
rect 9524 11488 9533 11528
rect 12067 11488 12076 11528
rect 12116 11488 13228 11528
rect 13268 11488 13277 11528
rect 17059 11488 17068 11528
rect 17108 11488 19180 11528
rect 19220 11488 19229 11528
rect 19747 11488 19756 11528
rect 19796 11488 20716 11528
rect 20756 11488 20765 11528
rect 24366 11488 24460 11528
rect 24500 11488 24509 11528
rect 27523 11488 27532 11528
rect 27572 11488 28396 11528
rect 28436 11488 28445 11528
rect 29155 11488 29164 11528
rect 29204 11488 29452 11528
rect 29492 11488 32428 11528
rect 32468 11488 32812 11528
rect 32852 11488 32861 11528
rect 33187 11488 33196 11528
rect 33236 11488 33676 11528
rect 33716 11488 33725 11528
rect 33859 11488 33868 11528
rect 33908 11488 34636 11528
rect 34676 11488 34685 11528
rect 35020 11488 35980 11528
rect 36020 11488 36268 11528
rect 36308 11488 36652 11528
rect 36692 11488 36701 11528
rect 40675 11488 40684 11528
rect 40724 11488 41548 11528
rect 41588 11488 41597 11528
rect 0 11468 80 11488
rect 24451 11487 24509 11488
rect 33187 11487 33245 11488
rect 30403 11444 30461 11445
rect 32899 11444 32957 11445
rect 35020 11444 35060 11488
rect 8227 11404 8236 11444
rect 8276 11404 9964 11444
rect 10004 11404 10013 11444
rect 11779 11404 11788 11444
rect 11828 11404 12268 11444
rect 12308 11404 14284 11444
rect 14324 11404 14333 11444
rect 17347 11404 17356 11444
rect 17396 11404 18164 11444
rect 20515 11404 20524 11444
rect 20564 11404 21484 11444
rect 21524 11404 21533 11444
rect 23920 11404 25036 11444
rect 25076 11404 25085 11444
rect 28960 11404 29740 11444
rect 29780 11404 29789 11444
rect 30403 11404 30412 11444
rect 30452 11404 30796 11444
rect 30836 11404 30845 11444
rect 31075 11404 31084 11444
rect 31124 11404 31564 11444
rect 31604 11404 32524 11444
rect 32564 11404 32573 11444
rect 32899 11404 32908 11444
rect 32948 11404 35060 11444
rect 35116 11404 36556 11444
rect 36596 11404 37076 11444
rect 42211 11404 42220 11444
rect 42260 11404 46444 11444
rect 46484 11404 47980 11444
rect 48020 11404 48364 11444
rect 48404 11404 48413 11444
rect 9388 11360 9428 11404
rect 18124 11360 18164 11404
rect 20419 11360 20477 11361
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 9187 11320 9196 11360
rect 9236 11320 9245 11360
rect 9348 11320 9388 11360
rect 9428 11320 9437 11360
rect 17220 11320 17260 11360
rect 17300 11320 17309 11360
rect 18115 11320 18124 11360
rect 18164 11320 18173 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 20334 11320 20428 11360
rect 20468 11320 20477 11360
rect 9196 11276 9236 11320
rect 17260 11276 17300 11320
rect 20419 11319 20477 11320
rect 23920 11276 23960 11404
rect 28960 11276 29000 11404
rect 30403 11403 30461 11404
rect 32899 11403 32957 11404
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 35116 11276 35156 11404
rect 36163 11360 36221 11361
rect 36078 11320 36172 11360
rect 36212 11320 36221 11360
rect 36163 11319 36221 11320
rect 8323 11236 8332 11276
rect 8372 11236 8716 11276
rect 8756 11236 8765 11276
rect 9196 11236 9580 11276
rect 9620 11236 9629 11276
rect 17260 11236 17644 11276
rect 17684 11236 19276 11276
rect 19316 11236 19325 11276
rect 21283 11236 21292 11276
rect 21332 11236 23500 11276
rect 23540 11236 23549 11276
rect 23596 11236 23960 11276
rect 24163 11236 24172 11276
rect 24212 11236 29000 11276
rect 29155 11236 29164 11276
rect 29204 11236 32332 11276
rect 32372 11236 33140 11276
rect 33187 11236 33196 11276
rect 33236 11236 33868 11276
rect 33908 11236 35156 11276
rect 18595 11192 18653 11193
rect 23596 11192 23636 11236
rect 33100 11192 33140 11236
rect 34243 11192 34301 11193
rect 3619 11152 3628 11192
rect 3668 11152 4684 11192
rect 4724 11152 5548 11192
rect 5588 11152 5597 11192
rect 7843 11152 7852 11192
rect 7892 11152 9100 11192
rect 9140 11152 9149 11192
rect 11299 11152 11308 11192
rect 11348 11152 12172 11192
rect 12212 11152 12221 11192
rect 16291 11152 16300 11192
rect 16340 11152 18604 11192
rect 18644 11152 18653 11192
rect 23395 11152 23404 11192
rect 23444 11152 23636 11192
rect 23875 11152 23884 11192
rect 23924 11152 24748 11192
rect 24788 11152 24797 11192
rect 31747 11152 31756 11192
rect 31796 11152 32428 11192
rect 32468 11152 32716 11192
rect 32756 11152 32765 11192
rect 33100 11152 34252 11192
rect 34292 11152 34301 11192
rect 18595 11151 18653 11152
rect 34243 11151 34301 11152
rect 32899 11108 32957 11109
rect 4003 11068 4012 11108
rect 4052 11068 5932 11108
rect 5972 11068 5981 11108
rect 7747 11068 7756 11108
rect 7796 11068 10156 11108
rect 10196 11068 10205 11108
rect 17923 11068 17932 11108
rect 17972 11068 19084 11108
rect 19124 11068 19564 11108
rect 19604 11068 20812 11108
rect 20852 11068 20861 11108
rect 31564 11068 32908 11108
rect 32948 11068 32957 11108
rect 31564 11024 31604 11068
rect 32899 11067 32957 11068
rect 32515 11024 32573 11025
rect 35116 11024 35156 11236
rect 36451 11276 36509 11277
rect 37036 11276 37076 11404
rect 42124 11320 42508 11360
rect 42548 11320 42557 11360
rect 42787 11320 42796 11360
rect 42836 11320 45100 11360
rect 45140 11320 45149 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 42124 11276 42164 11320
rect 36451 11236 36460 11276
rect 36500 11236 36652 11276
rect 36692 11236 36701 11276
rect 36941 11236 37036 11276
rect 37076 11236 37612 11276
rect 37652 11236 37661 11276
rect 42115 11236 42124 11276
rect 42164 11236 42173 11276
rect 36451 11235 36509 11236
rect 36067 11192 36125 11193
rect 36355 11192 36413 11193
rect 35203 11152 35212 11192
rect 35252 11152 35692 11192
rect 35732 11152 35741 11192
rect 35875 11152 35884 11192
rect 35924 11152 35933 11192
rect 36067 11152 36076 11192
rect 36116 11152 36172 11192
rect 36212 11152 36221 11192
rect 36355 11152 36364 11192
rect 36404 11152 36498 11192
rect 38947 11152 38956 11192
rect 38996 11152 39532 11192
rect 39572 11152 40012 11192
rect 40052 11152 40061 11192
rect 45379 11152 45388 11192
rect 45428 11152 45964 11192
rect 46004 11152 46636 11192
rect 46676 11152 48172 11192
rect 48212 11152 48221 11192
rect 35884 11108 35924 11152
rect 36067 11151 36125 11152
rect 36355 11151 36413 11152
rect 35299 11068 35308 11108
rect 35348 11068 36940 11108
rect 36980 11068 37132 11108
rect 37172 11068 37181 11108
rect 37987 11068 37996 11108
rect 38036 11068 38572 11108
rect 38612 11068 38621 11108
rect 41635 11068 41644 11108
rect 41684 11068 47308 11108
rect 47348 11068 47788 11108
rect 47828 11068 47837 11108
rect 48067 11068 48076 11108
rect 48116 11068 48460 11108
rect 48500 11068 48509 11108
rect 36172 11024 36212 11068
rect 2563 10984 2572 11024
rect 2612 10984 3436 11024
rect 3476 10984 3485 11024
rect 5251 10984 5260 11024
rect 5300 10984 7372 11024
rect 7412 10984 7421 11024
rect 8131 10984 8140 11024
rect 8180 10984 8908 11024
rect 8948 10984 8957 11024
rect 9283 10984 9292 11024
rect 9332 10984 9868 11024
rect 9908 10984 9917 11024
rect 13891 10984 13900 11024
rect 13940 10984 15140 11024
rect 16963 10984 16972 11024
rect 17012 10984 17548 11024
rect 17588 10984 17597 11024
rect 18019 10984 18028 11024
rect 18068 10984 19468 11024
rect 19508 10984 19517 11024
rect 19747 10984 19756 11024
rect 19796 10984 24076 11024
rect 24116 10984 24125 11024
rect 24355 10984 24364 11024
rect 24404 10984 24556 11024
rect 24596 10984 24605 11024
rect 24835 10984 24844 11024
rect 24884 10984 26956 11024
rect 26996 10984 27005 11024
rect 28099 10984 28108 11024
rect 28148 10984 28972 11024
rect 29012 10984 29021 11024
rect 30115 10984 30124 11024
rect 30164 10984 31564 11024
rect 31604 10984 31613 11024
rect 31948 10984 32524 11024
rect 32564 10984 32573 11024
rect 32707 10984 32716 11024
rect 32756 10984 33196 11024
rect 33236 10984 33245 11024
rect 34915 10984 34924 11024
rect 34964 10984 35156 11024
rect 36163 10984 36172 11024
rect 36212 10984 36221 11024
rect 36355 10984 36364 11024
rect 36404 10984 36844 11024
rect 36884 10984 36893 11024
rect 37507 10984 37516 11024
rect 37556 10984 38380 11024
rect 38420 10984 38429 11024
rect 40195 10984 40204 11024
rect 40244 10984 40684 11024
rect 40724 10984 40733 11024
rect 43651 10984 43660 11024
rect 43700 10984 45004 11024
rect 45044 10984 46156 11024
rect 46196 10984 46205 11024
rect 47683 10984 47692 11024
rect 47732 10984 48268 11024
rect 48308 10984 48317 11024
rect 15100 10940 15140 10984
rect 24364 10940 24404 10984
rect 30124 10940 30164 10984
rect 15100 10900 17740 10940
rect 17780 10900 17789 10940
rect 22339 10900 22348 10940
rect 22388 10900 24404 10940
rect 27235 10900 27244 10940
rect 27284 10900 30164 10940
rect 20899 10856 20957 10857
rect 31948 10856 31988 10984
rect 32515 10983 32573 10984
rect 36163 10940 36221 10941
rect 32035 10900 32044 10940
rect 32084 10900 34156 10940
rect 34196 10900 35020 10940
rect 35060 10900 35069 10940
rect 35587 10900 35596 10940
rect 35636 10900 35645 10940
rect 36163 10900 36172 10940
rect 36212 10900 36652 10940
rect 36692 10900 36701 10940
rect 1507 10816 1516 10856
rect 1556 10816 2572 10856
rect 2612 10816 2621 10856
rect 4099 10816 4108 10856
rect 4148 10816 5452 10856
rect 5492 10816 5501 10856
rect 8419 10816 8428 10856
rect 8468 10816 9676 10856
rect 9716 10816 9725 10856
rect 17443 10816 17452 10856
rect 17492 10816 18796 10856
rect 18836 10816 18845 10856
rect 19651 10816 19660 10856
rect 19700 10816 20908 10856
rect 20948 10816 23020 10856
rect 23060 10816 23692 10856
rect 23732 10816 23741 10856
rect 29059 10816 29068 10856
rect 29108 10816 31988 10856
rect 32131 10856 32189 10857
rect 35596 10856 35636 10900
rect 36163 10899 36221 10900
rect 32131 10816 32140 10856
rect 32180 10816 33772 10856
rect 33812 10816 33821 10856
rect 34339 10816 34348 10856
rect 34388 10816 36268 10856
rect 36308 10816 36748 10856
rect 36788 10816 37708 10856
rect 37748 10816 37757 10856
rect 45763 10816 45772 10856
rect 45812 10816 48364 10856
rect 48404 10816 48413 10856
rect 20899 10815 20957 10816
rect 32131 10815 32189 10816
rect 19363 10772 19421 10773
rect 9379 10732 9388 10772
rect 9428 10732 10060 10772
rect 10100 10732 10109 10772
rect 18403 10732 18412 10772
rect 18452 10732 18461 10772
rect 19363 10732 19372 10772
rect 19412 10732 19756 10772
rect 19796 10732 19805 10772
rect 37219 10732 37228 10772
rect 37268 10732 38188 10772
rect 38228 10732 38237 10772
rect 42883 10732 42892 10772
rect 42932 10732 43660 10772
rect 43700 10732 44428 10772
rect 44468 10732 44908 10772
rect 44948 10732 44957 10772
rect 48259 10732 48268 10772
rect 48308 10732 48556 10772
rect 48596 10732 48605 10772
rect 0 10688 80 10708
rect 18412 10688 18452 10732
rect 19363 10731 19421 10732
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 4771 10648 4780 10688
rect 4820 10648 5356 10688
rect 5396 10648 5405 10688
rect 5923 10648 5932 10688
rect 5972 10648 6316 10688
rect 6356 10648 9292 10688
rect 9332 10648 9341 10688
rect 18412 10648 20620 10688
rect 20660 10648 20669 10688
rect 27715 10648 27724 10688
rect 27764 10648 32908 10688
rect 32948 10648 32957 10688
rect 37507 10648 37516 10688
rect 37556 10648 38764 10688
rect 38804 10648 39820 10688
rect 39860 10648 39869 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 32227 10564 32236 10604
rect 32276 10564 33100 10604
rect 33140 10564 33149 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 37603 10564 37612 10604
rect 37652 10564 38228 10604
rect 46339 10564 46348 10604
rect 46388 10564 47212 10604
rect 47252 10564 47261 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 18115 10520 18173 10521
rect 20803 10520 20861 10521
rect 32131 10520 32189 10521
rect 38188 10520 38228 10564
rect 18115 10480 18124 10520
rect 18164 10480 19372 10520
rect 19412 10480 19421 10520
rect 20707 10480 20716 10520
rect 20756 10480 20812 10520
rect 20852 10480 20861 10520
rect 32046 10480 32140 10520
rect 32180 10480 32189 10520
rect 32803 10480 32812 10520
rect 32852 10480 34924 10520
rect 34964 10480 35308 10520
rect 35348 10480 35357 10520
rect 38179 10480 38188 10520
rect 38228 10480 38237 10520
rect 18115 10479 18173 10480
rect 19372 10436 19412 10480
rect 20803 10479 20861 10480
rect 32131 10479 32189 10480
rect 31651 10436 31709 10437
rect 3715 10396 3724 10436
rect 3764 10396 4204 10436
rect 4244 10396 4253 10436
rect 6979 10396 6988 10436
rect 7028 10396 7468 10436
rect 7508 10396 8428 10436
rect 8468 10396 8620 10436
rect 8660 10396 8669 10436
rect 8899 10396 8908 10436
rect 8948 10396 9772 10436
rect 9812 10396 10636 10436
rect 10676 10396 10685 10436
rect 16771 10396 16780 10436
rect 16820 10396 17644 10436
rect 17684 10396 18220 10436
rect 18260 10396 18269 10436
rect 18691 10396 18700 10436
rect 18740 10396 18988 10436
rect 19028 10396 19037 10436
rect 19372 10396 22636 10436
rect 22676 10396 22685 10436
rect 24547 10396 24556 10436
rect 24596 10396 24748 10436
rect 24788 10396 31660 10436
rect 31700 10396 31709 10436
rect 31651 10395 31709 10396
rect 31948 10396 33004 10436
rect 33044 10396 33484 10436
rect 33524 10396 33533 10436
rect 36547 10396 36556 10436
rect 36596 10396 37324 10436
rect 37364 10396 37373 10436
rect 37699 10396 37708 10436
rect 37748 10396 39148 10436
rect 39188 10396 39197 10436
rect 42883 10396 42892 10436
rect 42932 10396 48940 10436
rect 48980 10396 48989 10436
rect 17635 10352 17693 10353
rect 20323 10352 20381 10353
rect 21763 10352 21821 10353
rect 31948 10352 31988 10396
rect 43171 10352 43229 10353
rect 7555 10312 7564 10352
rect 7604 10312 8524 10352
rect 8564 10312 9100 10352
rect 9140 10312 9676 10352
rect 9716 10312 9725 10352
rect 9868 10312 11308 10352
rect 11348 10312 11357 10352
rect 17635 10312 17644 10352
rect 17684 10312 18604 10352
rect 18644 10312 18653 10352
rect 20238 10312 20332 10352
rect 20372 10312 21580 10352
rect 21620 10312 21629 10352
rect 21763 10312 21772 10352
rect 21812 10312 22156 10352
rect 22196 10312 25612 10352
rect 25652 10312 25661 10352
rect 29251 10312 29260 10352
rect 29300 10312 31372 10352
rect 31412 10312 31421 10352
rect 31747 10312 31756 10352
rect 31796 10312 31948 10352
rect 31988 10312 31997 10352
rect 32515 10312 32524 10352
rect 32564 10312 33100 10352
rect 33140 10312 33149 10352
rect 35011 10312 35020 10352
rect 35060 10312 36076 10352
rect 36116 10312 36125 10352
rect 36355 10312 36364 10352
rect 36404 10312 36844 10352
rect 36884 10312 36893 10352
rect 37411 10312 37420 10352
rect 37460 10312 37469 10352
rect 41635 10312 41644 10352
rect 41684 10312 42220 10352
rect 42260 10312 42269 10352
rect 43086 10312 43180 10352
rect 43220 10312 45676 10352
rect 45716 10312 45725 10352
rect 46636 10312 48076 10352
rect 48116 10312 48125 10352
rect 7564 10268 7604 10312
rect 3907 10228 3916 10268
rect 3956 10228 4876 10268
rect 4916 10228 7604 10268
rect 7651 10228 7660 10268
rect 7700 10228 9772 10268
rect 9812 10228 9821 10268
rect 9868 10184 9908 10312
rect 17635 10311 17693 10312
rect 20323 10311 20381 10312
rect 21763 10311 21821 10312
rect 36547 10268 36605 10269
rect 37420 10268 37460 10312
rect 43171 10311 43229 10312
rect 46636 10268 46676 10312
rect 11320 10228 15436 10268
rect 15476 10228 15485 10268
rect 17740 10228 22060 10268
rect 22100 10228 22109 10268
rect 22915 10228 22924 10268
rect 22964 10228 23697 10268
rect 23737 10228 25708 10268
rect 25748 10228 25757 10268
rect 26947 10228 26956 10268
rect 26996 10228 29452 10268
rect 29492 10228 29501 10268
rect 31651 10228 31660 10268
rect 31700 10228 32812 10268
rect 32852 10228 32861 10268
rect 34147 10228 34156 10268
rect 34196 10228 36404 10268
rect 11320 10184 11360 10228
rect 17740 10184 17780 10228
rect 24835 10184 24893 10185
rect 32899 10184 32957 10185
rect 35683 10184 35741 10185
rect 36364 10184 36404 10228
rect 36547 10228 36556 10268
rect 36596 10228 37460 10268
rect 37699 10228 37708 10268
rect 37748 10228 41600 10268
rect 42307 10228 42316 10268
rect 42356 10228 46636 10268
rect 46676 10228 46685 10268
rect 36547 10227 36605 10228
rect 36451 10184 36509 10185
rect 41560 10184 41600 10228
rect 2563 10144 2572 10184
rect 2612 10144 2764 10184
rect 2804 10144 4972 10184
rect 5012 10144 5356 10184
rect 5396 10144 6316 10184
rect 6356 10144 6892 10184
rect 6932 10144 6941 10184
rect 8227 10144 8236 10184
rect 8276 10144 8285 10184
rect 8707 10144 8716 10184
rect 8756 10144 9196 10184
rect 9236 10144 9868 10184
rect 9908 10144 9917 10184
rect 10531 10144 10540 10184
rect 10580 10144 10589 10184
rect 10723 10144 10732 10184
rect 10772 10144 11360 10184
rect 12163 10144 12172 10184
rect 12212 10144 13420 10184
rect 13460 10144 13469 10184
rect 17731 10144 17740 10184
rect 17780 10144 17789 10184
rect 19267 10144 19276 10184
rect 19316 10144 20236 10184
rect 20276 10144 20285 10184
rect 20515 10144 20524 10184
rect 20564 10144 21868 10184
rect 21908 10144 21917 10184
rect 22243 10144 22252 10184
rect 22292 10144 23404 10184
rect 23444 10144 23453 10184
rect 23587 10144 23596 10184
rect 23636 10144 24364 10184
rect 24404 10144 24844 10184
rect 24884 10144 24893 10184
rect 25603 10144 25612 10184
rect 25652 10144 27052 10184
rect 27092 10144 27101 10184
rect 27331 10144 27340 10184
rect 27380 10144 28012 10184
rect 28052 10144 28061 10184
rect 29635 10144 29644 10184
rect 29684 10144 30740 10184
rect 31555 10144 31564 10184
rect 31604 10144 32428 10184
rect 32468 10144 32477 10184
rect 32814 10144 32908 10184
rect 32948 10144 32957 10184
rect 34531 10144 34540 10184
rect 34580 10144 35404 10184
rect 35444 10144 35453 10184
rect 35598 10144 35692 10184
rect 35732 10144 35741 10184
rect 35784 10144 35793 10184
rect 35833 10144 35980 10184
rect 36020 10144 36029 10184
rect 36355 10144 36364 10184
rect 36404 10144 36460 10184
rect 36500 10144 36509 10184
rect 36739 10144 36748 10184
rect 36788 10144 37420 10184
rect 37460 10144 37469 10184
rect 38179 10144 38188 10184
rect 38228 10144 39628 10184
rect 39668 10144 41396 10184
rect 41560 10144 42604 10184
rect 42644 10144 42653 10184
rect 43555 10144 43564 10184
rect 43604 10144 44140 10184
rect 44180 10144 44189 10184
rect 44419 10144 44428 10184
rect 44468 10144 44477 10184
rect 47779 10144 47788 10184
rect 47828 10144 49036 10184
rect 49076 10144 49085 10184
rect 8236 10100 8276 10144
rect 10540 10100 10580 10144
rect 24835 10143 24893 10144
rect 17731 10100 17789 10101
rect 27340 10100 27380 10144
rect 30700 10100 30740 10144
rect 32899 10143 32957 10144
rect 35683 10143 35741 10144
rect 36451 10143 36509 10144
rect 4675 10060 4684 10100
rect 4724 10060 4916 10100
rect 8236 10060 8812 10100
rect 8852 10060 9964 10100
rect 10004 10060 10013 10100
rect 10540 10060 11692 10100
rect 11732 10060 13228 10100
rect 13268 10060 13277 10100
rect 17731 10060 17740 10100
rect 17780 10060 18508 10100
rect 18548 10060 18557 10100
rect 20611 10060 20620 10100
rect 20660 10060 20812 10100
rect 20852 10060 20861 10100
rect 20910 10060 20919 10100
rect 20959 10060 25324 10100
rect 25364 10060 25373 10100
rect 26851 10060 26860 10100
rect 26900 10060 27380 10100
rect 28387 10060 28396 10100
rect 28436 10060 29740 10100
rect 29780 10060 29789 10100
rect 30700 10060 32140 10100
rect 32180 10060 32189 10100
rect 32236 10060 33292 10100
rect 33332 10060 33341 10100
rect 34051 10060 34060 10100
rect 34100 10060 35308 10100
rect 35348 10060 35357 10100
rect 38659 10060 38668 10100
rect 38708 10060 39052 10100
rect 39092 10060 39101 10100
rect 4876 10016 4916 10060
rect 17731 10059 17789 10060
rect 24067 10016 24125 10017
rect 24259 10016 24317 10017
rect 32236 10016 32276 10060
rect 32620 10016 32660 10060
rect 41356 10016 41396 10144
rect 44428 10100 44468 10144
rect 43075 10060 43084 10100
rect 43124 10060 44468 10100
rect 44707 10060 44716 10100
rect 44756 10060 45484 10100
rect 45524 10060 46924 10100
rect 46964 10060 47692 10100
rect 47732 10060 47741 10100
rect 44716 10016 44756 10060
rect 3523 9976 3532 10016
rect 3572 9976 3916 10016
rect 3956 9976 3965 10016
rect 4867 9976 4876 10016
rect 4916 9976 4925 10016
rect 5827 9976 5836 10016
rect 5876 9976 9676 10016
rect 9716 9976 9725 10016
rect 11971 9976 11980 10016
rect 12020 9976 12460 10016
rect 12500 9976 12509 10016
rect 16579 9976 16588 10016
rect 16628 9976 16780 10016
rect 16820 9976 16829 10016
rect 23299 9976 23308 10016
rect 23348 9976 24076 10016
rect 24116 9976 24125 10016
rect 24174 9976 24268 10016
rect 24308 9976 24317 10016
rect 31555 9976 31564 10016
rect 31604 9976 32276 10016
rect 32611 9976 32620 10016
rect 32660 9976 32669 10016
rect 36643 9976 36652 10016
rect 36692 9976 37228 10016
rect 37268 9976 37277 10016
rect 41347 9976 41356 10016
rect 41396 9976 41405 10016
rect 43363 9976 43372 10016
rect 43412 9976 44756 10016
rect 24067 9975 24125 9976
rect 24259 9975 24317 9976
rect 32035 9932 32093 9933
rect 19075 9892 19084 9932
rect 19124 9892 24172 9932
rect 24212 9892 24221 9932
rect 28960 9892 29260 9932
rect 29300 9892 29309 9932
rect 31939 9892 31948 9932
rect 31988 9892 32044 9932
rect 32084 9892 32093 9932
rect 41059 9892 41068 9932
rect 41108 9892 41740 9932
rect 41780 9892 41789 9932
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 15523 9808 15532 9848
rect 15572 9808 15916 9848
rect 15956 9808 17068 9848
rect 17108 9808 17117 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 20323 9808 20332 9848
rect 20372 9808 25132 9848
rect 25172 9808 25181 9848
rect 0 9788 80 9808
rect 28960 9764 29000 9892
rect 32035 9891 32093 9892
rect 31651 9848 31709 9849
rect 36355 9848 36413 9849
rect 31651 9808 31660 9848
rect 31700 9808 32236 9848
rect 32276 9808 32285 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 35587 9808 35596 9848
rect 35636 9808 36364 9848
rect 36404 9808 36413 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 31651 9807 31709 9808
rect 36355 9807 36413 9808
rect 31843 9764 31901 9765
rect 16387 9724 16396 9764
rect 16436 9724 16972 9764
rect 17012 9724 17021 9764
rect 18787 9724 18796 9764
rect 18836 9724 29000 9764
rect 31747 9724 31756 9764
rect 31796 9724 31852 9764
rect 31892 9724 31901 9764
rect 31843 9723 31901 9724
rect 7171 9640 7180 9680
rect 7220 9640 9772 9680
rect 9812 9640 9821 9680
rect 15715 9640 15724 9680
rect 15764 9640 16012 9680
rect 16052 9640 17260 9680
rect 17300 9640 17309 9680
rect 20995 9640 21004 9680
rect 21044 9640 21964 9680
rect 22004 9640 22013 9680
rect 22723 9640 22732 9680
rect 22772 9640 23308 9680
rect 23348 9640 23357 9680
rect 25123 9640 25132 9680
rect 25172 9640 25516 9680
rect 25556 9640 25565 9680
rect 29827 9640 29836 9680
rect 29876 9640 30740 9680
rect 35875 9640 35884 9680
rect 35924 9640 36268 9680
rect 36308 9640 36317 9680
rect 41731 9640 41740 9680
rect 41780 9640 42988 9680
rect 43028 9640 43037 9680
rect 30700 9596 30740 9640
rect 32035 9596 32093 9597
rect 7651 9556 7660 9596
rect 7700 9556 8044 9596
rect 8084 9556 8093 9596
rect 10243 9556 10252 9596
rect 10292 9556 10924 9596
rect 10964 9556 10973 9596
rect 16483 9556 16492 9596
rect 16532 9556 17356 9596
rect 17396 9556 17405 9596
rect 22540 9556 30220 9596
rect 30260 9556 30269 9596
rect 30691 9556 30700 9596
rect 30740 9556 31276 9596
rect 31316 9556 32044 9596
rect 32084 9556 32093 9596
rect 21379 9512 21437 9513
rect 22540 9512 22580 9556
rect 32035 9555 32093 9556
rect 24931 9512 24989 9513
rect 27139 9512 27197 9513
rect 1603 9472 1612 9512
rect 1652 9472 3532 9512
rect 3572 9472 3581 9512
rect 4195 9472 4204 9512
rect 4244 9472 5260 9512
rect 5300 9472 5309 9512
rect 6979 9472 6988 9512
rect 7028 9472 8332 9512
rect 8372 9472 8381 9512
rect 15619 9472 15628 9512
rect 15668 9472 16780 9512
rect 16820 9472 16829 9512
rect 17059 9472 17068 9512
rect 17108 9472 17548 9512
rect 17588 9472 17740 9512
rect 17780 9472 18316 9512
rect 18356 9472 18365 9512
rect 20803 9472 20812 9512
rect 20852 9472 21388 9512
rect 21428 9472 21437 9512
rect 22531 9472 22540 9512
rect 22580 9472 22589 9512
rect 23683 9472 23692 9512
rect 23732 9472 24172 9512
rect 24212 9472 24556 9512
rect 24596 9472 24605 9512
rect 24931 9472 24940 9512
rect 24980 9472 25516 9512
rect 25556 9472 25565 9512
rect 27139 9472 27148 9512
rect 27188 9472 27436 9512
rect 27476 9472 27485 9512
rect 28579 9472 28588 9512
rect 28628 9472 32051 9512
rect 32091 9472 32100 9512
rect 35107 9472 35116 9512
rect 35156 9472 35788 9512
rect 35828 9472 35837 9512
rect 42403 9472 42412 9512
rect 42452 9472 42988 9512
rect 43028 9472 43037 9512
rect 44035 9472 44044 9512
rect 44084 9472 44428 9512
rect 44468 9472 44477 9512
rect 21379 9471 21437 9472
rect 24931 9471 24989 9472
rect 27139 9471 27197 9472
rect 21571 9428 21629 9429
rect 2500 9388 2860 9428
rect 2900 9388 4300 9428
rect 4340 9388 4588 9428
rect 4628 9388 6124 9428
rect 6164 9388 6173 9428
rect 21379 9388 21388 9428
rect 21428 9388 21580 9428
rect 21620 9388 21629 9428
rect 24067 9388 24076 9428
rect 24116 9388 24844 9428
rect 24884 9388 25324 9428
rect 25364 9388 25373 9428
rect 26947 9388 26956 9428
rect 26996 9388 27005 9428
rect 27907 9388 27916 9428
rect 27956 9388 28300 9428
rect 28340 9388 28349 9428
rect 29059 9388 29068 9428
rect 29108 9388 29644 9428
rect 29684 9388 30892 9428
rect 30932 9388 31660 9428
rect 31700 9388 31709 9428
rect 37795 9388 37804 9428
rect 37844 9388 38572 9428
rect 38612 9388 39244 9428
rect 39284 9388 39293 9428
rect 41347 9388 41356 9428
rect 41396 9388 43276 9428
rect 43316 9388 44620 9428
rect 44660 9388 44669 9428
rect 2500 9344 2540 9388
rect 21571 9387 21629 9388
rect 20803 9344 20861 9345
rect 26956 9344 26996 9388
rect 32035 9344 32093 9345
rect 1699 9304 1708 9344
rect 1748 9304 2540 9344
rect 4867 9304 4876 9344
rect 4916 9304 5740 9344
rect 5780 9304 5789 9344
rect 7267 9304 7276 9344
rect 7316 9304 9292 9344
rect 9332 9304 9341 9344
rect 13603 9304 13612 9344
rect 13652 9304 17644 9344
rect 17684 9304 17693 9344
rect 18019 9304 18028 9344
rect 18068 9304 18220 9344
rect 18260 9304 18269 9344
rect 20718 9304 20812 9344
rect 20852 9304 20861 9344
rect 21955 9304 21964 9344
rect 22004 9304 25364 9344
rect 26956 9304 28204 9344
rect 28244 9304 28253 9344
rect 29347 9304 29356 9344
rect 29396 9304 29932 9344
rect 29972 9304 31276 9344
rect 31316 9304 31325 9344
rect 31950 9304 32044 9344
rect 32084 9304 32093 9344
rect 35011 9304 35020 9344
rect 35060 9304 35884 9344
rect 35924 9304 35933 9344
rect 37987 9304 37996 9344
rect 38036 9304 38668 9344
rect 38708 9304 38717 9344
rect 42691 9304 42700 9344
rect 42740 9304 43180 9344
rect 43220 9304 43229 9344
rect 20803 9303 20861 9304
rect 25324 9260 25364 9304
rect 32035 9303 32093 9304
rect 1027 9220 1036 9260
rect 1076 9220 1900 9260
rect 1940 9220 1949 9260
rect 7660 9220 7852 9260
rect 7892 9220 7901 9260
rect 16675 9220 16684 9260
rect 16724 9220 17260 9260
rect 17300 9220 17309 9260
rect 23107 9220 23116 9260
rect 23156 9220 24172 9260
rect 24212 9220 24221 9260
rect 24643 9220 24652 9260
rect 24692 9220 25036 9260
rect 25076 9220 25085 9260
rect 25315 9220 25324 9260
rect 25364 9220 25373 9260
rect 31075 9220 31084 9260
rect 31124 9220 31372 9260
rect 31412 9220 31421 9260
rect 32236 9220 33580 9260
rect 33620 9220 33629 9260
rect 45859 9220 45868 9260
rect 45908 9220 47308 9260
rect 47348 9220 47357 9260
rect 7363 9136 7372 9176
rect 7412 9136 7564 9176
rect 7604 9136 7613 9176
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 1315 8884 1324 8924
rect 1364 8884 2284 8924
rect 2324 8884 4012 8924
rect 4052 8884 4061 8924
rect 7660 8840 7700 9220
rect 7747 9136 7756 9176
rect 7796 9136 9388 9176
rect 9428 9136 9437 9176
rect 20131 9136 20140 9176
rect 20180 9136 20332 9176
rect 20372 9136 20381 9176
rect 22819 9136 22828 9176
rect 22868 9136 23020 9176
rect 23060 9136 23069 9176
rect 2371 8800 2380 8840
rect 2420 8800 2540 8840
rect 2659 8800 2668 8840
rect 2708 8800 3724 8840
rect 3764 8800 3773 8840
rect 4099 8800 4108 8840
rect 4148 8800 5932 8840
rect 5972 8800 5981 8840
rect 7651 8800 7660 8840
rect 7700 8800 7709 8840
rect 2500 8756 2540 8800
rect 7756 8756 7796 9136
rect 32236 9093 32276 9220
rect 36067 9176 36125 9177
rect 35779 9136 35788 9176
rect 35828 9136 36076 9176
rect 36116 9136 36125 9176
rect 36067 9135 36125 9136
rect 26659 9092 26717 9093
rect 32227 9092 32285 9093
rect 14851 9052 14860 9092
rect 14900 9052 15148 9092
rect 15188 9052 16492 9092
rect 16532 9052 16541 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 20995 9052 21004 9092
rect 21044 9052 21292 9092
rect 21332 9052 22732 9092
rect 22772 9052 22781 9092
rect 26574 9052 26668 9092
rect 26708 9052 26717 9092
rect 31555 9052 31564 9092
rect 31604 9052 32236 9092
rect 32276 9052 32285 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 26659 9051 26717 9052
rect 32227 9051 32285 9052
rect 32323 9008 32381 9009
rect 20419 8968 20428 9008
rect 20468 8968 20477 9008
rect 30403 8968 30412 9008
rect 30452 8968 30461 9008
rect 32227 8968 32236 9008
rect 32276 8968 32332 9008
rect 32372 8968 32381 9008
rect 20428 8840 20468 8968
rect 24355 8924 24413 8925
rect 30307 8924 30365 8925
rect 20707 8884 20716 8924
rect 20756 8884 21964 8924
rect 22004 8884 22013 8924
rect 22819 8884 22828 8924
rect 22868 8884 23788 8924
rect 23828 8884 23837 8924
rect 24270 8884 24364 8924
rect 24404 8884 24884 8924
rect 30222 8884 30316 8924
rect 30356 8884 30365 8924
rect 24355 8883 24413 8884
rect 21475 8840 21533 8841
rect 24844 8840 24884 8884
rect 30307 8883 30365 8884
rect 27715 8840 27773 8841
rect 28003 8840 28061 8841
rect 30412 8840 30452 8968
rect 32323 8967 32381 8968
rect 34243 9008 34301 9009
rect 34243 8968 34252 9008
rect 34292 8968 34732 9008
rect 34772 8968 34781 9008
rect 34243 8967 34301 8968
rect 31555 8884 31564 8924
rect 31604 8884 32140 8924
rect 32180 8884 32189 8924
rect 33868 8884 34348 8924
rect 34388 8884 34397 8924
rect 30691 8840 30749 8841
rect 31459 8840 31517 8841
rect 33868 8840 33908 8884
rect 34051 8840 34109 8841
rect 8323 8800 8332 8840
rect 8372 8800 9004 8840
rect 9044 8800 9053 8840
rect 9475 8800 9484 8840
rect 9524 8800 10060 8840
rect 10100 8800 10109 8840
rect 17827 8800 17836 8840
rect 17876 8800 17885 8840
rect 18883 8800 18892 8840
rect 18932 8800 20468 8840
rect 20899 8800 20908 8840
rect 20948 8800 21484 8840
rect 21524 8800 21533 8840
rect 22435 8800 22444 8840
rect 22484 8800 23212 8840
rect 23252 8800 23261 8840
rect 23587 8800 23596 8840
rect 23636 8800 24748 8840
rect 24788 8800 24797 8840
rect 24844 8800 27239 8840
rect 27279 8800 27288 8840
rect 27630 8800 27724 8840
rect 27764 8800 27773 8840
rect 27918 8800 28012 8840
rect 28052 8800 28061 8840
rect 9484 8756 9524 8800
rect 17836 8756 17876 8800
rect 21475 8799 21533 8800
rect 27715 8799 27773 8800
rect 28003 8799 28061 8800
rect 29548 8800 30452 8840
rect 30606 8800 30700 8840
rect 30740 8800 30749 8840
rect 31344 8800 31372 8840
rect 31412 8800 31468 8840
rect 31508 8800 31948 8840
rect 31988 8800 31997 8840
rect 33571 8800 33580 8840
rect 33620 8800 33908 8840
rect 33966 8800 34060 8840
rect 34100 8800 34109 8840
rect 37891 8800 37900 8840
rect 37940 8800 38956 8840
rect 38996 8800 39005 8840
rect 41155 8800 41164 8840
rect 41204 8800 41548 8840
rect 41588 8800 41597 8840
rect 42787 8800 42796 8840
rect 42836 8800 44236 8840
rect 44276 8800 44285 8840
rect 46435 8800 46444 8840
rect 46484 8800 47116 8840
rect 47156 8800 47165 8840
rect 24643 8756 24701 8757
rect 24931 8756 24989 8757
rect 2500 8716 3628 8756
rect 3668 8716 3677 8756
rect 4963 8716 4972 8756
rect 5012 8716 7796 8756
rect 8035 8716 8044 8756
rect 8084 8716 9524 8756
rect 10243 8716 10252 8756
rect 10292 8716 10636 8756
rect 10676 8716 13900 8756
rect 13940 8716 13949 8756
rect 17836 8716 21868 8756
rect 21908 8716 24364 8756
rect 24404 8716 24413 8756
rect 24558 8716 24652 8756
rect 24692 8716 24701 8756
rect 24846 8716 24940 8756
rect 24980 8716 24989 8756
rect 28579 8716 28588 8756
rect 28628 8716 29164 8756
rect 29204 8716 29213 8756
rect 3523 8632 3532 8672
rect 3572 8632 3724 8672
rect 3764 8632 3773 8672
rect 6595 8632 6604 8672
rect 6644 8632 7468 8672
rect 7508 8632 7517 8672
rect 8044 8504 8084 8716
rect 24643 8715 24701 8716
rect 24931 8715 24989 8716
rect 23203 8672 23261 8673
rect 29548 8672 29588 8800
rect 30691 8799 30749 8800
rect 31459 8799 31517 8800
rect 34051 8799 34109 8800
rect 30595 8716 30604 8756
rect 30644 8716 30988 8756
rect 31028 8716 31037 8756
rect 33763 8716 33772 8756
rect 33812 8716 34252 8756
rect 34292 8716 34924 8756
rect 34964 8716 34973 8756
rect 41443 8716 41452 8756
rect 41492 8716 43468 8756
rect 43508 8716 43517 8756
rect 34147 8672 34205 8673
rect 8899 8632 8908 8672
rect 8948 8632 9868 8672
rect 9908 8632 9917 8672
rect 10723 8632 10732 8672
rect 10772 8632 11404 8672
rect 11444 8632 11453 8672
rect 11683 8632 11692 8672
rect 11732 8632 12268 8672
rect 12308 8632 12317 8672
rect 13987 8632 13996 8672
rect 14036 8632 14668 8672
rect 14708 8632 16012 8672
rect 16052 8632 16061 8672
rect 16387 8632 16396 8672
rect 16436 8632 17356 8672
rect 17396 8632 17405 8672
rect 18307 8632 18316 8672
rect 18356 8632 19084 8672
rect 19124 8632 19133 8672
rect 19747 8632 19756 8672
rect 19796 8632 21484 8672
rect 21524 8632 21533 8672
rect 22723 8632 22732 8672
rect 22772 8632 23212 8672
rect 23252 8632 23261 8672
rect 23395 8632 23404 8672
rect 23444 8632 23692 8672
rect 23732 8632 23741 8672
rect 23875 8632 23884 8672
rect 23924 8632 24076 8672
rect 24116 8632 24125 8672
rect 24259 8632 24268 8672
rect 24308 8632 27436 8672
rect 27476 8632 27485 8672
rect 27715 8632 27724 8672
rect 27764 8632 28012 8672
rect 28052 8632 28061 8672
rect 29539 8632 29548 8672
rect 29588 8632 29597 8672
rect 30307 8632 30316 8672
rect 30356 8632 31468 8672
rect 31508 8632 31517 8672
rect 34147 8632 34156 8672
rect 34196 8632 35020 8672
rect 35060 8632 35069 8672
rect 35203 8632 35212 8672
rect 35252 8632 35596 8672
rect 35636 8632 35645 8672
rect 40003 8632 40012 8672
rect 40052 8632 41356 8672
rect 41396 8632 41405 8672
rect 43363 8632 43372 8672
rect 43412 8632 45484 8672
rect 45524 8632 47116 8672
rect 47156 8632 48172 8672
rect 48212 8632 48221 8672
rect 9868 8588 9908 8632
rect 23203 8631 23261 8632
rect 20803 8588 20861 8589
rect 27436 8588 27476 8632
rect 34147 8631 34205 8632
rect 9868 8548 11596 8588
rect 11636 8548 11884 8588
rect 11924 8548 11933 8588
rect 18796 8548 20620 8588
rect 20660 8548 20669 8588
rect 20803 8548 20812 8588
rect 20852 8548 21140 8588
rect 22339 8548 22348 8588
rect 22388 8548 23308 8588
rect 23348 8548 23357 8588
rect 24355 8548 24364 8588
rect 24404 8548 25172 8588
rect 26563 8548 26572 8588
rect 26612 8548 26621 8588
rect 27436 8548 28588 8588
rect 28628 8548 28637 8588
rect 28867 8548 28876 8588
rect 28916 8548 29740 8588
rect 29780 8548 30065 8588
rect 30105 8548 30114 8588
rect 30220 8548 44812 8588
rect 44852 8548 45196 8588
rect 45236 8548 45245 8588
rect 18796 8504 18836 8548
rect 20803 8547 20861 8548
rect 19843 8504 19901 8505
rect 20899 8504 20957 8505
rect 21100 8504 21140 8548
rect 21475 8504 21533 8505
rect 25132 8504 25172 8548
rect 26572 8504 26612 8548
rect 28963 8504 29021 8505
rect 30220 8504 30260 8548
rect 33187 8504 33245 8505
rect 3523 8464 3532 8504
rect 3572 8464 8084 8504
rect 16963 8464 16972 8504
rect 17012 8464 18796 8504
rect 18836 8464 18845 8504
rect 19758 8464 19852 8504
rect 19892 8464 19901 8504
rect 19843 8463 19901 8464
rect 19948 8464 20332 8504
rect 20372 8464 20381 8504
rect 20814 8464 20908 8504
rect 20948 8464 20957 8504
rect 21091 8464 21100 8504
rect 21140 8464 21149 8504
rect 21475 8464 21484 8504
rect 21524 8464 21580 8504
rect 21620 8464 21629 8504
rect 22444 8464 22919 8504
rect 22959 8464 24596 8504
rect 24643 8464 24652 8504
rect 24692 8464 24701 8504
rect 25123 8464 25132 8504
rect 25172 8464 25181 8504
rect 25795 8464 25804 8504
rect 25844 8464 26476 8504
rect 26516 8464 26525 8504
rect 26572 8464 27628 8504
rect 27668 8464 28396 8504
rect 28436 8464 28445 8504
rect 28878 8464 28972 8504
rect 29012 8464 29021 8504
rect 29155 8464 29164 8504
rect 29204 8464 30260 8504
rect 30499 8464 30508 8504
rect 30548 8464 33196 8504
rect 33236 8464 33245 8504
rect 34435 8464 34444 8504
rect 34484 8464 35500 8504
rect 35540 8464 35549 8504
rect 38275 8464 38284 8504
rect 38324 8464 40204 8504
rect 40244 8464 40253 8504
rect 41731 8464 41740 8504
rect 41780 8464 43468 8504
rect 43508 8464 43517 8504
rect 19948 8420 19988 8464
rect 20899 8463 20957 8464
rect 21475 8463 21533 8464
rect 5059 8380 5068 8420
rect 5108 8380 6796 8420
rect 6836 8380 8620 8420
rect 8660 8380 9676 8420
rect 9716 8380 9725 8420
rect 15907 8380 15916 8420
rect 15956 8380 17260 8420
rect 17300 8380 19988 8420
rect 20035 8380 20044 8420
rect 20084 8380 20428 8420
rect 20468 8380 20477 8420
rect 20611 8380 20620 8420
rect 20660 8380 22348 8420
rect 22388 8380 22397 8420
rect 20515 8336 20573 8337
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 6019 8296 6028 8336
rect 6068 8296 10156 8336
rect 10196 8296 10828 8336
rect 10868 8296 10877 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 20227 8296 20236 8336
rect 20276 8296 20285 8336
rect 20515 8296 20524 8336
rect 20564 8296 22060 8336
rect 22100 8296 22109 8336
rect 20236 8252 20276 8296
rect 20515 8295 20573 8296
rect 22444 8252 22484 8464
rect 22531 8420 22589 8421
rect 22723 8420 22781 8421
rect 22531 8380 22540 8420
rect 22580 8380 22674 8420
rect 22723 8380 22732 8420
rect 22772 8380 23020 8420
rect 23060 8380 23069 8420
rect 22531 8379 22589 8380
rect 22723 8379 22781 8380
rect 24556 8336 24596 8464
rect 24652 8420 24692 8464
rect 28963 8463 29021 8464
rect 33187 8463 33245 8464
rect 30307 8420 30365 8421
rect 34243 8420 34301 8421
rect 24652 8380 30316 8420
rect 30356 8380 30365 8420
rect 34051 8380 34060 8420
rect 34100 8380 34252 8420
rect 34292 8380 34301 8420
rect 30307 8379 30365 8380
rect 34243 8379 34301 8380
rect 35596 8380 36076 8420
rect 36116 8380 36125 8420
rect 36547 8380 36556 8420
rect 36596 8380 42508 8420
rect 42548 8380 45772 8420
rect 45812 8380 45821 8420
rect 23107 8296 23116 8336
rect 23156 8296 23596 8336
rect 23636 8296 23645 8336
rect 23779 8296 23788 8336
rect 23828 8296 24500 8336
rect 24556 8296 24844 8336
rect 24884 8296 24893 8336
rect 25219 8296 25228 8336
rect 25268 8296 26284 8336
rect 26324 8296 26333 8336
rect 26659 8296 26668 8336
rect 26708 8296 27340 8336
rect 27380 8296 27389 8336
rect 27907 8296 27916 8336
rect 27956 8296 32812 8336
rect 32852 8296 32861 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 24460 8252 24500 8296
rect 25996 8252 26036 8296
rect 26659 8252 26717 8253
rect 35596 8252 35636 8380
rect 35779 8296 35788 8336
rect 35828 8296 38956 8336
rect 38996 8296 40876 8336
rect 40916 8296 40925 8336
rect 41059 8296 41068 8336
rect 41108 8296 43948 8336
rect 43988 8296 43997 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 16579 8212 16588 8252
rect 16628 8212 17068 8252
rect 17108 8212 17836 8252
rect 17876 8212 20276 8252
rect 20323 8212 20332 8252
rect 20372 8212 22484 8252
rect 23011 8212 23020 8252
rect 23060 8212 24364 8252
rect 24404 8212 24413 8252
rect 24460 8212 24596 8252
rect 24643 8212 24652 8252
rect 24692 8212 25420 8252
rect 25460 8212 25469 8252
rect 25987 8212 25996 8252
rect 26036 8212 26045 8252
rect 26659 8212 26668 8252
rect 26708 8212 31852 8252
rect 31892 8212 33868 8252
rect 33908 8212 33917 8252
rect 34828 8212 35636 8252
rect 38755 8212 38764 8252
rect 38804 8212 42700 8252
rect 42740 8212 42749 8252
rect 0 8168 80 8188
rect 9475 8168 9533 8169
rect 23203 8168 23261 8169
rect 24556 8168 24596 8212
rect 26659 8211 26717 8212
rect 27523 8168 27581 8169
rect 34828 8168 34868 8212
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 1027 8128 1036 8168
rect 1076 8128 2860 8168
rect 2900 8128 2909 8168
rect 7459 8128 7468 8168
rect 7508 8128 8140 8168
rect 8180 8128 8524 8168
rect 8564 8128 8573 8168
rect 9379 8128 9388 8168
rect 9428 8128 9484 8168
rect 9524 8128 9533 8168
rect 15811 8128 15820 8168
rect 15860 8128 21140 8168
rect 21187 8128 21196 8168
rect 21236 8128 21676 8168
rect 21716 8128 21725 8168
rect 23118 8128 23212 8168
rect 23252 8128 23261 8168
rect 23491 8128 23500 8168
rect 23540 8128 24172 8168
rect 24212 8128 24221 8168
rect 24547 8128 24556 8168
rect 24596 8128 24605 8168
rect 27438 8128 27532 8168
rect 27572 8128 27581 8168
rect 28099 8128 28108 8168
rect 28148 8128 28876 8168
rect 28916 8128 28925 8168
rect 29827 8128 29836 8168
rect 29876 8128 30988 8168
rect 31028 8128 31037 8168
rect 34819 8128 34828 8168
rect 34868 8128 34877 8168
rect 35299 8128 35308 8168
rect 35348 8128 35596 8168
rect 35636 8128 35645 8168
rect 35875 8128 35884 8168
rect 35924 8128 36212 8168
rect 36252 8128 36261 8168
rect 36355 8128 36364 8168
rect 36404 8128 36413 8168
rect 39427 8128 39436 8168
rect 39476 8128 41068 8168
rect 41108 8128 41117 8168
rect 46627 8128 46636 8168
rect 46676 8128 46924 8168
rect 46964 8128 46973 8168
rect 0 8108 80 8128
rect 9475 8127 9533 8128
rect 20515 8084 20573 8085
rect 21100 8084 21140 8128
rect 23203 8127 23261 8128
rect 27523 8127 27581 8128
rect 36364 8084 36404 8128
rect 1411 8044 1420 8084
rect 1460 8044 3436 8084
rect 3476 8044 4396 8084
rect 4436 8044 4972 8084
rect 5012 8044 5021 8084
rect 11107 8044 11116 8084
rect 11156 8044 11692 8084
rect 11732 8044 11741 8084
rect 18499 8044 18508 8084
rect 18548 8044 20332 8084
rect 20372 8044 20524 8084
rect 20564 8044 20573 8084
rect 21091 8044 21100 8084
rect 21140 8044 23308 8084
rect 23348 8044 23692 8084
rect 23732 8044 23741 8084
rect 24460 8044 26572 8084
rect 26612 8044 26621 8084
rect 27244 8044 36404 8084
rect 39619 8044 39628 8084
rect 39668 8044 41452 8084
rect 41492 8044 41501 8084
rect 20515 8043 20573 8044
rect 1603 7960 1612 8000
rect 1652 7960 2860 8000
rect 2900 7960 2909 8000
rect 4867 7960 4876 8000
rect 4916 7960 5356 8000
rect 5396 7960 5836 8000
rect 5876 7960 5885 8000
rect 7459 7960 7468 8000
rect 7508 7960 7852 8000
rect 7892 7960 7901 8000
rect 9763 7960 9772 8000
rect 9812 7960 9964 8000
rect 10004 7960 10540 8000
rect 10580 7960 10589 8000
rect 14371 7960 14380 8000
rect 14420 7960 17260 8000
rect 17300 7960 18892 8000
rect 18932 7960 18941 8000
rect 20419 7960 20428 8000
rect 20468 7960 21484 8000
rect 21524 7960 21533 8000
rect 22435 7960 22444 8000
rect 22484 7960 23884 8000
rect 23924 7960 23933 8000
rect 20803 7916 20861 7917
rect 24460 7916 24500 8044
rect 27244 8000 27284 8044
rect 29827 8000 29885 8001
rect 24739 7960 24748 8000
rect 24788 7960 25420 8000
rect 25460 7960 26092 8000
rect 26132 7960 26141 8000
rect 26371 7960 26380 8000
rect 26420 7960 27052 8000
rect 27092 7960 27101 8000
rect 27235 7960 27244 8000
rect 27284 7960 27293 8000
rect 27427 7960 27436 8000
rect 27476 7960 27764 8000
rect 27811 7960 27820 8000
rect 27860 7960 29452 8000
rect 29492 7960 29501 8000
rect 29742 7960 29836 8000
rect 29876 7960 29885 8000
rect 30019 7960 30028 8000
rect 30068 7960 30604 8000
rect 30644 7960 30653 8000
rect 31651 7960 31660 8000
rect 31700 7960 34828 8000
rect 34868 7960 34877 8000
rect 35971 7960 35980 8000
rect 36020 7960 36940 8000
rect 36980 7960 36989 8000
rect 37891 7960 37900 8000
rect 37940 7960 38284 8000
rect 38324 7960 38333 8000
rect 40195 7960 40204 8000
rect 40244 7960 41260 8000
rect 41300 7960 41309 8000
rect 41560 7960 41932 8000
rect 41972 7960 42796 8000
rect 42836 7960 42845 8000
rect 27724 7916 27764 7960
rect 29827 7959 29885 7960
rect 41560 7916 41600 7960
rect 835 7876 844 7916
rect 884 7876 1708 7916
rect 1748 7876 1996 7916
rect 2036 7876 2045 7916
rect 5251 7876 5260 7916
rect 5300 7876 6028 7916
rect 6068 7876 6077 7916
rect 20227 7876 20236 7916
rect 20276 7876 20620 7916
rect 20660 7876 20669 7916
rect 20718 7876 20812 7916
rect 20852 7876 20861 7916
rect 20803 7875 20861 7876
rect 21004 7876 24500 7916
rect 24547 7876 24556 7916
rect 24596 7876 25228 7916
rect 25268 7876 25277 7916
rect 27724 7876 29000 7916
rect 30403 7876 30412 7916
rect 30452 7876 32140 7916
rect 32180 7876 35884 7916
rect 35924 7876 35933 7916
rect 36355 7876 36364 7916
rect 36404 7876 37036 7916
rect 37076 7876 37085 7916
rect 37780 7876 41600 7916
rect 21004 7832 21044 7876
rect 1123 7792 1132 7832
rect 1172 7792 2476 7832
rect 2516 7792 2525 7832
rect 20419 7792 20428 7832
rect 20468 7792 21004 7832
rect 21044 7792 21053 7832
rect 21964 7792 22676 7832
rect 22723 7792 22732 7832
rect 22772 7792 23980 7832
rect 24020 7792 24029 7832
rect 835 7708 844 7748
rect 884 7708 1804 7748
rect 1844 7708 1853 7748
rect 2851 7708 2860 7748
rect 2900 7708 3628 7748
rect 3668 7708 3677 7748
rect 8035 7708 8044 7748
rect 8084 7708 8428 7748
rect 8468 7708 9292 7748
rect 9332 7708 9341 7748
rect 14371 7708 14380 7748
rect 14420 7708 16204 7748
rect 16244 7708 16253 7748
rect 8995 7664 9053 7665
rect 21964 7664 22004 7792
rect 22636 7748 22676 7792
rect 28960 7748 29000 7876
rect 33571 7792 33580 7832
rect 33620 7792 34060 7832
rect 34100 7792 34109 7832
rect 34339 7792 34348 7832
rect 34388 7792 35116 7832
rect 35156 7792 35165 7832
rect 36451 7792 36460 7832
rect 36500 7792 36940 7832
rect 36980 7792 36989 7832
rect 22636 7708 24460 7748
rect 24500 7708 24509 7748
rect 25132 7708 27820 7748
rect 27860 7708 27869 7748
rect 28960 7708 36556 7748
rect 36596 7708 36605 7748
rect 25132 7664 25172 7708
rect 26755 7664 26813 7665
rect 37780 7664 37820 7876
rect 42979 7792 42988 7832
rect 43028 7792 43468 7832
rect 43508 7792 43517 7832
rect 8910 7624 9004 7664
rect 9044 7624 9053 7664
rect 20515 7624 20524 7664
rect 20564 7624 22004 7664
rect 22147 7624 22156 7664
rect 22196 7624 23596 7664
rect 23636 7624 23645 7664
rect 24259 7624 24268 7664
rect 24308 7624 24317 7664
rect 24643 7624 24652 7664
rect 24692 7624 25132 7664
rect 25172 7624 25181 7664
rect 25315 7624 25324 7664
rect 25364 7624 26381 7664
rect 26421 7624 26430 7664
rect 26670 7624 26764 7664
rect 26804 7624 26813 7664
rect 30115 7624 30124 7664
rect 30164 7624 35116 7664
rect 35156 7624 35165 7664
rect 35875 7624 35884 7664
rect 35924 7624 37820 7664
rect 8995 7623 9053 7624
rect 24268 7580 24308 7624
rect 26755 7623 26813 7624
rect 32131 7580 32189 7581
rect 32515 7580 32573 7581
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 8707 7540 8716 7580
rect 8756 7540 9100 7580
rect 9140 7540 9149 7580
rect 11491 7540 11500 7580
rect 11540 7540 11692 7580
rect 11732 7540 12940 7580
rect 12980 7540 13132 7580
rect 13172 7540 13181 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 18691 7540 18700 7580
rect 18740 7540 18749 7580
rect 22051 7540 22060 7580
rect 22100 7540 22732 7580
rect 22772 7540 22781 7580
rect 23011 7540 23020 7580
rect 23060 7540 24308 7580
rect 24547 7540 24556 7580
rect 24596 7540 26284 7580
rect 26324 7540 27820 7580
rect 27860 7540 27869 7580
rect 29059 7540 29068 7580
rect 29108 7540 30028 7580
rect 30068 7540 30220 7580
rect 30260 7540 30269 7580
rect 31651 7540 31660 7580
rect 31700 7540 32140 7580
rect 32180 7540 32189 7580
rect 32430 7540 32524 7580
rect 32564 7540 32573 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 34243 7540 34252 7580
rect 34292 7540 35692 7580
rect 35732 7540 35741 7580
rect 37795 7540 37804 7580
rect 37844 7540 38092 7580
rect 38132 7540 38572 7580
rect 38612 7540 38621 7580
rect 44035 7540 44044 7580
rect 44084 7540 46732 7580
rect 46772 7540 46924 7580
rect 46964 7540 46973 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 18700 7496 18740 7540
rect 32131 7539 32189 7540
rect 32515 7539 32573 7540
rect 23971 7496 24029 7497
rect 27619 7496 27677 7497
rect 35683 7496 35741 7497
rect 16579 7456 16588 7496
rect 16628 7456 17644 7496
rect 17684 7456 17693 7496
rect 18508 7456 22636 7496
rect 22676 7456 22685 7496
rect 22732 7456 23980 7496
rect 24020 7456 24029 7496
rect 24451 7456 24460 7496
rect 24500 7456 25516 7496
rect 25556 7456 25565 7496
rect 27619 7456 27628 7496
rect 27668 7456 30124 7496
rect 30164 7456 30508 7496
rect 30548 7456 30557 7496
rect 31075 7456 31084 7496
rect 31124 7456 35692 7496
rect 35732 7456 35741 7496
rect 18508 7412 18548 7456
rect 22732 7412 22772 7456
rect 23971 7455 24029 7456
rect 27619 7455 27677 7456
rect 31084 7412 31124 7456
rect 35683 7455 35741 7456
rect 8803 7372 8812 7412
rect 8852 7372 9580 7412
rect 9620 7372 9629 7412
rect 18499 7372 18508 7412
rect 18548 7372 18557 7412
rect 20419 7372 20428 7412
rect 20468 7372 22772 7412
rect 22915 7372 22924 7412
rect 22964 7372 25132 7412
rect 25172 7372 25181 7412
rect 27139 7372 27148 7412
rect 27188 7372 27628 7412
rect 27668 7372 27677 7412
rect 29347 7372 29356 7412
rect 29396 7372 31124 7412
rect 31171 7372 31180 7412
rect 31220 7372 31700 7412
rect 31747 7372 31756 7412
rect 31796 7372 32524 7412
rect 32564 7372 32573 7412
rect 34339 7372 34348 7412
rect 34388 7372 34540 7412
rect 34580 7372 34589 7412
rect 37315 7372 37324 7412
rect 37364 7372 37996 7412
rect 38036 7372 38045 7412
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 1219 7288 1228 7328
rect 1268 7288 2764 7328
rect 2804 7288 4012 7328
rect 4052 7288 4061 7328
rect 9196 7288 9388 7328
rect 9428 7288 9437 7328
rect 0 7268 80 7288
rect 9196 7244 9236 7288
rect 9187 7204 9196 7244
rect 9236 7204 9245 7244
rect 9580 7160 9620 7372
rect 30595 7328 30653 7329
rect 31660 7328 31700 7372
rect 21667 7288 21676 7328
rect 21716 7288 23212 7328
rect 23252 7288 23261 7328
rect 23395 7288 23404 7328
rect 23444 7288 24172 7328
rect 24212 7288 24460 7328
rect 24500 7288 24509 7328
rect 30019 7288 30028 7328
rect 30068 7288 30412 7328
rect 30452 7288 30461 7328
rect 30595 7288 30604 7328
rect 30644 7288 30700 7328
rect 30740 7288 30749 7328
rect 31651 7288 31660 7328
rect 31700 7288 31709 7328
rect 32131 7288 32140 7328
rect 32180 7288 32332 7328
rect 32372 7288 35788 7328
rect 35828 7288 35837 7328
rect 37411 7288 37420 7328
rect 37460 7288 38764 7328
rect 38804 7288 38813 7328
rect 41635 7288 41644 7328
rect 41684 7288 42700 7328
rect 42740 7288 42892 7328
rect 42932 7288 42941 7328
rect 30595 7287 30653 7288
rect 16867 7204 16876 7244
rect 16916 7204 18508 7244
rect 18548 7204 18557 7244
rect 22339 7204 22348 7244
rect 22388 7204 23116 7244
rect 23156 7204 23165 7244
rect 23299 7204 23308 7244
rect 23348 7204 24556 7244
rect 24596 7204 24605 7244
rect 24652 7204 28204 7244
rect 28244 7204 28253 7244
rect 28771 7204 28780 7244
rect 28820 7204 29260 7244
rect 29300 7204 29740 7244
rect 29780 7204 34636 7244
rect 34676 7204 34685 7244
rect 19075 7160 19133 7161
rect 23779 7160 23837 7161
rect 23971 7160 24029 7161
rect 24652 7160 24692 7204
rect 27139 7160 27197 7161
rect 30403 7160 30461 7161
rect 34147 7160 34205 7161
rect 34732 7160 34772 7288
rect 35011 7204 35020 7244
rect 35060 7204 35404 7244
rect 35444 7204 35453 7244
rect 37602 7204 37611 7244
rect 37651 7204 37900 7244
rect 37940 7204 37949 7244
rect 38083 7204 38092 7244
rect 38132 7204 38668 7244
rect 38708 7204 40588 7244
rect 40628 7204 40637 7244
rect 9379 7120 9388 7160
rect 9428 7120 9620 7160
rect 9667 7120 9676 7160
rect 9716 7120 12076 7160
rect 12116 7120 12844 7160
rect 12884 7120 12893 7160
rect 17539 7120 17548 7160
rect 17588 7120 18700 7160
rect 18740 7120 18749 7160
rect 18979 7120 18988 7160
rect 19028 7120 19084 7160
rect 19124 7120 19133 7160
rect 20515 7120 20524 7160
rect 20564 7120 20812 7160
rect 20852 7120 20861 7160
rect 22243 7120 22252 7160
rect 22292 7120 23596 7160
rect 23636 7120 23645 7160
rect 23779 7120 23788 7160
rect 23828 7120 23922 7160
rect 23971 7120 23980 7160
rect 24020 7120 24692 7160
rect 24739 7120 24748 7160
rect 24788 7120 25036 7160
rect 25076 7120 25324 7160
rect 25364 7120 26380 7160
rect 26420 7120 26429 7160
rect 27054 7120 27148 7160
rect 27188 7120 27197 7160
rect 27427 7120 27436 7160
rect 27476 7120 29548 7160
rect 29588 7120 29597 7160
rect 29836 7120 30412 7160
rect 30452 7120 32044 7160
rect 32084 7120 32093 7160
rect 32227 7120 32236 7160
rect 32276 7120 33196 7160
rect 33236 7120 33245 7160
rect 34062 7120 34156 7160
rect 34196 7120 34205 7160
rect 34531 7120 34540 7160
rect 34580 7120 34772 7160
rect 35299 7120 35308 7160
rect 35348 7120 35357 7160
rect 36835 7120 36844 7160
rect 36884 7120 38188 7160
rect 38228 7120 39436 7160
rect 39476 7120 39485 7160
rect 41923 7120 41932 7160
rect 41972 7120 43756 7160
rect 43796 7120 43805 7160
rect 19075 7119 19133 7120
rect 23779 7119 23837 7120
rect 23971 7119 24029 7120
rect 27139 7119 27197 7120
rect 18787 7076 18845 7077
rect 29836 7076 29876 7120
rect 30403 7119 30461 7120
rect 34147 7119 34205 7120
rect 17347 7036 17356 7076
rect 17396 7036 17932 7076
rect 17972 7036 18796 7076
rect 18836 7036 18845 7076
rect 20611 7036 20620 7076
rect 20660 7036 21004 7076
rect 21044 7036 21388 7076
rect 21428 7036 26572 7076
rect 26612 7036 26621 7076
rect 29740 7036 29876 7076
rect 34243 7076 34301 7077
rect 35308 7076 35348 7120
rect 43171 7076 43229 7077
rect 34243 7036 34252 7076
rect 34292 7036 35116 7076
rect 35156 7036 35165 7076
rect 35308 7036 35980 7076
rect 36020 7036 41260 7076
rect 41300 7036 41309 7076
rect 43086 7036 43180 7076
rect 43220 7036 43229 7076
rect 18787 7035 18845 7036
rect 29740 6992 29780 7036
rect 34243 7035 34301 7036
rect 43171 7035 43229 7036
rect 3523 6952 3532 6992
rect 3572 6952 4204 6992
rect 4244 6952 4253 6992
rect 4579 6952 4588 6992
rect 4628 6952 4637 6992
rect 6019 6952 6028 6992
rect 6068 6952 7948 6992
rect 7988 6952 7997 6992
rect 8323 6952 8332 6992
rect 8372 6952 8716 6992
rect 8756 6952 8765 6992
rect 9763 6952 9772 6992
rect 9812 6952 11404 6992
rect 11444 6952 11453 6992
rect 14659 6952 14668 6992
rect 14708 6952 15628 6992
rect 15668 6952 15677 6992
rect 16867 6952 16876 6992
rect 16916 6952 18796 6992
rect 18836 6952 19180 6992
rect 19220 6952 19229 6992
rect 22819 6952 22828 6992
rect 22868 6952 24081 6992
rect 24121 6952 24460 6992
rect 24500 6952 24509 6992
rect 27235 6952 27244 6992
rect 27284 6952 29780 6992
rect 29836 6952 35308 6992
rect 35348 6952 36268 6992
rect 36308 6952 36317 6992
rect 37603 6952 37612 6992
rect 37652 6952 40972 6992
rect 41012 6952 41021 6992
rect 43459 6952 43468 6992
rect 43508 6952 46828 6992
rect 46868 6952 46877 6992
rect 4588 6908 4628 6952
rect 23683 6908 23741 6909
rect 29836 6908 29876 6952
rect 4588 6868 9484 6908
rect 9524 6868 9533 6908
rect 16099 6868 16108 6908
rect 16148 6868 17164 6908
rect 17204 6868 19276 6908
rect 19316 6868 19325 6908
rect 19372 6868 22540 6908
rect 22580 6868 22589 6908
rect 23598 6868 23692 6908
rect 23732 6868 23741 6908
rect 27811 6868 27820 6908
rect 27860 6868 29836 6908
rect 29876 6868 29885 6908
rect 30307 6868 30316 6908
rect 30356 6868 30796 6908
rect 30836 6868 30845 6908
rect 32803 6868 32812 6908
rect 32852 6868 34004 6908
rect 34051 6868 34060 6908
rect 34100 6868 36748 6908
rect 36788 6868 36797 6908
rect 5548 6824 5588 6868
rect 19372 6824 19412 6868
rect 23683 6867 23741 6868
rect 24643 6824 24701 6825
rect 33964 6824 34004 6868
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 5539 6784 5548 6824
rect 5588 6784 5597 6824
rect 8332 6784 10156 6824
rect 10196 6784 10205 6824
rect 17443 6784 17452 6824
rect 17492 6784 19412 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 23203 6784 23212 6824
rect 23252 6784 24652 6824
rect 24692 6784 24701 6824
rect 29443 6784 29452 6824
rect 29492 6784 30220 6824
rect 30260 6784 30269 6824
rect 30700 6784 32524 6824
rect 32564 6784 33196 6824
rect 33236 6784 33245 6824
rect 33964 6784 34156 6824
rect 34196 6784 34348 6824
rect 34388 6784 34397 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 35020 6784 35980 6824
rect 36020 6784 36029 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 8332 6656 8372 6784
rect 24643 6783 24701 6784
rect 30595 6740 30653 6741
rect 9571 6700 9580 6740
rect 9620 6700 10060 6740
rect 10100 6700 10109 6740
rect 17827 6700 17836 6740
rect 17876 6700 19796 6740
rect 28387 6700 28396 6740
rect 28436 6700 29356 6740
rect 29396 6700 29405 6740
rect 30115 6700 30124 6740
rect 30164 6700 30604 6740
rect 30644 6700 30653 6740
rect 19756 6656 19796 6700
rect 30595 6699 30653 6700
rect 24259 6656 24317 6657
rect 30700 6656 30740 6784
rect 35020 6740 35060 6784
rect 30787 6700 30796 6740
rect 30836 6700 31276 6740
rect 31316 6700 35060 6740
rect 37891 6700 37900 6740
rect 37940 6700 38572 6740
rect 38612 6700 38621 6740
rect 8323 6616 8332 6656
rect 8372 6616 8381 6656
rect 10147 6616 10156 6656
rect 10196 6616 11116 6656
rect 11156 6616 11165 6656
rect 16291 6616 16300 6656
rect 16340 6616 19468 6656
rect 19508 6616 19517 6656
rect 19747 6616 19756 6656
rect 19796 6616 19805 6656
rect 23107 6616 23116 6656
rect 23156 6616 23788 6656
rect 23828 6616 23837 6656
rect 24259 6616 24268 6656
rect 24308 6616 24940 6656
rect 24980 6616 30740 6656
rect 30883 6616 30892 6656
rect 30932 6616 34636 6656
rect 34676 6616 35020 6656
rect 35060 6616 35069 6656
rect 36067 6616 36076 6656
rect 36116 6616 36748 6656
rect 36788 6616 36797 6656
rect 24259 6615 24317 6616
rect 18883 6572 18941 6573
rect 24451 6572 24509 6573
rect 27715 6572 27773 6573
rect 32035 6572 32093 6573
rect 8803 6532 8812 6572
rect 8852 6532 9004 6572
rect 9044 6532 9053 6572
rect 18883 6532 18892 6572
rect 18932 6532 19026 6572
rect 22819 6532 22828 6572
rect 22868 6532 23500 6572
rect 23540 6532 24460 6572
rect 24500 6532 24509 6572
rect 27619 6532 27628 6572
rect 27668 6532 27724 6572
rect 27764 6532 27773 6572
rect 31363 6532 31372 6572
rect 31412 6532 31756 6572
rect 31796 6532 31805 6572
rect 31939 6532 31948 6572
rect 31988 6532 32044 6572
rect 32084 6532 32093 6572
rect 18883 6531 18941 6532
rect 24451 6531 24509 6532
rect 27715 6531 27773 6532
rect 32035 6531 32093 6532
rect 32227 6572 32285 6573
rect 34147 6572 34205 6573
rect 32227 6532 32236 6572
rect 32276 6532 32332 6572
rect 32372 6532 32381 6572
rect 34147 6532 34156 6572
rect 34196 6532 34732 6572
rect 34772 6532 34781 6572
rect 35587 6532 35596 6572
rect 35636 6532 35788 6572
rect 35828 6532 36884 6572
rect 37315 6532 37324 6572
rect 37364 6532 37516 6572
rect 37556 6532 37820 6572
rect 32227 6531 32285 6532
rect 34147 6531 34205 6532
rect 0 6488 80 6508
rect 9475 6488 9533 6489
rect 27619 6488 27677 6489
rect 35683 6488 35741 6489
rect 36844 6488 36884 6532
rect 37780 6488 37820 6532
rect 44716 6532 46252 6572
rect 46292 6532 46301 6572
rect 44716 6489 44756 6532
rect 44707 6488 44765 6489
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 2851 6448 2860 6488
rect 2900 6448 4012 6488
rect 4052 6448 4492 6488
rect 4532 6448 4541 6488
rect 7075 6448 7084 6488
rect 7124 6448 8372 6488
rect 8419 6448 8428 6488
rect 8468 6448 9100 6488
rect 9140 6448 9149 6488
rect 9390 6448 9484 6488
rect 9524 6448 9533 6488
rect 10243 6448 10252 6488
rect 10292 6448 11884 6488
rect 11924 6448 11933 6488
rect 12931 6448 12940 6488
rect 12980 6448 14668 6488
rect 14708 6448 14717 6488
rect 16387 6448 16396 6488
rect 16436 6448 16780 6488
rect 16820 6448 16829 6488
rect 19075 6448 19084 6488
rect 19124 6448 20524 6488
rect 20564 6448 20573 6488
rect 22723 6448 22732 6488
rect 22772 6448 23116 6488
rect 23156 6448 23165 6488
rect 23875 6448 23884 6488
rect 23924 6448 24268 6488
rect 24308 6448 24317 6488
rect 27523 6448 27532 6488
rect 27572 6448 27628 6488
rect 27668 6448 27677 6488
rect 28195 6448 28204 6488
rect 28244 6448 28588 6488
rect 28628 6448 28972 6488
rect 29012 6448 29021 6488
rect 29155 6448 29164 6488
rect 29204 6448 30892 6488
rect 30932 6448 30941 6488
rect 31459 6448 31468 6488
rect 31508 6448 32716 6488
rect 32756 6448 32765 6488
rect 35011 6448 35020 6488
rect 35060 6448 35692 6488
rect 35732 6448 35741 6488
rect 35875 6448 35884 6488
rect 35924 6448 35933 6488
rect 36835 6448 36844 6488
rect 36884 6448 37612 6488
rect 37652 6448 37661 6488
rect 37780 6448 38572 6488
rect 38612 6448 40684 6488
rect 40724 6448 40733 6488
rect 41251 6448 41260 6488
rect 41300 6448 41644 6488
rect 41684 6448 41693 6488
rect 44515 6448 44524 6488
rect 44564 6448 44573 6488
rect 44622 6448 44716 6488
rect 44756 6448 44765 6488
rect 45283 6448 45292 6488
rect 45332 6448 47116 6488
rect 47156 6448 47165 6488
rect 0 6428 80 6448
rect 8332 6404 8372 6448
rect 9475 6447 9533 6448
rect 27619 6447 27677 6448
rect 35683 6447 35741 6448
rect 22627 6404 22685 6405
rect 23395 6404 23453 6405
rect 35884 6404 35924 6448
rect 42211 6404 42269 6405
rect 5155 6364 5164 6404
rect 5204 6364 7468 6404
rect 7508 6364 7517 6404
rect 8323 6364 8332 6404
rect 8372 6364 8381 6404
rect 18115 6364 18124 6404
rect 18164 6364 19852 6404
rect 19892 6364 21484 6404
rect 21524 6364 21533 6404
rect 22542 6364 22636 6404
rect 22676 6364 23212 6404
rect 23252 6364 23261 6404
rect 23310 6364 23404 6404
rect 23444 6364 23453 6404
rect 23971 6364 23980 6404
rect 24020 6364 24748 6404
rect 24788 6364 24797 6404
rect 26563 6364 26572 6404
rect 26612 6364 29548 6404
rect 29588 6364 29597 6404
rect 29731 6364 29740 6404
rect 29780 6364 33908 6404
rect 35884 6364 37804 6404
rect 37844 6364 37853 6404
rect 42019 6364 42028 6404
rect 42068 6364 42220 6404
rect 42260 6364 42269 6404
rect 22627 6363 22685 6364
rect 23395 6363 23453 6364
rect 24259 6320 24317 6321
rect 33868 6320 33908 6364
rect 42211 6363 42269 6364
rect 43171 6404 43229 6405
rect 44524 6404 44564 6448
rect 44707 6447 44765 6448
rect 43171 6364 43180 6404
rect 43220 6364 44756 6404
rect 43171 6363 43229 6364
rect 44716 6320 44756 6364
rect 4195 6280 4204 6320
rect 4244 6280 4972 6320
rect 5012 6280 6028 6320
rect 6068 6280 6077 6320
rect 6595 6280 6604 6320
rect 6644 6280 6796 6320
rect 6836 6280 7372 6320
rect 7412 6280 7421 6320
rect 8227 6280 8236 6320
rect 8276 6280 8428 6320
rect 8468 6280 8477 6320
rect 9187 6280 9196 6320
rect 9236 6280 9676 6320
rect 9716 6280 10060 6320
rect 10100 6280 10109 6320
rect 22819 6280 22828 6320
rect 22868 6280 23692 6320
rect 23732 6280 23741 6320
rect 24163 6280 24172 6320
rect 24212 6280 24268 6320
rect 24308 6280 24317 6320
rect 24547 6280 24556 6320
rect 24596 6280 27436 6320
rect 27476 6280 27485 6320
rect 29635 6280 29644 6320
rect 29684 6280 31564 6320
rect 31604 6280 31613 6320
rect 32034 6280 32043 6320
rect 32083 6280 33196 6320
rect 33236 6280 33245 6320
rect 33859 6280 33868 6320
rect 33908 6280 35308 6320
rect 35348 6280 35788 6320
rect 35828 6280 35837 6320
rect 36067 6280 36076 6320
rect 36116 6280 37820 6320
rect 44707 6280 44716 6320
rect 44756 6280 44765 6320
rect 24259 6279 24317 6280
rect 32515 6236 32573 6237
rect 37780 6236 37820 6280
rect 7171 6196 7180 6236
rect 7220 6196 9292 6236
rect 9332 6196 9341 6236
rect 17923 6196 17932 6236
rect 17972 6196 22060 6236
rect 22100 6196 22109 6236
rect 23011 6196 23020 6236
rect 23060 6196 24268 6236
rect 24308 6196 24317 6236
rect 31651 6196 31660 6236
rect 31700 6196 32524 6236
rect 32564 6196 33004 6236
rect 33044 6196 33053 6236
rect 35395 6196 35404 6236
rect 35444 6196 36940 6236
rect 36980 6196 36989 6236
rect 37780 6196 37900 6236
rect 37940 6196 37949 6236
rect 32515 6195 32573 6196
rect 17251 6112 17260 6152
rect 17300 6112 19564 6152
rect 19604 6112 19613 6152
rect 19747 6112 19756 6152
rect 19796 6112 20812 6152
rect 20852 6112 20861 6152
rect 32044 6112 32428 6152
rect 32468 6112 32477 6152
rect 32611 6112 32620 6152
rect 32660 6112 32812 6152
rect 32852 6112 32861 6152
rect 33091 6112 33100 6152
rect 33140 6112 37820 6152
rect 18979 6068 19037 6069
rect 32044 6068 32084 6112
rect 32227 6068 32285 6069
rect 32899 6068 32957 6069
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 18979 6028 18988 6068
rect 19028 6028 19988 6068
rect 32035 6028 32044 6068
rect 32084 6028 32093 6068
rect 32227 6028 32236 6068
rect 32276 6028 32908 6068
rect 32948 6028 32957 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 18979 6027 19037 6028
rect 19363 5984 19421 5985
rect 19948 5984 19988 6028
rect 32227 6027 32285 6028
rect 32899 6027 32957 6028
rect 26563 5984 26621 5985
rect 17347 5944 17356 5984
rect 17396 5944 19372 5984
rect 19412 5944 19421 5984
rect 19939 5944 19948 5984
rect 19988 5944 26572 5984
rect 26612 5944 26621 5984
rect 30595 5944 30604 5984
rect 30644 5944 31084 5984
rect 31124 5944 31133 5984
rect 31939 5944 31948 5984
rect 31988 5944 32620 5984
rect 32660 5944 32669 5984
rect 34531 5944 34540 5984
rect 34580 5944 34828 5984
rect 34868 5944 35692 5984
rect 35732 5944 35741 5984
rect 19363 5943 19421 5944
rect 26563 5943 26621 5944
rect 37780 5900 37820 6112
rect 39907 6028 39916 6068
rect 39956 6028 42220 6068
rect 42260 6028 44236 6068
rect 44276 6028 45004 6068
rect 45044 6028 45053 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 15811 5860 15820 5900
rect 15860 5860 17452 5900
rect 17492 5860 17501 5900
rect 18883 5860 18892 5900
rect 18932 5860 19180 5900
rect 19220 5860 19229 5900
rect 26371 5860 26380 5900
rect 26420 5860 36308 5900
rect 37780 5860 39532 5900
rect 39572 5860 41644 5900
rect 41684 5860 41693 5900
rect 7747 5816 7805 5817
rect 7459 5776 7468 5816
rect 7508 5776 7756 5816
rect 7796 5776 7805 5816
rect 8995 5776 9004 5816
rect 9044 5776 9868 5816
rect 9908 5776 9917 5816
rect 16195 5776 16204 5816
rect 16244 5776 16340 5816
rect 16675 5776 16684 5816
rect 16724 5776 18988 5816
rect 19028 5776 19037 5816
rect 19267 5776 19276 5816
rect 19316 5776 19852 5816
rect 19892 5776 19901 5816
rect 20035 5776 20044 5816
rect 20084 5776 20093 5816
rect 21379 5776 21388 5816
rect 21428 5776 22732 5816
rect 22772 5776 22781 5816
rect 23971 5776 23980 5816
rect 24020 5776 29000 5816
rect 31171 5776 31180 5816
rect 31220 5776 31564 5816
rect 31604 5776 31613 5816
rect 31843 5776 31852 5816
rect 31892 5776 32524 5816
rect 32564 5776 33484 5816
rect 33524 5776 33533 5816
rect 35395 5776 35404 5816
rect 35444 5776 35453 5816
rect 7747 5775 7805 5776
rect 0 5648 80 5668
rect 0 5608 1036 5648
rect 1076 5608 1085 5648
rect 4771 5608 4780 5648
rect 4820 5608 5452 5648
rect 5492 5608 5501 5648
rect 7363 5608 7372 5648
rect 7412 5608 7660 5648
rect 7700 5608 7709 5648
rect 7939 5608 7948 5648
rect 7988 5608 8140 5648
rect 8180 5608 9393 5648
rect 9433 5608 9442 5648
rect 11971 5608 11980 5648
rect 12020 5608 13132 5648
rect 13172 5608 13181 5648
rect 0 5588 80 5608
rect 8899 5564 8957 5565
rect 16300 5564 16340 5776
rect 20044 5732 20084 5776
rect 28960 5732 29000 5776
rect 35404 5732 35444 5776
rect 16973 5692 16982 5732
rect 17022 5692 20084 5732
rect 22435 5692 22444 5732
rect 22484 5692 24844 5732
rect 24884 5692 24893 5732
rect 28960 5692 35444 5732
rect 26563 5648 26621 5649
rect 16771 5608 16780 5648
rect 16820 5608 17548 5648
rect 17588 5608 17597 5648
rect 19651 5608 19660 5648
rect 19700 5608 19709 5648
rect 23587 5608 23596 5648
rect 23636 5608 24076 5648
rect 24116 5608 24125 5648
rect 24355 5608 24364 5648
rect 24404 5608 24413 5648
rect 26563 5608 26572 5648
rect 26612 5608 26860 5648
rect 26900 5608 26909 5648
rect 27907 5608 27916 5648
rect 27956 5608 28492 5648
rect 28532 5608 28541 5648
rect 28963 5608 28972 5648
rect 29012 5608 29052 5648
rect 30211 5608 30220 5648
rect 30260 5608 31084 5648
rect 31124 5608 31133 5648
rect 31939 5608 31948 5648
rect 31988 5608 33004 5648
rect 33044 5608 33053 5648
rect 34915 5608 34924 5648
rect 34964 5608 35212 5648
rect 35252 5608 35261 5648
rect 35395 5608 35404 5648
rect 35444 5608 35980 5648
rect 36020 5608 36029 5648
rect 19660 5564 19700 5608
rect 24364 5564 24404 5608
rect 26563 5607 26621 5608
rect 28972 5565 29012 5608
rect 28963 5564 29021 5565
rect 32131 5564 32189 5565
rect 7459 5524 7468 5564
rect 7508 5524 7756 5564
rect 7796 5524 7805 5564
rect 8899 5524 8908 5564
rect 8948 5524 9042 5564
rect 12163 5524 12172 5564
rect 12212 5524 12940 5564
rect 12980 5524 15532 5564
rect 15572 5524 15581 5564
rect 16300 5524 19700 5564
rect 21571 5524 21580 5564
rect 21620 5524 22348 5564
rect 22388 5524 23788 5564
rect 23828 5524 24404 5564
rect 26440 5524 28972 5564
rect 29012 5524 29021 5564
rect 32046 5524 32140 5564
rect 32180 5524 35500 5564
rect 35540 5524 35549 5564
rect 8899 5523 8957 5524
rect 26440 5480 26480 5524
rect 28963 5523 29021 5524
rect 32131 5523 32189 5524
rect 36268 5480 36308 5860
rect 36355 5776 36364 5816
rect 36404 5776 38380 5816
rect 38420 5776 38429 5816
rect 38467 5692 38476 5732
rect 38516 5692 40780 5732
rect 40820 5692 40829 5732
rect 37123 5608 37132 5648
rect 37172 5608 37612 5648
rect 37652 5608 37661 5648
rect 38659 5608 38668 5648
rect 38708 5608 40876 5648
rect 40916 5608 40925 5648
rect 41827 5608 41836 5648
rect 41876 5608 42604 5648
rect 42644 5608 42653 5648
rect 43267 5608 43276 5648
rect 43316 5608 43948 5648
rect 43988 5608 44908 5648
rect 44948 5608 45580 5648
rect 45620 5608 45629 5648
rect 36643 5524 36652 5564
rect 36692 5524 38860 5564
rect 38900 5524 38909 5564
rect 43651 5524 43660 5564
rect 43700 5524 44812 5564
rect 44852 5524 44861 5564
rect 4195 5440 4204 5480
rect 4244 5440 5068 5480
rect 5108 5440 5117 5480
rect 7171 5440 7180 5480
rect 7220 5440 8428 5480
rect 8468 5440 8477 5480
rect 9091 5440 9100 5480
rect 9140 5440 9772 5480
rect 9812 5440 9821 5480
rect 14179 5440 14188 5480
rect 14228 5440 18508 5480
rect 18548 5440 18557 5480
rect 18883 5440 18892 5480
rect 18932 5440 23116 5480
rect 23156 5440 23165 5480
rect 26371 5440 26380 5480
rect 26420 5440 26480 5480
rect 27811 5440 27820 5480
rect 27860 5440 28780 5480
rect 28820 5440 28829 5480
rect 28963 5440 28972 5480
rect 29012 5440 29260 5480
rect 29300 5440 29740 5480
rect 29780 5440 29789 5480
rect 30499 5440 30508 5480
rect 30548 5440 32332 5480
rect 32372 5440 32381 5480
rect 35011 5440 35020 5480
rect 35060 5440 36172 5480
rect 36212 5440 36221 5480
rect 36268 5440 40492 5480
rect 40532 5440 40820 5480
rect 30691 5396 30749 5397
rect 40780 5396 40820 5440
rect 9379 5356 9388 5396
rect 9428 5356 9676 5396
rect 9716 5356 9725 5396
rect 16195 5356 16204 5396
rect 16244 5356 16972 5396
rect 17012 5356 19084 5396
rect 19124 5356 19133 5396
rect 23299 5356 23308 5396
rect 23348 5356 23596 5396
rect 23636 5356 26284 5396
rect 26324 5356 30700 5396
rect 30740 5356 32620 5396
rect 32660 5356 32669 5396
rect 38179 5356 38188 5396
rect 38228 5356 39820 5396
rect 39860 5356 39869 5396
rect 40771 5356 40780 5396
rect 40820 5356 40829 5396
rect 30691 5355 30749 5356
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 17923 5272 17932 5312
rect 17972 5272 19372 5312
rect 19412 5272 19421 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 23011 5272 23020 5312
rect 23060 5272 23692 5312
rect 23732 5272 23741 5312
rect 29539 5272 29548 5312
rect 29588 5272 32236 5312
rect 32276 5272 32285 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 4684 5188 5164 5228
rect 5204 5188 5213 5228
rect 16396 5188 18604 5228
rect 18644 5188 20908 5228
rect 20948 5188 20957 5228
rect 28771 5188 28780 5228
rect 28820 5188 29836 5228
rect 29876 5188 29885 5228
rect 4684 5144 4724 5188
rect 16396 5144 16436 5188
rect 4675 5104 4684 5144
rect 4724 5104 4733 5144
rect 8803 5104 8812 5144
rect 8852 5104 9196 5144
rect 9236 5104 9245 5144
rect 13027 5104 13036 5144
rect 13076 5104 16396 5144
rect 16436 5104 16445 5144
rect 17731 5104 17740 5144
rect 17780 5104 17789 5144
rect 21475 5104 21484 5144
rect 21524 5104 21533 5144
rect 28099 5104 28108 5144
rect 28148 5104 29164 5144
rect 29204 5104 29213 5144
rect 30403 5104 30412 5144
rect 30452 5104 30644 5144
rect 37795 5104 37804 5144
rect 37844 5104 38284 5144
rect 38324 5104 38333 5144
rect 17251 5060 17309 5061
rect 3715 5020 3724 5060
rect 3764 5020 5164 5060
rect 5204 5020 5213 5060
rect 9571 5020 9580 5060
rect 9620 5020 10348 5060
rect 10388 5020 10397 5060
rect 16003 5020 16012 5060
rect 16052 5020 17068 5060
rect 17108 5020 17117 5060
rect 17251 5020 17260 5060
rect 17300 5020 17394 5060
rect 17251 5019 17309 5020
rect 7747 4976 7805 4977
rect 17740 4976 17780 5104
rect 21484 5060 21524 5104
rect 21763 5060 21821 5061
rect 17827 5020 17836 5060
rect 17876 5020 18892 5060
rect 18932 5020 18941 5060
rect 21484 5020 21772 5060
rect 21812 5020 21821 5060
rect 21763 5019 21821 5020
rect 23011 5060 23069 5061
rect 24451 5060 24509 5061
rect 24643 5060 24701 5061
rect 28003 5060 28061 5061
rect 30604 5060 30644 5104
rect 23011 5020 23020 5060
rect 23060 5020 23299 5060
rect 23339 5020 23348 5060
rect 23395 5020 23404 5060
rect 23444 5020 23884 5060
rect 23924 5020 23933 5060
rect 24366 5020 24460 5060
rect 24500 5020 24509 5060
rect 24558 5020 24652 5060
rect 24692 5020 24701 5060
rect 24835 5020 24844 5060
rect 24884 5020 28012 5060
rect 28052 5020 28061 5060
rect 28291 5020 28300 5060
rect 28340 5020 29835 5060
rect 29875 5020 29884 5060
rect 30019 5020 30028 5060
rect 30068 5020 30508 5060
rect 30548 5020 30557 5060
rect 30604 5020 30988 5060
rect 31028 5020 31604 5060
rect 32707 5020 32716 5060
rect 32756 5020 34924 5060
rect 34964 5020 34973 5060
rect 35107 5020 35116 5060
rect 35156 5020 37420 5060
rect 37460 5020 38668 5060
rect 38708 5020 39628 5060
rect 39668 5020 39677 5060
rect 23011 5019 23069 5020
rect 24451 5019 24509 5020
rect 24643 5019 24701 5020
rect 28003 5019 28061 5020
rect 21571 4976 21629 4977
rect 31564 4976 31604 5020
rect 31939 4976 31997 4977
rect 34339 4976 34397 4977
rect 2947 4936 2956 4976
rect 2996 4936 5548 4976
rect 5588 4936 5597 4976
rect 6595 4936 6604 4976
rect 6644 4936 7372 4976
rect 7412 4936 7421 4976
rect 7662 4936 7756 4976
rect 7796 4936 7805 4976
rect 8707 4936 8716 4976
rect 8756 4936 9196 4976
rect 9236 4936 9245 4976
rect 9667 4936 9676 4976
rect 9716 4936 10156 4976
rect 10196 4936 10540 4976
rect 10580 4936 13324 4976
rect 13364 4936 13373 4976
rect 15100 4936 16108 4976
rect 16148 4936 18028 4976
rect 18068 4936 18077 4976
rect 19267 4936 19276 4976
rect 19316 4936 21388 4976
rect 21428 4936 21437 4976
rect 21571 4936 21580 4976
rect 21620 4936 21671 4976
rect 21711 4936 21720 4976
rect 21763 4936 21772 4976
rect 21812 4936 26476 4976
rect 26516 4936 26525 4976
rect 26851 4936 26860 4976
rect 26900 4936 27244 4976
rect 27284 4936 27293 4976
rect 28867 4936 28876 4976
rect 28916 4936 29260 4976
rect 29300 4936 29309 4976
rect 29443 4936 29452 4976
rect 29492 4936 29740 4976
rect 29780 4936 29789 4976
rect 29923 4936 29932 4976
rect 29972 4936 31084 4976
rect 31124 4936 31133 4976
rect 31555 4936 31564 4976
rect 31604 4936 31948 4976
rect 31988 4936 31997 4976
rect 34243 4936 34252 4976
rect 34292 4936 34348 4976
rect 34388 4936 34397 4976
rect 36355 4936 36364 4976
rect 36404 4936 38380 4976
rect 38420 4936 38429 4976
rect 38755 4936 38764 4976
rect 38804 4936 39244 4976
rect 39284 4936 39293 4976
rect 7747 4935 7805 4936
rect 4195 4852 4204 4892
rect 4244 4852 4684 4892
rect 4724 4852 4733 4892
rect 8803 4852 8812 4892
rect 8852 4852 10444 4892
rect 10484 4852 10493 4892
rect 0 4808 80 4828
rect 15100 4808 15140 4936
rect 21571 4935 21629 4936
rect 31939 4935 31997 4936
rect 18883 4892 18941 4893
rect 30307 4892 30365 4893
rect 34252 4892 34292 4936
rect 34339 4935 34397 4936
rect 16387 4852 16396 4892
rect 16436 4852 17548 4892
rect 17588 4852 17597 4892
rect 17731 4852 17740 4892
rect 17780 4852 18892 4892
rect 18932 4852 18988 4892
rect 19028 4852 19037 4892
rect 20131 4852 20140 4892
rect 20180 4852 20524 4892
rect 20564 4852 20573 4892
rect 20899 4852 20908 4892
rect 20948 4852 23116 4892
rect 23156 4852 24268 4892
rect 24308 4852 24317 4892
rect 25996 4852 26668 4892
rect 26708 4852 26717 4892
rect 28387 4852 28396 4892
rect 28436 4852 29356 4892
rect 29396 4852 29644 4892
rect 29684 4852 29693 4892
rect 30222 4852 30316 4892
rect 30356 4852 30365 4892
rect 31459 4852 31468 4892
rect 31508 4852 34292 4892
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 10051 4768 10060 4808
rect 10100 4768 10348 4808
rect 10388 4768 10397 4808
rect 11320 4768 11596 4808
rect 11636 4768 11645 4808
rect 14179 4768 14188 4808
rect 14228 4768 15140 4808
rect 17548 4808 17588 4852
rect 18883 4851 18941 4852
rect 25996 4808 26036 4852
rect 26668 4808 26708 4852
rect 30307 4851 30365 4852
rect 30883 4808 30941 4809
rect 17548 4768 17836 4808
rect 17876 4768 17885 4808
rect 19363 4768 19372 4808
rect 19412 4768 23212 4808
rect 23252 4768 23261 4808
rect 23788 4768 26036 4808
rect 26083 4768 26092 4808
rect 26132 4768 26284 4808
rect 26324 4768 26333 4808
rect 26668 4768 27148 4808
rect 27188 4768 27197 4808
rect 27331 4768 27340 4808
rect 27380 4768 29068 4808
rect 29108 4768 29117 4808
rect 30798 4768 30892 4808
rect 30932 4768 30941 4808
rect 32803 4768 32812 4808
rect 32852 4768 33676 4808
rect 33716 4768 33725 4808
rect 0 4748 80 4768
rect 4291 4684 4300 4724
rect 4340 4684 5932 4724
rect 5972 4684 5981 4724
rect 8995 4640 9053 4641
rect 11320 4640 11360 4768
rect 19372 4724 19412 4768
rect 23788 4724 23828 4768
rect 30883 4767 30941 4768
rect 25027 4724 25085 4725
rect 27619 4724 27677 4725
rect 28963 4724 29021 4725
rect 32899 4724 32957 4725
rect 18691 4684 18700 4724
rect 18740 4684 19412 4724
rect 20140 4684 23788 4724
rect 23828 4684 23837 4724
rect 24942 4684 25036 4724
rect 25076 4684 25085 4724
rect 8910 4600 9004 4640
rect 9044 4600 11360 4640
rect 17731 4640 17789 4641
rect 20140 4640 20180 4684
rect 25027 4683 25085 4684
rect 25132 4684 27628 4724
rect 27668 4684 28204 4724
rect 28244 4684 28253 4724
rect 28963 4684 28972 4724
rect 29012 4684 29106 4724
rect 32814 4684 32908 4724
rect 32948 4684 32957 4724
rect 25132 4640 25172 4684
rect 27619 4683 27677 4684
rect 28963 4683 29021 4684
rect 32899 4683 32957 4684
rect 17731 4600 17740 4640
rect 17780 4600 20180 4640
rect 23491 4600 23500 4640
rect 23540 4600 25172 4640
rect 25411 4600 25420 4640
rect 25460 4600 26516 4640
rect 27907 4600 27916 4640
rect 27956 4600 28780 4640
rect 28820 4600 29452 4640
rect 29492 4600 29501 4640
rect 8995 4599 9053 4600
rect 17731 4599 17789 4600
rect 26371 4556 26429 4557
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 20611 4516 20620 4556
rect 20660 4516 21100 4556
rect 21140 4516 23596 4556
rect 23636 4516 23645 4556
rect 24931 4516 24940 4556
rect 24980 4516 26380 4556
rect 26420 4516 26429 4556
rect 26476 4556 26516 4600
rect 31843 4556 31901 4557
rect 26476 4516 31700 4556
rect 31758 4516 31852 4556
rect 31892 4516 31901 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 26371 4515 26429 4516
rect 29539 4472 29597 4473
rect 16387 4432 16396 4472
rect 16436 4432 20236 4472
rect 20276 4432 20908 4472
rect 20948 4432 20957 4472
rect 27619 4432 27628 4472
rect 27668 4432 28108 4472
rect 28148 4432 28157 4472
rect 28960 4432 29548 4472
rect 29588 4432 29597 4472
rect 31660 4472 31700 4516
rect 31843 4515 31901 4516
rect 31660 4432 34540 4472
rect 34580 4432 34589 4472
rect 15811 4388 15869 4389
rect 28960 4388 29000 4432
rect 29539 4431 29597 4432
rect 11587 4348 11596 4388
rect 11636 4348 15820 4388
rect 15860 4348 15869 4388
rect 17251 4348 17260 4388
rect 17300 4348 17740 4388
rect 17780 4348 18508 4388
rect 18548 4348 18557 4388
rect 20140 4348 21196 4388
rect 21236 4348 22924 4388
rect 22964 4348 22973 4388
rect 23020 4348 25420 4388
rect 25460 4348 25469 4388
rect 26380 4348 28684 4388
rect 28724 4348 29000 4388
rect 33859 4348 33868 4388
rect 33908 4348 34252 4388
rect 34292 4348 34301 4388
rect 15811 4347 15869 4348
rect 19075 4304 19133 4305
rect 20140 4304 20180 4348
rect 9859 4264 9868 4304
rect 9908 4264 10252 4304
rect 10292 4264 10540 4304
rect 10580 4264 11020 4304
rect 11060 4264 11500 4304
rect 11540 4264 11788 4304
rect 11828 4264 11980 4304
rect 12020 4264 13420 4304
rect 13460 4264 13469 4304
rect 17155 4264 17164 4304
rect 17204 4264 17356 4304
rect 17396 4264 17644 4304
rect 17684 4264 17693 4304
rect 17827 4264 17836 4304
rect 17876 4264 19084 4304
rect 19124 4264 20180 4304
rect 20323 4304 20381 4305
rect 23020 4304 23060 4348
rect 25315 4304 25373 4305
rect 20323 4264 20332 4304
rect 20372 4264 20466 4304
rect 20899 4264 20908 4304
rect 20948 4264 23060 4304
rect 23587 4264 23596 4304
rect 23636 4264 24076 4304
rect 24116 4264 24844 4304
rect 24884 4264 24893 4304
rect 25230 4264 25324 4304
rect 25364 4264 25373 4304
rect 19075 4263 19133 4264
rect 20323 4263 20381 4264
rect 25315 4263 25373 4264
rect 26380 4220 26420 4348
rect 26467 4304 26525 4305
rect 26467 4264 26476 4304
rect 26516 4264 37228 4304
rect 37268 4264 37277 4304
rect 26467 4263 26525 4264
rect 10435 4180 10444 4220
rect 10484 4180 10924 4220
rect 10964 4180 11404 4220
rect 11444 4180 11884 4220
rect 11924 4180 11933 4220
rect 12163 4180 12172 4220
rect 12212 4180 16396 4220
rect 16436 4180 16445 4220
rect 16579 4180 16588 4220
rect 16628 4180 18220 4220
rect 18260 4180 18269 4220
rect 18403 4180 18412 4220
rect 18452 4180 19084 4220
rect 19124 4180 19133 4220
rect 20035 4180 20044 4220
rect 20084 4180 20372 4220
rect 22723 4180 22732 4220
rect 22772 4180 25900 4220
rect 25940 4180 25949 4220
rect 26371 4180 26380 4220
rect 26420 4180 26429 4220
rect 29539 4180 29548 4220
rect 29588 4180 30988 4220
rect 31028 4180 32716 4220
rect 32756 4180 32765 4220
rect 20332 4136 20372 4180
rect 5539 4096 5548 4136
rect 5588 4096 6604 4136
rect 6644 4096 6653 4136
rect 11779 4096 11788 4136
rect 11828 4096 13132 4136
rect 13172 4096 13181 4136
rect 13315 4096 13324 4136
rect 13364 4096 13612 4136
rect 13652 4096 13661 4136
rect 15331 4096 15340 4136
rect 15380 4096 16492 4136
rect 16532 4096 20180 4136
rect 20323 4096 20332 4136
rect 20372 4096 20812 4136
rect 20852 4096 20861 4136
rect 23971 4096 23980 4136
rect 24020 4096 25612 4136
rect 25652 4096 25661 4136
rect 26083 4096 26092 4136
rect 26132 4096 26668 4136
rect 26708 4096 27628 4136
rect 27668 4096 27677 4136
rect 28099 4096 28108 4136
rect 28148 4096 28396 4136
rect 28436 4096 28445 4136
rect 28579 4096 28588 4136
rect 28628 4096 29068 4136
rect 29108 4096 29117 4136
rect 31651 4096 31660 4136
rect 31700 4096 32908 4136
rect 32948 4096 32957 4136
rect 35875 4096 35884 4136
rect 35924 4096 36652 4136
rect 36692 4096 36701 4136
rect 38755 4096 38764 4136
rect 38804 4096 39244 4136
rect 39284 4096 39293 4136
rect 20140 4052 20180 4096
rect 6700 4012 7660 4052
rect 7700 4012 7709 4052
rect 15043 4012 15052 4052
rect 15092 4012 16108 4052
rect 16148 4012 16157 4052
rect 17539 4012 17548 4052
rect 17588 4012 18700 4052
rect 18740 4012 18749 4052
rect 20140 4012 20276 4052
rect 22051 4012 22060 4052
rect 22100 4012 24364 4052
rect 24404 4012 24413 4052
rect 26179 4012 26188 4052
rect 26228 4012 26476 4052
rect 26516 4012 28012 4052
rect 28052 4012 28061 4052
rect 36268 4012 37804 4052
rect 37844 4012 37853 4052
rect 0 3968 80 3988
rect 6700 3968 6740 4012
rect 8899 3968 8957 3969
rect 20236 3968 20276 4012
rect 36268 3968 36308 4012
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 6691 3928 6700 3968
rect 6740 3928 6749 3968
rect 7459 3928 7468 3968
rect 7508 3928 8140 3968
rect 8180 3928 8189 3968
rect 8803 3928 8812 3968
rect 8852 3928 8908 3968
rect 8948 3928 8957 3968
rect 9187 3928 9196 3968
rect 9236 3928 10252 3968
rect 10292 3928 10301 3968
rect 11107 3928 11116 3968
rect 11156 3928 15724 3968
rect 15764 3928 15773 3968
rect 17443 3928 17452 3968
rect 17492 3928 17836 3968
rect 17876 3928 17885 3968
rect 18499 3928 18508 3968
rect 18548 3928 20180 3968
rect 20227 3928 20236 3968
rect 20276 3928 20285 3968
rect 23779 3928 23788 3968
rect 23828 3928 26380 3968
rect 26420 3928 26429 3968
rect 27523 3928 27532 3968
rect 27572 3928 29740 3968
rect 29780 3928 29789 3968
rect 31459 3928 31468 3968
rect 31508 3928 34444 3968
rect 34484 3928 34493 3968
rect 34915 3928 34924 3968
rect 34964 3928 35308 3968
rect 35348 3928 35357 3968
rect 36259 3928 36268 3968
rect 36308 3928 36317 3968
rect 38371 3928 38380 3968
rect 38420 3928 39628 3968
rect 39668 3928 40492 3968
rect 40532 3928 40541 3968
rect 0 3908 80 3928
rect 8899 3927 8957 3928
rect 20140 3884 20180 3928
rect 27619 3884 27677 3885
rect 10627 3844 10636 3884
rect 10676 3844 16300 3884
rect 16340 3844 16349 3884
rect 17731 3844 17740 3884
rect 17780 3844 18892 3884
rect 18932 3844 18941 3884
rect 20140 3844 27436 3884
rect 27476 3844 27485 3884
rect 27619 3844 27628 3884
rect 27668 3844 27762 3884
rect 27820 3844 28052 3884
rect 28579 3844 28588 3884
rect 28628 3844 29068 3884
rect 29108 3844 29356 3884
rect 29396 3844 29644 3884
rect 29684 3844 29693 3884
rect 31267 3844 31276 3884
rect 31316 3844 31660 3884
rect 31700 3844 31709 3884
rect 37891 3844 37900 3884
rect 37940 3844 38284 3884
rect 38324 3844 38333 3884
rect 27619 3843 27677 3844
rect 27820 3800 27860 3844
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 5347 3760 5356 3800
rect 5396 3760 6796 3800
rect 6836 3760 6845 3800
rect 7939 3760 7948 3800
rect 7988 3760 9004 3800
rect 9044 3760 9053 3800
rect 9187 3760 9196 3800
rect 9236 3760 9676 3800
rect 9716 3760 9725 3800
rect 9955 3760 9964 3800
rect 10004 3760 10156 3800
rect 10196 3760 10205 3800
rect 12067 3760 12076 3800
rect 12116 3760 12748 3800
rect 12788 3760 12797 3800
rect 17539 3760 17548 3800
rect 17588 3760 18028 3800
rect 18068 3760 18077 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 20611 3760 20620 3800
rect 20660 3760 21580 3800
rect 21620 3760 21629 3800
rect 23299 3760 23308 3800
rect 23348 3760 26708 3800
rect 26755 3760 26764 3800
rect 26804 3760 27532 3800
rect 27572 3760 27860 3800
rect 27907 3760 27916 3800
rect 27956 3760 27965 3800
rect 26668 3716 26708 3760
rect 27811 3716 27869 3717
rect 17923 3676 17932 3716
rect 17972 3676 18124 3716
rect 18164 3676 18173 3716
rect 19939 3676 19948 3716
rect 19988 3676 20524 3716
rect 20564 3676 23500 3716
rect 23540 3676 24172 3716
rect 24212 3676 24221 3716
rect 26668 3676 27820 3716
rect 27860 3676 27869 3716
rect 27811 3675 27869 3676
rect 26659 3632 26717 3633
rect 7747 3592 7756 3632
rect 7796 3592 8716 3632
rect 8756 3592 8765 3632
rect 10051 3592 10060 3632
rect 10100 3592 11308 3632
rect 11348 3592 11357 3632
rect 14083 3592 14092 3632
rect 14132 3592 14668 3632
rect 14708 3592 14717 3632
rect 15907 3592 15916 3632
rect 15956 3592 16492 3632
rect 16532 3592 19372 3632
rect 19412 3592 19421 3632
rect 19468 3592 21100 3632
rect 21140 3592 21149 3632
rect 23779 3592 23788 3632
rect 23828 3592 24268 3632
rect 24308 3592 24317 3632
rect 25507 3592 25516 3632
rect 25556 3592 26668 3632
rect 26708 3592 26717 3632
rect 19468 3548 19508 3592
rect 26659 3591 26717 3592
rect 8227 3508 8236 3548
rect 8276 3508 10828 3548
rect 10868 3508 10877 3548
rect 17059 3508 17068 3548
rect 17108 3508 17836 3548
rect 17876 3508 17885 3548
rect 18019 3508 18028 3548
rect 18068 3508 19508 3548
rect 19747 3508 19756 3548
rect 19796 3508 20468 3548
rect 20899 3508 20908 3548
rect 20948 3508 21388 3548
rect 21428 3508 21437 3548
rect 24067 3508 24076 3548
rect 24116 3508 25420 3548
rect 25460 3508 25469 3548
rect 26563 3508 26572 3548
rect 26612 3508 27244 3548
rect 27284 3508 27436 3548
rect 27476 3508 27485 3548
rect 20428 3464 20468 3508
rect 22723 3464 22781 3465
rect 27916 3464 27956 3760
rect 28012 3716 28052 3844
rect 28099 3800 28157 3801
rect 28099 3760 28108 3800
rect 28148 3760 29164 3800
rect 29204 3760 29213 3800
rect 31075 3760 31084 3800
rect 31124 3760 31756 3800
rect 31796 3760 31805 3800
rect 31939 3760 31948 3800
rect 31988 3760 31997 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 37603 3760 37612 3800
rect 37652 3760 38092 3800
rect 38132 3760 38141 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 28099 3759 28157 3760
rect 31948 3716 31988 3760
rect 28012 3676 28492 3716
rect 28532 3676 29260 3716
rect 29300 3676 29309 3716
rect 30787 3676 30796 3716
rect 30836 3676 31180 3716
rect 31220 3676 31229 3716
rect 31363 3676 31372 3716
rect 31412 3676 31988 3716
rect 28963 3592 28972 3632
rect 29012 3592 33580 3632
rect 33620 3592 34060 3632
rect 34100 3592 34109 3632
rect 28675 3508 28684 3548
rect 28724 3508 29876 3548
rect 29836 3464 29876 3508
rect 6595 3424 6604 3464
rect 6644 3424 9388 3464
rect 9428 3424 9437 3464
rect 16291 3424 16300 3464
rect 16340 3424 19276 3464
rect 19316 3424 20140 3464
rect 20180 3424 20189 3464
rect 20419 3424 20428 3464
rect 20468 3424 20477 3464
rect 21091 3424 21100 3464
rect 21140 3424 21676 3464
rect 21716 3424 21725 3464
rect 22638 3424 22732 3464
rect 22772 3424 23692 3464
rect 23732 3424 23741 3464
rect 24259 3424 24268 3464
rect 24308 3424 26764 3464
rect 26804 3424 26813 3464
rect 27811 3424 27820 3464
rect 27860 3424 28108 3464
rect 28148 3424 28157 3464
rect 28387 3424 28396 3464
rect 28436 3424 29356 3464
rect 29396 3424 29405 3464
rect 29827 3424 29836 3464
rect 29876 3424 29885 3464
rect 30979 3424 30988 3464
rect 31028 3424 31276 3464
rect 31316 3424 31325 3464
rect 31555 3424 31564 3464
rect 31604 3424 32044 3464
rect 32084 3424 32093 3464
rect 36163 3424 36172 3464
rect 36212 3424 36652 3464
rect 36692 3424 36701 3464
rect 22723 3423 22781 3424
rect 8899 3340 8908 3380
rect 8948 3340 9772 3380
rect 9812 3340 9821 3380
rect 19171 3340 19180 3380
rect 19220 3340 21004 3380
rect 21044 3340 21484 3380
rect 21524 3340 21533 3380
rect 24451 3340 24460 3380
rect 24500 3340 25324 3380
rect 25364 3340 25373 3380
rect 28960 3340 29260 3380
rect 29300 3340 29932 3380
rect 29972 3340 31372 3380
rect 31412 3340 31421 3380
rect 15811 3296 15869 3297
rect 21283 3296 21341 3297
rect 28960 3296 29000 3340
rect 15726 3256 15820 3296
rect 15860 3256 15869 3296
rect 20131 3256 20140 3296
rect 20180 3256 20812 3296
rect 20852 3256 20861 3296
rect 21198 3256 21292 3296
rect 21332 3256 21341 3296
rect 24163 3256 24172 3296
rect 24212 3256 24364 3296
rect 24404 3256 29000 3296
rect 15811 3255 15869 3256
rect 21283 3255 21341 3256
rect 21292 3212 21332 3255
rect 27139 3212 27197 3213
rect 21292 3172 26572 3212
rect 26612 3172 27148 3212
rect 27188 3172 27197 3212
rect 27427 3172 27436 3212
rect 27476 3172 27820 3212
rect 27860 3172 27869 3212
rect 27139 3171 27197 3172
rect 0 3128 80 3148
rect 20323 3128 20381 3129
rect 0 3088 652 3128
rect 692 3088 701 3128
rect 15715 3088 15724 3128
rect 15764 3088 20332 3128
rect 20372 3088 21292 3128
rect 21332 3088 21341 3128
rect 27139 3088 27148 3128
rect 27188 3088 27916 3128
rect 27956 3088 29000 3128
rect 0 3068 80 3088
rect 20323 3087 20381 3088
rect 28960 3044 29000 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 17731 3004 17740 3044
rect 17780 3004 18028 3044
rect 18068 3004 18077 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 20803 3004 20812 3044
rect 20852 3004 25172 3044
rect 27235 3004 27244 3044
rect 27284 3004 28012 3044
rect 28052 3004 28061 3044
rect 28960 3004 29932 3044
rect 29972 3004 30124 3044
rect 30164 3004 30316 3044
rect 30356 3004 30365 3044
rect 31948 3004 32140 3044
rect 32180 3004 32189 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 25132 2960 25172 3004
rect 31948 2960 31988 3004
rect 16300 2920 18356 2960
rect 19363 2920 19372 2960
rect 19412 2920 20908 2960
rect 20948 2920 20957 2960
rect 25123 2920 25132 2960
rect 25172 2920 31988 2960
rect 32035 2920 32044 2960
rect 32084 2920 33332 2960
rect 16300 2876 16340 2920
rect 18316 2876 18356 2920
rect 33292 2876 33332 2920
rect 8227 2836 8236 2876
rect 8276 2836 9196 2876
rect 9236 2836 9245 2876
rect 16291 2836 16300 2876
rect 16340 2836 16349 2876
rect 16771 2836 16780 2876
rect 16820 2836 17932 2876
rect 17972 2836 17981 2876
rect 18307 2836 18316 2876
rect 18356 2836 18365 2876
rect 27619 2836 27628 2876
rect 27668 2836 28300 2876
rect 28340 2836 28349 2876
rect 33283 2836 33292 2876
rect 33332 2836 33341 2876
rect 37411 2836 37420 2876
rect 37460 2836 37996 2876
rect 38036 2836 38045 2876
rect 2500 2752 14284 2792
rect 14324 2752 14333 2792
rect 16579 2752 16588 2792
rect 16628 2752 17452 2792
rect 17492 2752 17836 2792
rect 17876 2752 17885 2792
rect 18019 2752 18028 2792
rect 18068 2752 22636 2792
rect 22676 2752 22685 2792
rect 25411 2752 25420 2792
rect 25460 2752 29740 2792
rect 29780 2752 31468 2792
rect 31508 2752 31517 2792
rect 2500 2708 2540 2752
rect 835 2668 844 2708
rect 884 2668 2540 2708
rect 7459 2668 7468 2708
rect 7508 2668 11404 2708
rect 11444 2668 11453 2708
rect 17251 2668 17260 2708
rect 17300 2668 19468 2708
rect 19508 2668 20620 2708
rect 20660 2668 20669 2708
rect 7171 2584 7180 2624
rect 7220 2584 7564 2624
rect 7604 2584 7613 2624
rect 16099 2584 16108 2624
rect 16148 2584 16876 2624
rect 16916 2584 16925 2624
rect 17155 2584 17164 2624
rect 17204 2584 17644 2624
rect 17684 2584 19660 2624
rect 19700 2584 19709 2624
rect 19843 2584 19852 2624
rect 19892 2584 20140 2624
rect 20180 2584 20189 2624
rect 20419 2584 20428 2624
rect 20468 2584 21196 2624
rect 21236 2584 21245 2624
rect 28099 2584 28108 2624
rect 28148 2584 28972 2624
rect 29012 2584 29021 2624
rect 29068 2584 29356 2624
rect 29396 2584 29405 2624
rect 31171 2584 31180 2624
rect 31220 2584 32276 2624
rect 32803 2584 32812 2624
rect 32852 2584 33100 2624
rect 33140 2584 34540 2624
rect 34580 2584 36460 2624
rect 36500 2584 36509 2624
rect 37987 2584 37996 2624
rect 38036 2584 38476 2624
rect 38516 2584 38525 2624
rect 17059 2540 17117 2541
rect 29068 2540 29108 2584
rect 32236 2540 32276 2584
rect 16387 2500 16396 2540
rect 16436 2500 17068 2540
rect 17108 2500 17117 2540
rect 17347 2500 17356 2540
rect 17396 2500 17780 2540
rect 18115 2500 18124 2540
rect 18164 2500 18316 2540
rect 18356 2500 18365 2540
rect 18595 2500 18604 2540
rect 18644 2500 18653 2540
rect 28867 2500 28876 2540
rect 28916 2500 29108 2540
rect 32227 2500 32236 2540
rect 32276 2500 32285 2540
rect 17059 2499 17117 2500
rect 17356 2456 17396 2500
rect 17740 2456 17780 2500
rect 18604 2456 18644 2500
rect 17155 2416 17164 2456
rect 17204 2416 17396 2456
rect 17539 2416 17548 2456
rect 17588 2416 17684 2456
rect 17740 2416 17932 2456
rect 17972 2416 18412 2456
rect 18452 2416 18461 2456
rect 18604 2416 19372 2456
rect 19412 2416 19421 2456
rect 20227 2416 20236 2456
rect 20276 2416 23020 2456
rect 23060 2416 24076 2456
rect 24116 2416 24125 2456
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 16675 2248 16684 2288
rect 16724 2248 17548 2288
rect 17588 2248 17597 2288
rect 0 2228 80 2248
rect 17644 2204 17684 2416
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 16483 2164 16492 2204
rect 16532 2164 17356 2204
rect 17396 2164 17684 2204
rect 16003 2080 16012 2120
rect 16052 2080 16532 2120
rect 21763 2080 21772 2120
rect 21812 2080 22444 2120
rect 22484 2080 22493 2120
rect 16492 2036 16532 2080
rect 16483 1996 16492 2036
rect 16532 1996 16876 2036
rect 16916 1996 16925 2036
rect 17059 1996 17068 2036
rect 17108 1996 17260 2036
rect 17300 1996 17309 2036
rect 22531 1996 22540 2036
rect 22580 1996 22924 2036
rect 22964 1996 22973 2036
rect 21571 1912 21580 1952
rect 21620 1912 22444 1952
rect 22484 1912 22493 1952
rect 26851 1912 26860 1952
rect 26900 1912 30124 1952
rect 30164 1912 32812 1952
rect 32852 1912 32861 1952
rect 18787 1744 18796 1784
rect 18836 1744 19372 1784
rect 19412 1744 19421 1784
rect 16483 1660 16492 1700
rect 16532 1660 16780 1700
rect 16820 1660 17452 1700
rect 17492 1660 17501 1700
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 25315 1240 25324 1280
rect 25364 1240 26284 1280
rect 26324 1240 26668 1280
rect 26708 1240 26717 1280
rect 17059 1112 17117 1113
rect 17059 1072 17068 1112
rect 17108 1072 17260 1112
rect 17300 1072 17309 1112
rect 19555 1072 19564 1112
rect 19604 1072 20716 1112
rect 20756 1072 20765 1112
rect 26851 1072 26860 1112
rect 26900 1072 27724 1112
rect 27764 1072 27773 1112
rect 17059 1071 17117 1072
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 76 36688 116 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 6796 35008 6836 35048
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 6796 34084 6836 34124
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4876 33244 4916 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 21292 32992 21332 33032
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 13612 32404 13652 32444
rect 4876 32320 4916 32360
rect 31756 31900 31796 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 13996 31564 14036 31604
rect 12844 31312 12884 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 13612 30976 13652 31016
rect 13996 30976 14036 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 12844 30556 12884 30596
rect 13900 30388 13940 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 11404 27448 11444 27488
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 30796 27028 30836 27068
rect 17164 26776 17204 26816
rect 13132 26692 13172 26732
rect 13804 26608 13844 26648
rect 14764 26608 14804 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 30796 26440 30836 26480
rect 31276 26440 31316 26480
rect 31756 26440 31796 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 14764 26272 14804 26312
rect 17644 26188 17684 26228
rect 13900 26104 13940 26144
rect 28492 26104 28532 26144
rect 30604 26104 30644 26144
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 13708 25516 13748 25556
rect 26476 25432 26516 25472
rect 45772 25180 45812 25220
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 11404 24508 11444 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 13132 23668 13172 23708
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 4876 22828 4916 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4780 22660 4820 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4780 21736 4820 21776
rect 5068 21736 5108 21776
rect 21484 21736 21524 21776
rect 23116 21736 23156 21776
rect 6028 21652 6068 21692
rect 5068 21232 5108 21272
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4876 20728 4916 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 21484 20224 21524 20264
rect 23116 20056 23156 20096
rect 26572 20056 26612 20096
rect 6028 19888 6068 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 6412 18880 6452 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 6412 18544 6452 18584
rect 20620 18544 20660 18584
rect 19372 18292 19412 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 5164 18124 5204 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 20332 17872 20372 17912
rect 28876 17788 28916 17828
rect 28876 17620 28916 17660
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 28012 17368 28052 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 19372 17284 19412 17324
rect 18124 16948 18164 16988
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 31660 16528 31700 16568
rect 28876 16276 28916 16316
rect 32140 16276 32180 16316
rect 34156 16276 34196 16316
rect 19948 16192 19988 16232
rect 31948 16024 31988 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4780 15856 4820 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 34348 15520 34388 15560
rect 5164 15352 5204 15392
rect 19084 15436 19124 15476
rect 6412 15352 6452 15392
rect 29740 15352 29780 15392
rect 19372 15268 19412 15308
rect 20140 15184 20180 15224
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 28876 15100 28916 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 20044 15016 20084 15056
rect 32908 14848 32948 14888
rect 23980 14764 24020 14804
rect 12844 14680 12884 14720
rect 22540 14596 22580 14636
rect 5164 14512 5204 14552
rect 23980 14512 24020 14552
rect 40876 14512 40916 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 28876 14344 28916 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 35020 14344 35060 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 4780 14176 4820 14216
rect 19372 14176 19412 14216
rect 21100 14176 21140 14216
rect 20044 14092 20084 14132
rect 22540 13924 22580 13964
rect 25516 14092 25556 14132
rect 31756 14008 31796 14048
rect 32716 14008 32756 14048
rect 30028 13840 30068 13880
rect 30700 13840 30740 13880
rect 30604 13672 30644 13712
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 32908 13588 32948 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 31660 13504 31700 13544
rect 18700 13168 18740 13208
rect 23980 13168 24020 13208
rect 30604 13168 30644 13208
rect 31852 13084 31892 13124
rect 29740 13000 29780 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 27628 12748 27668 12788
rect 18028 12580 18068 12620
rect 20236 12580 20276 12620
rect 23980 12580 24020 12620
rect 18700 12496 18740 12536
rect 21772 12496 21812 12536
rect 29548 12496 29588 12536
rect 11404 12328 11444 12368
rect 19084 12328 19124 12368
rect 23020 12244 23060 12284
rect 26188 12244 26228 12284
rect 18028 12160 18068 12200
rect 31852 12160 31892 12200
rect 34156 12160 34196 12200
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 30700 12076 30740 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 20236 11992 20276 12032
rect 31468 11908 31508 11948
rect 14476 11740 14516 11780
rect 11884 11656 11924 11696
rect 26572 11656 26612 11696
rect 28012 11656 28052 11696
rect 32332 11572 32372 11612
rect 24460 11488 24500 11528
rect 33196 11488 33236 11528
rect 30412 11404 30452 11444
rect 32908 11404 32948 11444
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 20428 11320 20468 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 36172 11320 36212 11360
rect 18604 11152 18644 11192
rect 34252 11152 34292 11192
rect 32908 11068 32948 11108
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 36460 11236 36500 11276
rect 36076 11152 36116 11192
rect 36364 11152 36404 11192
rect 32524 10984 32564 11024
rect 36172 10900 36212 10940
rect 20908 10816 20948 10856
rect 32140 10816 32180 10856
rect 19372 10732 19412 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 18124 10480 18164 10520
rect 20812 10480 20852 10520
rect 32140 10480 32180 10520
rect 31660 10396 31700 10436
rect 17644 10312 17684 10352
rect 20332 10312 20372 10352
rect 21772 10312 21812 10352
rect 43180 10312 43220 10352
rect 36556 10228 36596 10268
rect 24844 10144 24884 10184
rect 32908 10144 32948 10184
rect 35692 10144 35732 10184
rect 36460 10144 36500 10184
rect 17740 10060 17780 10100
rect 24076 9976 24116 10016
rect 24268 9976 24308 10016
rect 32044 9892 32084 9932
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 31660 9808 31700 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 36364 9808 36404 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 31852 9724 31892 9764
rect 32044 9556 32084 9596
rect 21388 9472 21428 9512
rect 24940 9472 24980 9512
rect 27148 9472 27188 9512
rect 21580 9388 21620 9428
rect 20812 9304 20852 9344
rect 32044 9304 32084 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 36076 9136 36116 9176
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 26668 9052 26708 9092
rect 32236 9052 32276 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 32332 8968 32372 9008
rect 24364 8884 24404 8924
rect 30316 8884 30356 8924
rect 34252 8968 34292 9008
rect 21484 8800 21524 8840
rect 27724 8800 27764 8840
rect 28012 8800 28052 8840
rect 30700 8800 30740 8840
rect 31468 8800 31508 8840
rect 34060 8800 34100 8840
rect 24652 8716 24692 8756
rect 24940 8716 24980 8756
rect 23212 8632 23252 8672
rect 34156 8632 34196 8672
rect 20812 8548 20852 8588
rect 19852 8464 19892 8504
rect 20908 8464 20948 8504
rect 21484 8464 21524 8504
rect 28972 8464 29012 8504
rect 33196 8464 33236 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 20524 8296 20564 8336
rect 22540 8380 22580 8420
rect 22732 8380 22772 8420
rect 30316 8380 30356 8420
rect 34252 8380 34292 8420
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 26668 8212 26708 8252
rect 9484 8128 9524 8168
rect 23212 8128 23252 8168
rect 27532 8128 27572 8168
rect 20524 8044 20564 8084
rect 29836 7960 29876 8000
rect 20812 7876 20852 7916
rect 9004 7624 9044 7664
rect 26764 7624 26804 7664
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 32140 7540 32180 7580
rect 32524 7540 32564 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 23980 7456 24020 7496
rect 27628 7456 27668 7496
rect 35692 7456 35732 7496
rect 30604 7288 30644 7328
rect 19084 7120 19124 7160
rect 23788 7120 23828 7160
rect 23980 7120 24020 7160
rect 27148 7120 27188 7160
rect 30412 7120 30452 7160
rect 34156 7120 34196 7160
rect 18796 7036 18836 7076
rect 34252 7036 34292 7076
rect 43180 7036 43220 7076
rect 23692 6868 23732 6908
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 24652 6784 24692 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 30604 6700 30644 6740
rect 24268 6616 24308 6656
rect 18892 6532 18932 6572
rect 24460 6532 24500 6572
rect 27724 6532 27764 6572
rect 32044 6532 32084 6572
rect 32236 6532 32276 6572
rect 34156 6532 34196 6572
rect 9484 6448 9524 6488
rect 27628 6448 27668 6488
rect 35692 6448 35732 6488
rect 44716 6448 44756 6488
rect 22636 6364 22676 6404
rect 23404 6364 23444 6404
rect 42220 6364 42260 6404
rect 43180 6364 43220 6404
rect 24268 6280 24308 6320
rect 32524 6196 32564 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 18988 6028 19028 6068
rect 32236 6028 32276 6068
rect 32908 6028 32948 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 19372 5944 19412 5984
rect 26572 5944 26612 5984
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 7756 5776 7796 5816
rect 26572 5608 26612 5648
rect 8908 5524 8948 5564
rect 28972 5524 29012 5564
rect 32140 5524 32180 5564
rect 30700 5356 30740 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 17260 5020 17300 5060
rect 21772 5020 21812 5060
rect 23020 5020 23060 5060
rect 24460 5020 24500 5060
rect 24652 5020 24692 5060
rect 28012 5020 28052 5060
rect 7756 4936 7796 4976
rect 21580 4936 21620 4976
rect 31948 4936 31988 4976
rect 34348 4936 34388 4976
rect 18892 4852 18932 4892
rect 30316 4852 30356 4892
rect 30892 4768 30932 4808
rect 25036 4684 25076 4724
rect 9004 4600 9044 4640
rect 27628 4684 27668 4724
rect 28972 4684 29012 4724
rect 32908 4684 32948 4724
rect 17740 4600 17780 4640
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 26380 4516 26420 4556
rect 31852 4516 31892 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 29548 4432 29588 4472
rect 15820 4348 15860 4388
rect 19084 4264 19124 4304
rect 20332 4264 20372 4304
rect 25324 4264 25364 4304
rect 26476 4264 26516 4304
rect 8908 3928 8948 3968
rect 27628 3844 27668 3884
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 27820 3676 27860 3716
rect 26668 3592 26708 3632
rect 28108 3760 28148 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 22732 3424 22772 3464
rect 15820 3256 15860 3296
rect 21292 3256 21332 3296
rect 27148 3172 27188 3212
rect 20332 3088 20372 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 17068 2500 17108 2540
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 17068 1072 17108 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 76 36728 116 36737
rect 76 20105 116 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 6796 35048 6836 35057
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 6796 34124 6836 35008
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 6796 34075 6836 34084
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4876 33284 4916 33293
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4876 32360 4916 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 21292 33032 21332 33041
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 4876 32311 4916 32320
rect 13612 32444 13652 32453
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 12844 31352 12884 31361
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 12844 30596 12884 31312
rect 13612 31016 13652 32404
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 13612 30967 13652 30976
rect 13996 31604 14036 31613
rect 13996 31016 14036 31564
rect 13996 30967 14036 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 12844 30547 12884 30556
rect 13900 30428 13940 30437
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 11404 27488 11444 27497
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 11404 24548 11444 27448
rect 11404 24499 11444 24508
rect 13132 26732 13172 26741
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 13132 23708 13172 26692
rect 13804 26648 13844 26657
rect 13804 26153 13844 26608
rect 13803 26144 13845 26153
rect 13803 26104 13804 26144
rect 13844 26104 13845 26144
rect 13803 26095 13845 26104
rect 13900 26144 13940 30388
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 21292 26825 21332 32992
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 31756 31940 31796 31949
rect 30796 27068 30836 27077
rect 17163 26816 17205 26825
rect 17163 26776 17164 26816
rect 17204 26776 17205 26816
rect 17163 26767 17205 26776
rect 21291 26816 21333 26825
rect 21291 26776 21292 26816
rect 21332 26776 21333 26816
rect 21291 26767 21333 26776
rect 17164 26682 17204 26767
rect 14764 26648 14804 26657
rect 14764 26312 14804 26608
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 30796 26480 30836 27028
rect 30796 26431 30836 26440
rect 31276 26480 31316 26489
rect 14764 26263 14804 26272
rect 13900 26095 13940 26104
rect 17644 26228 17684 26237
rect 17644 25901 17684 26188
rect 28492 26144 28532 26153
rect 28492 25901 28532 26104
rect 30603 26144 30645 26153
rect 30603 26104 30604 26144
rect 30644 26104 30645 26144
rect 30603 26095 30645 26104
rect 30604 26010 30644 26095
rect 17643 25892 17685 25901
rect 17643 25852 17644 25892
rect 17684 25852 17685 25892
rect 17643 25843 17685 25852
rect 28491 25892 28533 25901
rect 28491 25852 28492 25892
rect 28532 25852 28533 25892
rect 28491 25843 28533 25852
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 13708 25556 13748 25565
rect 13708 25229 13748 25516
rect 26476 25472 26516 25481
rect 26476 25229 26516 25432
rect 31276 25229 31316 26440
rect 31756 26480 31796 31900
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 31756 26431 31796 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 13707 25220 13749 25229
rect 13707 25180 13708 25220
rect 13748 25180 13749 25220
rect 13707 25171 13749 25180
rect 26475 25220 26517 25229
rect 26475 25180 26476 25220
rect 26516 25180 26517 25220
rect 26475 25171 26517 25180
rect 31275 25220 31317 25229
rect 31275 25180 31276 25220
rect 31316 25180 31317 25220
rect 31275 25171 31317 25180
rect 45771 25220 45813 25229
rect 45771 25180 45772 25220
rect 45812 25180 45813 25220
rect 45771 25171 45813 25180
rect 45772 25086 45812 25171
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 13132 23659 13172 23668
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 4876 22868 4916 22877
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4780 22700 4820 22709
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4780 21776 4820 22660
rect 4780 21727 4820 21736
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4876 20768 4916 22828
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 5068 21776 5108 21785
rect 5068 21272 5108 21736
rect 21484 21776 21524 21785
rect 5068 21223 5108 21232
rect 6028 21692 6068 21701
rect 4876 20719 4916 20728
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 75 20096 117 20105
rect 75 20056 76 20096
rect 116 20056 117 20096
rect 75 20047 117 20056
rect 6028 19928 6068 21652
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 21484 20264 21524 21736
rect 21484 20215 21524 20224
rect 23116 21776 23156 21785
rect 23116 20096 23156 21736
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 23116 20047 23156 20056
rect 26571 20096 26613 20105
rect 26571 20056 26572 20096
rect 26612 20056 26613 20096
rect 26571 20047 26613 20056
rect 26572 19962 26612 20047
rect 6028 19879 6068 19888
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 6412 18920 6452 18929
rect 6412 18584 6452 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 5164 18164 5204 18173
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4780 15896 4820 15905
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4780 14216 4820 15856
rect 5164 15392 5204 18124
rect 5164 14552 5204 15352
rect 6412 15392 6452 18544
rect 20620 18584 20660 18593
rect 19372 18332 19412 18341
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 19372 17324 19412 18292
rect 20332 17912 20372 17921
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 19372 17275 19412 17284
rect 6412 15343 6452 15352
rect 18124 16988 18164 16997
rect 12843 14720 12885 14729
rect 12843 14680 12844 14720
rect 12884 14680 12885 14720
rect 12843 14671 12885 14680
rect 12844 14586 12884 14671
rect 5164 14503 5204 14512
rect 4780 14167 4820 14176
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 18028 12620 18068 12629
rect 11403 12368 11445 12377
rect 11403 12328 11404 12368
rect 11444 12328 11445 12368
rect 11403 12319 11445 12328
rect 11404 12234 11444 12319
rect 18028 12200 18068 12580
rect 18028 12151 18068 12160
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 14475 11780 14517 11789
rect 14475 11740 14476 11780
rect 14516 11740 14517 11780
rect 14475 11731 14517 11740
rect 11883 11696 11925 11705
rect 11883 11656 11884 11696
rect 11924 11656 11925 11696
rect 11883 11647 11925 11656
rect 11884 11562 11924 11647
rect 14476 11646 14516 11731
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18124 10520 18164 16948
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 19948 16232 19988 16241
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 19084 15476 19124 15485
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18700 13208 18740 13217
rect 18700 12545 18740 13168
rect 18699 12536 18741 12545
rect 18699 12496 18700 12536
rect 18740 12496 18741 12536
rect 18699 12487 18741 12496
rect 18700 12401 18740 12487
rect 19084 12368 19124 15436
rect 19372 15308 19412 15317
rect 19372 14216 19412 15268
rect 19948 14561 19988 16192
rect 20139 15224 20181 15233
rect 20139 15184 20140 15224
rect 20180 15184 20181 15224
rect 20139 15175 20181 15184
rect 20140 15090 20180 15175
rect 20044 15056 20084 15065
rect 19947 14552 19989 14561
rect 19947 14512 19948 14552
rect 19988 14512 19989 14552
rect 19947 14503 19989 14512
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19372 14167 19412 14176
rect 20044 14132 20084 15016
rect 20044 14083 20084 14092
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 19084 12319 19124 12328
rect 20236 12620 20276 12629
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 20236 12032 20276 12580
rect 20236 11983 20276 11992
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 18603 11192 18645 11201
rect 18603 11152 18604 11192
rect 18644 11152 18645 11192
rect 18603 11143 18645 11152
rect 18604 11058 18644 11143
rect 19372 10772 19412 10781
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 18124 10471 18164 10480
rect 17644 10352 17684 10361
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 9484 8168 9524 8177
rect 9004 7664 9044 7673
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 7756 5816 7796 5825
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 7756 4976 7796 5776
rect 7756 4927 7796 4936
rect 8908 5564 8948 5573
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 8908 3968 8948 5524
rect 9004 4640 9044 7624
rect 9484 6488 9524 8128
rect 9484 6439 9524 6448
rect 17260 5060 17300 5071
rect 17260 4985 17300 5020
rect 17259 4976 17301 4985
rect 17259 4936 17260 4976
rect 17300 4936 17301 4976
rect 17259 4927 17301 4936
rect 9004 4591 9044 4600
rect 8908 3919 8948 3928
rect 15820 4388 15860 4397
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 15820 3305 15860 4348
rect 17644 3305 17684 10312
rect 17740 10100 17780 10109
rect 17740 4640 17780 10060
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 19084 7160 19124 7169
rect 18796 7076 18836 7085
rect 18836 7036 19028 7076
rect 18796 7027 18836 7036
rect 18892 6572 18932 6581
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18892 4892 18932 6532
rect 18988 6068 19028 7036
rect 18988 6019 19028 6028
rect 18892 4843 18932 4852
rect 17740 4591 17780 4600
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 19084 4304 19124 7120
rect 19372 5984 19412 10732
rect 20332 10352 20372 17872
rect 20332 10303 20372 10312
rect 20428 11360 20468 11369
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 19852 8513 19892 8598
rect 19851 8504 19893 8513
rect 19851 8464 19852 8504
rect 19892 8464 19893 8504
rect 19851 8455 19893 8464
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 19372 5935 19412 5944
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 20428 5069 20468 11320
rect 20620 11201 20660 18544
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 28876 17828 28916 17837
rect 28876 17660 28916 17788
rect 28012 17408 28052 17417
rect 22539 15224 22581 15233
rect 22539 15184 22540 15224
rect 22580 15184 22581 15224
rect 22539 15175 22581 15184
rect 22540 14636 22580 15175
rect 21100 14216 21140 14225
rect 21100 13889 21140 14176
rect 22540 13964 22580 14596
rect 23980 14804 24020 14813
rect 23980 14552 24020 14764
rect 23980 14503 24020 14512
rect 22540 13915 22580 13924
rect 25516 14132 25556 14141
rect 21099 13880 21141 13889
rect 21099 13840 21100 13880
rect 21140 13840 21141 13880
rect 21099 13831 21141 13840
rect 23980 13208 24020 13217
rect 23980 12620 24020 13168
rect 21771 12536 21813 12545
rect 21771 12496 21772 12536
rect 21812 12496 21813 12536
rect 21771 12487 21813 12496
rect 21772 12402 21812 12487
rect 23020 12284 23060 12293
rect 20619 11192 20661 11201
rect 20619 11152 20620 11192
rect 20660 11152 20661 11192
rect 20619 11143 20661 11152
rect 20908 10856 20948 10865
rect 20812 10520 20852 10529
rect 20812 9344 20852 10480
rect 20812 9295 20852 9304
rect 20812 8588 20852 8597
rect 20524 8336 20564 8345
rect 20524 8084 20564 8296
rect 20812 8261 20852 8548
rect 20908 8504 20948 10816
rect 21772 10352 21812 10361
rect 21388 9512 21428 9521
rect 21388 8849 21428 9472
rect 21580 9428 21620 9437
rect 21387 8840 21429 8849
rect 21387 8800 21388 8840
rect 21428 8800 21429 8840
rect 21387 8791 21429 8800
rect 21484 8840 21524 8849
rect 20908 8455 20948 8464
rect 21484 8504 21524 8800
rect 21484 8455 21524 8464
rect 20811 8252 20853 8261
rect 20811 8212 20812 8252
rect 20852 8212 20853 8252
rect 20811 8203 20853 8212
rect 20524 8035 20564 8044
rect 20812 7916 20852 8203
rect 20812 7867 20852 7876
rect 20427 5060 20469 5069
rect 20427 5020 20428 5060
rect 20468 5020 20469 5060
rect 20427 5011 20469 5020
rect 21580 4976 21620 9388
rect 21772 5060 21812 10312
rect 22635 8504 22677 8513
rect 22635 8464 22636 8504
rect 22676 8464 22677 8504
rect 22635 8455 22677 8464
rect 22539 8420 22581 8429
rect 22539 8380 22540 8420
rect 22580 8380 22581 8420
rect 22539 8371 22581 8380
rect 22540 8286 22580 8371
rect 22636 6404 22676 8455
rect 22636 6355 22676 6364
rect 22732 8420 22772 8429
rect 21772 4985 21812 5020
rect 21580 4901 21620 4936
rect 21771 4976 21813 4985
rect 21771 4936 21772 4976
rect 21812 4936 21813 4976
rect 21771 4927 21813 4936
rect 21579 4892 21621 4901
rect 21579 4852 21580 4892
rect 21620 4852 21621 4892
rect 21579 4843 21621 4852
rect 21772 4313 21812 4927
rect 19084 4255 19124 4264
rect 20332 4304 20372 4313
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 15819 3296 15861 3305
rect 15819 3256 15820 3296
rect 15860 3256 15861 3296
rect 15819 3247 15861 3256
rect 17643 3296 17685 3305
rect 17643 3256 17644 3296
rect 17684 3256 17685 3296
rect 17643 3247 17685 3256
rect 15820 3162 15860 3247
rect 20332 3128 20372 4264
rect 21771 4304 21813 4313
rect 21771 4264 21772 4304
rect 21812 4264 21813 4304
rect 21771 4255 21813 4264
rect 22732 3464 22772 8380
rect 23020 5060 23060 12244
rect 23212 8672 23252 8681
rect 23212 8177 23252 8632
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 23691 8168 23733 8177
rect 23691 8128 23692 8168
rect 23732 8128 23733 8168
rect 23691 8119 23733 8128
rect 23212 8034 23252 8119
rect 23692 6908 23732 8119
rect 23980 7496 24020 12580
rect 25516 11789 25556 14092
rect 27628 12788 27668 12797
rect 26187 12284 26229 12293
rect 26187 12244 26188 12284
rect 26228 12244 26229 12284
rect 26187 12235 26229 12244
rect 26188 12150 26228 12235
rect 25515 11780 25557 11789
rect 25515 11740 25516 11780
rect 25556 11740 25557 11780
rect 25515 11731 25557 11740
rect 26572 11696 26612 11705
rect 24460 11528 24500 11537
rect 24075 10016 24117 10025
rect 24075 9976 24076 10016
rect 24116 9976 24117 10016
rect 24075 9967 24117 9976
rect 24268 10016 24308 10025
rect 24076 9882 24116 9967
rect 23787 7160 23829 7169
rect 23787 7120 23788 7160
rect 23828 7120 23829 7160
rect 23787 7111 23829 7120
rect 23980 7160 24020 7456
rect 23980 7111 24020 7120
rect 23788 7026 23828 7111
rect 23692 6859 23732 6868
rect 24268 6656 24308 9976
rect 24364 8924 24404 8933
rect 24364 8177 24404 8884
rect 24363 8168 24405 8177
rect 24363 8128 24364 8168
rect 24404 8128 24405 8168
rect 24363 8119 24405 8128
rect 23403 6404 23445 6413
rect 23403 6364 23404 6404
rect 23444 6364 23445 6404
rect 23403 6355 23445 6364
rect 23404 6270 23444 6355
rect 24268 6320 24308 6616
rect 24460 6572 24500 11488
rect 24844 10184 24884 10195
rect 24844 10109 24884 10144
rect 24843 10100 24885 10109
rect 24843 10060 24844 10100
rect 24884 10060 24885 10100
rect 24843 10051 24885 10060
rect 24939 10016 24981 10025
rect 24939 9976 24940 10016
rect 24980 9976 24981 10016
rect 24939 9967 24981 9976
rect 24940 9512 24980 9967
rect 24652 8756 24692 8765
rect 24652 6824 24692 8716
rect 24940 8756 24980 9472
rect 24940 8429 24980 8716
rect 24939 8420 24981 8429
rect 24939 8380 24940 8420
rect 24980 8380 24981 8420
rect 24939 8371 24981 8380
rect 24652 6775 24692 6784
rect 24460 6523 24500 6532
rect 24268 6271 24308 6280
rect 26572 5984 26612 11656
rect 27148 9512 27188 9521
rect 26572 5648 26612 5944
rect 26572 5599 26612 5608
rect 26668 9092 26708 9101
rect 26668 8252 26708 9052
rect 23020 5011 23060 5020
rect 24459 5060 24501 5069
rect 24459 5020 24460 5060
rect 24500 5020 24501 5060
rect 24459 5011 24501 5020
rect 24652 5060 24692 5069
rect 24460 4817 24500 5011
rect 24459 4808 24501 4817
rect 24459 4768 24460 4808
rect 24500 4768 24501 4808
rect 24459 4759 24501 4768
rect 24652 4733 24692 5020
rect 24651 4724 24693 4733
rect 24651 4684 24652 4724
rect 24692 4684 24693 4724
rect 24651 4675 24693 4684
rect 25036 4724 25076 4733
rect 25036 4565 25076 4684
rect 25035 4556 25077 4565
rect 25035 4516 25036 4556
rect 25076 4516 25077 4556
rect 25035 4507 25077 4516
rect 26380 4556 26420 4565
rect 26420 4516 26516 4556
rect 26380 4507 26420 4516
rect 25323 4304 25365 4313
rect 25323 4264 25324 4304
rect 25364 4264 25365 4304
rect 25323 4255 25365 4264
rect 26476 4304 26516 4516
rect 26476 4255 26516 4264
rect 25324 4170 25364 4255
rect 26668 3632 26708 8212
rect 26763 8252 26805 8261
rect 26763 8212 26764 8252
rect 26804 8212 26805 8252
rect 26763 8203 26805 8212
rect 26764 7664 26804 8203
rect 26764 7615 26804 7624
rect 26668 3583 26708 3592
rect 27148 7160 27188 9472
rect 27531 8252 27573 8261
rect 27531 8212 27532 8252
rect 27572 8212 27573 8252
rect 27531 8203 27573 8212
rect 27532 8168 27572 8203
rect 27532 8117 27572 8128
rect 22732 3415 22772 3424
rect 21291 3296 21333 3305
rect 21291 3256 21292 3296
rect 21332 3256 21333 3296
rect 21291 3247 21333 3256
rect 21292 3162 21332 3247
rect 27148 3212 27188 7120
rect 27628 7496 27668 12748
rect 28012 11696 28052 17368
rect 28876 16316 28916 17620
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 28876 16267 28916 16276
rect 31660 16568 31700 16577
rect 29740 15392 29780 15401
rect 28876 15140 28916 15149
rect 28876 14384 28916 15100
rect 28876 14335 28916 14344
rect 29740 13040 29780 15352
rect 30027 13880 30069 13889
rect 30027 13840 30028 13880
rect 30068 13840 30069 13880
rect 30027 13831 30069 13840
rect 30700 13880 30740 13889
rect 30028 13746 30068 13831
rect 30604 13712 30644 13721
rect 30604 13208 30644 13672
rect 30604 13159 30644 13168
rect 29740 12991 29780 13000
rect 28012 11647 28052 11656
rect 29548 12536 29588 12545
rect 27724 8840 27764 8849
rect 27724 8765 27764 8800
rect 28012 8840 28052 8849
rect 27723 8756 27765 8765
rect 27723 8716 27724 8756
rect 27764 8716 27765 8756
rect 27723 8707 27765 8716
rect 27724 8705 27764 8707
rect 27628 6488 27668 7456
rect 27723 6572 27765 6581
rect 27723 6532 27724 6572
rect 27764 6532 27765 6572
rect 27723 6523 27765 6532
rect 27628 6439 27668 6448
rect 27724 6438 27764 6523
rect 28012 5060 28052 8800
rect 28971 8756 29013 8765
rect 28971 8716 28972 8756
rect 29012 8716 29013 8756
rect 28971 8707 29013 8716
rect 28972 8504 29012 8707
rect 28972 6581 29012 8464
rect 28971 6572 29013 6581
rect 28971 6532 28972 6572
rect 29012 6532 29013 6572
rect 28971 6523 29013 6532
rect 28012 5011 28052 5020
rect 28972 5564 29012 5573
rect 27628 4724 27668 4733
rect 27628 3884 27668 4684
rect 28972 4724 29012 5524
rect 28972 4675 29012 4684
rect 29548 4472 29588 12496
rect 30700 12116 30740 13840
rect 31660 13544 31700 16528
rect 32140 16316 32180 16325
rect 31948 16064 31988 16073
rect 31660 13495 31700 13504
rect 31756 14048 31796 14057
rect 31756 13376 31796 14008
rect 30700 12067 30740 12076
rect 31660 13336 31796 13376
rect 31468 11948 31508 11957
rect 30412 11444 30452 11453
rect 30316 8924 30356 8933
rect 30316 8420 30356 8884
rect 30316 8371 30356 8380
rect 29836 8000 29876 8009
rect 29836 7169 29876 7960
rect 29835 7160 29877 7169
rect 29835 7120 29836 7160
rect 29876 7120 29877 7160
rect 29835 7111 29877 7120
rect 30412 7160 30452 11404
rect 30700 8840 30740 8849
rect 30412 7111 30452 7120
rect 30604 7328 30644 7337
rect 30604 6740 30644 7288
rect 30604 6691 30644 6700
rect 30700 5396 30740 8800
rect 31468 8840 31508 11908
rect 31660 10436 31700 13336
rect 31660 9848 31700 10396
rect 31660 9799 31700 9808
rect 31852 13124 31892 13133
rect 31852 12200 31892 13084
rect 31852 9764 31892 12160
rect 31852 9715 31892 9724
rect 31468 8791 31508 8800
rect 30700 5347 30740 5356
rect 31948 4976 31988 16024
rect 32140 11705 32180 16276
rect 34156 16316 34196 16325
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 32908 14888 32948 14897
rect 32715 14636 32757 14645
rect 32715 14596 32716 14636
rect 32756 14596 32757 14636
rect 32715 14587 32757 14596
rect 32716 14048 32756 14587
rect 32716 13999 32756 14008
rect 32908 13628 32948 14848
rect 32908 13579 32948 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 34156 12200 34196 16276
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 34156 12151 34196 12160
rect 34348 15560 34388 15569
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 32139 11696 32181 11705
rect 32139 11656 32140 11696
rect 32180 11656 32181 11696
rect 32139 11647 32181 11656
rect 32332 11612 32372 11621
rect 32140 10856 32180 10865
rect 32140 10520 32180 10816
rect 32140 10471 32180 10480
rect 32044 9932 32084 9941
rect 32044 9596 32084 9892
rect 32044 9344 32084 9556
rect 32044 9295 32084 9304
rect 32236 9092 32276 9101
rect 32140 7580 32180 7589
rect 32043 6572 32085 6581
rect 32043 6532 32044 6572
rect 32084 6532 32085 6572
rect 32043 6523 32085 6532
rect 32044 6438 32084 6523
rect 32140 5564 32180 7540
rect 32236 6572 32276 9052
rect 32332 9008 32372 11572
rect 33196 11528 33236 11537
rect 32908 11444 32948 11453
rect 32908 11108 32948 11404
rect 32908 11059 32948 11068
rect 32523 11024 32565 11033
rect 32523 10984 32524 11024
rect 32564 10984 32565 11024
rect 32523 10975 32565 10984
rect 32524 10890 32564 10975
rect 32907 10184 32949 10193
rect 32907 10144 32908 10184
rect 32948 10144 32949 10184
rect 32907 10135 32949 10144
rect 32908 10050 32948 10135
rect 32332 8959 32372 8968
rect 33196 8504 33236 11488
rect 34252 11192 34292 11201
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 34252 9008 34292 11152
rect 34059 8840 34101 8849
rect 34059 8800 34060 8840
rect 34100 8800 34101 8840
rect 34059 8791 34101 8800
rect 34060 8706 34100 8791
rect 33196 8455 33236 8464
rect 34156 8672 34196 8681
rect 32236 6068 32276 6532
rect 32524 7580 32564 7589
rect 32524 6236 32564 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 34156 7160 34196 8632
rect 34156 6572 34196 7120
rect 34252 8420 34292 8968
rect 34252 7076 34292 8380
rect 34252 7027 34292 7036
rect 34156 6523 34196 6532
rect 32907 6320 32949 6329
rect 32907 6280 32908 6320
rect 32948 6280 32949 6320
rect 32907 6271 32949 6280
rect 32524 6187 32564 6196
rect 32236 6019 32276 6028
rect 32908 6068 32948 6271
rect 32908 6019 32948 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 32140 5515 32180 5524
rect 31948 4927 31988 4936
rect 34348 4976 34388 15520
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 35019 14636 35061 14645
rect 35019 14596 35020 14636
rect 35060 14596 35061 14636
rect 35019 14587 35061 14596
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 35020 14384 35060 14587
rect 40875 14552 40917 14561
rect 40875 14512 40876 14552
rect 40916 14512 40917 14552
rect 40875 14503 40917 14512
rect 40876 14418 40916 14503
rect 35020 14335 35060 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 36172 11360 36212 11369
rect 36076 11192 36116 11201
rect 35692 10184 35732 10193
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 35692 7496 35732 10144
rect 36076 9176 36116 11152
rect 36172 11033 36212 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 36460 11276 36500 11285
rect 36364 11192 36404 11201
rect 36171 11024 36213 11033
rect 36171 10984 36172 11024
rect 36212 10984 36213 11024
rect 36171 10975 36213 10984
rect 36172 10940 36212 10975
rect 36172 10860 36212 10900
rect 36364 9848 36404 11152
rect 36460 10184 36500 11236
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 43180 10352 43220 10361
rect 36556 10268 36596 10279
rect 36556 10193 36596 10228
rect 36460 10135 36500 10144
rect 36555 10184 36597 10193
rect 36555 10144 36556 10184
rect 36596 10144 36597 10184
rect 36555 10135 36597 10144
rect 43180 10109 43220 10312
rect 43179 10100 43221 10109
rect 43179 10060 43180 10100
rect 43220 10060 43221 10100
rect 43179 10051 43221 10060
rect 36364 9799 36404 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 36076 9127 36116 9136
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 35692 6488 35732 7456
rect 35692 6439 35732 6448
rect 43180 7076 43220 7085
rect 43180 6413 43220 7036
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 44715 6572 44757 6581
rect 44715 6532 44716 6572
rect 44756 6532 44757 6572
rect 44715 6523 44757 6532
rect 44716 6488 44756 6523
rect 44716 6437 44756 6448
rect 42220 6404 42260 6413
rect 42220 6245 42260 6364
rect 43179 6404 43221 6413
rect 43179 6364 43180 6404
rect 43220 6364 43221 6404
rect 43179 6355 43221 6364
rect 42219 6236 42261 6245
rect 42219 6196 42220 6236
rect 42260 6196 42261 6236
rect 42219 6187 42261 6196
rect 42220 6185 42260 6187
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 34348 4927 34388 4936
rect 30315 4892 30357 4901
rect 30315 4852 30316 4892
rect 30356 4852 30357 4892
rect 30315 4843 30357 4852
rect 30316 4758 30356 4843
rect 30891 4808 30933 4817
rect 30891 4768 30892 4808
rect 30932 4768 30933 4808
rect 30891 4759 30933 4768
rect 30892 4674 30932 4759
rect 32907 4724 32949 4733
rect 32907 4684 32908 4724
rect 32948 4684 32949 4724
rect 32907 4675 32949 4684
rect 32908 4590 32948 4675
rect 31851 4556 31893 4565
rect 31851 4516 31852 4556
rect 31892 4516 31893 4556
rect 31851 4507 31893 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 29548 4423 29588 4432
rect 31852 4422 31892 4507
rect 27628 3835 27668 3844
rect 28108 3800 28148 3809
rect 27820 3760 28108 3800
rect 27820 3716 27860 3760
rect 28108 3751 28148 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 27820 3667 27860 3676
rect 27148 3163 27188 3172
rect 20332 3079 20372 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 17068 2540 17108 2549
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 17068 1112 17108 2500
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 17068 1063 17108 1072
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 13804 26104 13844 26144
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 17164 26776 17204 26816
rect 21292 26776 21332 26816
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 30604 26104 30644 26144
rect 17644 25852 17684 25892
rect 28492 25852 28532 25892
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 13708 25180 13748 25220
rect 26476 25180 26516 25220
rect 31276 25180 31316 25220
rect 45772 25180 45812 25220
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 76 20056 116 20096
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 26572 20056 26612 20096
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 12844 14680 12884 14720
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 11404 12328 11444 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 14476 11740 14516 11780
rect 11884 11656 11924 11696
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18700 12496 18740 12536
rect 20140 15184 20180 15224
rect 19948 14512 19988 14552
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 18604 11152 18644 11192
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 17260 4936 17300 4976
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 19852 8464 19892 8504
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 22540 15184 22580 15224
rect 21100 13840 21140 13880
rect 21772 12496 21812 12536
rect 20620 11152 20660 11192
rect 21388 8800 21428 8840
rect 20812 8212 20852 8252
rect 20428 5020 20468 5060
rect 22636 8464 22676 8504
rect 22540 8380 22580 8420
rect 21772 4936 21812 4976
rect 21580 4852 21620 4892
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 15820 3256 15860 3296
rect 17644 3256 17684 3296
rect 21772 4264 21812 4304
rect 23212 8128 23252 8168
rect 23692 8128 23732 8168
rect 26188 12244 26228 12284
rect 25516 11740 25556 11780
rect 24076 9976 24116 10016
rect 23788 7120 23828 7160
rect 24364 8128 24404 8168
rect 23404 6364 23444 6404
rect 24844 10060 24884 10100
rect 24940 9976 24980 10016
rect 24940 8380 24980 8420
rect 24460 5020 24500 5060
rect 24460 4768 24500 4808
rect 24652 4684 24692 4724
rect 25036 4516 25076 4556
rect 25324 4264 25364 4304
rect 26764 8212 26804 8252
rect 27532 8212 27572 8252
rect 21292 3256 21332 3296
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 30028 13840 30068 13880
rect 27724 8716 27764 8756
rect 27724 6532 27764 6572
rect 28972 8716 29012 8756
rect 28972 6532 29012 6572
rect 29836 7120 29876 7160
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 32716 14596 32756 14636
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 32140 11656 32180 11696
rect 32044 6532 32084 6572
rect 32524 10984 32564 11024
rect 32908 10144 32948 10184
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 34060 8800 34100 8840
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 32908 6280 32948 6320
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 35020 14596 35060 14636
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 40876 14512 40916 14552
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 36172 10984 36212 11024
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 36556 10144 36596 10184
rect 43180 10060 43220 10100
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 44716 6532 44756 6572
rect 43180 6364 43220 6404
rect 42220 6196 42260 6236
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 30316 4852 30356 4892
rect 30892 4768 30932 4808
rect 32908 4684 32948 4724
rect 31852 4516 31892 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 17155 26776 17164 26816
rect 17204 26776 21292 26816
rect 21332 26776 21341 26816
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 13795 26104 13804 26144
rect 13844 26104 30604 26144
rect 30644 26104 30653 26144
rect 17635 25852 17644 25892
rect 17684 25852 28492 25892
rect 28532 25852 28541 25892
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 13699 25180 13708 25220
rect 13748 25180 26476 25220
rect 26516 25180 26525 25220
rect 31267 25180 31276 25220
rect 31316 25180 45772 25220
rect 45812 25180 45821 25220
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 67 20056 76 20096
rect 116 20056 26572 20096
rect 26612 20056 26621 20096
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 20131 15184 20140 15224
rect 20180 15184 22540 15224
rect 22580 15184 22589 15224
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 12835 14680 12844 14720
rect 12884 14680 20180 14720
rect 20140 14636 20180 14680
rect 20140 14596 32716 14636
rect 32756 14596 35020 14636
rect 35060 14596 35069 14636
rect 19939 14512 19948 14552
rect 19988 14512 40876 14552
rect 40916 14512 40925 14552
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 21091 13840 21100 13880
rect 21140 13840 30028 13880
rect 30068 13840 30077 13880
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 18691 12496 18700 12536
rect 18740 12496 21772 12536
rect 21812 12496 21821 12536
rect 11395 12328 11404 12368
rect 11444 12328 23960 12368
rect 23920 12284 23960 12328
rect 23920 12244 26188 12284
rect 26228 12244 26237 12284
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 14467 11740 14476 11780
rect 14516 11740 25516 11780
rect 25556 11740 25565 11780
rect 11875 11656 11884 11696
rect 11924 11656 32140 11696
rect 32180 11656 32189 11696
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 18595 11152 18604 11192
rect 18644 11152 20620 11192
rect 20660 11152 20669 11192
rect 32515 10984 32524 11024
rect 32564 10984 36172 11024
rect 36212 10984 36221 11024
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 32899 10144 32908 10184
rect 32948 10144 36556 10184
rect 36596 10144 36605 10184
rect 24835 10060 24844 10100
rect 24884 10060 43180 10100
rect 43220 10060 43229 10100
rect 24067 9976 24076 10016
rect 24116 9976 24940 10016
rect 24980 9976 24989 10016
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 21379 8800 21388 8840
rect 21428 8800 34060 8840
rect 34100 8800 34109 8840
rect 27715 8716 27724 8756
rect 27764 8716 28972 8756
rect 29012 8716 29021 8756
rect 19843 8464 19852 8504
rect 19892 8464 22636 8504
rect 22676 8464 22685 8504
rect 22531 8380 22540 8420
rect 22580 8380 24940 8420
rect 24980 8380 24989 8420
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 20803 8212 20812 8252
rect 20852 8212 26764 8252
rect 26804 8212 27532 8252
rect 27572 8212 27581 8252
rect 23203 8128 23212 8168
rect 23252 8128 23692 8168
rect 23732 8128 24364 8168
rect 24404 8128 24413 8168
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 23779 7120 23788 7160
rect 23828 7120 29836 7160
rect 29876 7120 29885 7160
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 27715 6532 27724 6572
rect 27764 6532 28972 6572
rect 29012 6532 32044 6572
rect 32084 6532 44716 6572
rect 44756 6532 44765 6572
rect 23395 6364 23404 6404
rect 23444 6364 43180 6404
rect 43220 6364 43229 6404
rect 32899 6280 32908 6320
rect 32948 6280 37820 6320
rect 37780 6236 37820 6280
rect 37780 6196 42220 6236
rect 42260 6196 42269 6236
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 20419 5020 20428 5060
rect 20468 5020 24460 5060
rect 24500 5020 24509 5060
rect 17251 4936 17260 4976
rect 17300 4936 21772 4976
rect 21812 4936 21821 4976
rect 21571 4852 21580 4892
rect 21620 4852 30316 4892
rect 30356 4852 30365 4892
rect 24451 4768 24460 4808
rect 24500 4768 30892 4808
rect 30932 4768 30941 4808
rect 24643 4684 24652 4724
rect 24692 4684 32908 4724
rect 32948 4684 32957 4724
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 25027 4516 25036 4556
rect 25076 4516 31852 4556
rect 31892 4516 31901 4556
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 21763 4264 21772 4304
rect 21812 4264 25324 4304
rect 25364 4264 25373 4304
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 15811 3256 15820 3296
rect 15860 3256 17644 3296
rect 17684 3256 21292 3296
rect 21332 3256 21341 3296
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 37843 94236 38600
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 38599 95476 38682
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676451365
transform 1 0 26400 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_0_0_clk
timestamp 1676451365
transform -1 0 8064 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk
timestamp 1676451365
transform -1 0 8256 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk
timestamp 1676451365
transform -1 0 15168 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk
timestamp 1676451365
transform 1 0 12960 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk
timestamp 1676451365
transform -1 0 7776 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk
timestamp 1676451365
transform -1 0 8640 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk
timestamp 1676451365
transform -1 0 16416 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk
timestamp 1676451365
transform -1 0 15936 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk
timestamp 1676451365
transform -1 0 38784 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk
timestamp 1676451365
transform 1 0 37728 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk
timestamp 1676451365
transform 1 0 44352 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk
timestamp 1676451365
transform -1 0 44352 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk
timestamp 1676451365
transform -1 0 33024 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk
timestamp 1676451365
transform -1 0 34272 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk
timestamp 1676451365
transform 1 0 40896 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk
timestamp 1676451365
transform -1 0 38400 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_0__f_clk
timestamp 1676451365
transform -1 0 5472 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_1__f_clk
timestamp 1676451365
transform -1 0 7776 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_2__f_clk
timestamp 1676451365
transform -1 0 5088 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_3__f_clk
timestamp 1676451365
transform 1 0 8640 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_4__f_clk
timestamp 1676451365
transform -1 0 14304 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_5__f_clk
timestamp 1676451365
transform 1 0 15840 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_6__f_clk
timestamp 1676451365
transform -1 0 12480 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_7__f_clk
timestamp 1676451365
transform 1 0 14592 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_8__f_clk
timestamp 1676451365
transform -1 0 4032 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_9__f_clk
timestamp 1676451365
transform -1 0 6816 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_10__f_clk
timestamp 1676451365
transform -1 0 5952 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_11__f_clk
timestamp 1676451365
transform 1 0 7872 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_12__f_clk
timestamp 1676451365
transform -1 0 13248 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_13__f_clk
timestamp 1676451365
transform 1 0 19392 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_14__f_clk
timestamp 1676451365
transform -1 0 14208 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_15__f_clk
timestamp 1676451365
transform 1 0 17280 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_16__f_clk
timestamp 1676451365
transform -1 0 37056 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_17__f_clk
timestamp 1676451365
transform 1 0 39264 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_18__f_clk
timestamp 1676451365
transform -1 0 38016 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_19__f_clk
timestamp 1676451365
transform 1 0 39360 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_20__f_clk
timestamp 1676451365
transform -1 0 43872 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_21__f_clk
timestamp 1676451365
transform 1 0 45984 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_22__f_clk
timestamp 1676451365
transform -1 0 43296 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_23__f_clk
timestamp 1676451365
transform 1 0 45216 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_24__f_clk
timestamp 1676451365
transform -1 0 28416 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_25__f_clk
timestamp 1676451365
transform -1 0 29472 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_26__f_clk
timestamp 1676451365
transform -1 0 30624 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_27__f_clk
timestamp 1676451365
transform -1 0 31872 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_28__f_clk
timestamp 1676451365
transform -1 0 45696 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_29__f_clk
timestamp 1676451365
transform 1 0 45696 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_30__f_clk
timestamp 1676451365
transform -1 0 35616 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_31__f_clk
timestamp 1676451365
transform 1 0 37920 0 -1 32508
box -48 -56 1296 834
use sg13g2_inv_1  clkload0
timestamp 1676382929
transform 1 0 6720 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  clkload1
timestamp 1676381911
transform 1 0 8640 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  clkload2
timestamp 1676381911
transform 1 0 9984 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  clkload3
timestamp 1676381911
transform 1 0 12672 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  clkload4
timestamp 1676381911
transform -1 0 35808 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  clkload5
timestamp 1676381911
transform -1 0 37536 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  clkload6
timestamp 1676381911
transform 1 0 41664 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  clkload7
timestamp 1676381911
transform 1 0 40320 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  clkload8
timestamp 1676381911
transform 1 0 26784 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  clkload9
timestamp 1676381911
transform 1 0 39552 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_8  fanout349
timestamp 1676451365
transform 1 0 31296 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout350
timestamp 1676451365
transform 1 0 31584 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout351
timestamp 1676451365
transform 1 0 25248 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout352
timestamp 1676451365
transform -1 0 17472 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout353
timestamp 1676451365
transform -1 0 26496 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout354
timestamp 1676451365
transform -1 0 27168 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout355
timestamp 1676451365
transform 1 0 32544 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  fanout356
timestamp 1676451365
transform 1 0 31776 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout357
timestamp 1676451365
transform -1 0 24000 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_8  fanout358
timestamp 1676451365
transform 1 0 22656 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout359
timestamp 1676451365
transform 1 0 30144 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_1  fanout360
timestamp 1676381911
transform 1 0 30624 0 1 14364
box -48 -56 432 834
use sg13g2_buf_8  fanout361
timestamp 1676451365
transform -1 0 25440 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout362
timestamp 1676451365
transform 1 0 31776 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  fanout363
timestamp 1676451365
transform 1 0 23808 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout364
timestamp 1676451365
transform 1 0 24096 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout365
timestamp 1676451365
transform 1 0 24480 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout366
timestamp 1676451365
transform -1 0 26784 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_2  fanout367
timestamp 1676381867
transform -1 0 27168 0 1 12852
box -48 -56 528 834
use sg13g2_buf_8  fanout368
timestamp 1676451365
transform -1 0 18912 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_1  fanout369
timestamp 1676381911
transform 1 0 16320 0 1 15876
box -48 -56 432 834
use sg13g2_buf_8  fanout370
timestamp 1676451365
transform 1 0 16800 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout371
timestamp 1676451365
transform -1 0 20544 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_2  fanout372
timestamp 1676381867
transform -1 0 20352 0 1 5292
box -48 -56 528 834
use sg13g2_buf_8  fanout373
timestamp 1676451365
transform 1 0 26688 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout374
timestamp 1676451365
transform -1 0 27744 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout375
timestamp 1676451365
transform 1 0 26688 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_1  fanout376
timestamp 1676381911
transform 1 0 27456 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_8  fanout377
timestamp 1676451365
transform -1 0 17952 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout378
timestamp 1676451365
transform -1 0 25440 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout379
timestamp 1676451365
transform -1 0 26304 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout380
timestamp 1676451365
transform 1 0 22080 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout381
timestamp 1676451365
transform -1 0 20352 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_1  fanout382
timestamp 1676381911
transform -1 0 24000 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_8  fanout383
timestamp 1676451365
transform -1 0 28896 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout384
timestamp 1676451365
transform -1 0 19392 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout385
timestamp 1676451365
transform -1 0 27648 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout386
timestamp 1676451365
transform -1 0 28224 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout387
timestamp 1676451365
transform 1 0 30048 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout388
timestamp 1676451365
transform -1 0 22368 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout389
timestamp 1676451365
transform 1 0 11424 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout390
timestamp 1676451365
transform 1 0 11520 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout391
timestamp 1676451365
transform 1 0 8064 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_2  fanout392
timestamp 1676381867
transform 1 0 38400 0 -1 8316
box -48 -56 528 834
use sg13g2_buf_8  fanout393
timestamp 1676451365
transform 1 0 26784 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout394
timestamp 1676451365
transform -1 0 26016 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_2  fanout395
timestamp 1676381867
transform 1 0 16416 0 1 26460
box -48 -56 528 834
use sg13g2_buf_1  fanout396
timestamp 1676381911
transform -1 0 28800 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_8  fanout397
timestamp 1676451365
transform 1 0 35904 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout398
timestamp 1676451365
transform 1 0 40416 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout399
timestamp 1676451365
transform 1 0 13920 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout400
timestamp 1676451365
transform -1 0 8064 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_1  fanout401
timestamp 1676381911
transform -1 0 6336 0 1 20412
box -48 -56 432 834
use sg13g2_buf_8  fanout402
timestamp 1676451365
transform 1 0 9984 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout403
timestamp 1676451365
transform -1 0 5760 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout404
timestamp 1676451365
transform -1 0 7776 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout405
timestamp 1676451365
transform -1 0 11520 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout406
timestamp 1676451365
transform -1 0 13056 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout407
timestamp 1676451365
transform 1 0 14976 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_1  fanout408
timestamp 1676381911
transform -1 0 16224 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout409
timestamp 1676381867
transform 1 0 3360 0 1 32508
box -48 -56 528 834
use sg13g2_buf_2  fanout410
timestamp 1676381867
transform 1 0 5664 0 -1 30996
box -48 -56 528 834
use sg13g2_buf_8  fanout411
timestamp 1676451365
transform -1 0 13344 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout412
timestamp 1676451365
transform -1 0 12576 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_2  fanout413
timestamp 1676381867
transform 1 0 11424 0 1 35532
box -48 -56 528 834
use sg13g2_buf_8  fanout414
timestamp 1676451365
transform -1 0 17760 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  fanout415
timestamp 1676451365
transform 1 0 15072 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_2  fanout416
timestamp 1676381867
transform -1 0 13824 0 -1 35532
box -48 -56 528 834
use sg13g2_buf_8  fanout417
timestamp 1676451365
transform 1 0 20352 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout418
timestamp 1676451365
transform -1 0 21312 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout419
timestamp 1676451365
transform 1 0 24192 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  fanout420
timestamp 1676451365
transform -1 0 22848 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_2  fanout421
timestamp 1676381867
transform 1 0 20544 0 1 30996
box -48 -56 528 834
use sg13g2_buf_8  fanout422
timestamp 1676451365
transform -1 0 21888 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout423
timestamp 1676451365
transform -1 0 41568 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout424
timestamp 1676451365
transform 1 0 35424 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout425
timestamp 1676451365
transform 1 0 32448 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout426
timestamp 1676451365
transform 1 0 34080 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout427
timestamp 1676451365
transform -1 0 33120 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_1  fanout428
timestamp 1676381911
transform -1 0 32736 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_8  fanout429
timestamp 1676451365
transform 1 0 34368 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_1  fanout430
timestamp 1676381911
transform 1 0 33408 0 1 32508
box -48 -56 432 834
use sg13g2_buf_2  fanout431
timestamp 1676381867
transform -1 0 34464 0 -1 30996
box -48 -56 528 834
use sg13g2_buf_8  fanout432
timestamp 1676451365
transform 1 0 38880 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout433
timestamp 1676451365
transform 1 0 48000 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout434
timestamp 1676451365
transform -1 0 48960 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout435
timestamp 1676451365
transform -1 0 44064 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout436
timestamp 1676451365
transform -1 0 45504 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_2  fanout437
timestamp 1676381867
transform -1 0 36096 0 1 27972
box -48 -56 528 834
use sg13g2_buf_1  fanout438
timestamp 1676381911
transform 1 0 32928 0 1 23436
box -48 -56 432 834
use sg13g2_buf_8  fanout439
timestamp 1676451365
transform -1 0 36864 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout440
timestamp 1676451365
transform -1 0 40032 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout441
timestamp 1676451365
transform -1 0 46848 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout442
timestamp 1676451365
transform 1 0 45312 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  fanout443
timestamp 1676451365
transform -1 0 44640 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout444
timestamp 1676451365
transform -1 0 43680 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout445
timestamp 1676451365
transform -1 0 46848 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout446
timestamp 1676451365
transform 1 0 19488 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_1  fanout447
timestamp 1676381911
transform 1 0 18720 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_8  fanout448
timestamp 1676451365
transform -1 0 31488 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_8  fanout449
timestamp 1676451365
transform -1 0 36384 0 -1 3780
box -48 -56 1296 834
use sg13g2_buf_8  fanout450
timestamp 1676451365
transform -1 0 36288 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout451
timestamp 1676451365
transform -1 0 38016 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_1  fanout452
timestamp 1676381911
transform -1 0 37152 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_8  fanout453
timestamp 1676451365
transform -1 0 36768 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout454
timestamp 1676451365
transform -1 0 16512 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout455
timestamp 1676451365
transform -1 0 16704 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  fanout456
timestamp 1676451365
transform 1 0 25728 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_2  fanout457
timestamp 1676381867
transform -1 0 27072 0 1 756
box -48 -56 528 834
use sg13g2_buf_8  fanout458
timestamp 1676451365
transform -1 0 25632 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_1  fanout459
timestamp 1676381911
transform 1 0 25248 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_8  fanout460
timestamp 1676451365
transform -1 0 35616 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_1  fanout461
timestamp 1676381911
transform -1 0 33984 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_8  fanout462
timestamp 1676451365
transform -1 0 31008 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout463
timestamp 1676451365
transform -1 0 38976 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout464
timestamp 1676451365
transform -1 0 39936 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout465
timestamp 1676451365
transform -1 0 42144 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout466
timestamp 1676451365
transform 1 0 37440 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout467
timestamp 1676451365
transform -1 0 22848 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_1  fanout468
timestamp 1676381911
transform -1 0 21984 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_8  fanout469
timestamp 1676451365
transform -1 0 25824 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout470
timestamp 1676451365
transform -1 0 24768 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout471
timestamp 1676451365
transform -1 0 9120 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout472
timestamp 1676451365
transform -1 0 28416 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout473
timestamp 1676451365
transform -1 0 31872 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_1  fanout474
timestamp 1676381911
transform -1 0 30240 0 1 26460
box -48 -56 432 834
use sg13g2_buf_8  fanout475
timestamp 1676451365
transform -1 0 29664 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout476
timestamp 1676451365
transform -1 0 14496 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout477
timestamp 1676451365
transform -1 0 14496 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout478
timestamp 1676451365
transform -1 0 17184 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout479
timestamp 1676451365
transform -1 0 23040 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout480
timestamp 1676451365
transform 1 0 22752 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout481
timestamp 1676451365
transform -1 0 24288 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout482
timestamp 1676451365
transform -1 0 32928 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout483
timestamp 1676451365
transform -1 0 31968 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout484
timestamp 1676451365
transform 1 0 37536 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout485
timestamp 1676451365
transform 1 0 38208 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout486
timestamp 1676451365
transform 1 0 28704 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout487
timestamp 1676451365
transform -1 0 29952 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout488
timestamp 1676451365
transform -1 0 11136 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout489
timestamp 1676451365
transform -1 0 12288 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout490
timestamp 1676451365
transform -1 0 14592 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_1  fanout491
timestamp 1676381911
transform 1 0 18816 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_8  fanout492
timestamp 1676451365
transform 1 0 13632 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout493
timestamp 1676451365
transform -1 0 15456 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout494
timestamp 1676451365
transform 1 0 4224 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout495
timestamp 1676451365
transform -1 0 12096 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout496
timestamp 1676451365
transform 1 0 9984 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_1  fanout497
timestamp 1676381911
transform -1 0 9504 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_8  fanout498
timestamp 1676451365
transform 1 0 11712 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  fanout499
timestamp 1676451365
transform -1 0 12384 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout500
timestamp 1676451365
transform -1 0 13920 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout501
timestamp 1676451365
transform 1 0 18048 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout502
timestamp 1676451365
transform 1 0 22944 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  fanout503
timestamp 1676451365
transform -1 0 24768 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout504
timestamp 1676451365
transform 1 0 14976 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout505
timestamp 1676451365
transform 1 0 33984 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout506
timestamp 1676451365
transform -1 0 35616 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout507
timestamp 1676451365
transform -1 0 48096 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout508
timestamp 1676451365
transform 1 0 43776 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout509
timestamp 1676451365
transform -1 0 43104 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout510
timestamp 1676451365
transform 1 0 33120 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout511
timestamp 1676451365
transform -1 0 33984 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout512
timestamp 1676451365
transform -1 0 36000 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout513
timestamp 1676451365
transform -1 0 45888 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_1  fanout514
timestamp 1676381911
transform -1 0 46464 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_8  fanout515
timestamp 1676451365
transform -1 0 45888 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_1  fanout516
timestamp 1676381911
transform 1 0 46464 0 1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout517
timestamp 1676381867
transform -1 0 45216 0 1 21924
box -48 -56 528 834
use sg13g2_buf_8  fanout518
timestamp 1676451365
transform 1 0 15456 0 -1 20412
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_168
timestamp 1679577901
transform 1 0 16704 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_172
timestamp 1677579658
transform 1 0 17088 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_177
timestamp 1679581782
transform 1 0 17568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_184
timestamp 1679581782
transform 1 0 18240 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_191
timestamp 1677580104
transform 1 0 18912 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_193
timestamp 1677579658
transform 1 0 19104 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_199
timestamp 1679581782
transform 1 0 19680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_206
timestamp 1679581782
transform 1 0 20352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_213
timestamp 1679581782
transform 1 0 21024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_220
timestamp 1679581782
transform 1 0 21696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_227
timestamp 1679581782
transform 1 0 22368 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_234
timestamp 1677580104
transform 1 0 23040 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_236
timestamp 1677579658
transform 1 0 23232 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_241
timestamp 1679581782
transform 1 0 23712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_248
timestamp 1679581782
transform 1 0 24384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_255
timestamp 1679581782
transform 1 0 25056 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_262
timestamp 1677580104
transform 1 0 25728 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_264
timestamp 1677579658
transform 1 0 25920 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_269
timestamp 1677580104
transform 1 0 26400 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_276
timestamp 1679581782
transform 1 0 27072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_283
timestamp 1679581782
transform 1 0 27744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_290
timestamp 1679581782
transform 1 0 28416 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_297
timestamp 1679577901
transform 1 0 29088 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_301
timestamp 1677579658
transform 1 0 29472 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_306
timestamp 1679581782
transform 1 0 29952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_313
timestamp 1679581782
transform 1 0 30624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_320
timestamp 1679581782
transform 1 0 31296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_327
timestamp 1679581782
transform 1 0 31968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_334
timestamp 1679581782
transform 1 0 32640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_341
timestamp 1679581782
transform 1 0 33312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_348
timestamp 1679581782
transform 1 0 33984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_355
timestamp 1679581782
transform 1 0 34656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_362
timestamp 1679581782
transform 1 0 35328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_369
timestamp 1679581782
transform 1 0 36000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_376
timestamp 1679581782
transform 1 0 36672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_383
timestamp 1679581782
transform 1 0 37344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_390
timestamp 1679581782
transform 1 0 38016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_397
timestamp 1679581782
transform 1 0 38688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_404
timestamp 1679581782
transform 1 0 39360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_411
timestamp 1679581782
transform 1 0 40032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_418
timestamp 1679581782
transform 1 0 40704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_425
timestamp 1679581782
transform 1 0 41376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_432
timestamp 1679581782
transform 1 0 42048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_439
timestamp 1679581782
transform 1 0 42720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_446
timestamp 1679581782
transform 1 0 43392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_453
timestamp 1679581782
transform 1 0 44064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_460
timestamp 1679581782
transform 1 0 44736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_467
timestamp 1679581782
transform 1 0 45408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_474
timestamp 1679581782
transform 1 0 46080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_481
timestamp 1679581782
transform 1 0 46752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_488
timestamp 1679581782
transform 1 0 47424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_495
timestamp 1679581782
transform 1 0 48096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_502
timestamp 1679581782
transform 1 0 48768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_509
timestamp 1679581782
transform 1 0 49440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_516
timestamp 1679581782
transform 1 0 50112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_523
timestamp 1679581782
transform 1 0 50784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_530
timestamp 1679581782
transform 1 0 51456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_537
timestamp 1679581782
transform 1 0 52128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_544
timestamp 1679581782
transform 1 0 52800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_551
timestamp 1679581782
transform 1 0 53472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_558
timestamp 1679581782
transform 1 0 54144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_565
timestamp 1679581782
transform 1 0 54816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_572
timestamp 1679581782
transform 1 0 55488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_579
timestamp 1679581782
transform 1 0 56160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_586
timestamp 1679581782
transform 1 0 56832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_593
timestamp 1679581782
transform 1 0 57504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_600
timestamp 1679581782
transform 1 0 58176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_607
timestamp 1679581782
transform 1 0 58848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_614
timestamp 1679581782
transform 1 0 59520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_621
timestamp 1679581782
transform 1 0 60192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_628
timestamp 1679581782
transform 1 0 60864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_635
timestamp 1679581782
transform 1 0 61536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_642
timestamp 1679581782
transform 1 0 62208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_649
timestamp 1679581782
transform 1 0 62880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_656
timestamp 1679581782
transform 1 0 63552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_663
timestamp 1679581782
transform 1 0 64224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_670
timestamp 1679581782
transform 1 0 64896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_677
timestamp 1679581782
transform 1 0 65568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_684
timestamp 1679581782
transform 1 0 66240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_691
timestamp 1679581782
transform 1 0 66912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_698
timestamp 1679581782
transform 1 0 67584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_705
timestamp 1679581782
transform 1 0 68256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_712
timestamp 1679581782
transform 1 0 68928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_719
timestamp 1679581782
transform 1 0 69600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_726
timestamp 1679581782
transform 1 0 70272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_733
timestamp 1679581782
transform 1 0 70944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_740
timestamp 1679581782
transform 1 0 71616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_747
timestamp 1679581782
transform 1 0 72288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_754
timestamp 1679581782
transform 1 0 72960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_761
timestamp 1679581782
transform 1 0 73632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_768
timestamp 1679581782
transform 1 0 74304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_775
timestamp 1679581782
transform 1 0 74976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_782
timestamp 1679581782
transform 1 0 75648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_789
timestamp 1679581782
transform 1 0 76320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_796
timestamp 1679581782
transform 1 0 76992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_803
timestamp 1679581782
transform 1 0 77664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_810
timestamp 1679581782
transform 1 0 78336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_817
timestamp 1679581782
transform 1 0 79008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_824
timestamp 1679581782
transform 1 0 79680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_831
timestamp 1679581782
transform 1 0 80352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_838
timestamp 1679581782
transform 1 0 81024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_845
timestamp 1679581782
transform 1 0 81696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_852
timestamp 1679581782
transform 1 0 82368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_859
timestamp 1679581782
transform 1 0 83040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_866
timestamp 1679581782
transform 1 0 83712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_873
timestamp 1679581782
transform 1 0 84384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_880
timestamp 1679581782
transform 1 0 85056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_887
timestamp 1679581782
transform 1 0 85728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_894
timestamp 1679581782
transform 1 0 86400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_901
timestamp 1679581782
transform 1 0 87072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_908
timestamp 1679581782
transform 1 0 87744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_915
timestamp 1679581782
transform 1 0 88416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_922
timestamp 1679581782
transform 1 0 89088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_929
timestamp 1679581782
transform 1 0 89760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_936
timestamp 1679581782
transform 1 0 90432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_943
timestamp 1679581782
transform 1 0 91104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_950
timestamp 1679581782
transform 1 0 91776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_957
timestamp 1679581782
transform 1 0 92448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_964
timestamp 1679581782
transform 1 0 93120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_971
timestamp 1679581782
transform 1 0 93792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_978
timestamp 1679581782
transform 1 0 94464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_985
timestamp 1679581782
transform 1 0 95136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_992
timestamp 1679581782
transform 1 0 95808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_999
timestamp 1679581782
transform 1 0 96480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1006
timestamp 1679581782
transform 1 0 97152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1013
timestamp 1679581782
transform 1 0 97824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1020
timestamp 1679581782
transform 1 0 98496 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_1027
timestamp 1677580104
transform 1 0 99168 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_161
timestamp 1677580104
transform 1 0 16032 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_185
timestamp 1677580104
transform 1 0 18336 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_224
timestamp 1677580104
transform 1 0 22080 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_226
timestamp 1677579658
transform 1 0 22272 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_231
timestamp 1677579658
transform 1 0 22752 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_259
timestamp 1677579658
transform 1 0 25440 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_288
timestamp 1679577901
transform 1 0 28224 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_292
timestamp 1677580104
transform 1 0 28608 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679581782
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679581782
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679581782
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679581782
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679581782
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679581782
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679581782
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679581782
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679581782
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679581782
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679581782
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679581782
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679581782
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679581782
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679581782
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_53
timestamp 1677579658
transform 1 0 5664 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_58
timestamp 1679581782
transform 1 0 6144 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_65
timestamp 1677580104
transform 1 0 6816 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_75
timestamp 1679577901
transform 1 0 7776 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_106
timestamp 1679581782
transform 1 0 10752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_113
timestamp 1679581782
transform 1 0 11424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_120
timestamp 1679581782
transform 1 0 12096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_127
timestamp 1679581782
transform 1 0 12768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_134
timestamp 1679581782
transform 1 0 13440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_141
timestamp 1679581782
transform 1 0 14112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_148
timestamp 1679581782
transform 1 0 14784 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_155
timestamp 1677580104
transform 1 0 15456 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_157
timestamp 1677579658
transform 1 0 15648 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_189
timestamp 1679577901
transform 1 0 18720 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_217
timestamp 1677580104
transform 1 0 21408 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_219
timestamp 1677579658
transform 1 0 21600 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_247
timestamp 1677579658
transform 1 0 24288 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_261
timestamp 1677579658
transform 1 0 25632 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_294
timestamp 1677580104
transform 1 0 28800 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_296
timestamp 1677579658
transform 1 0 28992 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_307
timestamp 1677580104
transform 1 0 30048 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_335
timestamp 1679577901
transform 1 0 32736 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_339
timestamp 1677579658
transform 1 0 33120 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_367
timestamp 1677579658
transform 1 0 35808 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_377
timestamp 1679581782
transform 1 0 36768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_394
timestamp 1679581782
transform 1 0 38400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_401
timestamp 1679581782
transform 1 0 39072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_408
timestamp 1679581782
transform 1 0 39744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_415
timestamp 1679581782
transform 1 0 40416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_422
timestamp 1679581782
transform 1 0 41088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_429
timestamp 1679581782
transform 1 0 41760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_436
timestamp 1679581782
transform 1 0 42432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_443
timestamp 1679581782
transform 1 0 43104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_450
timestamp 1679581782
transform 1 0 43776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_457
timestamp 1679581782
transform 1 0 44448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_464
timestamp 1679581782
transform 1 0 45120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_471
timestamp 1679581782
transform 1 0 45792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_478
timestamp 1679581782
transform 1 0 46464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_485
timestamp 1679581782
transform 1 0 47136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_492
timestamp 1679581782
transform 1 0 47808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_499
timestamp 1679581782
transform 1 0 48480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_506
timestamp 1679581782
transform 1 0 49152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_513
timestamp 1679581782
transform 1 0 49824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_520
timestamp 1679581782
transform 1 0 50496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_527
timestamp 1679581782
transform 1 0 51168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_534
timestamp 1679581782
transform 1 0 51840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_541
timestamp 1679581782
transform 1 0 52512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_548
timestamp 1679581782
transform 1 0 53184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_555
timestamp 1679581782
transform 1 0 53856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_562
timestamp 1679581782
transform 1 0 54528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_569
timestamp 1679581782
transform 1 0 55200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_576
timestamp 1679581782
transform 1 0 55872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_583
timestamp 1679581782
transform 1 0 56544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_590
timestamp 1679581782
transform 1 0 57216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_597
timestamp 1679581782
transform 1 0 57888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_604
timestamp 1679581782
transform 1 0 58560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_611
timestamp 1679581782
transform 1 0 59232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_618
timestamp 1679581782
transform 1 0 59904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_639
timestamp 1679581782
transform 1 0 61920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_646
timestamp 1679581782
transform 1 0 62592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_653
timestamp 1679581782
transform 1 0 63264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_660
timestamp 1679581782
transform 1 0 63936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_667
timestamp 1679581782
transform 1 0 64608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_674
timestamp 1679581782
transform 1 0 65280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_681
timestamp 1679581782
transform 1 0 65952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_688
timestamp 1679581782
transform 1 0 66624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_695
timestamp 1679581782
transform 1 0 67296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_702
timestamp 1679581782
transform 1 0 67968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_709
timestamp 1679581782
transform 1 0 68640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_730
timestamp 1679581782
transform 1 0 70656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_737
timestamp 1679581782
transform 1 0 71328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_744
timestamp 1679581782
transform 1 0 72000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_751
timestamp 1679581782
transform 1 0 72672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_758
timestamp 1679581782
transform 1 0 73344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_765
timestamp 1679581782
transform 1 0 74016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_772
timestamp 1679581782
transform 1 0 74688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_779
timestamp 1679581782
transform 1 0 75360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_786
timestamp 1679581782
transform 1 0 76032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_793
timestamp 1679581782
transform 1 0 76704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_800
timestamp 1679581782
transform 1 0 77376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_807
timestamp 1679581782
transform 1 0 78048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_814
timestamp 1679581782
transform 1 0 78720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_821
timestamp 1679581782
transform 1 0 79392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_828
timestamp 1679581782
transform 1 0 80064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_835
timestamp 1679581782
transform 1 0 80736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_842
timestamp 1679581782
transform 1 0 81408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_849
timestamp 1679581782
transform 1 0 82080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_856
timestamp 1679581782
transform 1 0 82752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_863
timestamp 1679581782
transform 1 0 83424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_870
timestamp 1679581782
transform 1 0 84096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_877
timestamp 1679581782
transform 1 0 84768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_884
timestamp 1679581782
transform 1 0 85440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_891
timestamp 1679581782
transform 1 0 86112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_898
timestamp 1679581782
transform 1 0 86784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_905
timestamp 1679581782
transform 1 0 87456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_912
timestamp 1679581782
transform 1 0 88128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_919
timestamp 1679581782
transform 1 0 88800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_926
timestamp 1679581782
transform 1 0 89472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_933
timestamp 1679581782
transform 1 0 90144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_940
timestamp 1679581782
transform 1 0 90816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_947
timestamp 1679581782
transform 1 0 91488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_954
timestamp 1679581782
transform 1 0 92160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_961
timestamp 1679581782
transform 1 0 92832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_968
timestamp 1679581782
transform 1 0 93504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_975
timestamp 1679581782
transform 1 0 94176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_982
timestamp 1679581782
transform 1 0 94848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_989
timestamp 1679581782
transform 1 0 95520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_996
timestamp 1679581782
transform 1 0 96192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1003
timestamp 1679581782
transform 1 0 96864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1010
timestamp 1679581782
transform 1 0 97536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1017
timestamp 1679581782
transform 1 0 98208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_1024
timestamp 1679577901
transform 1 0 98880 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_39
timestamp 1679577901
transform 1 0 4320 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_47
timestamp 1677580104
transform 1 0 5088 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_81
timestamp 1677580104
transform 1 0 8352 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_83
timestamp 1677579658
transform 1 0 8544 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_101
timestamp 1677580104
transform 1 0 10272 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_103
timestamp 1677579658
transform 1 0 10464 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_113
timestamp 1677580104
transform 1 0 11424 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_142
timestamp 1679581782
transform 1 0 14208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_149
timestamp 1679581782
transform 1 0 14880 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_156
timestamp 1677580104
transform 1 0 15552 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_183
timestamp 1679581782
transform 1 0 18144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_190
timestamp 1679577901
transform 1 0 18816 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_202
timestamp 1677580104
transform 1 0 19968 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_204
timestamp 1677579658
transform 1 0 20160 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_234
timestamp 1679577901
transform 1 0 23040 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_270
timestamp 1677580104
transform 1 0 26496 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_306
timestamp 1679581782
transform 1 0 29952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_313
timestamp 1679577901
transform 1 0 30624 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_317
timestamp 1677580104
transform 1 0 31008 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_329
timestamp 1677579658
transform 1 0 32160 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_334
timestamp 1677580104
transform 1 0 32640 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_349
timestamp 1677580104
transform 1 0 34080 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_373
timestamp 1679581782
transform 1 0 36384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_408
timestamp 1679581782
transform 1 0 39744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_415
timestamp 1679581782
transform 1 0 40416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_422
timestamp 1679581782
transform 1 0 41088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_429
timestamp 1679581782
transform 1 0 41760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_436
timestamp 1679581782
transform 1 0 42432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_443
timestamp 1679581782
transform 1 0 43104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_450
timestamp 1679581782
transform 1 0 43776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_457
timestamp 1679581782
transform 1 0 44448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_464
timestamp 1679581782
transform 1 0 45120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_471
timestamp 1679581782
transform 1 0 45792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_478
timestamp 1679581782
transform 1 0 46464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_485
timestamp 1679581782
transform 1 0 47136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_492
timestamp 1679581782
transform 1 0 47808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_499
timestamp 1679581782
transform 1 0 48480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_506
timestamp 1679581782
transform 1 0 49152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_513
timestamp 1679581782
transform 1 0 49824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_520
timestamp 1679581782
transform 1 0 50496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_527
timestamp 1679581782
transform 1 0 51168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_534
timestamp 1679581782
transform 1 0 51840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_541
timestamp 1679581782
transform 1 0 52512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_548
timestamp 1679581782
transform 1 0 53184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_555
timestamp 1679581782
transform 1 0 53856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_562
timestamp 1679581782
transform 1 0 54528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_569
timestamp 1679581782
transform 1 0 55200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_576
timestamp 1679581782
transform 1 0 55872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_583
timestamp 1679581782
transform 1 0 56544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_590
timestamp 1679581782
transform 1 0 57216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_597
timestamp 1679581782
transform 1 0 57888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_604
timestamp 1679581782
transform 1 0 58560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_611
timestamp 1679581782
transform 1 0 59232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_618
timestamp 1679581782
transform 1 0 59904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_625
timestamp 1679581782
transform 1 0 60576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_632
timestamp 1679581782
transform 1 0 61248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_639
timestamp 1679581782
transform 1 0 61920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_646
timestamp 1679581782
transform 1 0 62592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_653
timestamp 1679581782
transform 1 0 63264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_660
timestamp 1679581782
transform 1 0 63936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_667
timestamp 1679581782
transform 1 0 64608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_674
timestamp 1679581782
transform 1 0 65280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_681
timestamp 1679581782
transform 1 0 65952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_688
timestamp 1679581782
transform 1 0 66624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_695
timestamp 1679581782
transform 1 0 67296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_702
timestamp 1679581782
transform 1 0 67968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_709
timestamp 1679581782
transform 1 0 68640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_716
timestamp 1679581782
transform 1 0 69312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_723
timestamp 1679581782
transform 1 0 69984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_730
timestamp 1679581782
transform 1 0 70656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_737
timestamp 1679581782
transform 1 0 71328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_744
timestamp 1679581782
transform 1 0 72000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_751
timestamp 1679581782
transform 1 0 72672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_758
timestamp 1679581782
transform 1 0 73344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_765
timestamp 1679581782
transform 1 0 74016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_772
timestamp 1679581782
transform 1 0 74688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_779
timestamp 1679581782
transform 1 0 75360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_786
timestamp 1679581782
transform 1 0 76032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_793
timestamp 1679581782
transform 1 0 76704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_800
timestamp 1679581782
transform 1 0 77376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_807
timestamp 1679581782
transform 1 0 78048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_814
timestamp 1679581782
transform 1 0 78720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_821
timestamp 1679581782
transform 1 0 79392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_828
timestamp 1679581782
transform 1 0 80064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_835
timestamp 1679581782
transform 1 0 80736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_842
timestamp 1679581782
transform 1 0 81408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_849
timestamp 1679581782
transform 1 0 82080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_856
timestamp 1679581782
transform 1 0 82752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_863
timestamp 1679581782
transform 1 0 83424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_870
timestamp 1679581782
transform 1 0 84096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_877
timestamp 1679581782
transform 1 0 84768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_884
timestamp 1679581782
transform 1 0 85440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_891
timestamp 1679581782
transform 1 0 86112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_898
timestamp 1679581782
transform 1 0 86784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_905
timestamp 1679581782
transform 1 0 87456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_912
timestamp 1679581782
transform 1 0 88128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_919
timestamp 1679581782
transform 1 0 88800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_926
timestamp 1679581782
transform 1 0 89472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_933
timestamp 1679581782
transform 1 0 90144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_940
timestamp 1679581782
transform 1 0 90816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_947
timestamp 1679581782
transform 1 0 91488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_954
timestamp 1679581782
transform 1 0 92160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_961
timestamp 1679581782
transform 1 0 92832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_968
timestamp 1679581782
transform 1 0 93504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_975
timestamp 1679581782
transform 1 0 94176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_982
timestamp 1679581782
transform 1 0 94848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_989
timestamp 1679581782
transform 1 0 95520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_996
timestamp 1679581782
transform 1 0 96192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1003
timestamp 1679581782
transform 1 0 96864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1010
timestamp 1679581782
transform 1 0 97536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1017
timestamp 1679581782
transform 1 0 98208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_1024
timestamp 1679577901
transform 1 0 98880 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677579658
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_32
timestamp 1679577901
transform 1 0 3648 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_36
timestamp 1677580104
transform 1 0 4032 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_65
timestamp 1677579658
transform 1 0 6816 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_139
timestamp 1677579658
transform 1 0 13920 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_168
timestamp 1677580104
transform 1 0 16704 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_175
timestamp 1677580104
transform 1 0 17376 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_192
timestamp 1677580104
transform 1 0 19008 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_194
timestamp 1677579658
transform 1 0 19200 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_216
timestamp 1679581782
transform 1 0 21312 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_223
timestamp 1677580104
transform 1 0 21984 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_229
timestamp 1677580104
transform 1 0 22560 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_251
timestamp 1679577901
transform 1 0 24672 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_303
timestamp 1679581782
transform 1 0 29664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_310
timestamp 1679581782
transform 1 0 30336 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_317
timestamp 1677580104
transform 1 0 31008 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_319
timestamp 1677579658
transform 1 0 31200 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_365
timestamp 1677580104
transform 1 0 35616 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_421
timestamp 1679581782
transform 1 0 40992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_428
timestamp 1679581782
transform 1 0 41664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_435
timestamp 1679581782
transform 1 0 42336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_442
timestamp 1679581782
transform 1 0 43008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_449
timestamp 1679581782
transform 1 0 43680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_456
timestamp 1679581782
transform 1 0 44352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_463
timestamp 1679581782
transform 1 0 45024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_470
timestamp 1679581782
transform 1 0 45696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_477
timestamp 1679581782
transform 1 0 46368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_484
timestamp 1679581782
transform 1 0 47040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_491
timestamp 1679581782
transform 1 0 47712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_498
timestamp 1679581782
transform 1 0 48384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_505
timestamp 1679581782
transform 1 0 49056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_512
timestamp 1679581782
transform 1 0 49728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_519
timestamp 1679581782
transform 1 0 50400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_526
timestamp 1679581782
transform 1 0 51072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_533
timestamp 1679581782
transform 1 0 51744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_540
timestamp 1679581782
transform 1 0 52416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_547
timestamp 1679581782
transform 1 0 53088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_554
timestamp 1679581782
transform 1 0 53760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_561
timestamp 1679581782
transform 1 0 54432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_568
timestamp 1679581782
transform 1 0 55104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_575
timestamp 1679581782
transform 1 0 55776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_582
timestamp 1679581782
transform 1 0 56448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_589
timestamp 1679581782
transform 1 0 57120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_596
timestamp 1679581782
transform 1 0 57792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_603
timestamp 1679581782
transform 1 0 58464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_610
timestamp 1679581782
transform 1 0 59136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_617
timestamp 1679581782
transform 1 0 59808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_624
timestamp 1679581782
transform 1 0 60480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_631
timestamp 1679581782
transform 1 0 61152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_638
timestamp 1679581782
transform 1 0 61824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_645
timestamp 1679581782
transform 1 0 62496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_652
timestamp 1679581782
transform 1 0 63168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_659
timestamp 1679581782
transform 1 0 63840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_666
timestamp 1679581782
transform 1 0 64512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_673
timestamp 1679581782
transform 1 0 65184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_680
timestamp 1679581782
transform 1 0 65856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_687
timestamp 1679581782
transform 1 0 66528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_694
timestamp 1679581782
transform 1 0 67200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_701
timestamp 1679581782
transform 1 0 67872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_708
timestamp 1679581782
transform 1 0 68544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_715
timestamp 1679581782
transform 1 0 69216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_722
timestamp 1679581782
transform 1 0 69888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_729
timestamp 1679581782
transform 1 0 70560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_736
timestamp 1679581782
transform 1 0 71232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_743
timestamp 1679581782
transform 1 0 71904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_750
timestamp 1679581782
transform 1 0 72576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_757
timestamp 1679581782
transform 1 0 73248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_764
timestamp 1679581782
transform 1 0 73920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_771
timestamp 1679581782
transform 1 0 74592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_778
timestamp 1679581782
transform 1 0 75264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_785
timestamp 1679581782
transform 1 0 75936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_792
timestamp 1679581782
transform 1 0 76608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_799
timestamp 1679581782
transform 1 0 77280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_806
timestamp 1679581782
transform 1 0 77952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_813
timestamp 1679581782
transform 1 0 78624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_820
timestamp 1679581782
transform 1 0 79296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_827
timestamp 1679581782
transform 1 0 79968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_834
timestamp 1679581782
transform 1 0 80640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_841
timestamp 1679581782
transform 1 0 81312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_848
timestamp 1679581782
transform 1 0 81984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_855
timestamp 1679581782
transform 1 0 82656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_862
timestamp 1679581782
transform 1 0 83328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_869
timestamp 1679581782
transform 1 0 84000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_876
timestamp 1679581782
transform 1 0 84672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_883
timestamp 1679581782
transform 1 0 85344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_890
timestamp 1679581782
transform 1 0 86016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_897
timestamp 1679581782
transform 1 0 86688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_904
timestamp 1679581782
transform 1 0 87360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_911
timestamp 1679581782
transform 1 0 88032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_918
timestamp 1679581782
transform 1 0 88704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_925
timestamp 1679581782
transform 1 0 89376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_932
timestamp 1679581782
transform 1 0 90048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_939
timestamp 1679581782
transform 1 0 90720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_946
timestamp 1679581782
transform 1 0 91392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_953
timestamp 1679581782
transform 1 0 92064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_960
timestamp 1679581782
transform 1 0 92736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_967
timestamp 1679581782
transform 1 0 93408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_974
timestamp 1679581782
transform 1 0 94080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_981
timestamp 1679581782
transform 1 0 94752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_988
timestamp 1679581782
transform 1 0 95424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_995
timestamp 1679581782
transform 1 0 96096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1002
timestamp 1679581782
transform 1 0 96768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1009
timestamp 1679581782
transform 1 0 97440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1016
timestamp 1679581782
transform 1 0 98112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_1023
timestamp 1679577901
transform 1 0 98784 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_1027
timestamp 1677580104
transform 1 0 99168 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_39
timestamp 1677580104
transform 1 0 4320 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_54
timestamp 1677579658
transform 1 0 5760 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_78
timestamp 1679577901
transform 1 0 8064 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_82
timestamp 1677579658
transform 1 0 8448 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 10656 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_112
timestamp 1677579658
transform 1 0 11328 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_137
timestamp 1677580104
transform 1 0 13728 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_152
timestamp 1679581782
transform 1 0 15168 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_190
timestamp 1677580104
transform 1 0 18816 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_197
timestamp 1679577901
transform 1 0 19488 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_201
timestamp 1677579658
transform 1 0 19872 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_211
timestamp 1679577901
transform 1 0 20832 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_215
timestamp 1677579658
transform 1 0 21216 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_222
timestamp 1679581782
transform 1 0 21888 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_229
timestamp 1677579658
transform 1 0 22560 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_239
timestamp 1677579658
transform 1 0 23520 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_263
timestamp 1677580104
transform 1 0 25824 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_288
timestamp 1679577901
transform 1 0 28224 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_307
timestamp 1677579658
transform 1 0 30048 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_338
timestamp 1679577901
transform 1 0 33024 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_342
timestamp 1677580104
transform 1 0 33408 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_389
timestamp 1677579658
transform 1 0 37920 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_430
timestamp 1679581782
transform 1 0 41856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_437
timestamp 1679581782
transform 1 0 42528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_444
timestamp 1679581782
transform 1 0 43200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_451
timestamp 1679581782
transform 1 0 43872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_458
timestamp 1679581782
transform 1 0 44544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_465
timestamp 1679581782
transform 1 0 45216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_472
timestamp 1679581782
transform 1 0 45888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_479
timestamp 1679581782
transform 1 0 46560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_486
timestamp 1679581782
transform 1 0 47232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_493
timestamp 1679581782
transform 1 0 47904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_500
timestamp 1679581782
transform 1 0 48576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_507
timestamp 1679581782
transform 1 0 49248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_514
timestamp 1679581782
transform 1 0 49920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_521
timestamp 1679581782
transform 1 0 50592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_528
timestamp 1679581782
transform 1 0 51264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_535
timestamp 1679581782
transform 1 0 51936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_542
timestamp 1679581782
transform 1 0 52608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_549
timestamp 1679581782
transform 1 0 53280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_556
timestamp 1679581782
transform 1 0 53952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_563
timestamp 1679581782
transform 1 0 54624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_570
timestamp 1679581782
transform 1 0 55296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_577
timestamp 1679581782
transform 1 0 55968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_584
timestamp 1679581782
transform 1 0 56640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_591
timestamp 1679581782
transform 1 0 57312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_598
timestamp 1679581782
transform 1 0 57984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_605
timestamp 1679581782
transform 1 0 58656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_612
timestamp 1679581782
transform 1 0 59328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_619
timestamp 1679581782
transform 1 0 60000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_626
timestamp 1679581782
transform 1 0 60672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_633
timestamp 1679581782
transform 1 0 61344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_640
timestamp 1679581782
transform 1 0 62016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_647
timestamp 1679581782
transform 1 0 62688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_654
timestamp 1679581782
transform 1 0 63360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_661
timestamp 1679581782
transform 1 0 64032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_668
timestamp 1679581782
transform 1 0 64704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_675
timestamp 1679581782
transform 1 0 65376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_682
timestamp 1679581782
transform 1 0 66048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_689
timestamp 1679581782
transform 1 0 66720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_696
timestamp 1679581782
transform 1 0 67392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_703
timestamp 1679581782
transform 1 0 68064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_710
timestamp 1679581782
transform 1 0 68736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_717
timestamp 1679581782
transform 1 0 69408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_724
timestamp 1679581782
transform 1 0 70080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_731
timestamp 1679581782
transform 1 0 70752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_738
timestamp 1679581782
transform 1 0 71424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_745
timestamp 1679581782
transform 1 0 72096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_752
timestamp 1679581782
transform 1 0 72768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_759
timestamp 1679581782
transform 1 0 73440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_766
timestamp 1679581782
transform 1 0 74112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_773
timestamp 1679581782
transform 1 0 74784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_780
timestamp 1679581782
transform 1 0 75456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_787
timestamp 1679581782
transform 1 0 76128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_794
timestamp 1679581782
transform 1 0 76800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_801
timestamp 1679581782
transform 1 0 77472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679581782
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679581782
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_822
timestamp 1679581782
transform 1 0 79488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_829
timestamp 1679581782
transform 1 0 80160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_836
timestamp 1679581782
transform 1 0 80832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_843
timestamp 1679581782
transform 1 0 81504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_850
timestamp 1679581782
transform 1 0 82176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_857
timestamp 1679581782
transform 1 0 82848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_864
timestamp 1679581782
transform 1 0 83520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_871
timestamp 1679581782
transform 1 0 84192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_878
timestamp 1679581782
transform 1 0 84864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_885
timestamp 1679581782
transform 1 0 85536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_892
timestamp 1679581782
transform 1 0 86208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_899
timestamp 1679581782
transform 1 0 86880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_906
timestamp 1679581782
transform 1 0 87552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_913
timestamp 1679581782
transform 1 0 88224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_920
timestamp 1679581782
transform 1 0 88896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_927
timestamp 1679581782
transform 1 0 89568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_934
timestamp 1679581782
transform 1 0 90240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_941
timestamp 1679581782
transform 1 0 90912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_948
timestamp 1679581782
transform 1 0 91584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_955
timestamp 1679581782
transform 1 0 92256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_962
timestamp 1679581782
transform 1 0 92928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_969
timestamp 1679581782
transform 1 0 93600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_976
timestamp 1679581782
transform 1 0 94272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_983
timestamp 1679581782
transform 1 0 94944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_990
timestamp 1679581782
transform 1 0 95616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_997
timestamp 1679581782
transform 1 0 96288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1004
timestamp 1679581782
transform 1 0 96960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1011
timestamp 1679581782
transform 1 0 97632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1018
timestamp 1679581782
transform 1 0 98304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_1025
timestamp 1679577901
transform 1 0 98976 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_8
timestamp 1679581782
transform 1 0 1344 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_15
timestamp 1677580104
transform 1 0 2016 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 2592 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_28
timestamp 1677580104
transform 1 0 3264 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_67
timestamp 1677579658
transform 1 0 7008 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_84
timestamp 1677580104
transform 1 0 8640 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 9984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 10656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_112
timestamp 1679577901
transform 1 0 11328 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_116
timestamp 1677579658
transform 1 0 11712 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_122
timestamp 1679577901
transform 1 0 12288 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_126
timestamp 1677580104
transform 1 0 12672 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_184
timestamp 1677580104
transform 1 0 18240 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_200
timestamp 1677579658
transform 1 0 19776 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_206
timestamp 1677579658
transform 1 0 20352 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_214
timestamp 1677579658
transform 1 0 21120 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_219
timestamp 1679577901
transform 1 0 21600 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_230
timestamp 1677580104
transform 1 0 22656 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_232
timestamp 1677579658
transform 1 0 22848 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_255
timestamp 1679581782
transform 1 0 25056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_262
timestamp 1679577901
transform 1 0 25728 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_266
timestamp 1677579658
transform 1 0 26112 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_285
timestamp 1677580104
transform 1 0 27936 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_300
timestamp 1677580104
transform 1 0 29376 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_307
timestamp 1679581782
transform 1 0 30048 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_314
timestamp 1677580104
transform 1 0 30720 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_316
timestamp 1677579658
transform 1 0 30912 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_344
timestamp 1679581782
transform 1 0 33600 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_351
timestamp 1677579658
transform 1 0 34272 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_384
timestamp 1677579658
transform 1 0 37440 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_394
timestamp 1677579658
transform 1 0 38400 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_407
timestamp 1677579658
transform 1 0 39648 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_422
timestamp 1679581782
transform 1 0 41088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_429
timestamp 1679577901
transform 1 0 41760 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_442
timestamp 1679581782
transform 1 0 43008 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_449
timestamp 1677580104
transform 1 0 43680 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_464
timestamp 1679581782
transform 1 0 45120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_471
timestamp 1679581782
transform 1 0 45792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_478
timestamp 1679581782
transform 1 0 46464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_485
timestamp 1679581782
transform 1 0 47136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_492
timestamp 1679581782
transform 1 0 47808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_499
timestamp 1679581782
transform 1 0 48480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_506
timestamp 1679581782
transform 1 0 49152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_513
timestamp 1679581782
transform 1 0 49824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_520
timestamp 1679581782
transform 1 0 50496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_527
timestamp 1679581782
transform 1 0 51168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_534
timestamp 1679581782
transform 1 0 51840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_541
timestamp 1679581782
transform 1 0 52512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_548
timestamp 1679581782
transform 1 0 53184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_555
timestamp 1679581782
transform 1 0 53856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_562
timestamp 1679581782
transform 1 0 54528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_569
timestamp 1679581782
transform 1 0 55200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_576
timestamp 1679581782
transform 1 0 55872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_583
timestamp 1679581782
transform 1 0 56544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_590
timestamp 1679581782
transform 1 0 57216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_597
timestamp 1679581782
transform 1 0 57888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_604
timestamp 1679581782
transform 1 0 58560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_611
timestamp 1679581782
transform 1 0 59232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_618
timestamp 1679581782
transform 1 0 59904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_625
timestamp 1679581782
transform 1 0 60576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_632
timestamp 1679581782
transform 1 0 61248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_639
timestamp 1679581782
transform 1 0 61920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_646
timestamp 1679581782
transform 1 0 62592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_653
timestamp 1679581782
transform 1 0 63264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_660
timestamp 1679581782
transform 1 0 63936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_667
timestamp 1679581782
transform 1 0 64608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_674
timestamp 1679581782
transform 1 0 65280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_681
timestamp 1679581782
transform 1 0 65952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_688
timestamp 1679581782
transform 1 0 66624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_695
timestamp 1679581782
transform 1 0 67296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_702
timestamp 1679581782
transform 1 0 67968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_709
timestamp 1679581782
transform 1 0 68640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_716
timestamp 1679581782
transform 1 0 69312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_723
timestamp 1679581782
transform 1 0 69984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_730
timestamp 1679581782
transform 1 0 70656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_737
timestamp 1679581782
transform 1 0 71328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_744
timestamp 1679581782
transform 1 0 72000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_751
timestamp 1679581782
transform 1 0 72672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_758
timestamp 1679581782
transform 1 0 73344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_765
timestamp 1679581782
transform 1 0 74016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_772
timestamp 1679581782
transform 1 0 74688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_779
timestamp 1679581782
transform 1 0 75360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_786
timestamp 1679581782
transform 1 0 76032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_793
timestamp 1679581782
transform 1 0 76704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_800
timestamp 1679581782
transform 1 0 77376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_807
timestamp 1679581782
transform 1 0 78048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_814
timestamp 1679581782
transform 1 0 78720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_821
timestamp 1679581782
transform 1 0 79392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_828
timestamp 1679581782
transform 1 0 80064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_835
timestamp 1679581782
transform 1 0 80736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_842
timestamp 1679581782
transform 1 0 81408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_849
timestamp 1679581782
transform 1 0 82080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_856
timestamp 1679581782
transform 1 0 82752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_863
timestamp 1679581782
transform 1 0 83424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_870
timestamp 1679581782
transform 1 0 84096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_877
timestamp 1679581782
transform 1 0 84768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_884
timestamp 1679581782
transform 1 0 85440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_891
timestamp 1679581782
transform 1 0 86112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_898
timestamp 1679581782
transform 1 0 86784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_905
timestamp 1679581782
transform 1 0 87456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_912
timestamp 1679581782
transform 1 0 88128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_919
timestamp 1679581782
transform 1 0 88800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_926
timestamp 1679581782
transform 1 0 89472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_933
timestamp 1679581782
transform 1 0 90144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_940
timestamp 1679581782
transform 1 0 90816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_947
timestamp 1679581782
transform 1 0 91488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_954
timestamp 1679581782
transform 1 0 92160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_961
timestamp 1679581782
transform 1 0 92832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_968
timestamp 1679581782
transform 1 0 93504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_975
timestamp 1679581782
transform 1 0 94176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_982
timestamp 1679581782
transform 1 0 94848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_989
timestamp 1679581782
transform 1 0 95520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_996
timestamp 1679581782
transform 1 0 96192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1003
timestamp 1679581782
transform 1 0 96864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1010
timestamp 1679581782
transform 1 0 97536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1017
timestamp 1679581782
transform 1 0 98208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_1024
timestamp 1679577901
transform 1 0 98880 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677579658
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_4
timestamp 1677580104
transform 1 0 960 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_6
timestamp 1677579658
transform 1 0 1152 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_11
timestamp 1679577901
transform 1 0 1632 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_15
timestamp 1677579658
transform 1 0 2016 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_28
timestamp 1677580104
transform 1 0 3264 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_30
timestamp 1677579658
transform 1 0 3456 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_49
timestamp 1677579658
transform 1 0 5280 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_76
timestamp 1677580104
transform 1 0 7872 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_78
timestamp 1677579658
transform 1 0 8064 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_129
timestamp 1679577901
transform 1 0 12960 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_133
timestamp 1677580104
transform 1 0 13344 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_144
timestamp 1679581782
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_151
timestamp 1679577901
transform 1 0 15072 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_177
timestamp 1677580104
transform 1 0 17568 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_179
timestamp 1677579658
transform 1 0 17760 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_186
timestamp 1677580104
transform 1 0 18432 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_188
timestamp 1677579658
transform 1 0 18624 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_204
timestamp 1679581782
transform 1 0 20160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_211
timestamp 1679581782
transform 1 0 20832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_218
timestamp 1679581782
transform 1 0 21504 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_225
timestamp 1677580104
transform 1 0 22176 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_227
timestamp 1677579658
transform 1 0 22368 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_250
timestamp 1679581782
transform 1 0 24576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_257
timestamp 1679581782
transform 1 0 25248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_264
timestamp 1679581782
transform 1 0 25920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_271
timestamp 1679577901
transform 1 0 26592 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_275
timestamp 1677580104
transform 1 0 26976 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_283
timestamp 1679577901
transform 1 0 27744 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_309
timestamp 1679581782
transform 1 0 30240 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_316
timestamp 1677580104
transform 1 0 30912 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_318
timestamp 1677579658
transform 1 0 31104 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_383
timestamp 1677579658
transform 1 0 37344 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_400
timestamp 1677580104
transform 1 0 38976 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_486
timestamp 1679581782
transform 1 0 47232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_493
timestamp 1679581782
transform 1 0 47904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_500
timestamp 1679581782
transform 1 0 48576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_507
timestamp 1679581782
transform 1 0 49248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_514
timestamp 1679581782
transform 1 0 49920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_521
timestamp 1679581782
transform 1 0 50592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_528
timestamp 1679581782
transform 1 0 51264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_535
timestamp 1679581782
transform 1 0 51936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_542
timestamp 1679581782
transform 1 0 52608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_549
timestamp 1679581782
transform 1 0 53280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_556
timestamp 1679581782
transform 1 0 53952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_563
timestamp 1679581782
transform 1 0 54624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_570
timestamp 1679581782
transform 1 0 55296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_577
timestamp 1679581782
transform 1 0 55968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_584
timestamp 1679581782
transform 1 0 56640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_591
timestamp 1679581782
transform 1 0 57312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_598
timestamp 1679581782
transform 1 0 57984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_605
timestamp 1679581782
transform 1 0 58656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_612
timestamp 1679581782
transform 1 0 59328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_619
timestamp 1679581782
transform 1 0 60000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_626
timestamp 1679581782
transform 1 0 60672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_633
timestamp 1679581782
transform 1 0 61344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_640
timestamp 1679581782
transform 1 0 62016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_647
timestamp 1679581782
transform 1 0 62688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_654
timestamp 1679581782
transform 1 0 63360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_661
timestamp 1679581782
transform 1 0 64032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_668
timestamp 1679581782
transform 1 0 64704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_675
timestamp 1679581782
transform 1 0 65376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_682
timestamp 1679581782
transform 1 0 66048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_689
timestamp 1679581782
transform 1 0 66720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_696
timestamp 1679581782
transform 1 0 67392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_703
timestamp 1679581782
transform 1 0 68064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_710
timestamp 1679581782
transform 1 0 68736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_717
timestamp 1679581782
transform 1 0 69408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_724
timestamp 1679581782
transform 1 0 70080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_731
timestamp 1679581782
transform 1 0 70752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_738
timestamp 1679581782
transform 1 0 71424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_745
timestamp 1679581782
transform 1 0 72096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_752
timestamp 1679581782
transform 1 0 72768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_759
timestamp 1679581782
transform 1 0 73440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_766
timestamp 1679581782
transform 1 0 74112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_773
timestamp 1679581782
transform 1 0 74784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_780
timestamp 1679581782
transform 1 0 75456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_787
timestamp 1679581782
transform 1 0 76128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_794
timestamp 1679581782
transform 1 0 76800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_801
timestamp 1679581782
transform 1 0 77472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_808
timestamp 1679581782
transform 1 0 78144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_815
timestamp 1679581782
transform 1 0 78816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_822
timestamp 1679581782
transform 1 0 79488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_829
timestamp 1679581782
transform 1 0 80160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_836
timestamp 1679581782
transform 1 0 80832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_843
timestamp 1679581782
transform 1 0 81504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_850
timestamp 1679581782
transform 1 0 82176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_857
timestamp 1679581782
transform 1 0 82848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_864
timestamp 1679581782
transform 1 0 83520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_871
timestamp 1679581782
transform 1 0 84192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_878
timestamp 1679581782
transform 1 0 84864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_885
timestamp 1679581782
transform 1 0 85536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_892
timestamp 1679581782
transform 1 0 86208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_899
timestamp 1679581782
transform 1 0 86880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_906
timestamp 1679581782
transform 1 0 87552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_913
timestamp 1679581782
transform 1 0 88224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_920
timestamp 1679581782
transform 1 0 88896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_927
timestamp 1679581782
transform 1 0 89568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_934
timestamp 1679581782
transform 1 0 90240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_941
timestamp 1679581782
transform 1 0 90912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_948
timestamp 1679581782
transform 1 0 91584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_955
timestamp 1679581782
transform 1 0 92256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_962
timestamp 1679581782
transform 1 0 92928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_969
timestamp 1679581782
transform 1 0 93600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_976
timestamp 1679581782
transform 1 0 94272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_983
timestamp 1679581782
transform 1 0 94944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_990
timestamp 1679581782
transform 1 0 95616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_997
timestamp 1679581782
transform 1 0 96288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1004
timestamp 1679581782
transform 1 0 96960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1011
timestamp 1679581782
transform 1 0 97632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1018
timestamp 1679581782
transform 1 0 98304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_1025
timestamp 1679577901
transform 1 0 98976 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_0
timestamp 1677580104
transform 1 0 576 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_82
timestamp 1677579658
transform 1 0 8448 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_96
timestamp 1677580104
transform 1 0 9792 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_111
timestamp 1677579658
transform 1 0 11232 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_121
timestamp 1679581782
transform 1 0 12192 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_128
timestamp 1677580104
transform 1 0 12864 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_200
timestamp 1679577901
transform 1 0 19776 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_204
timestamp 1677580104
transform 1 0 20160 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_221
timestamp 1679577901
transform 1 0 21792 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1679581782
transform 1 0 25440 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_266
timestamp 1677580104
transform 1 0 26112 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_272
timestamp 1679577901
transform 1 0 26688 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_285
timestamp 1679581782
transform 1 0 27936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_292
timestamp 1679577901
transform 1 0 28608 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_317
timestamp 1677580104
transform 1 0 31008 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_319
timestamp 1677579658
transform 1 0 31200 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_327
timestamp 1677580104
transform 1 0 31968 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_341
timestamp 1679581782
transform 1 0 33312 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_348
timestamp 1677579658
transform 1 0 33984 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_356
timestamp 1677579658
transform 1 0 34752 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_380
timestamp 1677580104
transform 1 0 37056 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_442
timestamp 1677579658
transform 1 0 43008 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_467
timestamp 1677579658
transform 1 0 45408 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_485
timestamp 1679581782
transform 1 0 47136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_492
timestamp 1679581782
transform 1 0 47808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_499
timestamp 1679581782
transform 1 0 48480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_506
timestamp 1679581782
transform 1 0 49152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_513
timestamp 1679581782
transform 1 0 49824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_520
timestamp 1679581782
transform 1 0 50496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_527
timestamp 1679581782
transform 1 0 51168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_534
timestamp 1679581782
transform 1 0 51840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_541
timestamp 1679581782
transform 1 0 52512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_548
timestamp 1679581782
transform 1 0 53184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_555
timestamp 1679581782
transform 1 0 53856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_562
timestamp 1679581782
transform 1 0 54528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_569
timestamp 1679581782
transform 1 0 55200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_576
timestamp 1679581782
transform 1 0 55872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_583
timestamp 1679581782
transform 1 0 56544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_590
timestamp 1679581782
transform 1 0 57216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_597
timestamp 1679581782
transform 1 0 57888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_604
timestamp 1679581782
transform 1 0 58560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_611
timestamp 1679581782
transform 1 0 59232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_618
timestamp 1679581782
transform 1 0 59904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_625
timestamp 1679581782
transform 1 0 60576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_632
timestamp 1679581782
transform 1 0 61248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_639
timestamp 1679581782
transform 1 0 61920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_646
timestamp 1679581782
transform 1 0 62592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_653
timestamp 1679581782
transform 1 0 63264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_660
timestamp 1679581782
transform 1 0 63936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_667
timestamp 1679581782
transform 1 0 64608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_674
timestamp 1679581782
transform 1 0 65280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_681
timestamp 1679581782
transform 1 0 65952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_688
timestamp 1679581782
transform 1 0 66624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_695
timestamp 1679581782
transform 1 0 67296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_702
timestamp 1679581782
transform 1 0 67968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_709
timestamp 1679581782
transform 1 0 68640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_716
timestamp 1679581782
transform 1 0 69312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_723
timestamp 1679581782
transform 1 0 69984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_730
timestamp 1679581782
transform 1 0 70656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_737
timestamp 1679581782
transform 1 0 71328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_744
timestamp 1679581782
transform 1 0 72000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_751
timestamp 1679581782
transform 1 0 72672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_758
timestamp 1679581782
transform 1 0 73344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679581782
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679581782
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_779
timestamp 1679581782
transform 1 0 75360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_786
timestamp 1679581782
transform 1 0 76032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_793
timestamp 1679581782
transform 1 0 76704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_800
timestamp 1679581782
transform 1 0 77376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_807
timestamp 1679581782
transform 1 0 78048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_814
timestamp 1679581782
transform 1 0 78720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_821
timestamp 1679581782
transform 1 0 79392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_828
timestamp 1679581782
transform 1 0 80064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_835
timestamp 1679581782
transform 1 0 80736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_842
timestamp 1679581782
transform 1 0 81408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_849
timestamp 1679581782
transform 1 0 82080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_856
timestamp 1679581782
transform 1 0 82752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_863
timestamp 1679581782
transform 1 0 83424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_870
timestamp 1679581782
transform 1 0 84096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_877
timestamp 1679581782
transform 1 0 84768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_884
timestamp 1679581782
transform 1 0 85440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_891
timestamp 1679581782
transform 1 0 86112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_898
timestamp 1679581782
transform 1 0 86784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_905
timestamp 1679581782
transform 1 0 87456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_912
timestamp 1679581782
transform 1 0 88128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_919
timestamp 1679581782
transform 1 0 88800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_926
timestamp 1679581782
transform 1 0 89472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_933
timestamp 1679581782
transform 1 0 90144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_940
timestamp 1679581782
transform 1 0 90816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_947
timestamp 1679581782
transform 1 0 91488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_954
timestamp 1679581782
transform 1 0 92160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_961
timestamp 1679581782
transform 1 0 92832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_968
timestamp 1679581782
transform 1 0 93504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_975
timestamp 1679581782
transform 1 0 94176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_982
timestamp 1679581782
transform 1 0 94848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_989
timestamp 1679581782
transform 1 0 95520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_996
timestamp 1679581782
transform 1 0 96192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1003
timestamp 1679581782
transform 1 0 96864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1010
timestamp 1679581782
transform 1 0 97536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1017
timestamp 1679581782
transform 1 0 98208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_1024
timestamp 1679577901
transform 1 0 98880 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_1028
timestamp 1677579658
transform 1 0 99264 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1677580104
transform 1 0 576 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_21
timestamp 1677580104
transform 1 0 2592 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_90
timestamp 1677580104
transform 1 0 9216 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_111
timestamp 1679577901
transform 1 0 11232 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_142
timestamp 1679577901
transform 1 0 14208 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_146
timestamp 1677580104
transform 1 0 14592 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_152
timestamp 1679577901
transform 1 0 15168 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_156
timestamp 1677580104
transform 1 0 15552 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_184
timestamp 1679577901
transform 1 0 18240 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_188
timestamp 1677580104
transform 1 0 18624 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_194
timestamp 1679581782
transform 1 0 19200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_201
timestamp 1679577901
transform 1 0 19872 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_221
timestamp 1679577901
transform 1 0 21792 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_225
timestamp 1677579658
transform 1 0 22176 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_245
timestamp 1677580104
transform 1 0 24096 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_247
timestamp 1677579658
transform 1 0 24288 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_271
timestamp 1679577901
transform 1 0 26592 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_286
timestamp 1679581782
transform 1 0 28032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_293
timestamp 1679581782
transform 1 0 28704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_300
timestamp 1679577901
transform 1 0 29376 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_309
timestamp 1679581782
transform 1 0 30240 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_316
timestamp 1677580104
transform 1 0 30912 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_324
timestamp 1677579658
transform 1 0 31680 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_331
timestamp 1679581782
transform 1 0 32352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_338
timestamp 1679581782
transform 1 0 33024 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_345
timestamp 1677580104
transform 1 0 33696 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_347
timestamp 1677579658
transform 1 0 33888 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_383
timestamp 1677579658
transform 1 0 37344 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_427
timestamp 1677580104
transform 1 0 41568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_457
timestamp 1677580104
transform 1 0 44448 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_459
timestamp 1677579658
transform 1 0 44640 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_488
timestamp 1679581782
transform 1 0 47424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_495
timestamp 1679581782
transform 1 0 48096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_502
timestamp 1679581782
transform 1 0 48768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_509
timestamp 1679581782
transform 1 0 49440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_516
timestamp 1679581782
transform 1 0 50112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_523
timestamp 1679581782
transform 1 0 50784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_530
timestamp 1679581782
transform 1 0 51456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_537
timestamp 1679581782
transform 1 0 52128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_544
timestamp 1679581782
transform 1 0 52800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_551
timestamp 1679581782
transform 1 0 53472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_558
timestamp 1679581782
transform 1 0 54144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_565
timestamp 1679581782
transform 1 0 54816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_572
timestamp 1679581782
transform 1 0 55488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_579
timestamp 1679581782
transform 1 0 56160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_586
timestamp 1679581782
transform 1 0 56832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_593
timestamp 1679581782
transform 1 0 57504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_600
timestamp 1679581782
transform 1 0 58176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_607
timestamp 1679581782
transform 1 0 58848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_614
timestamp 1679581782
transform 1 0 59520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_621
timestamp 1679581782
transform 1 0 60192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_628
timestamp 1679581782
transform 1 0 60864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_635
timestamp 1679581782
transform 1 0 61536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_642
timestamp 1679581782
transform 1 0 62208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_649
timestamp 1679581782
transform 1 0 62880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_656
timestamp 1679581782
transform 1 0 63552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_663
timestamp 1679581782
transform 1 0 64224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_670
timestamp 1679581782
transform 1 0 64896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_677
timestamp 1679581782
transform 1 0 65568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_684
timestamp 1679581782
transform 1 0 66240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_691
timestamp 1679581782
transform 1 0 66912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_698
timestamp 1679581782
transform 1 0 67584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_705
timestamp 1679581782
transform 1 0 68256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_712
timestamp 1679581782
transform 1 0 68928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_719
timestamp 1679581782
transform 1 0 69600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_726
timestamp 1679581782
transform 1 0 70272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_733
timestamp 1679581782
transform 1 0 70944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_740
timestamp 1679581782
transform 1 0 71616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_747
timestamp 1679581782
transform 1 0 72288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_754
timestamp 1679581782
transform 1 0 72960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_761
timestamp 1679581782
transform 1 0 73632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_768
timestamp 1679581782
transform 1 0 74304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_775
timestamp 1679581782
transform 1 0 74976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_782
timestamp 1679581782
transform 1 0 75648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_789
timestamp 1679581782
transform 1 0 76320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_796
timestamp 1679581782
transform 1 0 76992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_803
timestamp 1679581782
transform 1 0 77664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_810
timestamp 1679581782
transform 1 0 78336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_817
timestamp 1679581782
transform 1 0 79008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_824
timestamp 1679581782
transform 1 0 79680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_831
timestamp 1679581782
transform 1 0 80352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_838
timestamp 1679581782
transform 1 0 81024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_845
timestamp 1679581782
transform 1 0 81696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_852
timestamp 1679581782
transform 1 0 82368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_859
timestamp 1679581782
transform 1 0 83040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_866
timestamp 1679581782
transform 1 0 83712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_873
timestamp 1679581782
transform 1 0 84384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_880
timestamp 1679581782
transform 1 0 85056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_887
timestamp 1679581782
transform 1 0 85728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_894
timestamp 1679581782
transform 1 0 86400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_901
timestamp 1679581782
transform 1 0 87072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_908
timestamp 1679581782
transform 1 0 87744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_915
timestamp 1679581782
transform 1 0 88416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_922
timestamp 1679581782
transform 1 0 89088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_929
timestamp 1679581782
transform 1 0 89760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_936
timestamp 1679581782
transform 1 0 90432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_943
timestamp 1679581782
transform 1 0 91104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_950
timestamp 1679581782
transform 1 0 91776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_957
timestamp 1679581782
transform 1 0 92448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_964
timestamp 1679581782
transform 1 0 93120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_971
timestamp 1679581782
transform 1 0 93792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_978
timestamp 1679581782
transform 1 0 94464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_985
timestamp 1679581782
transform 1 0 95136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_992
timestamp 1679581782
transform 1 0 95808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_999
timestamp 1679581782
transform 1 0 96480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1006
timestamp 1679581782
transform 1 0 97152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1013
timestamp 1679581782
transform 1 0 97824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1020
timestamp 1679581782
transform 1 0 98496 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_1027
timestamp 1677580104
transform 1 0 99168 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_91
timestamp 1677580104
transform 1 0 9312 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_93
timestamp 1677579658
transform 1 0 9504 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_98
timestamp 1679577901
transform 1 0 9984 0 1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_10_107
timestamp 1679577901
transform 1 0 10848 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_111
timestamp 1677579658
transform 1 0 11232 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_124
timestamp 1679581782
transform 1 0 12480 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_131
timestamp 1677580104
transform 1 0 13152 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_146
timestamp 1679581782
transform 1 0 14592 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_153
timestamp 1677580104
transform 1 0 15264 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_181
timestamp 1677580104
transform 1 0 17952 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_183
timestamp 1677579658
transform 1 0 18144 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_192
timestamp 1679581782
transform 1 0 19008 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_210
timestamp 1677579658
transform 1 0 20736 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_225
timestamp 1679577901
transform 1 0 22176 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_229
timestamp 1677579658
transform 1 0 22560 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_256
timestamp 1679577901
transform 1 0 25152 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_260
timestamp 1677579658
transform 1 0 25536 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_264
timestamp 1677580104
transform 1 0 25920 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_271
timestamp 1679577901
transform 1 0 26592 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_275
timestamp 1677579658
transform 1 0 26976 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_293
timestamp 1677579658
transform 1 0 28704 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_314
timestamp 1679581782
transform 1 0 30720 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_321
timestamp 1677579658
transform 1 0 31392 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_338
timestamp 1679577901
transform 1 0 33024 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_342
timestamp 1677579658
transform 1 0 33408 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_373
timestamp 1679581782
transform 1 0 36384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_380
timestamp 1679577901
transform 1 0 37056 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_384
timestamp 1677579658
transform 1 0 37440 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_507
timestamp 1679581782
transform 1 0 49248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_514
timestamp 1679581782
transform 1 0 49920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_521
timestamp 1679581782
transform 1 0 50592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_528
timestamp 1679581782
transform 1 0 51264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_535
timestamp 1679581782
transform 1 0 51936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_542
timestamp 1679581782
transform 1 0 52608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_549
timestamp 1679581782
transform 1 0 53280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_556
timestamp 1679581782
transform 1 0 53952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_563
timestamp 1679581782
transform 1 0 54624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_570
timestamp 1679581782
transform 1 0 55296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_577
timestamp 1679581782
transform 1 0 55968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_584
timestamp 1679581782
transform 1 0 56640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_591
timestamp 1679581782
transform 1 0 57312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_598
timestamp 1679581782
transform 1 0 57984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_605
timestamp 1679581782
transform 1 0 58656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_612
timestamp 1679581782
transform 1 0 59328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_619
timestamp 1679581782
transform 1 0 60000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_626
timestamp 1679581782
transform 1 0 60672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_633
timestamp 1679581782
transform 1 0 61344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_640
timestamp 1679581782
transform 1 0 62016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_647
timestamp 1679581782
transform 1 0 62688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_654
timestamp 1679581782
transform 1 0 63360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_661
timestamp 1679581782
transform 1 0 64032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_668
timestamp 1679581782
transform 1 0 64704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_675
timestamp 1679581782
transform 1 0 65376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_682
timestamp 1679581782
transform 1 0 66048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_689
timestamp 1679581782
transform 1 0 66720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_696
timestamp 1679581782
transform 1 0 67392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_703
timestamp 1679581782
transform 1 0 68064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_710
timestamp 1679581782
transform 1 0 68736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_717
timestamp 1679581782
transform 1 0 69408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_724
timestamp 1679581782
transform 1 0 70080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_731
timestamp 1679581782
transform 1 0 70752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_738
timestamp 1679581782
transform 1 0 71424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_745
timestamp 1679581782
transform 1 0 72096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_752
timestamp 1679581782
transform 1 0 72768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_759
timestamp 1679581782
transform 1 0 73440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_766
timestamp 1679581782
transform 1 0 74112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_773
timestamp 1679581782
transform 1 0 74784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_780
timestamp 1679581782
transform 1 0 75456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_787
timestamp 1679581782
transform 1 0 76128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_794
timestamp 1679581782
transform 1 0 76800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_801
timestamp 1679581782
transform 1 0 77472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_808
timestamp 1679581782
transform 1 0 78144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_815
timestamp 1679581782
transform 1 0 78816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_822
timestamp 1679581782
transform 1 0 79488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_829
timestamp 1679581782
transform 1 0 80160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_836
timestamp 1679581782
transform 1 0 80832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_843
timestamp 1679581782
transform 1 0 81504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_850
timestamp 1679581782
transform 1 0 82176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_857
timestamp 1679581782
transform 1 0 82848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_864
timestamp 1679581782
transform 1 0 83520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_871
timestamp 1679581782
transform 1 0 84192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_878
timestamp 1679581782
transform 1 0 84864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_885
timestamp 1679581782
transform 1 0 85536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_892
timestamp 1679581782
transform 1 0 86208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_899
timestamp 1679581782
transform 1 0 86880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_906
timestamp 1679581782
transform 1 0 87552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_913
timestamp 1679581782
transform 1 0 88224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_920
timestamp 1679581782
transform 1 0 88896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_927
timestamp 1679581782
transform 1 0 89568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_934
timestamp 1679581782
transform 1 0 90240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_941
timestamp 1679581782
transform 1 0 90912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_948
timestamp 1679581782
transform 1 0 91584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_955
timestamp 1679581782
transform 1 0 92256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_962
timestamp 1679581782
transform 1 0 92928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_969
timestamp 1679581782
transform 1 0 93600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_976
timestamp 1679581782
transform 1 0 94272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_983
timestamp 1679581782
transform 1 0 94944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_990
timestamp 1679581782
transform 1 0 95616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_997
timestamp 1679581782
transform 1 0 96288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1004
timestamp 1679581782
transform 1 0 96960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1011
timestamp 1679581782
transform 1 0 97632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1018
timestamp 1679581782
transform 1 0 98304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_1025
timestamp 1679577901
transform 1 0 98976 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_4
timestamp 1677580104
transform 1 0 960 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_6
timestamp 1677579658
transform 1 0 1152 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_32
timestamp 1677579658
transform 1 0 3648 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_59
timestamp 1679581782
transform 1 0 6240 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_77
timestamp 1677580104
transform 1 0 7968 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_79
timestamp 1677579658
transform 1 0 8160 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_127
timestamp 1679581782
transform 1 0 12768 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_134
timestamp 1677579658
transform 1 0 13440 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_162
timestamp 1677580104
transform 1 0 16128 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679581782
transform 1 0 19392 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_203
timestamp 1677580104
transform 1 0 20064 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_214
timestamp 1679577901
transform 1 0 21120 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_218
timestamp 1677579658
transform 1 0 21504 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_233
timestamp 1677580104
transform 1 0 22944 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_261
timestamp 1679581782
transform 1 0 25632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_268
timestamp 1679577901
transform 1 0 26304 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_272
timestamp 1677580104
transform 1 0 26688 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_293
timestamp 1679577901
transform 1 0 28704 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_297
timestamp 1677579658
transform 1 0 29088 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_317
timestamp 1677580104
transform 1 0 31008 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_338
timestamp 1679581782
transform 1 0 33024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_345
timestamp 1679577901
transform 1 0 33696 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_354
timestamp 1677580104
transform 1 0 34560 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_372
timestamp 1679581782
transform 1 0 36288 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_379
timestamp 1677580104
transform 1 0 36960 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_381
timestamp 1677579658
transform 1 0 37152 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_385
timestamp 1679577901
transform 1 0 37536 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_389
timestamp 1677580104
transform 1 0 37920 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679581782
transform 1 0 48960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679581782
transform 1 0 49632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_518
timestamp 1679581782
transform 1 0 50304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_525
timestamp 1679581782
transform 1 0 50976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_532
timestamp 1679581782
transform 1 0 51648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_539
timestamp 1679581782
transform 1 0 52320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_546
timestamp 1679581782
transform 1 0 52992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_553
timestamp 1679581782
transform 1 0 53664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_560
timestamp 1679581782
transform 1 0 54336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_567
timestamp 1679581782
transform 1 0 55008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_574
timestamp 1679581782
transform 1 0 55680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_581
timestamp 1679581782
transform 1 0 56352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_588
timestamp 1679581782
transform 1 0 57024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_595
timestamp 1679581782
transform 1 0 57696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_602
timestamp 1679581782
transform 1 0 58368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_609
timestamp 1679581782
transform 1 0 59040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_616
timestamp 1679581782
transform 1 0 59712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679581782
transform 1 0 60384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_630
timestamp 1679581782
transform 1 0 61056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_637
timestamp 1679581782
transform 1 0 61728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_644
timestamp 1679581782
transform 1 0 62400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_651
timestamp 1679581782
transform 1 0 63072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_658
timestamp 1679581782
transform 1 0 63744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_665
timestamp 1679581782
transform 1 0 64416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_672
timestamp 1679581782
transform 1 0 65088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_679
timestamp 1679581782
transform 1 0 65760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_686
timestamp 1679581782
transform 1 0 66432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_693
timestamp 1679581782
transform 1 0 67104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_700
timestamp 1679581782
transform 1 0 67776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_707
timestamp 1679581782
transform 1 0 68448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_714
timestamp 1679581782
transform 1 0 69120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_721
timestamp 1679581782
transform 1 0 69792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_728
timestamp 1679581782
transform 1 0 70464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_735
timestamp 1679581782
transform 1 0 71136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_742
timestamp 1679581782
transform 1 0 71808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679581782
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679581782
transform 1 0 73152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_763
timestamp 1679581782
transform 1 0 73824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_770
timestamp 1679581782
transform 1 0 74496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_777
timestamp 1679581782
transform 1 0 75168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_784
timestamp 1679581782
transform 1 0 75840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_791
timestamp 1679581782
transform 1 0 76512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_798
timestamp 1679581782
transform 1 0 77184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_805
timestamp 1679581782
transform 1 0 77856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_812
timestamp 1679581782
transform 1 0 78528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_819
timestamp 1679581782
transform 1 0 79200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_826
timestamp 1679581782
transform 1 0 79872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_833
timestamp 1679581782
transform 1 0 80544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_840
timestamp 1679581782
transform 1 0 81216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_847
timestamp 1679581782
transform 1 0 81888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_854
timestamp 1679581782
transform 1 0 82560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_861
timestamp 1679581782
transform 1 0 83232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_868
timestamp 1679581782
transform 1 0 83904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_875
timestamp 1679581782
transform 1 0 84576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_882
timestamp 1679581782
transform 1 0 85248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_889
timestamp 1679581782
transform 1 0 85920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_896
timestamp 1679581782
transform 1 0 86592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_903
timestamp 1679581782
transform 1 0 87264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_910
timestamp 1679581782
transform 1 0 87936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_917
timestamp 1679581782
transform 1 0 88608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_924
timestamp 1679581782
transform 1 0 89280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_931
timestamp 1679581782
transform 1 0 89952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_938
timestamp 1679581782
transform 1 0 90624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_945
timestamp 1679581782
transform 1 0 91296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_952
timestamp 1679581782
transform 1 0 91968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_959
timestamp 1679581782
transform 1 0 92640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_966
timestamp 1679581782
transform 1 0 93312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_973
timestamp 1679581782
transform 1 0 93984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_980
timestamp 1679581782
transform 1 0 94656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_987
timestamp 1679581782
transform 1 0 95328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_994
timestamp 1679581782
transform 1 0 96000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1001
timestamp 1679581782
transform 1 0 96672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1008
timestamp 1679581782
transform 1 0 97344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1015
timestamp 1679581782
transform 1 0 98016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1022
timestamp 1679581782
transform 1 0 98688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_4
timestamp 1679577901
transform 1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_8
timestamp 1677579658
transform 1 0 1344 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_74
timestamp 1679577901
transform 1 0 7680 0 1 9828
box -48 -56 432 834
use sg13g2_decap_4  FILLER_12_84
timestamp 1679577901
transform 1 0 8640 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_116
timestamp 1677580104
transform 1 0 11712 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_135
timestamp 1679577901
transform 1 0 13536 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_139
timestamp 1677579658
transform 1 0 13920 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679581782
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_151
timestamp 1677580104
transform 1 0 15072 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_175
timestamp 1677580104
transform 1 0 17376 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_177
timestamp 1677579658
transform 1 0 17568 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_200
timestamp 1679577901
transform 1 0 19776 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_228
timestamp 1677580104
transform 1 0 22464 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_251
timestamp 1677579658
transform 1 0 24672 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_262
timestamp 1679577901
transform 1 0 25728 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_266
timestamp 1677579658
transform 1 0 26112 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_277
timestamp 1679577901
transform 1 0 27168 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_281
timestamp 1677579658
transform 1 0 27552 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_290
timestamp 1679581782
transform 1 0 28416 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_297
timestamp 1677579658
transform 1 0 29088 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_306
timestamp 1677579658
transform 1 0 29952 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_316
timestamp 1679577901
transform 1 0 30912 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_345
timestamp 1677579658
transform 1 0 33696 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_439
timestamp 1677579658
transform 1 0 42720 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_510
timestamp 1679581782
transform 1 0 49536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_517
timestamp 1679581782
transform 1 0 50208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_524
timestamp 1679581782
transform 1 0 50880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_531
timestamp 1679581782
transform 1 0 51552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_538
timestamp 1679581782
transform 1 0 52224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_545
timestamp 1679581782
transform 1 0 52896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_552
timestamp 1679581782
transform 1 0 53568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_559
timestamp 1679581782
transform 1 0 54240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_566
timestamp 1679581782
transform 1 0 54912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_573
timestamp 1679581782
transform 1 0 55584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_580
timestamp 1679581782
transform 1 0 56256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_587
timestamp 1679581782
transform 1 0 56928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_594
timestamp 1679581782
transform 1 0 57600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_601
timestamp 1679581782
transform 1 0 58272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_608
timestamp 1679581782
transform 1 0 58944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_615
timestamp 1679581782
transform 1 0 59616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_622
timestamp 1679581782
transform 1 0 60288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_629
timestamp 1679581782
transform 1 0 60960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_636
timestamp 1679581782
transform 1 0 61632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_643
timestamp 1679581782
transform 1 0 62304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_650
timestamp 1679581782
transform 1 0 62976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_657
timestamp 1679581782
transform 1 0 63648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_664
timestamp 1679581782
transform 1 0 64320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_671
timestamp 1679581782
transform 1 0 64992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_678
timestamp 1679581782
transform 1 0 65664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_685
timestamp 1679581782
transform 1 0 66336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_692
timestamp 1679581782
transform 1 0 67008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_699
timestamp 1679581782
transform 1 0 67680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_706
timestamp 1679581782
transform 1 0 68352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_713
timestamp 1679581782
transform 1 0 69024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_720
timestamp 1679581782
transform 1 0 69696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_727
timestamp 1679581782
transform 1 0 70368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_734
timestamp 1679581782
transform 1 0 71040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_741
timestamp 1679581782
transform 1 0 71712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_748
timestamp 1679581782
transform 1 0 72384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_755
timestamp 1679581782
transform 1 0 73056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_762
timestamp 1679581782
transform 1 0 73728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_769
timestamp 1679581782
transform 1 0 74400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_776
timestamp 1679581782
transform 1 0 75072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_783
timestamp 1679581782
transform 1 0 75744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_790
timestamp 1679581782
transform 1 0 76416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_797
timestamp 1679581782
transform 1 0 77088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_804
timestamp 1679581782
transform 1 0 77760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_811
timestamp 1679581782
transform 1 0 78432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_818
timestamp 1679581782
transform 1 0 79104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_825
timestamp 1679581782
transform 1 0 79776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_832
timestamp 1679581782
transform 1 0 80448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_839
timestamp 1679581782
transform 1 0 81120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_846
timestamp 1679581782
transform 1 0 81792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_853
timestamp 1679581782
transform 1 0 82464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_860
timestamp 1679581782
transform 1 0 83136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_867
timestamp 1679581782
transform 1 0 83808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_874
timestamp 1679581782
transform 1 0 84480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_881
timestamp 1679581782
transform 1 0 85152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_888
timestamp 1679581782
transform 1 0 85824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_895
timestamp 1679581782
transform 1 0 86496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_902
timestamp 1679581782
transform 1 0 87168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_909
timestamp 1679581782
transform 1 0 87840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_916
timestamp 1679581782
transform 1 0 88512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_923
timestamp 1679581782
transform 1 0 89184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_930
timestamp 1679581782
transform 1 0 89856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_937
timestamp 1679581782
transform 1 0 90528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_944
timestamp 1679581782
transform 1 0 91200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_951
timestamp 1679581782
transform 1 0 91872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_958
timestamp 1679581782
transform 1 0 92544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_965
timestamp 1679581782
transform 1 0 93216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_972
timestamp 1679581782
transform 1 0 93888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_979
timestamp 1679581782
transform 1 0 94560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_986
timestamp 1679581782
transform 1 0 95232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_993
timestamp 1679581782
transform 1 0 95904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1000
timestamp 1679581782
transform 1 0 96576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1007
timestamp 1679581782
transform 1 0 97248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1014
timestamp 1679581782
transform 1 0 97920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1021
timestamp 1679581782
transform 1 0 98592 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_1028
timestamp 1677579658
transform 1 0 99264 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_11
timestamp 1677580104
transform 1 0 1632 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_13
timestamp 1677579658
transform 1 0 1824 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_18
timestamp 1677580104
transform 1 0 2304 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_25
timestamp 1679577901
transform 1 0 2976 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_68
timestamp 1679577901
transform 1 0 7104 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_72
timestamp 1677579658
transform 1 0 7488 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_101
timestamp 1679581782
transform 1 0 10272 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_108
timestamp 1677580104
transform 1 0 10944 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_110
timestamp 1677579658
transform 1 0 11136 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_165
timestamp 1677580104
transform 1 0 16416 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_167
timestamp 1677579658
transform 1 0 16608 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_201
timestamp 1679577901
transform 1 0 19872 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_205
timestamp 1677580104
transform 1 0 20256 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_213
timestamp 1679581782
transform 1 0 21024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_220
timestamp 1679581782
transform 1 0 21696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_227
timestamp 1679581782
transform 1 0 22368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_234
timestamp 1679577901
transform 1 0 23040 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_238
timestamp 1677579658
transform 1 0 23424 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_249
timestamp 1677580104
transform 1 0 24480 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_257
timestamp 1679581782
transform 1 0 25248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_264
timestamp 1679581782
transform 1 0 25920 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_271
timestamp 1677580104
transform 1 0 26592 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_273
timestamp 1677579658
transform 1 0 26784 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_288
timestamp 1679577901
transform 1 0 28224 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_292
timestamp 1677580104
transform 1 0 28608 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_317
timestamp 1679577901
transform 1 0 31008 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_343
timestamp 1679581782
transform 1 0 33504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_350
timestamp 1679581782
transform 1 0 34176 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_362
timestamp 1677579658
transform 1 0 35328 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_368
timestamp 1677580104
transform 1 0 35904 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_472
timestamp 1677579658
transform 1 0 45888 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_486
timestamp 1677579658
transform 1 0 47232 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_507
timestamp 1679581782
transform 1 0 49248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_514
timestamp 1679581782
transform 1 0 49920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_521
timestamp 1679581782
transform 1 0 50592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_528
timestamp 1679581782
transform 1 0 51264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_535
timestamp 1679581782
transform 1 0 51936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_542
timestamp 1679581782
transform 1 0 52608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_549
timestamp 1679581782
transform 1 0 53280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_556
timestamp 1679581782
transform 1 0 53952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_563
timestamp 1679581782
transform 1 0 54624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_570
timestamp 1679581782
transform 1 0 55296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_577
timestamp 1679581782
transform 1 0 55968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_584
timestamp 1679581782
transform 1 0 56640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_591
timestamp 1679581782
transform 1 0 57312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_598
timestamp 1679581782
transform 1 0 57984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_605
timestamp 1679581782
transform 1 0 58656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_612
timestamp 1679581782
transform 1 0 59328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_619
timestamp 1679581782
transform 1 0 60000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_626
timestamp 1679581782
transform 1 0 60672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_633
timestamp 1679581782
transform 1 0 61344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_640
timestamp 1679581782
transform 1 0 62016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_647
timestamp 1679581782
transform 1 0 62688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_654
timestamp 1679581782
transform 1 0 63360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_661
timestamp 1679581782
transform 1 0 64032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_668
timestamp 1679581782
transform 1 0 64704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_675
timestamp 1679581782
transform 1 0 65376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_682
timestamp 1679581782
transform 1 0 66048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_689
timestamp 1679581782
transform 1 0 66720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_696
timestamp 1679581782
transform 1 0 67392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_703
timestamp 1679581782
transform 1 0 68064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_710
timestamp 1679581782
transform 1 0 68736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_717
timestamp 1679581782
transform 1 0 69408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_724
timestamp 1679581782
transform 1 0 70080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_731
timestamp 1679581782
transform 1 0 70752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_738
timestamp 1679581782
transform 1 0 71424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_745
timestamp 1679581782
transform 1 0 72096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_752
timestamp 1679581782
transform 1 0 72768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_759
timestamp 1679581782
transform 1 0 73440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_766
timestamp 1679581782
transform 1 0 74112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_773
timestamp 1679581782
transform 1 0 74784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_780
timestamp 1679581782
transform 1 0 75456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_787
timestamp 1679581782
transform 1 0 76128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_794
timestamp 1679581782
transform 1 0 76800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_801
timestamp 1679581782
transform 1 0 77472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_808
timestamp 1679581782
transform 1 0 78144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_815
timestamp 1679581782
transform 1 0 78816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_822
timestamp 1679581782
transform 1 0 79488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_829
timestamp 1679581782
transform 1 0 80160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_836
timestamp 1679581782
transform 1 0 80832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_843
timestamp 1679581782
transform 1 0 81504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_850
timestamp 1679581782
transform 1 0 82176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_857
timestamp 1679581782
transform 1 0 82848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_864
timestamp 1679581782
transform 1 0 83520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_871
timestamp 1679581782
transform 1 0 84192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_878
timestamp 1679581782
transform 1 0 84864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_885
timestamp 1679581782
transform 1 0 85536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_892
timestamp 1679581782
transform 1 0 86208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_899
timestamp 1679581782
transform 1 0 86880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_906
timestamp 1679581782
transform 1 0 87552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_913
timestamp 1679581782
transform 1 0 88224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_920
timestamp 1679581782
transform 1 0 88896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_927
timestamp 1679581782
transform 1 0 89568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_934
timestamp 1679581782
transform 1 0 90240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_941
timestamp 1679581782
transform 1 0 90912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_948
timestamp 1679581782
transform 1 0 91584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_955
timestamp 1679581782
transform 1 0 92256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_962
timestamp 1679581782
transform 1 0 92928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_969
timestamp 1679581782
transform 1 0 93600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_976
timestamp 1679581782
transform 1 0 94272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_983
timestamp 1679581782
transform 1 0 94944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_990
timestamp 1679581782
transform 1 0 95616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_997
timestamp 1679581782
transform 1 0 96288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1004
timestamp 1679581782
transform 1 0 96960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1011
timestamp 1679581782
transform 1 0 97632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1018
timestamp 1679581782
transform 1 0 98304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_1025
timestamp 1679577901
transform 1 0 98976 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_65
timestamp 1679581782
transform 1 0 6816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_72
timestamp 1679577901
transform 1 0 7488 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_101
timestamp 1679581782
transform 1 0 10272 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_108
timestamp 1677580104
transform 1 0 10944 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_153
timestamp 1679581782
transform 1 0 15264 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_180
timestamp 1677580104
transform 1 0 17856 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_187
timestamp 1677580104
transform 1 0 18528 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_195
timestamp 1679577901
transform 1 0 19296 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_212
timestamp 1677579658
transform 1 0 20928 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_221
timestamp 1679581782
transform 1 0 21792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_228
timestamp 1679581782
transform 1 0 22464 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_235
timestamp 1677580104
transform 1 0 23136 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_237
timestamp 1677579658
transform 1 0 23328 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_255
timestamp 1679581782
transform 1 0 25056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_262
timestamp 1679577901
transform 1 0 25728 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_266
timestamp 1677579658
transform 1 0 26112 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_292
timestamp 1677580104
transform 1 0 28608 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_299
timestamp 1679581782
transform 1 0 29280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_306
timestamp 1679581782
transform 1 0 29952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_313
timestamp 1679581782
transform 1 0 30624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_339
timestamp 1679577901
transform 1 0 33120 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_343
timestamp 1677579658
transform 1 0 33504 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_359
timestamp 1677579658
transform 1 0 35040 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_363
timestamp 1679581782
transform 1 0 35424 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_373
timestamp 1677579658
transform 1 0 36384 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_398
timestamp 1679577901
transform 1 0 38784 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_409
timestamp 1677580104
transform 1 0 39840 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_462
timestamp 1677579658
transform 1 0 44928 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_472
timestamp 1677580104
transform 1 0 45888 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_510
timestamp 1679581782
transform 1 0 49536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_517
timestamp 1679581782
transform 1 0 50208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_524
timestamp 1679581782
transform 1 0 50880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_531
timestamp 1679581782
transform 1 0 51552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_538
timestamp 1679581782
transform 1 0 52224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_545
timestamp 1679581782
transform 1 0 52896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_552
timestamp 1679581782
transform 1 0 53568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_559
timestamp 1679581782
transform 1 0 54240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_566
timestamp 1679581782
transform 1 0 54912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_573
timestamp 1679581782
transform 1 0 55584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_580
timestamp 1679581782
transform 1 0 56256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_587
timestamp 1679581782
transform 1 0 56928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_594
timestamp 1679581782
transform 1 0 57600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_601
timestamp 1679581782
transform 1 0 58272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_608
timestamp 1679581782
transform 1 0 58944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_615
timestamp 1679581782
transform 1 0 59616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_622
timestamp 1679581782
transform 1 0 60288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_629
timestamp 1679581782
transform 1 0 60960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_636
timestamp 1679581782
transform 1 0 61632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_643
timestamp 1679581782
transform 1 0 62304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_650
timestamp 1679581782
transform 1 0 62976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_657
timestamp 1679581782
transform 1 0 63648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_664
timestamp 1679581782
transform 1 0 64320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_671
timestamp 1679581782
transform 1 0 64992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_678
timestamp 1679581782
transform 1 0 65664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_685
timestamp 1679581782
transform 1 0 66336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_692
timestamp 1679581782
transform 1 0 67008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_699
timestamp 1679581782
transform 1 0 67680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_706
timestamp 1679581782
transform 1 0 68352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_713
timestamp 1679581782
transform 1 0 69024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_720
timestamp 1679581782
transform 1 0 69696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_727
timestamp 1679581782
transform 1 0 70368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_734
timestamp 1679581782
transform 1 0 71040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_741
timestamp 1679581782
transform 1 0 71712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_748
timestamp 1679581782
transform 1 0 72384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_755
timestamp 1679581782
transform 1 0 73056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_762
timestamp 1679581782
transform 1 0 73728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_769
timestamp 1679581782
transform 1 0 74400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_776
timestamp 1679581782
transform 1 0 75072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_783
timestamp 1679581782
transform 1 0 75744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_790
timestamp 1679581782
transform 1 0 76416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_797
timestamp 1679581782
transform 1 0 77088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_804
timestamp 1679581782
transform 1 0 77760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_811
timestamp 1679581782
transform 1 0 78432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_818
timestamp 1679581782
transform 1 0 79104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_825
timestamp 1679581782
transform 1 0 79776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_832
timestamp 1679581782
transform 1 0 80448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_839
timestamp 1679581782
transform 1 0 81120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_846
timestamp 1679581782
transform 1 0 81792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_853
timestamp 1679581782
transform 1 0 82464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_860
timestamp 1679581782
transform 1 0 83136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_867
timestamp 1679581782
transform 1 0 83808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_874
timestamp 1679581782
transform 1 0 84480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_881
timestamp 1679581782
transform 1 0 85152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_888
timestamp 1679581782
transform 1 0 85824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_895
timestamp 1679581782
transform 1 0 86496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_902
timestamp 1679581782
transform 1 0 87168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_909
timestamp 1679581782
transform 1 0 87840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_916
timestamp 1679581782
transform 1 0 88512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_923
timestamp 1679581782
transform 1 0 89184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_930
timestamp 1679581782
transform 1 0 89856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_937
timestamp 1679581782
transform 1 0 90528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_944
timestamp 1679581782
transform 1 0 91200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_951
timestamp 1679581782
transform 1 0 91872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_958
timestamp 1679581782
transform 1 0 92544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_965
timestamp 1679581782
transform 1 0 93216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_972
timestamp 1679581782
transform 1 0 93888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_979
timestamp 1679581782
transform 1 0 94560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_986
timestamp 1679581782
transform 1 0 95232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_993
timestamp 1679581782
transform 1 0 95904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1000
timestamp 1679581782
transform 1 0 96576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1007
timestamp 1679581782
transform 1 0 97248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1014
timestamp 1679581782
transform 1 0 97920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1021
timestamp 1679581782
transform 1 0 98592 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_1028
timestamp 1677579658
transform 1 0 99264 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_18
timestamp 1679577901
transform 1 0 2304 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_22
timestamp 1677580104
transform 1 0 2688 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_80
timestamp 1677580104
transform 1 0 8256 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_108
timestamp 1677579658
transform 1 0 10944 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_127
timestamp 1677579658
transform 1 0 12768 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_137
timestamp 1677580104
transform 1 0 13728 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_152
timestamp 1679581782
transform 1 0 15168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_159
timestamp 1679581782
transform 1 0 15840 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_191
timestamp 1677580104
transform 1 0 18912 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_199
timestamp 1677580104
transform 1 0 19680 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_232
timestamp 1679581782
transform 1 0 22848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_239
timestamp 1679581782
transform 1 0 23520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_246
timestamp 1679581782
transform 1 0 24192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_253
timestamp 1679577901
transform 1 0 24864 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_15_270
timestamp 1679577901
transform 1 0 26496 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_282
timestamp 1677579658
transform 1 0 27648 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_302
timestamp 1679581782
transform 1 0 29568 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_309
timestamp 1677579658
transform 1 0 30240 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_334
timestamp 1679581782
transform 1 0 32640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_341
timestamp 1679581782
transform 1 0 33312 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_359
timestamp 1677580104
transform 1 0 35040 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_366
timestamp 1679581782
transform 1 0 35712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_373
timestamp 1679577901
transform 1 0 36384 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_377
timestamp 1677580104
transform 1 0 36768 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_426
timestamp 1677580104
transform 1 0 41472 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_428
timestamp 1677579658
transform 1 0 41664 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_480
timestamp 1677580104
transform 1 0 46656 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_491
timestamp 1677580104
transform 1 0 47712 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_502
timestamp 1679581782
transform 1 0 48768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_509
timestamp 1679581782
transform 1 0 49440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_516
timestamp 1679581782
transform 1 0 50112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_523
timestamp 1679581782
transform 1 0 50784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_530
timestamp 1679581782
transform 1 0 51456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_537
timestamp 1679581782
transform 1 0 52128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_544
timestamp 1679581782
transform 1 0 52800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_551
timestamp 1679581782
transform 1 0 53472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_558
timestamp 1679581782
transform 1 0 54144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_565
timestamp 1679581782
transform 1 0 54816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_572
timestamp 1679581782
transform 1 0 55488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_579
timestamp 1679581782
transform 1 0 56160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_586
timestamp 1679581782
transform 1 0 56832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_593
timestamp 1679581782
transform 1 0 57504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_600
timestamp 1679581782
transform 1 0 58176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_607
timestamp 1679581782
transform 1 0 58848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_614
timestamp 1679581782
transform 1 0 59520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_621
timestamp 1679581782
transform 1 0 60192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_628
timestamp 1679581782
transform 1 0 60864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_635
timestamp 1679581782
transform 1 0 61536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_642
timestamp 1679581782
transform 1 0 62208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_649
timestamp 1679581782
transform 1 0 62880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_656
timestamp 1679581782
transform 1 0 63552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_663
timestamp 1679581782
transform 1 0 64224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_670
timestamp 1679581782
transform 1 0 64896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_677
timestamp 1679581782
transform 1 0 65568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_684
timestamp 1679581782
transform 1 0 66240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_691
timestamp 1679581782
transform 1 0 66912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_698
timestamp 1679581782
transform 1 0 67584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_705
timestamp 1679581782
transform 1 0 68256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_712
timestamp 1679581782
transform 1 0 68928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_719
timestamp 1679581782
transform 1 0 69600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_726
timestamp 1679581782
transform 1 0 70272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_733
timestamp 1679581782
transform 1 0 70944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_740
timestamp 1679581782
transform 1 0 71616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_747
timestamp 1679581782
transform 1 0 72288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_754
timestamp 1679581782
transform 1 0 72960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_761
timestamp 1679581782
transform 1 0 73632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_768
timestamp 1679581782
transform 1 0 74304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_775
timestamp 1679581782
transform 1 0 74976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_782
timestamp 1679581782
transform 1 0 75648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_789
timestamp 1679581782
transform 1 0 76320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_796
timestamp 1679581782
transform 1 0 76992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_803
timestamp 1679581782
transform 1 0 77664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_810
timestamp 1679581782
transform 1 0 78336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_817
timestamp 1679581782
transform 1 0 79008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_824
timestamp 1679581782
transform 1 0 79680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_831
timestamp 1679581782
transform 1 0 80352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_838
timestamp 1679581782
transform 1 0 81024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_845
timestamp 1679581782
transform 1 0 81696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_852
timestamp 1679581782
transform 1 0 82368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_859
timestamp 1679581782
transform 1 0 83040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_866
timestamp 1679581782
transform 1 0 83712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_873
timestamp 1679581782
transform 1 0 84384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_880
timestamp 1679581782
transform 1 0 85056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_887
timestamp 1679581782
transform 1 0 85728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_894
timestamp 1679581782
transform 1 0 86400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_901
timestamp 1679581782
transform 1 0 87072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_908
timestamp 1679581782
transform 1 0 87744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_915
timestamp 1679581782
transform 1 0 88416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_922
timestamp 1679581782
transform 1 0 89088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_929
timestamp 1679581782
transform 1 0 89760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_936
timestamp 1679581782
transform 1 0 90432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_943
timestamp 1679581782
transform 1 0 91104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_950
timestamp 1679581782
transform 1 0 91776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_957
timestamp 1679581782
transform 1 0 92448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_964
timestamp 1679581782
transform 1 0 93120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_971
timestamp 1679581782
transform 1 0 93792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_978
timestamp 1679581782
transform 1 0 94464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_985
timestamp 1679581782
transform 1 0 95136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_992
timestamp 1679581782
transform 1 0 95808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_999
timestamp 1679581782
transform 1 0 96480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1006
timestamp 1679581782
transform 1 0 97152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1013
timestamp 1679581782
transform 1 0 97824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1020
timestamp 1679581782
transform 1 0 98496 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_1027
timestamp 1677580104
transform 1 0 99168 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679581782
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_18
timestamp 1679581782
transform 1 0 2304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_25
timestamp 1679577901
transform 1 0 2976 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_114
timestamp 1677580104
transform 1 0 11520 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_116
timestamp 1677579658
transform 1 0 11712 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_127
timestamp 1677579658
transform 1 0 12768 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_164
timestamp 1679581782
transform 1 0 16320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_171
timestamp 1679577901
transform 1 0 16992 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_175
timestamp 1677580104
transform 1 0 17376 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_183
timestamp 1677579658
transform 1 0 18144 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_204
timestamp 1677579658
transform 1 0 20160 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_222
timestamp 1677580104
transform 1 0 21888 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_224
timestamp 1677579658
transform 1 0 22080 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_234
timestamp 1677580104
transform 1 0 23040 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_240
timestamp 1679581782
transform 1 0 23616 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_247
timestamp 1677580104
transform 1 0 24288 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_277
timestamp 1679577901
transform 1 0 27168 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_281
timestamp 1677579658
transform 1 0 27552 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_294
timestamp 1677580104
transform 1 0 28800 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_317
timestamp 1679577901
transform 1 0 31008 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_321
timestamp 1677579658
transform 1 0 31392 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_326
timestamp 1677579658
transform 1 0 31872 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_333
timestamp 1677580104
transform 1 0 32544 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_339
timestamp 1679577901
transform 1 0 33120 0 1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_16_353
timestamp 1679577901
transform 1 0 34464 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_375
timestamp 1679581782
transform 1 0 36576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_489
timestamp 1679581782
transform 1 0 47520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_496
timestamp 1679581782
transform 1 0 48192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_503
timestamp 1679581782
transform 1 0 48864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_510
timestamp 1679581782
transform 1 0 49536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_517
timestamp 1679581782
transform 1 0 50208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_524
timestamp 1679581782
transform 1 0 50880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_531
timestamp 1679581782
transform 1 0 51552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_538
timestamp 1679581782
transform 1 0 52224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_545
timestamp 1679581782
transform 1 0 52896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_552
timestamp 1679581782
transform 1 0 53568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_559
timestamp 1679581782
transform 1 0 54240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_566
timestamp 1679581782
transform 1 0 54912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_573
timestamp 1679581782
transform 1 0 55584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_580
timestamp 1679581782
transform 1 0 56256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_587
timestamp 1679581782
transform 1 0 56928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_594
timestamp 1679581782
transform 1 0 57600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_601
timestamp 1679581782
transform 1 0 58272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_608
timestamp 1679581782
transform 1 0 58944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_615
timestamp 1679581782
transform 1 0 59616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_622
timestamp 1679581782
transform 1 0 60288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_629
timestamp 1679581782
transform 1 0 60960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_636
timestamp 1679581782
transform 1 0 61632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_643
timestamp 1679581782
transform 1 0 62304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_650
timestamp 1679581782
transform 1 0 62976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_657
timestamp 1679581782
transform 1 0 63648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_664
timestamp 1679581782
transform 1 0 64320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_671
timestamp 1679581782
transform 1 0 64992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_678
timestamp 1679581782
transform 1 0 65664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_685
timestamp 1679581782
transform 1 0 66336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_692
timestamp 1679581782
transform 1 0 67008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_699
timestamp 1679581782
transform 1 0 67680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_706
timestamp 1679581782
transform 1 0 68352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_713
timestamp 1679581782
transform 1 0 69024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_720
timestamp 1679581782
transform 1 0 69696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_727
timestamp 1679581782
transform 1 0 70368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_734
timestamp 1679581782
transform 1 0 71040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_741
timestamp 1679581782
transform 1 0 71712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_748
timestamp 1679581782
transform 1 0 72384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_755
timestamp 1679581782
transform 1 0 73056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_762
timestamp 1679581782
transform 1 0 73728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_769
timestamp 1679581782
transform 1 0 74400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_776
timestamp 1679581782
transform 1 0 75072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_783
timestamp 1679581782
transform 1 0 75744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_790
timestamp 1679581782
transform 1 0 76416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_797
timestamp 1679581782
transform 1 0 77088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_804
timestamp 1679581782
transform 1 0 77760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679581782
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_818
timestamp 1679581782
transform 1 0 79104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_825
timestamp 1679581782
transform 1 0 79776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_832
timestamp 1679581782
transform 1 0 80448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_839
timestamp 1679581782
transform 1 0 81120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_846
timestamp 1679581782
transform 1 0 81792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_853
timestamp 1679581782
transform 1 0 82464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_860
timestamp 1679581782
transform 1 0 83136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_867
timestamp 1679581782
transform 1 0 83808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_874
timestamp 1679581782
transform 1 0 84480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_881
timestamp 1679581782
transform 1 0 85152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_888
timestamp 1679581782
transform 1 0 85824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_895
timestamp 1679581782
transform 1 0 86496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_902
timestamp 1679581782
transform 1 0 87168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_909
timestamp 1679581782
transform 1 0 87840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_916
timestamp 1679581782
transform 1 0 88512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_923
timestamp 1679581782
transform 1 0 89184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_930
timestamp 1679581782
transform 1 0 89856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_937
timestamp 1679581782
transform 1 0 90528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_944
timestamp 1679581782
transform 1 0 91200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_951
timestamp 1679581782
transform 1 0 91872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_958
timestamp 1679581782
transform 1 0 92544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_965
timestamp 1679581782
transform 1 0 93216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_972
timestamp 1679581782
transform 1 0 93888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_979
timestamp 1679581782
transform 1 0 94560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_986
timestamp 1679581782
transform 1 0 95232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_993
timestamp 1679581782
transform 1 0 95904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1000
timestamp 1679581782
transform 1 0 96576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1007
timestamp 1679581782
transform 1 0 97248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1014
timestamp 1679581782
transform 1 0 97920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1021
timestamp 1679581782
transform 1 0 98592 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_1028
timestamp 1677579658
transform 1 0 99264 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_4
timestamp 1679581782
transform 1 0 960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_11
timestamp 1679581782
transform 1 0 1632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_18
timestamp 1679581782
transform 1 0 2304 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_25
timestamp 1677580104
transform 1 0 2976 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_40
timestamp 1677579658
transform 1 0 4416 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_65
timestamp 1677580104
transform 1 0 6816 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_80
timestamp 1677580104
transform 1 0 8256 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_82
timestamp 1677579658
transform 1 0 8448 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_87
timestamp 1679581782
transform 1 0 8928 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_94
timestamp 1677579658
transform 1 0 9600 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_122
timestamp 1677579658
transform 1 0 12288 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_132
timestamp 1679577901
transform 1 0 13248 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_153
timestamp 1677580104
transform 1 0 15264 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_155
timestamp 1677579658
transform 1 0 15456 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_161
timestamp 1679581782
transform 1 0 16032 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_168
timestamp 1677579658
transform 1 0 16704 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_180
timestamp 1677580104
transform 1 0 17856 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_195
timestamp 1677580104
transform 1 0 19296 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_207
timestamp 1677579658
transform 1 0 20448 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_236
timestamp 1679581782
transform 1 0 23232 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_243
timestamp 1677580104
transform 1 0 23904 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_258
timestamp 1677580104
transform 1 0 25344 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_273
timestamp 1677580104
transform 1 0 26784 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_275
timestamp 1677579658
transform 1 0 26976 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_286
timestamp 1677579658
transform 1 0 28032 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_292
timestamp 1679581782
transform 1 0 28608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_299
timestamp 1679581782
transform 1 0 29280 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_306
timestamp 1677580104
transform 1 0 29952 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_313
timestamp 1679581782
transform 1 0 30624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_320
timestamp 1679577901
transform 1 0 31296 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_17_351
timestamp 1679577901
transform 1 0 34272 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_355
timestamp 1677580104
transform 1 0 34656 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_400
timestamp 1679577901
transform 1 0 38976 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_404
timestamp 1677579658
transform 1 0 39360 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_409
timestamp 1679577901
transform 1 0 39840 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_413
timestamp 1677580104
transform 1 0 40224 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_433
timestamp 1677580104
transform 1 0 42144 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_435
timestamp 1677579658
transform 1 0 42336 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_449
timestamp 1679577901
transform 1 0 43680 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_481
timestamp 1679581782
transform 1 0 46752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_488
timestamp 1679581782
transform 1 0 47424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_495
timestamp 1679581782
transform 1 0 48096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_502
timestamp 1679581782
transform 1 0 48768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_509
timestamp 1679581782
transform 1 0 49440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_516
timestamp 1679581782
transform 1 0 50112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_523
timestamp 1679581782
transform 1 0 50784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_530
timestamp 1679581782
transform 1 0 51456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_537
timestamp 1679581782
transform 1 0 52128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_544
timestamp 1679581782
transform 1 0 52800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_551
timestamp 1679581782
transform 1 0 53472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_558
timestamp 1679581782
transform 1 0 54144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_565
timestamp 1679581782
transform 1 0 54816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_572
timestamp 1679581782
transform 1 0 55488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_579
timestamp 1679581782
transform 1 0 56160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_586
timestamp 1679581782
transform 1 0 56832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_593
timestamp 1679581782
transform 1 0 57504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_600
timestamp 1679581782
transform 1 0 58176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_607
timestamp 1679581782
transform 1 0 58848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_614
timestamp 1679581782
transform 1 0 59520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_621
timestamp 1679581782
transform 1 0 60192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_628
timestamp 1679581782
transform 1 0 60864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_635
timestamp 1679581782
transform 1 0 61536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_642
timestamp 1679581782
transform 1 0 62208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_649
timestamp 1679581782
transform 1 0 62880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_656
timestamp 1679581782
transform 1 0 63552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_663
timestamp 1679581782
transform 1 0 64224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_670
timestamp 1679581782
transform 1 0 64896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_677
timestamp 1679581782
transform 1 0 65568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_684
timestamp 1679581782
transform 1 0 66240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_691
timestamp 1679581782
transform 1 0 66912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_698
timestamp 1679581782
transform 1 0 67584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_705
timestamp 1679581782
transform 1 0 68256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_712
timestamp 1679581782
transform 1 0 68928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_719
timestamp 1679581782
transform 1 0 69600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_726
timestamp 1679581782
transform 1 0 70272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_733
timestamp 1679581782
transform 1 0 70944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_740
timestamp 1679581782
transform 1 0 71616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_747
timestamp 1679581782
transform 1 0 72288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_754
timestamp 1679581782
transform 1 0 72960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_761
timestamp 1679581782
transform 1 0 73632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_768
timestamp 1679581782
transform 1 0 74304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_775
timestamp 1679581782
transform 1 0 74976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_782
timestamp 1679581782
transform 1 0 75648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_789
timestamp 1679581782
transform 1 0 76320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_796
timestamp 1679581782
transform 1 0 76992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_803
timestamp 1679581782
transform 1 0 77664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_810
timestamp 1679581782
transform 1 0 78336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_817
timestamp 1679581782
transform 1 0 79008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_824
timestamp 1679581782
transform 1 0 79680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_831
timestamp 1679581782
transform 1 0 80352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_838
timestamp 1679581782
transform 1 0 81024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_845
timestamp 1679581782
transform 1 0 81696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_852
timestamp 1679581782
transform 1 0 82368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_859
timestamp 1679581782
transform 1 0 83040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_866
timestamp 1679581782
transform 1 0 83712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_873
timestamp 1679581782
transform 1 0 84384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_880
timestamp 1679581782
transform 1 0 85056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_887
timestamp 1679581782
transform 1 0 85728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_894
timestamp 1679581782
transform 1 0 86400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_901
timestamp 1679581782
transform 1 0 87072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_908
timestamp 1679581782
transform 1 0 87744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_915
timestamp 1679581782
transform 1 0 88416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_922
timestamp 1679581782
transform 1 0 89088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_929
timestamp 1679581782
transform 1 0 89760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_936
timestamp 1679581782
transform 1 0 90432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_943
timestamp 1679581782
transform 1 0 91104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_950
timestamp 1679581782
transform 1 0 91776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_957
timestamp 1679581782
transform 1 0 92448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_964
timestamp 1679581782
transform 1 0 93120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_971
timestamp 1679581782
transform 1 0 93792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_978
timestamp 1679581782
transform 1 0 94464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_985
timestamp 1679581782
transform 1 0 95136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_992
timestamp 1679581782
transform 1 0 95808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_999
timestamp 1679581782
transform 1 0 96480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1006
timestamp 1679581782
transform 1 0 97152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1013
timestamp 1679581782
transform 1 0 97824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1020
timestamp 1679581782
transform 1 0 98496 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_1027
timestamp 1677580104
transform 1 0 99168 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_8
timestamp 1677580104
transform 1 0 1344 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_10
timestamp 1677579658
transform 1 0 1536 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_15
timestamp 1677580104
transform 1 0 2016 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_17
timestamp 1677579658
transform 1 0 2208 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_45
timestamp 1677579658
transform 1 0 4896 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_90
timestamp 1679577901
transform 1 0 9216 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_151
timestamp 1677579658
transform 1 0 15072 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_160
timestamp 1677580104
transform 1 0 15936 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_196
timestamp 1677580104
transform 1 0 19392 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_198
timestamp 1677579658
transform 1 0 19584 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_204
timestamp 1677579658
transform 1 0 20160 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_220
timestamp 1677580104
transform 1 0 21696 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_222
timestamp 1677579658
transform 1 0 21888 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_229
timestamp 1679581782
transform 1 0 22560 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_236
timestamp 1677580104
transform 1 0 23232 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_254
timestamp 1677579658
transform 1 0 24960 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_270
timestamp 1677580104
transform 1 0 26496 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_307
timestamp 1679577901
transform 1 0 30048 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_311
timestamp 1677580104
transform 1 0 30432 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_358
timestamp 1679581782
transform 1 0 34944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_365
timestamp 1679581782
transform 1 0 35616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_372
timestamp 1679581782
transform 1 0 36288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_379
timestamp 1679577901
transform 1 0 36960 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_383
timestamp 1677579658
transform 1 0 37344 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_410
timestamp 1679581782
transform 1 0 39936 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_417
timestamp 1677580104
transform 1 0 40608 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_426
timestamp 1677580104
transform 1 0 41472 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_491
timestamp 1679581782
transform 1 0 47712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_498
timestamp 1679581782
transform 1 0 48384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_505
timestamp 1679581782
transform 1 0 49056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_512
timestamp 1679581782
transform 1 0 49728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_519
timestamp 1679581782
transform 1 0 50400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_526
timestamp 1679581782
transform 1 0 51072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_533
timestamp 1679581782
transform 1 0 51744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_540
timestamp 1679581782
transform 1 0 52416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_547
timestamp 1679581782
transform 1 0 53088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_554
timestamp 1679581782
transform 1 0 53760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_561
timestamp 1679581782
transform 1 0 54432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_568
timestamp 1679581782
transform 1 0 55104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_575
timestamp 1679581782
transform 1 0 55776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_582
timestamp 1679581782
transform 1 0 56448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_589
timestamp 1679581782
transform 1 0 57120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_596
timestamp 1679581782
transform 1 0 57792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_603
timestamp 1679581782
transform 1 0 58464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_610
timestamp 1679581782
transform 1 0 59136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_617
timestamp 1679581782
transform 1 0 59808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_624
timestamp 1679581782
transform 1 0 60480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_631
timestamp 1679581782
transform 1 0 61152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_638
timestamp 1679581782
transform 1 0 61824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_645
timestamp 1679581782
transform 1 0 62496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_652
timestamp 1679581782
transform 1 0 63168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_659
timestamp 1679581782
transform 1 0 63840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_666
timestamp 1679581782
transform 1 0 64512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_673
timestamp 1679581782
transform 1 0 65184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_680
timestamp 1679581782
transform 1 0 65856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_687
timestamp 1679581782
transform 1 0 66528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_694
timestamp 1679581782
transform 1 0 67200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_701
timestamp 1679581782
transform 1 0 67872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_708
timestamp 1679581782
transform 1 0 68544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_715
timestamp 1679581782
transform 1 0 69216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_722
timestamp 1679581782
transform 1 0 69888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_729
timestamp 1679581782
transform 1 0 70560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_736
timestamp 1679581782
transform 1 0 71232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_743
timestamp 1679581782
transform 1 0 71904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_750
timestamp 1679581782
transform 1 0 72576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_757
timestamp 1679581782
transform 1 0 73248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_764
timestamp 1679581782
transform 1 0 73920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_771
timestamp 1679581782
transform 1 0 74592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_778
timestamp 1679581782
transform 1 0 75264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_785
timestamp 1679581782
transform 1 0 75936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_792
timestamp 1679581782
transform 1 0 76608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_799
timestamp 1679581782
transform 1 0 77280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_806
timestamp 1679581782
transform 1 0 77952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_813
timestamp 1679581782
transform 1 0 78624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_820
timestamp 1679581782
transform 1 0 79296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_827
timestamp 1679581782
transform 1 0 79968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_834
timestamp 1679581782
transform 1 0 80640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_841
timestamp 1679581782
transform 1 0 81312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_848
timestamp 1679581782
transform 1 0 81984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_855
timestamp 1679581782
transform 1 0 82656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_862
timestamp 1679581782
transform 1 0 83328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_869
timestamp 1679581782
transform 1 0 84000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_876
timestamp 1679581782
transform 1 0 84672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_883
timestamp 1679581782
transform 1 0 85344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_890
timestamp 1679581782
transform 1 0 86016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_897
timestamp 1679581782
transform 1 0 86688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_904
timestamp 1679581782
transform 1 0 87360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_911
timestamp 1679581782
transform 1 0 88032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_918
timestamp 1679581782
transform 1 0 88704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_925
timestamp 1679581782
transform 1 0 89376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_932
timestamp 1679581782
transform 1 0 90048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_939
timestamp 1679581782
transform 1 0 90720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_946
timestamp 1679581782
transform 1 0 91392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_953
timestamp 1679581782
transform 1 0 92064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_960
timestamp 1679581782
transform 1 0 92736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_967
timestamp 1679581782
transform 1 0 93408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_974
timestamp 1679581782
transform 1 0 94080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_981
timestamp 1679581782
transform 1 0 94752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_988
timestamp 1679581782
transform 1 0 95424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_995
timestamp 1679581782
transform 1 0 96096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1002
timestamp 1679581782
transform 1 0 96768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1009
timestamp 1679581782
transform 1 0 97440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1016
timestamp 1679581782
transform 1 0 98112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_1023
timestamp 1679577901
transform 1 0 98784 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_1027
timestamp 1677580104
transform 1 0 99168 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_0
timestamp 1677579658
transform 1 0 576 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_46
timestamp 1677579658
transform 1 0 4992 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_103
timestamp 1679577901
transform 1 0 10464 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_107
timestamp 1677580104
transform 1 0 10848 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_122
timestamp 1677580104
transform 1 0 12288 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_127
timestamp 1677580104
transform 1 0 12768 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_129
timestamp 1677579658
transform 1 0 12960 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_167
timestamp 1677579658
transform 1 0 16608 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_181
timestamp 1679577901
transform 1 0 17952 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_213
timestamp 1679581782
transform 1 0 21024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_227
timestamp 1679581782
transform 1 0 22368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_234
timestamp 1679577901
transform 1 0 23040 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_238
timestamp 1677580104
transform 1 0 23424 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_244
timestamp 1677580104
transform 1 0 24000 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_259
timestamp 1679577901
transform 1 0 25440 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_263
timestamp 1677579658
transform 1 0 25824 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_285
timestamp 1679577901
transform 1 0 27936 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_300
timestamp 1677580104
transform 1 0 29376 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_326
timestamp 1679577901
transform 1 0 31872 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_335
timestamp 1677580104
transform 1 0 32736 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_337
timestamp 1677579658
transform 1 0 32928 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_395
timestamp 1679581782
transform 1 0 38496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_402
timestamp 1679577901
transform 1 0 39168 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_406
timestamp 1677579658
transform 1 0 39552 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_411
timestamp 1679581782
transform 1 0 40032 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_418
timestamp 1677580104
transform 1 0 40704 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_433
timestamp 1679581782
transform 1 0 42144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_440
timestamp 1679581782
transform 1 0 42816 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_447
timestamp 1677580104
transform 1 0 43488 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_449
timestamp 1677579658
transform 1 0 43680 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_463
timestamp 1679581782
transform 1 0 45024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_470
timestamp 1679581782
transform 1 0 45696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_477
timestamp 1679581782
transform 1 0 46368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_484
timestamp 1679581782
transform 1 0 47040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_491
timestamp 1679581782
transform 1 0 47712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_498
timestamp 1679581782
transform 1 0 48384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_505
timestamp 1679581782
transform 1 0 49056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_512
timestamp 1679581782
transform 1 0 49728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_519
timestamp 1679581782
transform 1 0 50400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_526
timestamp 1679581782
transform 1 0 51072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_533
timestamp 1679581782
transform 1 0 51744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_540
timestamp 1679581782
transform 1 0 52416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_547
timestamp 1679581782
transform 1 0 53088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_554
timestamp 1679581782
transform 1 0 53760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_561
timestamp 1679581782
transform 1 0 54432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_568
timestamp 1679581782
transform 1 0 55104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_575
timestamp 1679581782
transform 1 0 55776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_582
timestamp 1679581782
transform 1 0 56448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_589
timestamp 1679581782
transform 1 0 57120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_596
timestamp 1679581782
transform 1 0 57792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_603
timestamp 1679581782
transform 1 0 58464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_610
timestamp 1679581782
transform 1 0 59136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_617
timestamp 1679581782
transform 1 0 59808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_624
timestamp 1679581782
transform 1 0 60480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_631
timestamp 1679581782
transform 1 0 61152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_638
timestamp 1679581782
transform 1 0 61824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_645
timestamp 1679581782
transform 1 0 62496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_652
timestamp 1679581782
transform 1 0 63168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_659
timestamp 1679581782
transform 1 0 63840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_666
timestamp 1679581782
transform 1 0 64512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_673
timestamp 1679581782
transform 1 0 65184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_680
timestamp 1679581782
transform 1 0 65856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_687
timestamp 1679581782
transform 1 0 66528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_694
timestamp 1679581782
transform 1 0 67200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_701
timestamp 1679581782
transform 1 0 67872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_708
timestamp 1679581782
transform 1 0 68544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_715
timestamp 1679581782
transform 1 0 69216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_722
timestamp 1679581782
transform 1 0 69888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_729
timestamp 1679581782
transform 1 0 70560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_736
timestamp 1679581782
transform 1 0 71232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_743
timestamp 1679581782
transform 1 0 71904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_750
timestamp 1679581782
transform 1 0 72576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_757
timestamp 1679581782
transform 1 0 73248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_764
timestamp 1679581782
transform 1 0 73920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_771
timestamp 1679581782
transform 1 0 74592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_778
timestamp 1679581782
transform 1 0 75264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_785
timestamp 1679581782
transform 1 0 75936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_792
timestamp 1679581782
transform 1 0 76608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_799
timestamp 1679581782
transform 1 0 77280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_806
timestamp 1679581782
transform 1 0 77952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_813
timestamp 1679581782
transform 1 0 78624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_820
timestamp 1679581782
transform 1 0 79296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_827
timestamp 1679581782
transform 1 0 79968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_834
timestamp 1679581782
transform 1 0 80640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_841
timestamp 1679581782
transform 1 0 81312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_848
timestamp 1679581782
transform 1 0 81984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_855
timestamp 1679581782
transform 1 0 82656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_862
timestamp 1679581782
transform 1 0 83328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_869
timestamp 1679581782
transform 1 0 84000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_876
timestamp 1679581782
transform 1 0 84672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_883
timestamp 1679581782
transform 1 0 85344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_890
timestamp 1679581782
transform 1 0 86016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_897
timestamp 1679581782
transform 1 0 86688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_904
timestamp 1679581782
transform 1 0 87360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_911
timestamp 1679581782
transform 1 0 88032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_918
timestamp 1679581782
transform 1 0 88704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_925
timestamp 1679581782
transform 1 0 89376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_932
timestamp 1679581782
transform 1 0 90048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_939
timestamp 1679581782
transform 1 0 90720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_946
timestamp 1679581782
transform 1 0 91392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_953
timestamp 1679581782
transform 1 0 92064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_960
timestamp 1679581782
transform 1 0 92736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_967
timestamp 1679581782
transform 1 0 93408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_974
timestamp 1679581782
transform 1 0 94080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_981
timestamp 1679581782
transform 1 0 94752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_988
timestamp 1679581782
transform 1 0 95424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_995
timestamp 1679581782
transform 1 0 96096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1002
timestamp 1679581782
transform 1 0 96768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1009
timestamp 1679581782
transform 1 0 97440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1016
timestamp 1679581782
transform 1 0 98112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_1023
timestamp 1679577901
transform 1 0 98784 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_1027
timestamp 1677580104
transform 1 0 99168 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_0
timestamp 1677579658
transform 1 0 576 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_85
timestamp 1677579658
transform 1 0 8736 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_95
timestamp 1677580104
transform 1 0 9696 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_137
timestamp 1677580104
transform 1 0 13728 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_152
timestamp 1679581782
transform 1 0 15168 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_159
timestamp 1677579658
transform 1 0 15840 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_191
timestamp 1679581782
transform 1 0 18912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_198
timestamp 1679577901
transform 1 0 19584 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_202
timestamp 1677579658
transform 1 0 19968 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_215
timestamp 1677580104
transform 1 0 21216 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_223
timestamp 1679581782
transform 1 0 21984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_230
timestamp 1679581782
transform 1 0 22656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_237
timestamp 1679577901
transform 1 0 23328 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_241
timestamp 1677579658
transform 1 0 23712 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679581782
transform 1 0 26112 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_273
timestamp 1677580104
transform 1 0 26784 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_281
timestamp 1677580104
transform 1 0 27552 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_283
timestamp 1677579658
transform 1 0 27744 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_288
timestamp 1679581782
transform 1 0 28224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_295
timestamp 1679577901
transform 1 0 28896 0 1 15876
box -48 -56 432 834
use sg13g2_decap_4  FILLER_20_304
timestamp 1679577901
transform 1 0 29760 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_308
timestamp 1677580104
transform 1 0 30144 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_315
timestamp 1677580104
transform 1 0 30816 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_336
timestamp 1679581782
transform 1 0 32832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_343
timestamp 1679577901
transform 1 0 33504 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_347
timestamp 1677579658
transform 1 0 33888 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_352
timestamp 1679581782
transform 1 0 34368 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_372
timestamp 1677580104
transform 1 0 36288 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_374
timestamp 1677579658
transform 1 0 36480 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_438
timestamp 1679581782
transform 1 0 42624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_445
timestamp 1679581782
transform 1 0 43296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_452
timestamp 1679581782
transform 1 0 43968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_459
timestamp 1679581782
transform 1 0 44640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_466
timestamp 1679581782
transform 1 0 45312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_473
timestamp 1679581782
transform 1 0 45984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_480
timestamp 1679581782
transform 1 0 46656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_487
timestamp 1679581782
transform 1 0 47328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_494
timestamp 1679581782
transform 1 0 48000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_501
timestamp 1679581782
transform 1 0 48672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_508
timestamp 1679581782
transform 1 0 49344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_515
timestamp 1679581782
transform 1 0 50016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_522
timestamp 1679581782
transform 1 0 50688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_529
timestamp 1679581782
transform 1 0 51360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_536
timestamp 1679581782
transform 1 0 52032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_543
timestamp 1679581782
transform 1 0 52704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_550
timestamp 1679581782
transform 1 0 53376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_557
timestamp 1679581782
transform 1 0 54048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_564
timestamp 1679581782
transform 1 0 54720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_571
timestamp 1679581782
transform 1 0 55392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_578
timestamp 1679581782
transform 1 0 56064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_585
timestamp 1679581782
transform 1 0 56736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_592
timestamp 1679581782
transform 1 0 57408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_599
timestamp 1679581782
transform 1 0 58080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_606
timestamp 1679581782
transform 1 0 58752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_613
timestamp 1679581782
transform 1 0 59424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_620
timestamp 1679581782
transform 1 0 60096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_627
timestamp 1679581782
transform 1 0 60768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_634
timestamp 1679581782
transform 1 0 61440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_641
timestamp 1679581782
transform 1 0 62112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_648
timestamp 1679581782
transform 1 0 62784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_655
timestamp 1679581782
transform 1 0 63456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_662
timestamp 1679581782
transform 1 0 64128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_669
timestamp 1679581782
transform 1 0 64800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_676
timestamp 1679581782
transform 1 0 65472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_683
timestamp 1679581782
transform 1 0 66144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_690
timestamp 1679581782
transform 1 0 66816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_697
timestamp 1679581782
transform 1 0 67488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_704
timestamp 1679581782
transform 1 0 68160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_711
timestamp 1679581782
transform 1 0 68832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_718
timestamp 1679581782
transform 1 0 69504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_725
timestamp 1679581782
transform 1 0 70176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_732
timestamp 1679581782
transform 1 0 70848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_739
timestamp 1679581782
transform 1 0 71520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_746
timestamp 1679581782
transform 1 0 72192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_753
timestamp 1679581782
transform 1 0 72864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_760
timestamp 1679581782
transform 1 0 73536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_767
timestamp 1679581782
transform 1 0 74208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_774
timestamp 1679581782
transform 1 0 74880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_781
timestamp 1679581782
transform 1 0 75552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_788
timestamp 1679581782
transform 1 0 76224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_795
timestamp 1679581782
transform 1 0 76896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_802
timestamp 1679581782
transform 1 0 77568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_809
timestamp 1679581782
transform 1 0 78240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_816
timestamp 1679581782
transform 1 0 78912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_823
timestamp 1679581782
transform 1 0 79584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_830
timestamp 1679581782
transform 1 0 80256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_837
timestamp 1679581782
transform 1 0 80928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_844
timestamp 1679581782
transform 1 0 81600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_851
timestamp 1679581782
transform 1 0 82272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_858
timestamp 1679581782
transform 1 0 82944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_865
timestamp 1679581782
transform 1 0 83616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_872
timestamp 1679581782
transform 1 0 84288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_879
timestamp 1679581782
transform 1 0 84960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_886
timestamp 1679581782
transform 1 0 85632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_893
timestamp 1679581782
transform 1 0 86304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_900
timestamp 1679581782
transform 1 0 86976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_907
timestamp 1679581782
transform 1 0 87648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_914
timestamp 1679581782
transform 1 0 88320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_921
timestamp 1679581782
transform 1 0 88992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_928
timestamp 1679581782
transform 1 0 89664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_935
timestamp 1679581782
transform 1 0 90336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_942
timestamp 1679581782
transform 1 0 91008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_949
timestamp 1679581782
transform 1 0 91680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_956
timestamp 1679581782
transform 1 0 92352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_963
timestamp 1679581782
transform 1 0 93024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_970
timestamp 1679581782
transform 1 0 93696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_977
timestamp 1679581782
transform 1 0 94368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_984
timestamp 1679581782
transform 1 0 95040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_991
timestamp 1679581782
transform 1 0 95712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_998
timestamp 1679581782
transform 1 0 96384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1005
timestamp 1679581782
transform 1 0 97056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1012
timestamp 1679581782
transform 1 0 97728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1019
timestamp 1679581782
transform 1 0 98400 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_1026
timestamp 1677580104
transform 1 0 99072 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_1028
timestamp 1677579658
transform 1 0 99264 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_4
timestamp 1677580104
transform 1 0 960 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_6
timestamp 1677579658
transform 1 0 1152 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_47
timestamp 1677579658
transform 1 0 5088 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_123
timestamp 1679581782
transform 1 0 12384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13056 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_137
timestamp 1677580104
transform 1 0 13728 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_148
timestamp 1677580104
transform 1 0 14784 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_154
timestamp 1679577901
transform 1 0 15360 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_158
timestamp 1677579658
transform 1 0 15744 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_206
timestamp 1679577901
transform 1 0 20352 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_210
timestamp 1677580104
transform 1 0 20736 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_216
timestamp 1679577901
transform 1 0 21312 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_220
timestamp 1677579658
transform 1 0 21696 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_233
timestamp 1679581782
transform 1 0 22944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_240
timestamp 1679577901
transform 1 0 23616 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_244
timestamp 1677579658
transform 1 0 24000 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_265
timestamp 1677580104
transform 1 0 26016 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_273
timestamp 1679581782
transform 1 0 26784 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_307
timestamp 1677580104
transform 1 0 30048 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_309
timestamp 1677579658
transform 1 0 30240 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_335
timestamp 1679577901
transform 1 0 32736 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_339
timestamp 1677579658
transform 1 0 33120 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_381
timestamp 1677579658
transform 1 0 37152 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_409
timestamp 1679581782
transform 1 0 39840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_416
timestamp 1679581782
transform 1 0 40512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_423
timestamp 1679581782
transform 1 0 41184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_456
timestamp 1679581782
transform 1 0 44352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_463
timestamp 1679581782
transform 1 0 45024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_470
timestamp 1679581782
transform 1 0 45696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_477
timestamp 1679581782
transform 1 0 46368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_484
timestamp 1679581782
transform 1 0 47040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_491
timestamp 1679581782
transform 1 0 47712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_498
timestamp 1679581782
transform 1 0 48384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_505
timestamp 1679581782
transform 1 0 49056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_512
timestamp 1679581782
transform 1 0 49728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_519
timestamp 1679581782
transform 1 0 50400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_526
timestamp 1679581782
transform 1 0 51072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_533
timestamp 1679581782
transform 1 0 51744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_540
timestamp 1679581782
transform 1 0 52416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_547
timestamp 1679581782
transform 1 0 53088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_554
timestamp 1679581782
transform 1 0 53760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_561
timestamp 1679581782
transform 1 0 54432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_568
timestamp 1679581782
transform 1 0 55104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_575
timestamp 1679581782
transform 1 0 55776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_582
timestamp 1679581782
transform 1 0 56448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_589
timestamp 1679581782
transform 1 0 57120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_596
timestamp 1679581782
transform 1 0 57792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_603
timestamp 1679581782
transform 1 0 58464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_610
timestamp 1679581782
transform 1 0 59136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_617
timestamp 1679581782
transform 1 0 59808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_624
timestamp 1679581782
transform 1 0 60480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_631
timestamp 1679581782
transform 1 0 61152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_638
timestamp 1679581782
transform 1 0 61824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_645
timestamp 1679581782
transform 1 0 62496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_652
timestamp 1679581782
transform 1 0 63168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_659
timestamp 1679581782
transform 1 0 63840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_666
timestamp 1679581782
transform 1 0 64512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_673
timestamp 1679581782
transform 1 0 65184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_680
timestamp 1679581782
transform 1 0 65856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_687
timestamp 1679581782
transform 1 0 66528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_694
timestamp 1679581782
transform 1 0 67200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_701
timestamp 1679581782
transform 1 0 67872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_708
timestamp 1679581782
transform 1 0 68544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_715
timestamp 1679581782
transform 1 0 69216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_722
timestamp 1679581782
transform 1 0 69888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_729
timestamp 1679581782
transform 1 0 70560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_736
timestamp 1679581782
transform 1 0 71232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_743
timestamp 1679581782
transform 1 0 71904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_750
timestamp 1679581782
transform 1 0 72576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_757
timestamp 1679581782
transform 1 0 73248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_764
timestamp 1679581782
transform 1 0 73920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_771
timestamp 1679581782
transform 1 0 74592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_778
timestamp 1679581782
transform 1 0 75264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_785
timestamp 1679581782
transform 1 0 75936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_792
timestamp 1679581782
transform 1 0 76608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_799
timestamp 1679581782
transform 1 0 77280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_806
timestamp 1679581782
transform 1 0 77952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_813
timestamp 1679581782
transform 1 0 78624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_820
timestamp 1679581782
transform 1 0 79296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_827
timestamp 1679581782
transform 1 0 79968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_834
timestamp 1679581782
transform 1 0 80640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_841
timestamp 1679581782
transform 1 0 81312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_848
timestamp 1679581782
transform 1 0 81984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_855
timestamp 1679581782
transform 1 0 82656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_862
timestamp 1679581782
transform 1 0 83328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_869
timestamp 1679581782
transform 1 0 84000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_876
timestamp 1679581782
transform 1 0 84672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_883
timestamp 1679581782
transform 1 0 85344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_890
timestamp 1679581782
transform 1 0 86016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_897
timestamp 1679581782
transform 1 0 86688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_904
timestamp 1679581782
transform 1 0 87360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_911
timestamp 1679581782
transform 1 0 88032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_918
timestamp 1679581782
transform 1 0 88704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_925
timestamp 1679581782
transform 1 0 89376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_932
timestamp 1679581782
transform 1 0 90048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_939
timestamp 1679581782
transform 1 0 90720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_946
timestamp 1679581782
transform 1 0 91392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_953
timestamp 1679581782
transform 1 0 92064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_960
timestamp 1679581782
transform 1 0 92736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_967
timestamp 1679581782
transform 1 0 93408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_974
timestamp 1679581782
transform 1 0 94080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_981
timestamp 1679581782
transform 1 0 94752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_988
timestamp 1679581782
transform 1 0 95424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_995
timestamp 1679581782
transform 1 0 96096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1002
timestamp 1679581782
transform 1 0 96768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1009
timestamp 1679581782
transform 1 0 97440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1016
timestamp 1679581782
transform 1 0 98112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1023
timestamp 1679577901
transform 1 0 98784 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_1027
timestamp 1677580104
transform 1 0 99168 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_0
timestamp 1677580104
transform 1 0 576 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_33
timestamp 1677579658
transform 1 0 3744 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_60
timestamp 1677579658
transform 1 0 6336 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_74
timestamp 1677579658
transform 1 0 7680 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_111
timestamp 1679581782
transform 1 0 11232 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_118
timestamp 1677579658
transform 1 0 11904 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_201
timestamp 1679581782
transform 1 0 19872 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_228
timestamp 1677580104
transform 1 0 22464 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_243
timestamp 1677580104
transform 1 0 23904 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_256
timestamp 1677579658
transform 1 0 25152 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_283
timestamp 1677579658
transform 1 0 27744 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_297
timestamp 1677579658
transform 1 0 29088 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_308
timestamp 1677580104
transform 1 0 30144 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_310
timestamp 1677579658
transform 1 0 30336 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_320
timestamp 1677580104
transform 1 0 31296 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_322
timestamp 1677579658
transform 1 0 31488 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_336
timestamp 1677580104
transform 1 0 32832 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_365
timestamp 1677580104
transform 1 0 35616 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_367
timestamp 1677579658
transform 1 0 35808 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_372
timestamp 1679577901
transform 1 0 36288 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_376
timestamp 1677579658
transform 1 0 36672 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_390
timestamp 1679581782
transform 1 0 38016 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_397
timestamp 1677579658
transform 1 0 38688 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_407
timestamp 1679577901
transform 1 0 39648 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_411
timestamp 1677579658
transform 1 0 40032 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_430
timestamp 1679581782
transform 1 0 41856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_437
timestamp 1679581782
transform 1 0 42528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_444
timestamp 1679581782
transform 1 0 43200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_451
timestamp 1679581782
transform 1 0 43872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_458
timestamp 1679581782
transform 1 0 44544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_465
timestamp 1679581782
transform 1 0 45216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_472
timestamp 1679581782
transform 1 0 45888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_479
timestamp 1679581782
transform 1 0 46560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_486
timestamp 1679581782
transform 1 0 47232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_493
timestamp 1679581782
transform 1 0 47904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_500
timestamp 1679581782
transform 1 0 48576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_507
timestamp 1679581782
transform 1 0 49248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_514
timestamp 1679581782
transform 1 0 49920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_521
timestamp 1679581782
transform 1 0 50592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_528
timestamp 1679581782
transform 1 0 51264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_535
timestamp 1679581782
transform 1 0 51936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_542
timestamp 1679581782
transform 1 0 52608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_549
timestamp 1679581782
transform 1 0 53280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_556
timestamp 1679581782
transform 1 0 53952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_563
timestamp 1679581782
transform 1 0 54624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_570
timestamp 1679581782
transform 1 0 55296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_577
timestamp 1679581782
transform 1 0 55968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_584
timestamp 1679581782
transform 1 0 56640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_591
timestamp 1679581782
transform 1 0 57312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_598
timestamp 1679581782
transform 1 0 57984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_605
timestamp 1679581782
transform 1 0 58656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_612
timestamp 1679581782
transform 1 0 59328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_619
timestamp 1679581782
transform 1 0 60000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_626
timestamp 1679581782
transform 1 0 60672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_633
timestamp 1679581782
transform 1 0 61344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_640
timestamp 1679581782
transform 1 0 62016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_647
timestamp 1679581782
transform 1 0 62688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_654
timestamp 1679581782
transform 1 0 63360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_661
timestamp 1679581782
transform 1 0 64032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_668
timestamp 1679581782
transform 1 0 64704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_675
timestamp 1679581782
transform 1 0 65376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_682
timestamp 1679581782
transform 1 0 66048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_689
timestamp 1679581782
transform 1 0 66720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_696
timestamp 1679581782
transform 1 0 67392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_703
timestamp 1679581782
transform 1 0 68064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_710
timestamp 1679581782
transform 1 0 68736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_717
timestamp 1679581782
transform 1 0 69408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_724
timestamp 1679581782
transform 1 0 70080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_731
timestamp 1679581782
transform 1 0 70752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_738
timestamp 1679581782
transform 1 0 71424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_745
timestamp 1679581782
transform 1 0 72096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_752
timestamp 1679581782
transform 1 0 72768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_759
timestamp 1679581782
transform 1 0 73440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_766
timestamp 1679581782
transform 1 0 74112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_773
timestamp 1679581782
transform 1 0 74784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_780
timestamp 1679581782
transform 1 0 75456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_787
timestamp 1679581782
transform 1 0 76128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_794
timestamp 1679581782
transform 1 0 76800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_801
timestamp 1679581782
transform 1 0 77472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_808
timestamp 1679581782
transform 1 0 78144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_815
timestamp 1679581782
transform 1 0 78816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_822
timestamp 1679581782
transform 1 0 79488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_829
timestamp 1679581782
transform 1 0 80160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_836
timestamp 1679581782
transform 1 0 80832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_843
timestamp 1679581782
transform 1 0 81504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_850
timestamp 1679581782
transform 1 0 82176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_857
timestamp 1679581782
transform 1 0 82848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_864
timestamp 1679581782
transform 1 0 83520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_871
timestamp 1679581782
transform 1 0 84192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_878
timestamp 1679581782
transform 1 0 84864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_885
timestamp 1679581782
transform 1 0 85536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_892
timestamp 1679581782
transform 1 0 86208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_899
timestamp 1679581782
transform 1 0 86880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_906
timestamp 1679581782
transform 1 0 87552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_913
timestamp 1679581782
transform 1 0 88224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_920
timestamp 1679581782
transform 1 0 88896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_927
timestamp 1679581782
transform 1 0 89568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_934
timestamp 1679581782
transform 1 0 90240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_941
timestamp 1679581782
transform 1 0 90912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_948
timestamp 1679581782
transform 1 0 91584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_955
timestamp 1679581782
transform 1 0 92256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_962
timestamp 1679581782
transform 1 0 92928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_969
timestamp 1679581782
transform 1 0 93600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_976
timestamp 1679581782
transform 1 0 94272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_983
timestamp 1679581782
transform 1 0 94944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_990
timestamp 1679581782
transform 1 0 95616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_997
timestamp 1679581782
transform 1 0 96288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1004
timestamp 1679581782
transform 1 0 96960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1011
timestamp 1679581782
transform 1 0 97632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1018
timestamp 1679581782
transform 1 0 98304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_1025
timestamp 1679577901
transform 1 0 98976 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_15
timestamp 1679581782
transform 1 0 2016 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_50
timestamp 1677579658
transform 1 0 5376 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_57
timestamp 1677579658
transform 1 0 6048 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_82
timestamp 1677580104
transform 1 0 8448 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_110
timestamp 1679581782
transform 1 0 11136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_117
timestamp 1679581782
transform 1 0 11808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_128
timestamp 1679581782
transform 1 0 12864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_135
timestamp 1679581782
transform 1 0 13536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_142
timestamp 1679577901
transform 1 0 14208 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_146
timestamp 1677579658
transform 1 0 14592 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_201
timestamp 1679581782
transform 1 0 19872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_220
timestamp 1679577901
transform 1 0 21696 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_224
timestamp 1677580104
transform 1 0 22080 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_232
timestamp 1679581782
transform 1 0 22848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_239
timestamp 1679577901
transform 1 0 23520 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_243
timestamp 1677580104
transform 1 0 23904 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_254
timestamp 1677579658
transform 1 0 24960 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_268
timestamp 1679581782
transform 1 0 26304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_275
timestamp 1679577901
transform 1 0 26976 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_279
timestamp 1677579658
transform 1 0 27360 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_297
timestamp 1677580104
transform 1 0 29088 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_308
timestamp 1677579658
transform 1 0 30144 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_313
timestamp 1679581782
transform 1 0 30624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_320
timestamp 1679581782
transform 1 0 31296 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_327
timestamp 1677579658
transform 1 0 31968 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_334
timestamp 1677580104
transform 1 0 32640 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_341
timestamp 1677580104
transform 1 0 33312 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_343
timestamp 1677579658
transform 1 0 33504 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_385
timestamp 1677580104
transform 1 0 37536 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_387
timestamp 1677579658
transform 1 0 37728 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_442
timestamp 1679581782
transform 1 0 43008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_449
timestamp 1679577901
transform 1 0 43680 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_453
timestamp 1677579658
transform 1 0 44064 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_482
timestamp 1679581782
transform 1 0 46848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_489
timestamp 1679581782
transform 1 0 47520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_496
timestamp 1679581782
transform 1 0 48192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_503
timestamp 1679581782
transform 1 0 48864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_510
timestamp 1679581782
transform 1 0 49536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_517
timestamp 1679581782
transform 1 0 50208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_524
timestamp 1679581782
transform 1 0 50880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_531
timestamp 1679581782
transform 1 0 51552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_538
timestamp 1679581782
transform 1 0 52224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_545
timestamp 1679581782
transform 1 0 52896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_552
timestamp 1679581782
transform 1 0 53568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_559
timestamp 1679581782
transform 1 0 54240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_566
timestamp 1679581782
transform 1 0 54912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_573
timestamp 1679581782
transform 1 0 55584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_580
timestamp 1679581782
transform 1 0 56256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_587
timestamp 1679581782
transform 1 0 56928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_594
timestamp 1679581782
transform 1 0 57600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_601
timestamp 1679581782
transform 1 0 58272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_608
timestamp 1679581782
transform 1 0 58944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_615
timestamp 1679581782
transform 1 0 59616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_622
timestamp 1679581782
transform 1 0 60288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_629
timestamp 1679581782
transform 1 0 60960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_636
timestamp 1679581782
transform 1 0 61632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_643
timestamp 1679581782
transform 1 0 62304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_650
timestamp 1679581782
transform 1 0 62976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_657
timestamp 1679581782
transform 1 0 63648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_664
timestamp 1679581782
transform 1 0 64320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_671
timestamp 1679581782
transform 1 0 64992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_678
timestamp 1679581782
transform 1 0 65664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_685
timestamp 1679581782
transform 1 0 66336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_692
timestamp 1679581782
transform 1 0 67008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_699
timestamp 1679581782
transform 1 0 67680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_706
timestamp 1679581782
transform 1 0 68352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_713
timestamp 1679581782
transform 1 0 69024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_720
timestamp 1679581782
transform 1 0 69696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_727
timestamp 1679581782
transform 1 0 70368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_734
timestamp 1679581782
transform 1 0 71040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_741
timestamp 1679581782
transform 1 0 71712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_748
timestamp 1679581782
transform 1 0 72384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_755
timestamp 1679581782
transform 1 0 73056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_762
timestamp 1679581782
transform 1 0 73728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_769
timestamp 1679581782
transform 1 0 74400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_776
timestamp 1679581782
transform 1 0 75072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_783
timestamp 1679581782
transform 1 0 75744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_790
timestamp 1679581782
transform 1 0 76416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_797
timestamp 1679581782
transform 1 0 77088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_804
timestamp 1679581782
transform 1 0 77760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_811
timestamp 1679581782
transform 1 0 78432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_818
timestamp 1679581782
transform 1 0 79104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_825
timestamp 1679581782
transform 1 0 79776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_832
timestamp 1679581782
transform 1 0 80448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_839
timestamp 1679581782
transform 1 0 81120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_846
timestamp 1679581782
transform 1 0 81792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_853
timestamp 1679581782
transform 1 0 82464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_860
timestamp 1679581782
transform 1 0 83136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_867
timestamp 1679581782
transform 1 0 83808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_874
timestamp 1679581782
transform 1 0 84480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_881
timestamp 1679581782
transform 1 0 85152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_888
timestamp 1679581782
transform 1 0 85824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_895
timestamp 1679581782
transform 1 0 86496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_902
timestamp 1679581782
transform 1 0 87168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_909
timestamp 1679581782
transform 1 0 87840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_916
timestamp 1679581782
transform 1 0 88512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_923
timestamp 1679581782
transform 1 0 89184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_930
timestamp 1679581782
transform 1 0 89856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_937
timestamp 1679581782
transform 1 0 90528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_944
timestamp 1679581782
transform 1 0 91200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_951
timestamp 1679581782
transform 1 0 91872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_958
timestamp 1679581782
transform 1 0 92544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_965
timestamp 1679581782
transform 1 0 93216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_972
timestamp 1679581782
transform 1 0 93888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_979
timestamp 1679581782
transform 1 0 94560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_986
timestamp 1679581782
transform 1 0 95232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_993
timestamp 1679581782
transform 1 0 95904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1000
timestamp 1679581782
transform 1 0 96576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1007
timestamp 1679581782
transform 1 0 97248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1014
timestamp 1679581782
transform 1 0 97920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1021
timestamp 1679581782
transform 1 0 98592 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677579658
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_11
timestamp 1677580104
transform 1 0 1632 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_40
timestamp 1677580104
transform 1 0 4416 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_70
timestamp 1679577901
transform 1 0 7296 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_74
timestamp 1677579658
transform 1 0 7680 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_79
timestamp 1677579658
transform 1 0 8160 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_88
timestamp 1677580104
transform 1 0 9024 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_94
timestamp 1677580104
transform 1 0 9600 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_96
timestamp 1677579658
transform 1 0 9792 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_106
timestamp 1677580104
transform 1 0 10752 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_113
timestamp 1679577901
transform 1 0 11424 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_144
timestamp 1677580104
transform 1 0 14400 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_159
timestamp 1677580104
transform 1 0 15840 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_232
timestamp 1677580104
transform 1 0 22848 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_234
timestamp 1677579658
transform 1 0 23040 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_245
timestamp 1679581782
transform 1 0 24096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_252
timestamp 1679577901
transform 1 0 24768 0 1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_24_266
timestamp 1679577901
transform 1 0 26112 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_270
timestamp 1677580104
transform 1 0 26496 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_313
timestamp 1679581782
transform 1 0 30624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_320
timestamp 1679581782
transform 1 0 31296 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_327
timestamp 1677579658
transform 1 0 31968 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_390
timestamp 1677579658
transform 1 0 38016 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_405
timestamp 1677579658
transform 1 0 39456 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_423
timestamp 1679581782
transform 1 0 41184 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_430
timestamp 1677580104
transform 1 0 41856 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_432
timestamp 1677579658
transform 1 0 42048 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_442
timestamp 1677579658
transform 1 0 43008 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_465
timestamp 1679581782
transform 1 0 45216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_472
timestamp 1679581782
transform 1 0 45888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_479
timestamp 1679581782
transform 1 0 46560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_486
timestamp 1679581782
transform 1 0 47232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_493
timestamp 1679581782
transform 1 0 47904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_500
timestamp 1679581782
transform 1 0 48576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_507
timestamp 1679581782
transform 1 0 49248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_514
timestamp 1679581782
transform 1 0 49920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_521
timestamp 1679581782
transform 1 0 50592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_528
timestamp 1679581782
transform 1 0 51264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_535
timestamp 1679581782
transform 1 0 51936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_542
timestamp 1679581782
transform 1 0 52608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_549
timestamp 1679581782
transform 1 0 53280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_556
timestamp 1679581782
transform 1 0 53952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_563
timestamp 1679581782
transform 1 0 54624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_570
timestamp 1679581782
transform 1 0 55296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_577
timestamp 1679581782
transform 1 0 55968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_584
timestamp 1679581782
transform 1 0 56640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_591
timestamp 1679581782
transform 1 0 57312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_598
timestamp 1679581782
transform 1 0 57984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_605
timestamp 1679581782
transform 1 0 58656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_612
timestamp 1679581782
transform 1 0 59328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_619
timestamp 1679581782
transform 1 0 60000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_626
timestamp 1679581782
transform 1 0 60672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_633
timestamp 1679581782
transform 1 0 61344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_640
timestamp 1679581782
transform 1 0 62016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_647
timestamp 1679581782
transform 1 0 62688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_654
timestamp 1679581782
transform 1 0 63360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_661
timestamp 1679581782
transform 1 0 64032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_668
timestamp 1679581782
transform 1 0 64704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_675
timestamp 1679581782
transform 1 0 65376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_682
timestamp 1679581782
transform 1 0 66048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_689
timestamp 1679581782
transform 1 0 66720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_696
timestamp 1679581782
transform 1 0 67392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_703
timestamp 1679581782
transform 1 0 68064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_710
timestamp 1679581782
transform 1 0 68736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_717
timestamp 1679581782
transform 1 0 69408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_724
timestamp 1679581782
transform 1 0 70080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_731
timestamp 1679581782
transform 1 0 70752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_738
timestamp 1679581782
transform 1 0 71424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_745
timestamp 1679581782
transform 1 0 72096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_752
timestamp 1679581782
transform 1 0 72768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_759
timestamp 1679581782
transform 1 0 73440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_766
timestamp 1679581782
transform 1 0 74112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_773
timestamp 1679581782
transform 1 0 74784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_780
timestamp 1679581782
transform 1 0 75456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_787
timestamp 1679581782
transform 1 0 76128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_794
timestamp 1679581782
transform 1 0 76800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_801
timestamp 1679581782
transform 1 0 77472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_808
timestamp 1679581782
transform 1 0 78144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_815
timestamp 1679581782
transform 1 0 78816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_822
timestamp 1679581782
transform 1 0 79488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_829
timestamp 1679581782
transform 1 0 80160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_836
timestamp 1679581782
transform 1 0 80832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_843
timestamp 1679581782
transform 1 0 81504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_850
timestamp 1679581782
transform 1 0 82176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_857
timestamp 1679581782
transform 1 0 82848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_864
timestamp 1679581782
transform 1 0 83520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_871
timestamp 1679581782
transform 1 0 84192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_878
timestamp 1679581782
transform 1 0 84864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_885
timestamp 1679581782
transform 1 0 85536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_892
timestamp 1679581782
transform 1 0 86208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_899
timestamp 1679581782
transform 1 0 86880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_906
timestamp 1679581782
transform 1 0 87552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_913
timestamp 1679581782
transform 1 0 88224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_920
timestamp 1679581782
transform 1 0 88896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_927
timestamp 1679581782
transform 1 0 89568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_934
timestamp 1679581782
transform 1 0 90240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_941
timestamp 1679581782
transform 1 0 90912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_948
timestamp 1679581782
transform 1 0 91584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_955
timestamp 1679581782
transform 1 0 92256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_962
timestamp 1679581782
transform 1 0 92928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_969
timestamp 1679581782
transform 1 0 93600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_976
timestamp 1679581782
transform 1 0 94272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_983
timestamp 1679581782
transform 1 0 94944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_990
timestamp 1679581782
transform 1 0 95616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_997
timestamp 1679581782
transform 1 0 96288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1004
timestamp 1679581782
transform 1 0 96960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1011
timestamp 1679581782
transform 1 0 97632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1018
timestamp 1679581782
transform 1 0 98304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_1025
timestamp 1679577901
transform 1 0 98976 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_22
timestamp 1679581782
transform 1 0 2688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_29
timestamp 1679577901
transform 1 0 3360 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_38
timestamp 1679577901
transform 1 0 4224 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_42
timestamp 1677580104
transform 1 0 4608 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_79
timestamp 1677580104
transform 1 0 8160 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_84
timestamp 1677579658
transform 1 0 8640 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_186
timestamp 1677580104
transform 1 0 18432 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_188
timestamp 1677579658
transform 1 0 18624 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_207
timestamp 1679577901
transform 1 0 20448 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_211
timestamp 1677579658
transform 1 0 20832 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_225
timestamp 1677579658
transform 1 0 22176 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_266
timestamp 1677580104
transform 1 0 26112 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_268
timestamp 1677579658
transform 1 0 26304 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_295
timestamp 1677579658
transform 1 0 28896 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_329
timestamp 1679581782
transform 1 0 32160 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_336
timestamp 1677579658
transform 1 0 32832 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_341
timestamp 1679577901
transform 1 0 33312 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_349
timestamp 1679581782
transform 1 0 34080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_356
timestamp 1679581782
transform 1 0 34752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_363
timestamp 1679577901
transform 1 0 35424 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_367
timestamp 1677580104
transform 1 0 35808 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_373
timestamp 1677579658
transform 1 0 36384 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_386
timestamp 1677579658
transform 1 0 37632 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_401
timestamp 1677579658
transform 1 0 39072 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_408
timestamp 1679577901
transform 1 0 39744 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_412
timestamp 1677580104
transform 1 0 40128 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_427
timestamp 1677579658
transform 1 0 41568 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_460
timestamp 1679577901
transform 1 0 44736 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_491
timestamp 1679581782
transform 1 0 47712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_498
timestamp 1679581782
transform 1 0 48384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_505
timestamp 1679581782
transform 1 0 49056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_512
timestamp 1679581782
transform 1 0 49728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_519
timestamp 1679581782
transform 1 0 50400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_526
timestamp 1679581782
transform 1 0 51072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_533
timestamp 1679581782
transform 1 0 51744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_540
timestamp 1679581782
transform 1 0 52416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_547
timestamp 1679581782
transform 1 0 53088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_554
timestamp 1679581782
transform 1 0 53760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_561
timestamp 1679581782
transform 1 0 54432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_568
timestamp 1679581782
transform 1 0 55104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_575
timestamp 1679581782
transform 1 0 55776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_582
timestamp 1679581782
transform 1 0 56448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_589
timestamp 1679581782
transform 1 0 57120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_596
timestamp 1679581782
transform 1 0 57792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_603
timestamp 1679581782
transform 1 0 58464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_610
timestamp 1679581782
transform 1 0 59136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_617
timestamp 1679581782
transform 1 0 59808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_624
timestamp 1679581782
transform 1 0 60480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_631
timestamp 1679581782
transform 1 0 61152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_638
timestamp 1679581782
transform 1 0 61824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_645
timestamp 1679581782
transform 1 0 62496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_652
timestamp 1679581782
transform 1 0 63168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_659
timestamp 1679581782
transform 1 0 63840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_666
timestamp 1679581782
transform 1 0 64512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_673
timestamp 1679581782
transform 1 0 65184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_680
timestamp 1679581782
transform 1 0 65856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_687
timestamp 1679581782
transform 1 0 66528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_694
timestamp 1679581782
transform 1 0 67200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_701
timestamp 1679581782
transform 1 0 67872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_708
timestamp 1679581782
transform 1 0 68544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_715
timestamp 1679581782
transform 1 0 69216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_722
timestamp 1679581782
transform 1 0 69888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_729
timestamp 1679581782
transform 1 0 70560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_736
timestamp 1679581782
transform 1 0 71232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_743
timestamp 1679581782
transform 1 0 71904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_750
timestamp 1679581782
transform 1 0 72576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_757
timestamp 1679581782
transform 1 0 73248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_764
timestamp 1679581782
transform 1 0 73920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_771
timestamp 1679581782
transform 1 0 74592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_778
timestamp 1679581782
transform 1 0 75264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_785
timestamp 1679581782
transform 1 0 75936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_792
timestamp 1679581782
transform 1 0 76608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_799
timestamp 1679581782
transform 1 0 77280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_806
timestamp 1679581782
transform 1 0 77952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_813
timestamp 1679581782
transform 1 0 78624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_820
timestamp 1679581782
transform 1 0 79296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_827
timestamp 1679581782
transform 1 0 79968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_834
timestamp 1679581782
transform 1 0 80640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_841
timestamp 1679581782
transform 1 0 81312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_848
timestamp 1679581782
transform 1 0 81984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_855
timestamp 1679581782
transform 1 0 82656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_862
timestamp 1679581782
transform 1 0 83328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_869
timestamp 1679581782
transform 1 0 84000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_876
timestamp 1679581782
transform 1 0 84672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_883
timestamp 1679581782
transform 1 0 85344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_890
timestamp 1679581782
transform 1 0 86016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_897
timestamp 1679581782
transform 1 0 86688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_904
timestamp 1679581782
transform 1 0 87360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_911
timestamp 1679581782
transform 1 0 88032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_918
timestamp 1679581782
transform 1 0 88704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_925
timestamp 1679581782
transform 1 0 89376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_932
timestamp 1679581782
transform 1 0 90048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_939
timestamp 1679581782
transform 1 0 90720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_946
timestamp 1679581782
transform 1 0 91392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_953
timestamp 1679581782
transform 1 0 92064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_960
timestamp 1679581782
transform 1 0 92736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_967
timestamp 1679581782
transform 1 0 93408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_974
timestamp 1679581782
transform 1 0 94080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_981
timestamp 1679581782
transform 1 0 94752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_988
timestamp 1679581782
transform 1 0 95424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_995
timestamp 1679581782
transform 1 0 96096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1002
timestamp 1679581782
transform 1 0 96768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1009
timestamp 1679581782
transform 1 0 97440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1016
timestamp 1679581782
transform 1 0 98112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_1023
timestamp 1679577901
transform 1 0 98784 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_1027
timestamp 1677580104
transform 1 0 99168 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679581782
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679581782
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_47
timestamp 1679577901
transform 1 0 5088 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_55
timestamp 1677579658
transform 1 0 5856 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_78
timestamp 1679581782
transform 1 0 8064 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_99
timestamp 1677580104
transform 1 0 10080 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_142
timestamp 1677580104
transform 1 0 14208 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_144
timestamp 1677579658
transform 1 0 14400 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_148
timestamp 1677580104
transform 1 0 14784 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_167
timestamp 1679577901
transform 1 0 16608 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_175
timestamp 1679581782
transform 1 0 17376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_182
timestamp 1679581782
transform 1 0 18048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_189
timestamp 1679581782
transform 1 0 18720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_196
timestamp 1679577901
transform 1 0 19392 0 1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_26_212
timestamp 1679577901
transform 1 0 20928 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_226
timestamp 1677580104
transform 1 0 22272 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_248
timestamp 1679577901
transform 1 0 24384 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_252
timestamp 1677580104
transform 1 0 24768 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_282
timestamp 1679581782
transform 1 0 27648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_289
timestamp 1679581782
transform 1 0 28320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_296
timestamp 1679581782
transform 1 0 28992 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_303
timestamp 1677580104
transform 1 0 29664 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_305
timestamp 1677579658
transform 1 0 29856 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_310
timestamp 1677580104
transform 1 0 30336 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_312
timestamp 1677579658
transform 1 0 30528 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_326
timestamp 1677580104
transform 1 0 31872 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_328
timestamp 1677579658
transform 1 0 32064 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_345
timestamp 1679581782
transform 1 0 33696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_352
timestamp 1679581782
transform 1 0 34368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_359
timestamp 1679577901
transform 1 0 35040 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_363
timestamp 1677579658
transform 1 0 35424 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_412
timestamp 1677580104
transform 1 0 40128 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_414
timestamp 1677579658
transform 1 0 40320 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_463
timestamp 1677580104
transform 1 0 45024 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_487
timestamp 1679577901
transform 1 0 47328 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_491
timestamp 1677579658
transform 1 0 47712 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_519
timestamp 1679581782
transform 1 0 50400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_526
timestamp 1679581782
transform 1 0 51072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_533
timestamp 1679581782
transform 1 0 51744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_540
timestamp 1679581782
transform 1 0 52416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_547
timestamp 1679581782
transform 1 0 53088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_554
timestamp 1679581782
transform 1 0 53760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_561
timestamp 1679581782
transform 1 0 54432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_568
timestamp 1679581782
transform 1 0 55104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_575
timestamp 1679581782
transform 1 0 55776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_582
timestamp 1679581782
transform 1 0 56448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_589
timestamp 1679581782
transform 1 0 57120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_596
timestamp 1679581782
transform 1 0 57792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_603
timestamp 1679581782
transform 1 0 58464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_610
timestamp 1679581782
transform 1 0 59136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_617
timestamp 1679581782
transform 1 0 59808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_624
timestamp 1679581782
transform 1 0 60480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_631
timestamp 1679581782
transform 1 0 61152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_638
timestamp 1679581782
transform 1 0 61824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_645
timestamp 1679581782
transform 1 0 62496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_652
timestamp 1679581782
transform 1 0 63168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_659
timestamp 1679581782
transform 1 0 63840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_666
timestamp 1679581782
transform 1 0 64512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_673
timestamp 1679581782
transform 1 0 65184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_680
timestamp 1679581782
transform 1 0 65856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_687
timestamp 1679581782
transform 1 0 66528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_694
timestamp 1679581782
transform 1 0 67200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_701
timestamp 1679581782
transform 1 0 67872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_708
timestamp 1679581782
transform 1 0 68544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_715
timestamp 1679581782
transform 1 0 69216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_722
timestamp 1679581782
transform 1 0 69888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_729
timestamp 1679581782
transform 1 0 70560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_736
timestamp 1679581782
transform 1 0 71232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_743
timestamp 1679581782
transform 1 0 71904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_750
timestamp 1679581782
transform 1 0 72576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_757
timestamp 1679581782
transform 1 0 73248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_764
timestamp 1679581782
transform 1 0 73920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_771
timestamp 1679581782
transform 1 0 74592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_778
timestamp 1679581782
transform 1 0 75264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_785
timestamp 1679581782
transform 1 0 75936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_792
timestamp 1679581782
transform 1 0 76608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_799
timestamp 1679581782
transform 1 0 77280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_806
timestamp 1679581782
transform 1 0 77952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_813
timestamp 1679581782
transform 1 0 78624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_820
timestamp 1679581782
transform 1 0 79296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_827
timestamp 1679581782
transform 1 0 79968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_834
timestamp 1679581782
transform 1 0 80640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_841
timestamp 1679581782
transform 1 0 81312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_848
timestamp 1679581782
transform 1 0 81984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_855
timestamp 1679581782
transform 1 0 82656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_862
timestamp 1679581782
transform 1 0 83328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_869
timestamp 1679581782
transform 1 0 84000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_876
timestamp 1679581782
transform 1 0 84672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_883
timestamp 1679581782
transform 1 0 85344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_890
timestamp 1679581782
transform 1 0 86016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_897
timestamp 1679581782
transform 1 0 86688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_904
timestamp 1679581782
transform 1 0 87360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_911
timestamp 1679581782
transform 1 0 88032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_918
timestamp 1679581782
transform 1 0 88704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_925
timestamp 1679581782
transform 1 0 89376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_932
timestamp 1679581782
transform 1 0 90048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_939
timestamp 1679581782
transform 1 0 90720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_946
timestamp 1679581782
transform 1 0 91392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_953
timestamp 1679581782
transform 1 0 92064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_960
timestamp 1679581782
transform 1 0 92736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_967
timestamp 1679581782
transform 1 0 93408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_974
timestamp 1679581782
transform 1 0 94080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_981
timestamp 1679581782
transform 1 0 94752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_988
timestamp 1679581782
transform 1 0 95424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_995
timestamp 1679581782
transform 1 0 96096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1002
timestamp 1679581782
transform 1 0 96768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1009
timestamp 1679581782
transform 1 0 97440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1016
timestamp 1679581782
transform 1 0 98112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_1023
timestamp 1679577901
transform 1 0 98784 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_1027
timestamp 1677580104
transform 1 0 99168 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_7
timestamp 1679577901
transform 1 0 1248 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_42
timestamp 1677579658
transform 1 0 4608 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_56
timestamp 1677579658
transform 1 0 5952 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 8640 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_91
timestamp 1677580104
transform 1 0 9312 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_132
timestamp 1679581782
transform 1 0 13248 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_193
timestamp 1677580104
transform 1 0 19104 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_195
timestamp 1677579658
transform 1 0 19296 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_223
timestamp 1679577901
transform 1 0 21984 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_227
timestamp 1677579658
transform 1 0 22368 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 24096 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_267
timestamp 1677579658
transform 1 0 26208 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_299
timestamp 1677580104
transform 1 0 29280 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_301
timestamp 1677579658
transform 1 0 29472 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_306
timestamp 1679581782
transform 1 0 29952 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_313
timestamp 1677580104
transform 1 0 30624 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_315
timestamp 1677579658
transform 1 0 30816 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_362
timestamp 1677579658
transform 1 0 35328 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_385
timestamp 1677580104
transform 1 0 37536 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_387
timestamp 1677579658
transform 1 0 37728 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_407
timestamp 1677580104
transform 1 0 39648 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_472
timestamp 1677580104
transform 1 0 45888 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_482
timestamp 1677579658
transform 1 0 46848 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_506
timestamp 1679577901
transform 1 0 49152 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_510
timestamp 1677579658
transform 1 0 49536 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_515
timestamp 1679581782
transform 1 0 50016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_522
timestamp 1679581782
transform 1 0 50688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_529
timestamp 1679581782
transform 1 0 51360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_536
timestamp 1679581782
transform 1 0 52032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_543
timestamp 1679581782
transform 1 0 52704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_550
timestamp 1679581782
transform 1 0 53376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_557
timestamp 1679581782
transform 1 0 54048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_564
timestamp 1679581782
transform 1 0 54720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_571
timestamp 1679581782
transform 1 0 55392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_578
timestamp 1679581782
transform 1 0 56064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_585
timestamp 1679581782
transform 1 0 56736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_592
timestamp 1679581782
transform 1 0 57408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_599
timestamp 1679581782
transform 1 0 58080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_606
timestamp 1679581782
transform 1 0 58752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_613
timestamp 1679581782
transform 1 0 59424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_620
timestamp 1679581782
transform 1 0 60096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_627
timestamp 1679581782
transform 1 0 60768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_634
timestamp 1679581782
transform 1 0 61440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_641
timestamp 1679581782
transform 1 0 62112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_648
timestamp 1679581782
transform 1 0 62784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_655
timestamp 1679581782
transform 1 0 63456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_662
timestamp 1679581782
transform 1 0 64128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_669
timestamp 1679581782
transform 1 0 64800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_676
timestamp 1679581782
transform 1 0 65472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_683
timestamp 1679581782
transform 1 0 66144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_690
timestamp 1679581782
transform 1 0 66816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_697
timestamp 1679581782
transform 1 0 67488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_704
timestamp 1679581782
transform 1 0 68160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_711
timestamp 1679581782
transform 1 0 68832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_718
timestamp 1679581782
transform 1 0 69504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_725
timestamp 1679581782
transform 1 0 70176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_732
timestamp 1679581782
transform 1 0 70848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_739
timestamp 1679581782
transform 1 0 71520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_746
timestamp 1679581782
transform 1 0 72192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_753
timestamp 1679581782
transform 1 0 72864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_760
timestamp 1679581782
transform 1 0 73536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_767
timestamp 1679581782
transform 1 0 74208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_774
timestamp 1679581782
transform 1 0 74880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_781
timestamp 1679581782
transform 1 0 75552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_788
timestamp 1679581782
transform 1 0 76224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_795
timestamp 1679581782
transform 1 0 76896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_802
timestamp 1679581782
transform 1 0 77568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_809
timestamp 1679581782
transform 1 0 78240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_816
timestamp 1679581782
transform 1 0 78912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_823
timestamp 1679581782
transform 1 0 79584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_830
timestamp 1679581782
transform 1 0 80256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_837
timestamp 1679581782
transform 1 0 80928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_844
timestamp 1679581782
transform 1 0 81600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_851
timestamp 1679581782
transform 1 0 82272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_858
timestamp 1679581782
transform 1 0 82944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_865
timestamp 1679581782
transform 1 0 83616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_872
timestamp 1679581782
transform 1 0 84288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_879
timestamp 1679581782
transform 1 0 84960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_886
timestamp 1679581782
transform 1 0 85632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_893
timestamp 1679581782
transform 1 0 86304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_900
timestamp 1679581782
transform 1 0 86976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_907
timestamp 1679581782
transform 1 0 87648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_914
timestamp 1679581782
transform 1 0 88320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_921
timestamp 1679581782
transform 1 0 88992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_928
timestamp 1679581782
transform 1 0 89664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_935
timestamp 1679581782
transform 1 0 90336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_942
timestamp 1679581782
transform 1 0 91008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_949
timestamp 1679581782
transform 1 0 91680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_956
timestamp 1679581782
transform 1 0 92352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_963
timestamp 1679581782
transform 1 0 93024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_970
timestamp 1679581782
transform 1 0 93696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_977
timestamp 1679581782
transform 1 0 94368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_984
timestamp 1679581782
transform 1 0 95040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_991
timestamp 1679581782
transform 1 0 95712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_998
timestamp 1679581782
transform 1 0 96384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1005
timestamp 1679581782
transform 1 0 97056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1012
timestamp 1679581782
transform 1 0 97728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1019
timestamp 1679581782
transform 1 0 98400 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_1026
timestamp 1677580104
transform 1 0 99072 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_1028
timestamp 1677579658
transform 1 0 99264 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_4
timestamp 1677580104
transform 1 0 960 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_6
timestamp 1677579658
transform 1 0 1152 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_48
timestamp 1677580104
transform 1 0 5184 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_28_84
timestamp 1679577901
transform 1 0 8640 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_88
timestamp 1677580104
transform 1 0 9024 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_130
timestamp 1677580104
transform 1 0 13056 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_132
timestamp 1677579658
transform 1 0 13248 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_143
timestamp 1677580104
transform 1 0 14304 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_180
timestamp 1677580104
transform 1 0 17856 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_195
timestamp 1677580104
transform 1 0 19296 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_28_241
timestamp 1679577901
transform 1 0 23712 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_250
timestamp 1679581782
transform 1 0 24576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_257
timestamp 1679581782
transform 1 0 25248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_264
timestamp 1679581782
transform 1 0 25920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_271
timestamp 1679577901
transform 1 0 26592 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_275
timestamp 1677580104
transform 1 0 26976 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_281
timestamp 1679581782
transform 1 0 27552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_288
timestamp 1679581782
transform 1 0 28224 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_295
timestamp 1677580104
transform 1 0 28896 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_347
timestamp 1677580104
transform 1 0 33888 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_355
timestamp 1677579658
transform 1 0 34656 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_369
timestamp 1679581782
transform 1 0 36000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_376
timestamp 1679577901
transform 1 0 36672 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_380
timestamp 1677580104
transform 1 0 37056 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_409
timestamp 1677580104
transform 1 0 39840 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_496
timestamp 1677579658
transform 1 0 48192 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_533
timestamp 1679581782
transform 1 0 51744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_540
timestamp 1679581782
transform 1 0 52416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_547
timestamp 1679581782
transform 1 0 53088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_554
timestamp 1679581782
transform 1 0 53760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_561
timestamp 1679581782
transform 1 0 54432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_568
timestamp 1679581782
transform 1 0 55104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_575
timestamp 1679581782
transform 1 0 55776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_582
timestamp 1679581782
transform 1 0 56448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_589
timestamp 1679581782
transform 1 0 57120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_596
timestamp 1679581782
transform 1 0 57792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_603
timestamp 1679581782
transform 1 0 58464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_610
timestamp 1679581782
transform 1 0 59136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_617
timestamp 1679581782
transform 1 0 59808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_624
timestamp 1679581782
transform 1 0 60480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_631
timestamp 1679581782
transform 1 0 61152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_638
timestamp 1679581782
transform 1 0 61824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_645
timestamp 1679581782
transform 1 0 62496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_652
timestamp 1679581782
transform 1 0 63168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_659
timestamp 1679581782
transform 1 0 63840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_666
timestamp 1679581782
transform 1 0 64512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_673
timestamp 1679581782
transform 1 0 65184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_680
timestamp 1679581782
transform 1 0 65856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_687
timestamp 1679581782
transform 1 0 66528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_694
timestamp 1679581782
transform 1 0 67200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_701
timestamp 1679581782
transform 1 0 67872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_708
timestamp 1679581782
transform 1 0 68544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_715
timestamp 1679581782
transform 1 0 69216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_722
timestamp 1679581782
transform 1 0 69888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_729
timestamp 1679581782
transform 1 0 70560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_736
timestamp 1679581782
transform 1 0 71232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_743
timestamp 1679581782
transform 1 0 71904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_750
timestamp 1679581782
transform 1 0 72576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_757
timestamp 1679581782
transform 1 0 73248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_764
timestamp 1679581782
transform 1 0 73920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_771
timestamp 1679581782
transform 1 0 74592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_778
timestamp 1679581782
transform 1 0 75264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_785
timestamp 1679581782
transform 1 0 75936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_792
timestamp 1679581782
transform 1 0 76608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_799
timestamp 1679581782
transform 1 0 77280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_806
timestamp 1679581782
transform 1 0 77952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_813
timestamp 1679581782
transform 1 0 78624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_820
timestamp 1679581782
transform 1 0 79296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_827
timestamp 1679581782
transform 1 0 79968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_834
timestamp 1679581782
transform 1 0 80640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_841
timestamp 1679581782
transform 1 0 81312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_848
timestamp 1679581782
transform 1 0 81984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_855
timestamp 1679581782
transform 1 0 82656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_862
timestamp 1679581782
transform 1 0 83328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_869
timestamp 1679581782
transform 1 0 84000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_876
timestamp 1679581782
transform 1 0 84672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_883
timestamp 1679581782
transform 1 0 85344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_890
timestamp 1679581782
transform 1 0 86016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_897
timestamp 1679581782
transform 1 0 86688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_904
timestamp 1679581782
transform 1 0 87360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_911
timestamp 1679581782
transform 1 0 88032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_918
timestamp 1679581782
transform 1 0 88704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_925
timestamp 1679581782
transform 1 0 89376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_932
timestamp 1679581782
transform 1 0 90048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_939
timestamp 1679581782
transform 1 0 90720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_946
timestamp 1679581782
transform 1 0 91392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_953
timestamp 1679581782
transform 1 0 92064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_960
timestamp 1679581782
transform 1 0 92736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_967
timestamp 1679581782
transform 1 0 93408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_974
timestamp 1679581782
transform 1 0 94080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_981
timestamp 1679581782
transform 1 0 94752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_988
timestamp 1679581782
transform 1 0 95424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_995
timestamp 1679581782
transform 1 0 96096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1002
timestamp 1679581782
transform 1 0 96768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1009
timestamp 1679581782
transform 1 0 97440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1016
timestamp 1679581782
transform 1 0 98112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_1023
timestamp 1679577901
transform 1 0 98784 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_1027
timestamp 1677580104
transform 1 0 99168 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_4
timestamp 1679577901
transform 1 0 960 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_35
timestamp 1677579658
transform 1 0 3936 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_59
timestamp 1677580104
transform 1 0 6240 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_79
timestamp 1679577901
transform 1 0 8160 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_83
timestamp 1677579658
transform 1 0 8544 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_116
timestamp 1677579658
transform 1 0 11712 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_139
timestamp 1677579658
transform 1 0 13920 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_153
timestamp 1677579658
transform 1 0 15264 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_163
timestamp 1677579658
transform 1 0 16224 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_173
timestamp 1677580104
transform 1 0 17184 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_212
timestamp 1679581782
transform 1 0 20928 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_260
timestamp 1677580104
transform 1 0 25536 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_290
timestamp 1677580104
transform 1 0 28416 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_292
timestamp 1677579658
transform 1 0 28608 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_316
timestamp 1677579658
transform 1 0 30912 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_384
timestamp 1677580104
transform 1 0 37440 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_386
timestamp 1677579658
transform 1 0 37632 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_391
timestamp 1679577901
transform 1 0 38112 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_398
timestamp 1677579658
transform 1 0 38784 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_416
timestamp 1677579658
transform 1 0 40512 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_444
timestamp 1677579658
transform 1 0 43200 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_483
timestamp 1677580104
transform 1 0 46944 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_490
timestamp 1677579658
transform 1 0 47616 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_518
timestamp 1679581782
transform 1 0 50304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_525
timestamp 1679581782
transform 1 0 50976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_532
timestamp 1679581782
transform 1 0 51648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_539
timestamp 1679581782
transform 1 0 52320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_546
timestamp 1679581782
transform 1 0 52992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_553
timestamp 1679581782
transform 1 0 53664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_560
timestamp 1679581782
transform 1 0 54336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_567
timestamp 1679581782
transform 1 0 55008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_574
timestamp 1679581782
transform 1 0 55680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_581
timestamp 1679581782
transform 1 0 56352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_588
timestamp 1679581782
transform 1 0 57024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_595
timestamp 1679581782
transform 1 0 57696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_602
timestamp 1679581782
transform 1 0 58368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_609
timestamp 1679581782
transform 1 0 59040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_616
timestamp 1679581782
transform 1 0 59712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_623
timestamp 1679581782
transform 1 0 60384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_630
timestamp 1679581782
transform 1 0 61056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_637
timestamp 1679581782
transform 1 0 61728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_644
timestamp 1679581782
transform 1 0 62400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_651
timestamp 1679581782
transform 1 0 63072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_658
timestamp 1679581782
transform 1 0 63744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_665
timestamp 1679581782
transform 1 0 64416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_672
timestamp 1679581782
transform 1 0 65088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_679
timestamp 1679581782
transform 1 0 65760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_686
timestamp 1679581782
transform 1 0 66432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_693
timestamp 1679581782
transform 1 0 67104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_700
timestamp 1679581782
transform 1 0 67776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_707
timestamp 1679581782
transform 1 0 68448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_714
timestamp 1679581782
transform 1 0 69120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_721
timestamp 1679581782
transform 1 0 69792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_728
timestamp 1679581782
transform 1 0 70464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_735
timestamp 1679581782
transform 1 0 71136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_742
timestamp 1679581782
transform 1 0 71808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_749
timestamp 1679581782
transform 1 0 72480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_756
timestamp 1679581782
transform 1 0 73152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_763
timestamp 1679581782
transform 1 0 73824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_770
timestamp 1679581782
transform 1 0 74496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_777
timestamp 1679581782
transform 1 0 75168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_784
timestamp 1679581782
transform 1 0 75840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_791
timestamp 1679581782
transform 1 0 76512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_798
timestamp 1679581782
transform 1 0 77184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_805
timestamp 1679581782
transform 1 0 77856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_812
timestamp 1679581782
transform 1 0 78528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_819
timestamp 1679581782
transform 1 0 79200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_826
timestamp 1679581782
transform 1 0 79872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_833
timestamp 1679581782
transform 1 0 80544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_840
timestamp 1679581782
transform 1 0 81216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_847
timestamp 1679581782
transform 1 0 81888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_854
timestamp 1679581782
transform 1 0 82560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_861
timestamp 1679581782
transform 1 0 83232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_868
timestamp 1679581782
transform 1 0 83904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_875
timestamp 1679581782
transform 1 0 84576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_882
timestamp 1679581782
transform 1 0 85248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_889
timestamp 1679581782
transform 1 0 85920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_896
timestamp 1679581782
transform 1 0 86592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_903
timestamp 1679581782
transform 1 0 87264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_910
timestamp 1679581782
transform 1 0 87936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_917
timestamp 1679581782
transform 1 0 88608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_924
timestamp 1679581782
transform 1 0 89280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_931
timestamp 1679581782
transform 1 0 89952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_938
timestamp 1679581782
transform 1 0 90624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_945
timestamp 1679581782
transform 1 0 91296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_952
timestamp 1679581782
transform 1 0 91968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_959
timestamp 1679581782
transform 1 0 92640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_966
timestamp 1679581782
transform 1 0 93312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_973
timestamp 1679581782
transform 1 0 93984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_980
timestamp 1679581782
transform 1 0 94656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_987
timestamp 1679581782
transform 1 0 95328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_994
timestamp 1679581782
transform 1 0 96000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1001
timestamp 1679581782
transform 1 0 96672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1008
timestamp 1679581782
transform 1 0 97344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1015
timestamp 1679581782
transform 1 0 98016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1022
timestamp 1679581782
transform 1 0 98688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_0
timestamp 1679577901
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_4
timestamp 1677579658
transform 1 0 960 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_40
timestamp 1677579658
transform 1 0 4416 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_46
timestamp 1677579658
transform 1 0 4992 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_114
timestamp 1677580104
transform 1 0 11520 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_116
timestamp 1677579658
transform 1 0 11712 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_130
timestamp 1679581782
transform 1 0 13056 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_169
timestamp 1677579658
transform 1 0 16800 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_198
timestamp 1679581782
transform 1 0 19584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_205
timestamp 1679577901
transform 1 0 20256 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_222
timestamp 1679581782
transform 1 0 21888 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_229
timestamp 1677580104
transform 1 0 22560 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_244
timestamp 1677579658
transform 1 0 24000 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_276
timestamp 1677579658
transform 1 0 27072 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_335
timestamp 1677580104
transform 1 0 32736 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_404
timestamp 1679577901
transform 1 0 39360 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_408
timestamp 1677580104
transform 1 0 39744 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_417
timestamp 1677579658
transform 1 0 40608 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_435
timestamp 1677580104
transform 1 0 42336 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_450
timestamp 1679581782
transform 1 0 43776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_457
timestamp 1679577901
transform 1 0 44448 0 1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_30_465
timestamp 1679577901
transform 1 0 45216 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_507
timestamp 1677579658
transform 1 0 49248 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_525
timestamp 1679581782
transform 1 0 50976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_532
timestamp 1679581782
transform 1 0 51648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679581782
transform 1 0 52320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_546
timestamp 1679581782
transform 1 0 52992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_553
timestamp 1679581782
transform 1 0 53664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_560
timestamp 1679581782
transform 1 0 54336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_567
timestamp 1679581782
transform 1 0 55008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_574
timestamp 1679581782
transform 1 0 55680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_581
timestamp 1679581782
transform 1 0 56352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_588
timestamp 1679581782
transform 1 0 57024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_595
timestamp 1679581782
transform 1 0 57696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_602
timestamp 1679581782
transform 1 0 58368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_609
timestamp 1679581782
transform 1 0 59040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_616
timestamp 1679581782
transform 1 0 59712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_623
timestamp 1679581782
transform 1 0 60384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_630
timestamp 1679581782
transform 1 0 61056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_637
timestamp 1679581782
transform 1 0 61728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_644
timestamp 1679581782
transform 1 0 62400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_651
timestamp 1679581782
transform 1 0 63072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_658
timestamp 1679581782
transform 1 0 63744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_665
timestamp 1679581782
transform 1 0 64416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_672
timestamp 1679581782
transform 1 0 65088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_679
timestamp 1679581782
transform 1 0 65760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_686
timestamp 1679581782
transform 1 0 66432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_693
timestamp 1679581782
transform 1 0 67104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_700
timestamp 1679581782
transform 1 0 67776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_707
timestamp 1679581782
transform 1 0 68448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_714
timestamp 1679581782
transform 1 0 69120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_721
timestamp 1679581782
transform 1 0 69792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_728
timestamp 1679581782
transform 1 0 70464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_735
timestamp 1679581782
transform 1 0 71136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_742
timestamp 1679581782
transform 1 0 71808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_749
timestamp 1679581782
transform 1 0 72480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_756
timestamp 1679581782
transform 1 0 73152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_763
timestamp 1679581782
transform 1 0 73824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_770
timestamp 1679581782
transform 1 0 74496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_777
timestamp 1679581782
transform 1 0 75168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_784
timestamp 1679581782
transform 1 0 75840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_791
timestamp 1679581782
transform 1 0 76512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_798
timestamp 1679581782
transform 1 0 77184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_805
timestamp 1679581782
transform 1 0 77856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_812
timestamp 1679581782
transform 1 0 78528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_819
timestamp 1679581782
transform 1 0 79200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_826
timestamp 1679581782
transform 1 0 79872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_833
timestamp 1679581782
transform 1 0 80544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_840
timestamp 1679581782
transform 1 0 81216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_847
timestamp 1679581782
transform 1 0 81888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_854
timestamp 1679581782
transform 1 0 82560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_861
timestamp 1679581782
transform 1 0 83232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_868
timestamp 1679581782
transform 1 0 83904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_875
timestamp 1679581782
transform 1 0 84576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_882
timestamp 1679581782
transform 1 0 85248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_889
timestamp 1679581782
transform 1 0 85920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_896
timestamp 1679581782
transform 1 0 86592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_903
timestamp 1679581782
transform 1 0 87264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_910
timestamp 1679581782
transform 1 0 87936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_917
timestamp 1679581782
transform 1 0 88608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_924
timestamp 1679581782
transform 1 0 89280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_931
timestamp 1679581782
transform 1 0 89952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_938
timestamp 1679581782
transform 1 0 90624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_945
timestamp 1679581782
transform 1 0 91296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_952
timestamp 1679581782
transform 1 0 91968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_959
timestamp 1679581782
transform 1 0 92640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_966
timestamp 1679581782
transform 1 0 93312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_973
timestamp 1679581782
transform 1 0 93984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_980
timestamp 1679581782
transform 1 0 94656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_987
timestamp 1679581782
transform 1 0 95328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_994
timestamp 1679581782
transform 1 0 96000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1001
timestamp 1679581782
transform 1 0 96672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1008
timestamp 1679581782
transform 1 0 97344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1015
timestamp 1679581782
transform 1 0 98016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1022
timestamp 1679581782
transform 1 0 98688 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_0
timestamp 1677580104
transform 1 0 576 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_32
timestamp 1677580104
transform 1 0 3648 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_48
timestamp 1677580104
transform 1 0 5184 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_82
timestamp 1677579658
transform 1 0 8448 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_146
timestamp 1677579658
transform 1 0 14592 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_151
timestamp 1677580104
transform 1 0 15072 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_153
timestamp 1677579658
transform 1 0 15264 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_164
timestamp 1679577901
transform 1 0 16320 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_168
timestamp 1677580104
transform 1 0 16704 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_198
timestamp 1679581782
transform 1 0 19584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_205
timestamp 1679577901
transform 1 0 20256 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_209
timestamp 1677580104
transform 1 0 20640 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_237
timestamp 1677580104
transform 1 0 23328 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_271
timestamp 1677580104
transform 1 0 26592 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_273
timestamp 1677579658
transform 1 0 26784 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_301
timestamp 1677579658
transform 1 0 29472 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_311
timestamp 1677580104
transform 1 0 30432 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_313
timestamp 1677579658
transform 1 0 30624 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_330
timestamp 1677580104
transform 1 0 32256 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679581782
transform 1 0 36192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679581782
transform 1 0 36864 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_419
timestamp 1677579658
transform 1 0 40800 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_457
timestamp 1677580104
transform 1 0 44448 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_472
timestamp 1677580104
transform 1 0 45888 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_474
timestamp 1677579658
transform 1 0 46080 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_534
timestamp 1679581782
transform 1 0 51840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_541
timestamp 1679581782
transform 1 0 52512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_548
timestamp 1679581782
transform 1 0 53184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_555
timestamp 1679581782
transform 1 0 53856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_562
timestamp 1679581782
transform 1 0 54528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_569
timestamp 1679581782
transform 1 0 55200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_576
timestamp 1679581782
transform 1 0 55872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_583
timestamp 1679581782
transform 1 0 56544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_590
timestamp 1679581782
transform 1 0 57216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_597
timestamp 1679581782
transform 1 0 57888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_604
timestamp 1679581782
transform 1 0 58560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_611
timestamp 1679581782
transform 1 0 59232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_618
timestamp 1679581782
transform 1 0 59904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_625
timestamp 1679581782
transform 1 0 60576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_632
timestamp 1679581782
transform 1 0 61248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_639
timestamp 1679581782
transform 1 0 61920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_646
timestamp 1679581782
transform 1 0 62592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_653
timestamp 1679581782
transform 1 0 63264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_660
timestamp 1679581782
transform 1 0 63936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_667
timestamp 1679581782
transform 1 0 64608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_674
timestamp 1679581782
transform 1 0 65280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_681
timestamp 1679581782
transform 1 0 65952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_688
timestamp 1679581782
transform 1 0 66624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_695
timestamp 1679581782
transform 1 0 67296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_702
timestamp 1679581782
transform 1 0 67968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_709
timestamp 1679581782
transform 1 0 68640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_716
timestamp 1679581782
transform 1 0 69312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_723
timestamp 1679581782
transform 1 0 69984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_730
timestamp 1679581782
transform 1 0 70656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_737
timestamp 1679581782
transform 1 0 71328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_744
timestamp 1679581782
transform 1 0 72000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_751
timestamp 1679581782
transform 1 0 72672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_758
timestamp 1679581782
transform 1 0 73344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_765
timestamp 1679581782
transform 1 0 74016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_772
timestamp 1679581782
transform 1 0 74688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_779
timestamp 1679581782
transform 1 0 75360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_786
timestamp 1679581782
transform 1 0 76032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_793
timestamp 1679581782
transform 1 0 76704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_800
timestamp 1679581782
transform 1 0 77376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_807
timestamp 1679581782
transform 1 0 78048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_814
timestamp 1679581782
transform 1 0 78720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_821
timestamp 1679581782
transform 1 0 79392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_828
timestamp 1679581782
transform 1 0 80064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_835
timestamp 1679581782
transform 1 0 80736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_842
timestamp 1679581782
transform 1 0 81408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_849
timestamp 1679581782
transform 1 0 82080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_856
timestamp 1679581782
transform 1 0 82752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_863
timestamp 1679581782
transform 1 0 83424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_870
timestamp 1679581782
transform 1 0 84096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_877
timestamp 1679581782
transform 1 0 84768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_884
timestamp 1679581782
transform 1 0 85440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_891
timestamp 1679581782
transform 1 0 86112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_898
timestamp 1679581782
transform 1 0 86784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_905
timestamp 1679581782
transform 1 0 87456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_912
timestamp 1679581782
transform 1 0 88128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_919
timestamp 1679581782
transform 1 0 88800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_926
timestamp 1679581782
transform 1 0 89472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_933
timestamp 1679581782
transform 1 0 90144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_940
timestamp 1679581782
transform 1 0 90816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_947
timestamp 1679581782
transform 1 0 91488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_954
timestamp 1679581782
transform 1 0 92160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_961
timestamp 1679581782
transform 1 0 92832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_968
timestamp 1679581782
transform 1 0 93504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_975
timestamp 1679581782
transform 1 0 94176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_982
timestamp 1679581782
transform 1 0 94848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_989
timestamp 1679581782
transform 1 0 95520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_996
timestamp 1679581782
transform 1 0 96192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1003
timestamp 1679581782
transform 1 0 96864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1010
timestamp 1679581782
transform 1 0 97536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1017
timestamp 1679581782
transform 1 0 98208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_1024
timestamp 1679577901
transform 1 0 98880 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_1028
timestamp 1677579658
transform 1 0 99264 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_0
timestamp 1679577901
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_40
timestamp 1677579658
transform 1 0 4416 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_61
timestamp 1677580104
transform 1 0 6432 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_101
timestamp 1677580104
transform 1 0 10272 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_122
timestamp 1677580104
transform 1 0 12288 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_128
timestamp 1677580104
transform 1 0 12864 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_147
timestamp 1677580104
transform 1 0 14688 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_154
timestamp 1679581782
transform 1 0 15360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_166
timestamp 1679581782
transform 1 0 16512 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_173
timestamp 1677580104
transform 1 0 17184 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_175
timestamp 1677579658
transform 1 0 17376 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_249
timestamp 1677579658
transform 1 0 24480 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_255
timestamp 1679581782
transform 1 0 25056 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_262
timestamp 1677580104
transform 1 0 25728 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_264
timestamp 1677579658
transform 1 0 25920 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_290
timestamp 1677580104
transform 1 0 28416 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_292
timestamp 1677579658
transform 1 0 28608 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_306
timestamp 1677579658
transform 1 0 29952 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_320
timestamp 1679577901
transform 1 0 31296 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_369
timestamp 1677579658
transform 1 0 36000 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_394
timestamp 1679577901
transform 1 0 38400 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_398
timestamp 1677579658
transform 1 0 38784 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_412
timestamp 1677579658
transform 1 0 40128 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_452
timestamp 1679577901
transform 1 0 43968 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_456
timestamp 1677579658
transform 1 0 44352 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_462
timestamp 1677579658
transform 1 0 44928 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_535
timestamp 1679581782
transform 1 0 51936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_542
timestamp 1679581782
transform 1 0 52608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_549
timestamp 1679581782
transform 1 0 53280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_556
timestamp 1679581782
transform 1 0 53952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_563
timestamp 1679581782
transform 1 0 54624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_570
timestamp 1679581782
transform 1 0 55296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_577
timestamp 1679581782
transform 1 0 55968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_584
timestamp 1679581782
transform 1 0 56640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_591
timestamp 1679581782
transform 1 0 57312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_598
timestamp 1679581782
transform 1 0 57984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_605
timestamp 1679581782
transform 1 0 58656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_612
timestamp 1679581782
transform 1 0 59328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_619
timestamp 1679581782
transform 1 0 60000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_626
timestamp 1679581782
transform 1 0 60672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_633
timestamp 1679581782
transform 1 0 61344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_640
timestamp 1679581782
transform 1 0 62016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_647
timestamp 1679581782
transform 1 0 62688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_654
timestamp 1679581782
transform 1 0 63360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_661
timestamp 1679581782
transform 1 0 64032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_668
timestamp 1679581782
transform 1 0 64704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_675
timestamp 1679581782
transform 1 0 65376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_682
timestamp 1679581782
transform 1 0 66048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_689
timestamp 1679581782
transform 1 0 66720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_696
timestamp 1679581782
transform 1 0 67392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_703
timestamp 1679581782
transform 1 0 68064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_710
timestamp 1679581782
transform 1 0 68736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_717
timestamp 1679581782
transform 1 0 69408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_724
timestamp 1679581782
transform 1 0 70080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_731
timestamp 1679581782
transform 1 0 70752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_738
timestamp 1679581782
transform 1 0 71424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_745
timestamp 1679581782
transform 1 0 72096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_752
timestamp 1679581782
transform 1 0 72768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_759
timestamp 1679581782
transform 1 0 73440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_766
timestamp 1679581782
transform 1 0 74112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_773
timestamp 1679581782
transform 1 0 74784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_780
timestamp 1679581782
transform 1 0 75456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_787
timestamp 1679581782
transform 1 0 76128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_794
timestamp 1679581782
transform 1 0 76800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_801
timestamp 1679581782
transform 1 0 77472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_808
timestamp 1679581782
transform 1 0 78144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_815
timestamp 1679581782
transform 1 0 78816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_822
timestamp 1679581782
transform 1 0 79488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_829
timestamp 1679581782
transform 1 0 80160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_836
timestamp 1679581782
transform 1 0 80832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_843
timestamp 1679581782
transform 1 0 81504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_850
timestamp 1679581782
transform 1 0 82176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_857
timestamp 1679581782
transform 1 0 82848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_864
timestamp 1679581782
transform 1 0 83520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_871
timestamp 1679581782
transform 1 0 84192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_878
timestamp 1679581782
transform 1 0 84864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_885
timestamp 1679581782
transform 1 0 85536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_892
timestamp 1679581782
transform 1 0 86208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_899
timestamp 1679581782
transform 1 0 86880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_906
timestamp 1679581782
transform 1 0 87552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_913
timestamp 1679581782
transform 1 0 88224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_920
timestamp 1679581782
transform 1 0 88896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_927
timestamp 1679581782
transform 1 0 89568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_934
timestamp 1679581782
transform 1 0 90240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_941
timestamp 1679581782
transform 1 0 90912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_948
timestamp 1679581782
transform 1 0 91584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_955
timestamp 1679581782
transform 1 0 92256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_962
timestamp 1679581782
transform 1 0 92928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_969
timestamp 1679581782
transform 1 0 93600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_976
timestamp 1679581782
transform 1 0 94272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_983
timestamp 1679581782
transform 1 0 94944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_990
timestamp 1679581782
transform 1 0 95616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_997
timestamp 1679581782
transform 1 0 96288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1004
timestamp 1679581782
transform 1 0 96960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1011
timestamp 1679581782
transform 1 0 97632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1018
timestamp 1679581782
transform 1 0 98304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_1025
timestamp 1679577901
transform 1 0 98976 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_38
timestamp 1677579658
transform 1 0 4224 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_51
timestamp 1677580104
transform 1 0 5472 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_63
timestamp 1677580104
transform 1 0 6624 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_83
timestamp 1677580104
transform 1 0 8544 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_125
timestamp 1679581782
transform 1 0 12576 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_132
timestamp 1677580104
transform 1 0 13248 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_134
timestamp 1677579658
transform 1 0 13440 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_150
timestamp 1677580104
transform 1 0 14976 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_156
timestamp 1677579658
transform 1 0 15552 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_165
timestamp 1677579658
transform 1 0 16416 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_190
timestamp 1677579658
transform 1 0 18816 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_219
timestamp 1677580104
transform 1 0 21600 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_221
timestamp 1677579658
transform 1 0 21792 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_226
timestamp 1679581782
transform 1 0 22272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_233
timestamp 1679577901
transform 1 0 22944 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_237
timestamp 1677580104
transform 1 0 23328 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_266
timestamp 1677580104
transform 1 0 26112 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_294
timestamp 1677580104
transform 1 0 28800 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_301
timestamp 1677579658
transform 1 0 29472 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_307
timestamp 1677580104
transform 1 0 30048 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_316
timestamp 1679577901
transform 1 0 30912 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_365
timestamp 1677580104
transform 1 0 35616 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_367
timestamp 1677579658
transform 1 0 35808 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_385
timestamp 1677580104
transform 1 0 37536 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_402
timestamp 1679581782
transform 1 0 39168 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_409
timestamp 1677580104
transform 1 0 39840 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_420
timestamp 1677580104
transform 1 0 40896 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_437
timestamp 1677580104
transform 1 0 42528 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_461
timestamp 1677579658
transform 1 0 44832 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_489
timestamp 1677580104
transform 1 0 47520 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_514
timestamp 1677579658
transform 1 0 49920 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_533
timestamp 1679581782
transform 1 0 51744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_540
timestamp 1679581782
transform 1 0 52416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_547
timestamp 1679581782
transform 1 0 53088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_554
timestamp 1679581782
transform 1 0 53760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_561
timestamp 1679581782
transform 1 0 54432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_568
timestamp 1679581782
transform 1 0 55104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_575
timestamp 1679581782
transform 1 0 55776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_582
timestamp 1679581782
transform 1 0 56448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_589
timestamp 1679581782
transform 1 0 57120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_596
timestamp 1679581782
transform 1 0 57792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_603
timestamp 1679581782
transform 1 0 58464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_610
timestamp 1679581782
transform 1 0 59136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_617
timestamp 1679581782
transform 1 0 59808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_624
timestamp 1679581782
transform 1 0 60480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_631
timestamp 1679581782
transform 1 0 61152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_638
timestamp 1679581782
transform 1 0 61824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_645
timestamp 1679581782
transform 1 0 62496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_652
timestamp 1679581782
transform 1 0 63168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_659
timestamp 1679581782
transform 1 0 63840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_666
timestamp 1679581782
transform 1 0 64512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_673
timestamp 1679581782
transform 1 0 65184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_680
timestamp 1679581782
transform 1 0 65856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_687
timestamp 1679581782
transform 1 0 66528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_694
timestamp 1679581782
transform 1 0 67200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_701
timestamp 1679581782
transform 1 0 67872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_708
timestamp 1679581782
transform 1 0 68544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_715
timestamp 1679581782
transform 1 0 69216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_722
timestamp 1679581782
transform 1 0 69888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_729
timestamp 1679581782
transform 1 0 70560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_736
timestamp 1679581782
transform 1 0 71232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_743
timestamp 1679581782
transform 1 0 71904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_750
timestamp 1679581782
transform 1 0 72576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_757
timestamp 1679581782
transform 1 0 73248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_764
timestamp 1679581782
transform 1 0 73920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_771
timestamp 1679581782
transform 1 0 74592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_778
timestamp 1679581782
transform 1 0 75264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_785
timestamp 1679581782
transform 1 0 75936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_792
timestamp 1679581782
transform 1 0 76608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_799
timestamp 1679581782
transform 1 0 77280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_806
timestamp 1679581782
transform 1 0 77952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_813
timestamp 1679581782
transform 1 0 78624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_820
timestamp 1679581782
transform 1 0 79296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_827
timestamp 1679581782
transform 1 0 79968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_834
timestamp 1679581782
transform 1 0 80640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_841
timestamp 1679581782
transform 1 0 81312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_848
timestamp 1679581782
transform 1 0 81984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_855
timestamp 1679581782
transform 1 0 82656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_862
timestamp 1679581782
transform 1 0 83328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_869
timestamp 1679581782
transform 1 0 84000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_876
timestamp 1679581782
transform 1 0 84672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_883
timestamp 1679581782
transform 1 0 85344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_890
timestamp 1679581782
transform 1 0 86016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_897
timestamp 1679581782
transform 1 0 86688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_904
timestamp 1679581782
transform 1 0 87360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_911
timestamp 1679581782
transform 1 0 88032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_918
timestamp 1679581782
transform 1 0 88704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_925
timestamp 1679581782
transform 1 0 89376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_932
timestamp 1679581782
transform 1 0 90048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_939
timestamp 1679581782
transform 1 0 90720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_946
timestamp 1679581782
transform 1 0 91392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_953
timestamp 1679581782
transform 1 0 92064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_960
timestamp 1679581782
transform 1 0 92736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_967
timestamp 1679581782
transform 1 0 93408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_974
timestamp 1679581782
transform 1 0 94080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_981
timestamp 1679581782
transform 1 0 94752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_988
timestamp 1679581782
transform 1 0 95424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_995
timestamp 1679581782
transform 1 0 96096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1002
timestamp 1679581782
transform 1 0 96768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1009
timestamp 1679581782
transform 1 0 97440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1016
timestamp 1679581782
transform 1 0 98112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_1023
timestamp 1679577901
transform 1 0 98784 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_1027
timestamp 1677580104
transform 1 0 99168 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_14
timestamp 1677580104
transform 1 0 1920 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_20
timestamp 1677580104
transform 1 0 2496 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_38
timestamp 1677579658
transform 1 0 4224 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_84
timestamp 1677580104
transform 1 0 8640 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_118
timestamp 1679577901
transform 1 0 11904 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_122
timestamp 1677579658
transform 1 0 12288 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_158
timestamp 1677580104
transform 1 0 15744 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_174
timestamp 1679577901
transform 1 0 17280 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_186
timestamp 1677579658
transform 1 0 18432 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_206
timestamp 1677579658
transform 1 0 20352 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_234
timestamp 1677579658
transform 1 0 23040 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_257
timestamp 1677579658
transform 1 0 25248 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_272
timestamp 1677579658
transform 1 0 26688 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_304
timestamp 1677579658
transform 1 0 29760 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_309
timestamp 1677580104
transform 1 0 30240 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_321
timestamp 1679577901
transform 1 0 31392 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_352
timestamp 1677580104
transform 1 0 34368 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_359
timestamp 1677580104
transform 1 0 35040 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_368
timestamp 1679581782
transform 1 0 35904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_375
timestamp 1679577901
transform 1 0 36576 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_379
timestamp 1677580104
transform 1 0 36960 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_409
timestamp 1677579658
transform 1 0 39840 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_417
timestamp 1677580104
transform 1 0 40608 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_419
timestamp 1677579658
transform 1 0 40800 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_433
timestamp 1679577901
transform 1 0 42144 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_437
timestamp 1677579658
transform 1 0 42528 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_483
timestamp 1677580104
transform 1 0 46944 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_534
timestamp 1679581782
transform 1 0 51840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_541
timestamp 1679581782
transform 1 0 52512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_548
timestamp 1679581782
transform 1 0 53184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_555
timestamp 1679581782
transform 1 0 53856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_562
timestamp 1679581782
transform 1 0 54528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_569
timestamp 1679581782
transform 1 0 55200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_576
timestamp 1679581782
transform 1 0 55872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_583
timestamp 1679581782
transform 1 0 56544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_590
timestamp 1679581782
transform 1 0 57216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_597
timestamp 1679581782
transform 1 0 57888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_604
timestamp 1679581782
transform 1 0 58560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_611
timestamp 1679581782
transform 1 0 59232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_618
timestamp 1679581782
transform 1 0 59904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_625
timestamp 1679581782
transform 1 0 60576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_632
timestamp 1679581782
transform 1 0 61248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_639
timestamp 1679581782
transform 1 0 61920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_646
timestamp 1679581782
transform 1 0 62592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_653
timestamp 1679581782
transform 1 0 63264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_660
timestamp 1679581782
transform 1 0 63936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_667
timestamp 1679581782
transform 1 0 64608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_674
timestamp 1679581782
transform 1 0 65280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_681
timestamp 1679581782
transform 1 0 65952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_688
timestamp 1679581782
transform 1 0 66624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_695
timestamp 1679581782
transform 1 0 67296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_702
timestamp 1679581782
transform 1 0 67968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_709
timestamp 1679581782
transform 1 0 68640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_716
timestamp 1679581782
transform 1 0 69312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_723
timestamp 1679581782
transform 1 0 69984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_730
timestamp 1679581782
transform 1 0 70656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_737
timestamp 1679581782
transform 1 0 71328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_744
timestamp 1679581782
transform 1 0 72000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_751
timestamp 1679581782
transform 1 0 72672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_758
timestamp 1679581782
transform 1 0 73344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_765
timestamp 1679581782
transform 1 0 74016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_772
timestamp 1679581782
transform 1 0 74688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_779
timestamp 1679581782
transform 1 0 75360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_786
timestamp 1679581782
transform 1 0 76032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_793
timestamp 1679581782
transform 1 0 76704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_800
timestamp 1679581782
transform 1 0 77376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_807
timestamp 1679581782
transform 1 0 78048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_814
timestamp 1679581782
transform 1 0 78720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_821
timestamp 1679581782
transform 1 0 79392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_828
timestamp 1679581782
transform 1 0 80064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_835
timestamp 1679581782
transform 1 0 80736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_842
timestamp 1679581782
transform 1 0 81408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_849
timestamp 1679581782
transform 1 0 82080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_856
timestamp 1679581782
transform 1 0 82752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_863
timestamp 1679581782
transform 1 0 83424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_870
timestamp 1679581782
transform 1 0 84096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_877
timestamp 1679581782
transform 1 0 84768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_884
timestamp 1679581782
transform 1 0 85440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_891
timestamp 1679581782
transform 1 0 86112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_898
timestamp 1679581782
transform 1 0 86784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_905
timestamp 1679581782
transform 1 0 87456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_912
timestamp 1679581782
transform 1 0 88128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_919
timestamp 1679581782
transform 1 0 88800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_926
timestamp 1679581782
transform 1 0 89472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_933
timestamp 1679581782
transform 1 0 90144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_940
timestamp 1679581782
transform 1 0 90816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_947
timestamp 1679581782
transform 1 0 91488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_954
timestamp 1679581782
transform 1 0 92160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_961
timestamp 1679581782
transform 1 0 92832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_968
timestamp 1679581782
transform 1 0 93504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_975
timestamp 1679581782
transform 1 0 94176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_982
timestamp 1679581782
transform 1 0 94848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_989
timestamp 1679581782
transform 1 0 95520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_996
timestamp 1679581782
transform 1 0 96192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1003
timestamp 1679581782
transform 1 0 96864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1010
timestamp 1679581782
transform 1 0 97536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1017
timestamp 1679581782
transform 1 0 98208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_1024
timestamp 1679577901
transform 1 0 98880 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_1028
timestamp 1677579658
transform 1 0 99264 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_0
timestamp 1679577901
transform 1 0 576 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_4
timestamp 1677580104
transform 1 0 960 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_160
timestamp 1679577901
transform 1 0 15936 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_164
timestamp 1677579658
transform 1 0 16320 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_169
timestamp 1679577901
transform 1 0 16800 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_173
timestamp 1677579658
transform 1 0 17184 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_194
timestamp 1677580104
transform 1 0 19200 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_247
timestamp 1679577901
transform 1 0 24288 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_269
timestamp 1679581782
transform 1 0 26400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_276
timestamp 1679581782
transform 1 0 27072 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_288
timestamp 1677580104
transform 1 0 28224 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_298
timestamp 1679577901
transform 1 0 29184 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_302
timestamp 1677579658
transform 1 0 29568 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_339
timestamp 1677579658
transform 1 0 33120 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_343
timestamp 1677579658
transform 1 0 33504 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_376
timestamp 1677580104
transform 1 0 36672 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_435
timestamp 1679577901
transform 1 0 42336 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_439
timestamp 1677579658
transform 1 0 42720 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_528
timestamp 1679581782
transform 1 0 51264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_535
timestamp 1679581782
transform 1 0 51936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_542
timestamp 1679581782
transform 1 0 52608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_549
timestamp 1679581782
transform 1 0 53280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_556
timestamp 1679581782
transform 1 0 53952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_563
timestamp 1679581782
transform 1 0 54624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_570
timestamp 1679581782
transform 1 0 55296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_577
timestamp 1679581782
transform 1 0 55968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_584
timestamp 1679581782
transform 1 0 56640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_591
timestamp 1679581782
transform 1 0 57312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_598
timestamp 1679581782
transform 1 0 57984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_605
timestamp 1679581782
transform 1 0 58656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_612
timestamp 1679581782
transform 1 0 59328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_619
timestamp 1679581782
transform 1 0 60000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_626
timestamp 1679581782
transform 1 0 60672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_633
timestamp 1679581782
transform 1 0 61344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_640
timestamp 1679581782
transform 1 0 62016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_647
timestamp 1679581782
transform 1 0 62688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_654
timestamp 1679581782
transform 1 0 63360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_661
timestamp 1679581782
transform 1 0 64032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_668
timestamp 1679581782
transform 1 0 64704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_675
timestamp 1679581782
transform 1 0 65376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_682
timestamp 1679581782
transform 1 0 66048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_689
timestamp 1679581782
transform 1 0 66720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_696
timestamp 1679581782
transform 1 0 67392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_703
timestamp 1679581782
transform 1 0 68064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_710
timestamp 1679581782
transform 1 0 68736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_717
timestamp 1679581782
transform 1 0 69408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_724
timestamp 1679581782
transform 1 0 70080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_731
timestamp 1679581782
transform 1 0 70752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_738
timestamp 1679581782
transform 1 0 71424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_745
timestamp 1679581782
transform 1 0 72096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_752
timestamp 1679581782
transform 1 0 72768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_759
timestamp 1679581782
transform 1 0 73440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_766
timestamp 1679581782
transform 1 0 74112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_773
timestamp 1679581782
transform 1 0 74784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_780
timestamp 1679581782
transform 1 0 75456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_787
timestamp 1679581782
transform 1 0 76128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_794
timestamp 1679581782
transform 1 0 76800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_801
timestamp 1679581782
transform 1 0 77472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_808
timestamp 1679581782
transform 1 0 78144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_815
timestamp 1679581782
transform 1 0 78816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_822
timestamp 1679581782
transform 1 0 79488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_829
timestamp 1679581782
transform 1 0 80160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_836
timestamp 1679581782
transform 1 0 80832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_843
timestamp 1679581782
transform 1 0 81504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_850
timestamp 1679581782
transform 1 0 82176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_857
timestamp 1679581782
transform 1 0 82848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_864
timestamp 1679581782
transform 1 0 83520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_871
timestamp 1679581782
transform 1 0 84192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_878
timestamp 1679581782
transform 1 0 84864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_885
timestamp 1679581782
transform 1 0 85536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_892
timestamp 1679581782
transform 1 0 86208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_899
timestamp 1679581782
transform 1 0 86880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_906
timestamp 1679581782
transform 1 0 87552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_913
timestamp 1679581782
transform 1 0 88224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_920
timestamp 1679581782
transform 1 0 88896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_927
timestamp 1679581782
transform 1 0 89568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_934
timestamp 1679581782
transform 1 0 90240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_941
timestamp 1679581782
transform 1 0 90912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_948
timestamp 1679581782
transform 1 0 91584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_955
timestamp 1679581782
transform 1 0 92256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_962
timestamp 1679581782
transform 1 0 92928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_969
timestamp 1679581782
transform 1 0 93600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_976
timestamp 1679581782
transform 1 0 94272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_983
timestamp 1679581782
transform 1 0 94944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_990
timestamp 1679581782
transform 1 0 95616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_997
timestamp 1679581782
transform 1 0 96288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1004
timestamp 1679581782
transform 1 0 96960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1011
timestamp 1679581782
transform 1 0 97632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1018
timestamp 1679581782
transform 1 0 98304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_1025
timestamp 1679577901
transform 1 0 98976 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_7
timestamp 1679577901
transform 1 0 1248 0 1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_36_15
timestamp 1679577901
transform 1 0 2016 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_19
timestamp 1677579658
transform 1 0 2400 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_56
timestamp 1677579658
transform 1 0 5952 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_93
timestamp 1677579658
transform 1 0 9504 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_130
timestamp 1677580104
transform 1 0 13056 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_145
timestamp 1677580104
transform 1 0 14496 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_190
timestamp 1677579658
transform 1 0 18816 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_227
timestamp 1679581782
transform 1 0 22368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_234
timestamp 1679577901
transform 1 0 23040 0 1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_36_242
timestamp 1679577901
transform 1 0 23808 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_246
timestamp 1677580104
transform 1 0 24192 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_275
timestamp 1677580104
transform 1 0 26976 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_277
timestamp 1677579658
transform 1 0 27168 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_310
timestamp 1677580104
transform 1 0 30336 0 1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_382
timestamp 1679577901
transform 1 0 37248 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_390
timestamp 1677580104
transform 1 0 38016 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_405
timestamp 1677579658
transform 1 0 39456 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_439
timestamp 1677579658
transform 1 0 42720 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_472
timestamp 1677579658
transform 1 0 45888 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_476
timestamp 1677579658
transform 1 0 46272 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_486
timestamp 1677579658
transform 1 0 47232 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_510
timestamp 1677580104
transform 1 0 49536 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_512
timestamp 1677579658
transform 1 0 49728 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_522
timestamp 1679581782
transform 1 0 50688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_529
timestamp 1679581782
transform 1 0 51360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_536
timestamp 1679581782
transform 1 0 52032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_543
timestamp 1679581782
transform 1 0 52704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_550
timestamp 1679581782
transform 1 0 53376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_557
timestamp 1679581782
transform 1 0 54048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_564
timestamp 1679581782
transform 1 0 54720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_571
timestamp 1679581782
transform 1 0 55392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_578
timestamp 1679581782
transform 1 0 56064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_585
timestamp 1679581782
transform 1 0 56736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_592
timestamp 1679581782
transform 1 0 57408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_599
timestamp 1679581782
transform 1 0 58080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_606
timestamp 1679581782
transform 1 0 58752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_613
timestamp 1679581782
transform 1 0 59424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_620
timestamp 1679581782
transform 1 0 60096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_627
timestamp 1679581782
transform 1 0 60768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_634
timestamp 1679581782
transform 1 0 61440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_641
timestamp 1679581782
transform 1 0 62112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_648
timestamp 1679581782
transform 1 0 62784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_655
timestamp 1679581782
transform 1 0 63456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_662
timestamp 1679581782
transform 1 0 64128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_669
timestamp 1679581782
transform 1 0 64800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_676
timestamp 1679581782
transform 1 0 65472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_683
timestamp 1679581782
transform 1 0 66144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_690
timestamp 1679581782
transform 1 0 66816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_697
timestamp 1679581782
transform 1 0 67488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_704
timestamp 1679581782
transform 1 0 68160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_711
timestamp 1679581782
transform 1 0 68832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_718
timestamp 1679581782
transform 1 0 69504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_725
timestamp 1679581782
transform 1 0 70176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_732
timestamp 1679581782
transform 1 0 70848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_739
timestamp 1679581782
transform 1 0 71520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_746
timestamp 1679581782
transform 1 0 72192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_753
timestamp 1679581782
transform 1 0 72864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_760
timestamp 1679581782
transform 1 0 73536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_767
timestamp 1679581782
transform 1 0 74208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_774
timestamp 1679581782
transform 1 0 74880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_781
timestamp 1679581782
transform 1 0 75552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_788
timestamp 1679581782
transform 1 0 76224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_795
timestamp 1679581782
transform 1 0 76896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_802
timestamp 1679581782
transform 1 0 77568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_809
timestamp 1679581782
transform 1 0 78240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_816
timestamp 1679581782
transform 1 0 78912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_823
timestamp 1679581782
transform 1 0 79584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_830
timestamp 1679581782
transform 1 0 80256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_837
timestamp 1679581782
transform 1 0 80928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_844
timestamp 1679581782
transform 1 0 81600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_851
timestamp 1679581782
transform 1 0 82272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_858
timestamp 1679581782
transform 1 0 82944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_865
timestamp 1679581782
transform 1 0 83616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_872
timestamp 1679581782
transform 1 0 84288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_879
timestamp 1679581782
transform 1 0 84960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_886
timestamp 1679581782
transform 1 0 85632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_893
timestamp 1679581782
transform 1 0 86304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_900
timestamp 1679581782
transform 1 0 86976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_907
timestamp 1679581782
transform 1 0 87648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_914
timestamp 1679581782
transform 1 0 88320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_921
timestamp 1679581782
transform 1 0 88992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_928
timestamp 1679581782
transform 1 0 89664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_935
timestamp 1679581782
transform 1 0 90336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_942
timestamp 1679581782
transform 1 0 91008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_949
timestamp 1679581782
transform 1 0 91680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_956
timestamp 1679581782
transform 1 0 92352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_963
timestamp 1679581782
transform 1 0 93024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_970
timestamp 1679581782
transform 1 0 93696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_977
timestamp 1679581782
transform 1 0 94368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_984
timestamp 1679581782
transform 1 0 95040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_991
timestamp 1679581782
transform 1 0 95712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_998
timestamp 1679581782
transform 1 0 96384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1005
timestamp 1679581782
transform 1 0 97056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1012
timestamp 1679581782
transform 1 0 97728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1019
timestamp 1679581782
transform 1 0 98400 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_1026
timestamp 1677580104
transform 1 0 99072 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_1028
timestamp 1677579658
transform 1 0 99264 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_0
timestamp 1677580104
transform 1 0 576 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_2
timestamp 1677579658
transform 1 0 768 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_43
timestamp 1677579658
transform 1 0 4704 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_111
timestamp 1679577901
transform 1 0 11232 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_115
timestamp 1677579658
transform 1 0 11616 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_125
timestamp 1679581782
transform 1 0 12576 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_132
timestamp 1677580104
transform 1 0 13248 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_138
timestamp 1679577901
transform 1 0 13824 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_142
timestamp 1677580104
transform 1 0 14208 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_150
timestamp 1677580104
transform 1 0 14976 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_202
timestamp 1679577901
transform 1 0 19968 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_219
timestamp 1679581782
transform 1 0 21600 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_226
timestamp 1677580104
transform 1 0 22272 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_247
timestamp 1677580104
transform 1 0 24288 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_268
timestamp 1677580104
transform 1 0 26304 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_285
timestamp 1677579658
transform 1 0 27936 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_291
timestamp 1679577901
transform 1 0 28512 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_295
timestamp 1677580104
transform 1 0 28896 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_323
timestamp 1677580104
transform 1 0 31584 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_380
timestamp 1677579658
transform 1 0 37056 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_386
timestamp 1677580104
transform 1 0 37632 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_399
timestamp 1679577901
transform 1 0 38880 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_403
timestamp 1677580104
transform 1 0 39264 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_441
timestamp 1677579658
transform 1 0 42912 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_451
timestamp 1677579658
transform 1 0 43872 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_470
timestamp 1677579658
transform 1 0 45696 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_507
timestamp 1679581782
transform 1 0 49248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_514
timestamp 1679581782
transform 1 0 49920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_521
timestamp 1679581782
transform 1 0 50592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_528
timestamp 1679581782
transform 1 0 51264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_535
timestamp 1679581782
transform 1 0 51936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_542
timestamp 1679581782
transform 1 0 52608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_549
timestamp 1679581782
transform 1 0 53280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_556
timestamp 1679581782
transform 1 0 53952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_563
timestamp 1679581782
transform 1 0 54624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_570
timestamp 1679581782
transform 1 0 55296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_577
timestamp 1679581782
transform 1 0 55968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_584
timestamp 1679581782
transform 1 0 56640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_591
timestamp 1679581782
transform 1 0 57312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_598
timestamp 1679581782
transform 1 0 57984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_605
timestamp 1679581782
transform 1 0 58656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_612
timestamp 1679581782
transform 1 0 59328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_619
timestamp 1679581782
transform 1 0 60000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_626
timestamp 1679581782
transform 1 0 60672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_633
timestamp 1679581782
transform 1 0 61344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_640
timestamp 1679581782
transform 1 0 62016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_647
timestamp 1679581782
transform 1 0 62688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_654
timestamp 1679581782
transform 1 0 63360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_661
timestamp 1679581782
transform 1 0 64032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_668
timestamp 1679581782
transform 1 0 64704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_675
timestamp 1679581782
transform 1 0 65376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_682
timestamp 1679581782
transform 1 0 66048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_689
timestamp 1679581782
transform 1 0 66720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_696
timestamp 1679581782
transform 1 0 67392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_703
timestamp 1679581782
transform 1 0 68064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_710
timestamp 1679581782
transform 1 0 68736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_717
timestamp 1679581782
transform 1 0 69408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_724
timestamp 1679581782
transform 1 0 70080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_731
timestamp 1679581782
transform 1 0 70752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_738
timestamp 1679581782
transform 1 0 71424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_745
timestamp 1679581782
transform 1 0 72096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_752
timestamp 1679581782
transform 1 0 72768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_759
timestamp 1679581782
transform 1 0 73440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_766
timestamp 1679581782
transform 1 0 74112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_773
timestamp 1679581782
transform 1 0 74784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_780
timestamp 1679581782
transform 1 0 75456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_787
timestamp 1679581782
transform 1 0 76128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_794
timestamp 1679581782
transform 1 0 76800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_801
timestamp 1679581782
transform 1 0 77472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_808
timestamp 1679581782
transform 1 0 78144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_815
timestamp 1679581782
transform 1 0 78816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_822
timestamp 1679581782
transform 1 0 79488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_829
timestamp 1679581782
transform 1 0 80160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_836
timestamp 1679581782
transform 1 0 80832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_843
timestamp 1679581782
transform 1 0 81504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_850
timestamp 1679581782
transform 1 0 82176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_857
timestamp 1679581782
transform 1 0 82848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_864
timestamp 1679581782
transform 1 0 83520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_871
timestamp 1679581782
transform 1 0 84192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_878
timestamp 1679581782
transform 1 0 84864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_885
timestamp 1679581782
transform 1 0 85536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_892
timestamp 1679581782
transform 1 0 86208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_899
timestamp 1679581782
transform 1 0 86880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_906
timestamp 1679581782
transform 1 0 87552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_913
timestamp 1679581782
transform 1 0 88224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_920
timestamp 1679581782
transform 1 0 88896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_927
timestamp 1679581782
transform 1 0 89568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_934
timestamp 1679581782
transform 1 0 90240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_941
timestamp 1679581782
transform 1 0 90912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_948
timestamp 1679581782
transform 1 0 91584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_955
timestamp 1679581782
transform 1 0 92256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_962
timestamp 1679581782
transform 1 0 92928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_969
timestamp 1679581782
transform 1 0 93600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_976
timestamp 1679581782
transform 1 0 94272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_983
timestamp 1679581782
transform 1 0 94944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_990
timestamp 1679581782
transform 1 0 95616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_997
timestamp 1679581782
transform 1 0 96288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1004
timestamp 1679581782
transform 1 0 96960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1011
timestamp 1679581782
transform 1 0 97632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1018
timestamp 1679581782
transform 1 0 98304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_1025
timestamp 1679577901
transform 1 0 98976 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_34
timestamp 1677580104
transform 1 0 3840 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_51
timestamp 1677579658
transform 1 0 5472 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_100
timestamp 1679581782
transform 1 0 10176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_213
timestamp 1679577901
transform 1 0 21024 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_217
timestamp 1677580104
transform 1 0 21408 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_227
timestamp 1677579658
transform 1 0 22368 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_255
timestamp 1677579658
transform 1 0 25056 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_270
timestamp 1677579658
transform 1 0 26496 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_284
timestamp 1679581782
transform 1 0 27840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_291
timestamp 1679577901
transform 1 0 28512 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_295
timestamp 1677579658
transform 1 0 28896 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_345
timestamp 1677580104
transform 1 0 33696 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_356
timestamp 1677580104
transform 1 0 34752 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_363
timestamp 1677580104
transform 1 0 35424 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_410
timestamp 1677580104
transform 1 0 39936 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_412
timestamp 1677579658
transform 1 0 40128 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_441
timestamp 1677580104
transform 1 0 42912 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679581782
transform 1 0 46944 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_490
timestamp 1677579658
transform 1 0 47616 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_494
timestamp 1679581782
transform 1 0 48000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_501
timestamp 1679581782
transform 1 0 48672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_508
timestamp 1679581782
transform 1 0 49344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_515
timestamp 1679581782
transform 1 0 50016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_522
timestamp 1679581782
transform 1 0 50688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_529
timestamp 1679581782
transform 1 0 51360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_536
timestamp 1679581782
transform 1 0 52032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_543
timestamp 1679581782
transform 1 0 52704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_550
timestamp 1679581782
transform 1 0 53376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_557
timestamp 1679581782
transform 1 0 54048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_564
timestamp 1679581782
transform 1 0 54720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_571
timestamp 1679581782
transform 1 0 55392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_578
timestamp 1679581782
transform 1 0 56064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_585
timestamp 1679581782
transform 1 0 56736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_592
timestamp 1679581782
transform 1 0 57408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_599
timestamp 1679581782
transform 1 0 58080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_606
timestamp 1679581782
transform 1 0 58752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_613
timestamp 1679581782
transform 1 0 59424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_620
timestamp 1679581782
transform 1 0 60096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_627
timestamp 1679581782
transform 1 0 60768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_634
timestamp 1679581782
transform 1 0 61440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_641
timestamp 1679581782
transform 1 0 62112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_648
timestamp 1679581782
transform 1 0 62784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_655
timestamp 1679581782
transform 1 0 63456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_662
timestamp 1679581782
transform 1 0 64128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_669
timestamp 1679581782
transform 1 0 64800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_676
timestamp 1679581782
transform 1 0 65472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_683
timestamp 1679581782
transform 1 0 66144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_690
timestamp 1679581782
transform 1 0 66816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_697
timestamp 1679581782
transform 1 0 67488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_704
timestamp 1679581782
transform 1 0 68160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_711
timestamp 1679581782
transform 1 0 68832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_718
timestamp 1679581782
transform 1 0 69504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_725
timestamp 1679581782
transform 1 0 70176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_732
timestamp 1679581782
transform 1 0 70848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_739
timestamp 1679581782
transform 1 0 71520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_746
timestamp 1679581782
transform 1 0 72192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_753
timestamp 1679581782
transform 1 0 72864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_760
timestamp 1679581782
transform 1 0 73536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_767
timestamp 1679581782
transform 1 0 74208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_774
timestamp 1679581782
transform 1 0 74880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_781
timestamp 1679581782
transform 1 0 75552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_788
timestamp 1679581782
transform 1 0 76224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_795
timestamp 1679581782
transform 1 0 76896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_802
timestamp 1679581782
transform 1 0 77568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_809
timestamp 1679581782
transform 1 0 78240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_816
timestamp 1679581782
transform 1 0 78912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_823
timestamp 1679581782
transform 1 0 79584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_830
timestamp 1679581782
transform 1 0 80256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_837
timestamp 1679581782
transform 1 0 80928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_844
timestamp 1679581782
transform 1 0 81600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_851
timestamp 1679581782
transform 1 0 82272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_858
timestamp 1679581782
transform 1 0 82944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_865
timestamp 1679581782
transform 1 0 83616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_872
timestamp 1679581782
transform 1 0 84288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_879
timestamp 1679581782
transform 1 0 84960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_886
timestamp 1679581782
transform 1 0 85632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_893
timestamp 1679581782
transform 1 0 86304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_900
timestamp 1679581782
transform 1 0 86976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_907
timestamp 1679581782
transform 1 0 87648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_914
timestamp 1679581782
transform 1 0 88320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_921
timestamp 1679581782
transform 1 0 88992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_928
timestamp 1679581782
transform 1 0 89664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_935
timestamp 1679581782
transform 1 0 90336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_942
timestamp 1679581782
transform 1 0 91008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_949
timestamp 1679581782
transform 1 0 91680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_956
timestamp 1679581782
transform 1 0 92352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_963
timestamp 1679581782
transform 1 0 93024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_970
timestamp 1679581782
transform 1 0 93696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_977
timestamp 1679581782
transform 1 0 94368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_984
timestamp 1679581782
transform 1 0 95040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_991
timestamp 1679581782
transform 1 0 95712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_998
timestamp 1679581782
transform 1 0 96384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1005
timestamp 1679581782
transform 1 0 97056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1012
timestamp 1679581782
transform 1 0 97728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1019
timestamp 1679581782
transform 1 0 98400 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_1026
timestamp 1677580104
transform 1 0 99072 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_1028
timestamp 1677579658
transform 1 0 99264 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_7
timestamp 1679577901
transform 1 0 1248 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_11
timestamp 1677579658
transform 1 0 1632 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_16
timestamp 1679581782
transform 1 0 2112 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_23
timestamp 1677580104
transform 1 0 2784 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_48
timestamp 1677579658
transform 1 0 5184 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_70
timestamp 1677580104
transform 1 0 7296 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_99
timestamp 1679577901
transform 1 0 10080 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_103
timestamp 1677580104
transform 1 0 10464 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_123
timestamp 1677579658
transform 1 0 12384 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_152
timestamp 1677580104
transform 1 0 15168 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_164
timestamp 1677579658
transform 1 0 16320 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_197
timestamp 1677579658
transform 1 0 19488 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_243
timestamp 1679581782
transform 1 0 23904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_250
timestamp 1679577901
transform 1 0 24576 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_334
timestamp 1677579658
transform 1 0 32640 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_372
timestamp 1677579658
transform 1 0 36288 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_420
timestamp 1679577901
transform 1 0 40896 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_424
timestamp 1677579658
transform 1 0 41280 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_452
timestamp 1679577901
transform 1 0 43968 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_472
timestamp 1679581782
transform 1 0 45888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_479
timestamp 1679581782
transform 1 0 46560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_486
timestamp 1679581782
transform 1 0 47232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_493
timestamp 1679581782
transform 1 0 47904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_500
timestamp 1679581782
transform 1 0 48576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_507
timestamp 1679581782
transform 1 0 49248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_514
timestamp 1679581782
transform 1 0 49920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_521
timestamp 1679581782
transform 1 0 50592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_528
timestamp 1679581782
transform 1 0 51264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_535
timestamp 1679581782
transform 1 0 51936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_542
timestamp 1679581782
transform 1 0 52608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_549
timestamp 1679581782
transform 1 0 53280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_556
timestamp 1679581782
transform 1 0 53952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_563
timestamp 1679581782
transform 1 0 54624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_570
timestamp 1679581782
transform 1 0 55296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_577
timestamp 1679581782
transform 1 0 55968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_584
timestamp 1679581782
transform 1 0 56640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_591
timestamp 1679581782
transform 1 0 57312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_598
timestamp 1679581782
transform 1 0 57984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_605
timestamp 1679581782
transform 1 0 58656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_612
timestamp 1679581782
transform 1 0 59328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_619
timestamp 1679581782
transform 1 0 60000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_626
timestamp 1679581782
transform 1 0 60672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_633
timestamp 1679581782
transform 1 0 61344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_640
timestamp 1679581782
transform 1 0 62016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_647
timestamp 1679581782
transform 1 0 62688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_654
timestamp 1679581782
transform 1 0 63360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_661
timestamp 1679581782
transform 1 0 64032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_668
timestamp 1679581782
transform 1 0 64704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_675
timestamp 1679581782
transform 1 0 65376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_682
timestamp 1679581782
transform 1 0 66048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_689
timestamp 1679581782
transform 1 0 66720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_696
timestamp 1679581782
transform 1 0 67392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_703
timestamp 1679581782
transform 1 0 68064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_710
timestamp 1679581782
transform 1 0 68736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_717
timestamp 1679581782
transform 1 0 69408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_724
timestamp 1679581782
transform 1 0 70080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_731
timestamp 1679581782
transform 1 0 70752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_738
timestamp 1679581782
transform 1 0 71424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_745
timestamp 1679581782
transform 1 0 72096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_752
timestamp 1679581782
transform 1 0 72768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_759
timestamp 1679581782
transform 1 0 73440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_766
timestamp 1679581782
transform 1 0 74112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_773
timestamp 1679581782
transform 1 0 74784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_780
timestamp 1679581782
transform 1 0 75456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_787
timestamp 1679581782
transform 1 0 76128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_794
timestamp 1679581782
transform 1 0 76800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_801
timestamp 1679581782
transform 1 0 77472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_808
timestamp 1679581782
transform 1 0 78144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_815
timestamp 1679581782
transform 1 0 78816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_822
timestamp 1679581782
transform 1 0 79488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_829
timestamp 1679581782
transform 1 0 80160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_836
timestamp 1679581782
transform 1 0 80832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_843
timestamp 1679581782
transform 1 0 81504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_850
timestamp 1679581782
transform 1 0 82176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_857
timestamp 1679581782
transform 1 0 82848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_864
timestamp 1679581782
transform 1 0 83520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_871
timestamp 1679581782
transform 1 0 84192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_878
timestamp 1679581782
transform 1 0 84864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_885
timestamp 1679581782
transform 1 0 85536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_892
timestamp 1679581782
transform 1 0 86208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_899
timestamp 1679581782
transform 1 0 86880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_906
timestamp 1679581782
transform 1 0 87552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_913
timestamp 1679581782
transform 1 0 88224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_920
timestamp 1679581782
transform 1 0 88896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_927
timestamp 1679581782
transform 1 0 89568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_934
timestamp 1679581782
transform 1 0 90240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_941
timestamp 1679581782
transform 1 0 90912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_948
timestamp 1679581782
transform 1 0 91584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_955
timestamp 1679581782
transform 1 0 92256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_962
timestamp 1679581782
transform 1 0 92928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_969
timestamp 1679581782
transform 1 0 93600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_976
timestamp 1679581782
transform 1 0 94272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_983
timestamp 1679581782
transform 1 0 94944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_990
timestamp 1679581782
transform 1 0 95616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_997
timestamp 1679581782
transform 1 0 96288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1004
timestamp 1679581782
transform 1 0 96960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1011
timestamp 1679581782
transform 1 0 97632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1018
timestamp 1679581782
transform 1 0 98304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_1025
timestamp 1679577901
transform 1 0 98976 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_40_0
timestamp 1679577901
transform 1 0 576 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_4
timestamp 1677579658
transform 1 0 960 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_36
timestamp 1677580104
transform 1 0 4032 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_62
timestamp 1677579658
transform 1 0 6528 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_89
timestamp 1679577901
transform 1 0 9120 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_93
timestamp 1677579658
transform 1 0 9504 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_129
timestamp 1677580104
transform 1 0 12960 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_144
timestamp 1677579658
transform 1 0 14400 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_203
timestamp 1679577901
transform 1 0 20064 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_207
timestamp 1677579658
transform 1 0 20448 0 1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_213
timestamp 1679577901
transform 1 0 21024 0 1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_40_235
timestamp 1679577901
transform 1 0 23136 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_239
timestamp 1677580104
transform 1 0 23520 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_271
timestamp 1679581782
transform 1 0 26592 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_278
timestamp 1677579658
transform 1 0 27264 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_292
timestamp 1679581782
transform 1 0 28608 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_352
timestamp 1677580104
transform 1 0 34368 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_354
timestamp 1677579658
transform 1 0 34560 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_382
timestamp 1677580104
transform 1 0 37248 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_427
timestamp 1677580104
transform 1 0 41568 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_429
timestamp 1677579658
transform 1 0 41760 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_441
timestamp 1677580104
transform 1 0 42912 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_446
timestamp 1679581782
transform 1 0 43392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_453
timestamp 1679581782
transform 1 0 44064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_460
timestamp 1679581782
transform 1 0 44736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_467
timestamp 1679581782
transform 1 0 45408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_474
timestamp 1679581782
transform 1 0 46080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_481
timestamp 1679581782
transform 1 0 46752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_488
timestamp 1679581782
transform 1 0 47424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_495
timestamp 1679581782
transform 1 0 48096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_502
timestamp 1679581782
transform 1 0 48768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_509
timestamp 1679581782
transform 1 0 49440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_516
timestamp 1679581782
transform 1 0 50112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_523
timestamp 1679581782
transform 1 0 50784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_530
timestamp 1679581782
transform 1 0 51456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_537
timestamp 1679581782
transform 1 0 52128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_544
timestamp 1679581782
transform 1 0 52800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_551
timestamp 1679581782
transform 1 0 53472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_558
timestamp 1679581782
transform 1 0 54144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_565
timestamp 1679581782
transform 1 0 54816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_572
timestamp 1679581782
transform 1 0 55488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_579
timestamp 1679581782
transform 1 0 56160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_586
timestamp 1679581782
transform 1 0 56832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_593
timestamp 1679581782
transform 1 0 57504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_600
timestamp 1679581782
transform 1 0 58176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_607
timestamp 1679581782
transform 1 0 58848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_614
timestamp 1679581782
transform 1 0 59520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_621
timestamp 1679581782
transform 1 0 60192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_628
timestamp 1679581782
transform 1 0 60864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_635
timestamp 1679581782
transform 1 0 61536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_642
timestamp 1679581782
transform 1 0 62208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_649
timestamp 1679581782
transform 1 0 62880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_656
timestamp 1679581782
transform 1 0 63552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_663
timestamp 1679581782
transform 1 0 64224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_670
timestamp 1679581782
transform 1 0 64896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_677
timestamp 1679581782
transform 1 0 65568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_684
timestamp 1679581782
transform 1 0 66240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_691
timestamp 1679581782
transform 1 0 66912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_698
timestamp 1679581782
transform 1 0 67584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_705
timestamp 1679581782
transform 1 0 68256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_712
timestamp 1679581782
transform 1 0 68928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_719
timestamp 1679581782
transform 1 0 69600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_726
timestamp 1679581782
transform 1 0 70272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_733
timestamp 1679581782
transform 1 0 70944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_740
timestamp 1679581782
transform 1 0 71616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_747
timestamp 1679581782
transform 1 0 72288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_754
timestamp 1679581782
transform 1 0 72960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_761
timestamp 1679581782
transform 1 0 73632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_768
timestamp 1679581782
transform 1 0 74304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_775
timestamp 1679581782
transform 1 0 74976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_782
timestamp 1679581782
transform 1 0 75648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_789
timestamp 1679581782
transform 1 0 76320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_796
timestamp 1679581782
transform 1 0 76992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_803
timestamp 1679581782
transform 1 0 77664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_810
timestamp 1679581782
transform 1 0 78336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_817
timestamp 1679581782
transform 1 0 79008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_824
timestamp 1679581782
transform 1 0 79680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_831
timestamp 1679581782
transform 1 0 80352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_838
timestamp 1679581782
transform 1 0 81024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_845
timestamp 1679581782
transform 1 0 81696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_852
timestamp 1679581782
transform 1 0 82368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_859
timestamp 1679581782
transform 1 0 83040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_866
timestamp 1679581782
transform 1 0 83712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_873
timestamp 1679581782
transform 1 0 84384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_880
timestamp 1679581782
transform 1 0 85056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_887
timestamp 1679581782
transform 1 0 85728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_894
timestamp 1679581782
transform 1 0 86400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_901
timestamp 1679581782
transform 1 0 87072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_908
timestamp 1679581782
transform 1 0 87744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_915
timestamp 1679581782
transform 1 0 88416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_922
timestamp 1679581782
transform 1 0 89088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_929
timestamp 1679581782
transform 1 0 89760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_936
timestamp 1679581782
transform 1 0 90432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_943
timestamp 1679581782
transform 1 0 91104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_950
timestamp 1679581782
transform 1 0 91776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_957
timestamp 1679581782
transform 1 0 92448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_964
timestamp 1679581782
transform 1 0 93120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_971
timestamp 1679581782
transform 1 0 93792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_978
timestamp 1679581782
transform 1 0 94464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_985
timestamp 1679581782
transform 1 0 95136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_992
timestamp 1679581782
transform 1 0 95808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_999
timestamp 1679581782
transform 1 0 96480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1006
timestamp 1679581782
transform 1 0 97152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1013
timestamp 1679581782
transform 1 0 97824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1020
timestamp 1679581782
transform 1 0 98496 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_1027
timestamp 1677580104
transform 1 0 99168 0 1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_0
timestamp 1679577901
transform 1 0 576 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_4
timestamp 1677579658
transform 1 0 960 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_41
timestamp 1677580104
transform 1 0 4512 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_62
timestamp 1677579658
transform 1 0 6528 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_66
timestamp 1677580104
transform 1 0 6912 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_73
timestamp 1677580104
transform 1 0 7584 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_75
timestamp 1677579658
transform 1 0 7776 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_81
timestamp 1679581782
transform 1 0 8352 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_88
timestamp 1677579658
transform 1 0 9024 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_124
timestamp 1677579658
transform 1 0 12480 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_162
timestamp 1677579658
transform 1 0 16128 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_184
timestamp 1677579658
transform 1 0 18240 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_213
timestamp 1679577901
transform 1 0 21024 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_217
timestamp 1677580104
transform 1 0 21408 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_232
timestamp 1677579658
transform 1 0 22848 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_250
timestamp 1677580104
transform 1 0 24576 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_252
timestamp 1677579658
transform 1 0 24768 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_262
timestamp 1677579658
transform 1 0 25728 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_286
timestamp 1679577901
transform 1 0 28032 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_290
timestamp 1677580104
transform 1 0 28416 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_304
timestamp 1677580104
transform 1 0 29760 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_341
timestamp 1679577901
transform 1 0 33312 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_387
timestamp 1677580104
transform 1 0 37728 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_418
timestamp 1679581782
transform 1 0 40704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_425
timestamp 1679581782
transform 1 0 41376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_432
timestamp 1679581782
transform 1 0 42048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_439
timestamp 1679581782
transform 1 0 42720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_446
timestamp 1679581782
transform 1 0 43392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_453
timestamp 1679581782
transform 1 0 44064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_460
timestamp 1679581782
transform 1 0 44736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_467
timestamp 1679581782
transform 1 0 45408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_474
timestamp 1679581782
transform 1 0 46080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_481
timestamp 1679581782
transform 1 0 46752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_488
timestamp 1679581782
transform 1 0 47424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_495
timestamp 1679581782
transform 1 0 48096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_502
timestamp 1679581782
transform 1 0 48768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_509
timestamp 1679581782
transform 1 0 49440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_516
timestamp 1679581782
transform 1 0 50112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_523
timestamp 1679581782
transform 1 0 50784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_530
timestamp 1679581782
transform 1 0 51456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_537
timestamp 1679581782
transform 1 0 52128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_544
timestamp 1679581782
transform 1 0 52800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_551
timestamp 1679581782
transform 1 0 53472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_558
timestamp 1679581782
transform 1 0 54144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_565
timestamp 1679581782
transform 1 0 54816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_572
timestamp 1679581782
transform 1 0 55488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_579
timestamp 1679581782
transform 1 0 56160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_586
timestamp 1679581782
transform 1 0 56832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_593
timestamp 1679581782
transform 1 0 57504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_600
timestamp 1679581782
transform 1 0 58176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_607
timestamp 1679581782
transform 1 0 58848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_614
timestamp 1679581782
transform 1 0 59520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_621
timestamp 1679581782
transform 1 0 60192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_628
timestamp 1679581782
transform 1 0 60864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_635
timestamp 1679581782
transform 1 0 61536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_642
timestamp 1679581782
transform 1 0 62208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_649
timestamp 1679581782
transform 1 0 62880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_656
timestamp 1679581782
transform 1 0 63552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_663
timestamp 1679581782
transform 1 0 64224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_670
timestamp 1679581782
transform 1 0 64896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_677
timestamp 1679581782
transform 1 0 65568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_684
timestamp 1679581782
transform 1 0 66240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_691
timestamp 1679581782
transform 1 0 66912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_698
timestamp 1679581782
transform 1 0 67584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_705
timestamp 1679581782
transform 1 0 68256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_712
timestamp 1679581782
transform 1 0 68928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_719
timestamp 1679581782
transform 1 0 69600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_726
timestamp 1679581782
transform 1 0 70272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_733
timestamp 1679581782
transform 1 0 70944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_740
timestamp 1679581782
transform 1 0 71616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_747
timestamp 1679581782
transform 1 0 72288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_754
timestamp 1679581782
transform 1 0 72960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_761
timestamp 1679581782
transform 1 0 73632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_768
timestamp 1679581782
transform 1 0 74304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_775
timestamp 1679581782
transform 1 0 74976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_782
timestamp 1679581782
transform 1 0 75648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_789
timestamp 1679581782
transform 1 0 76320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_796
timestamp 1679581782
transform 1 0 76992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_803
timestamp 1679581782
transform 1 0 77664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_810
timestamp 1679581782
transform 1 0 78336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_817
timestamp 1679581782
transform 1 0 79008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_824
timestamp 1679581782
transform 1 0 79680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_831
timestamp 1679581782
transform 1 0 80352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_838
timestamp 1679581782
transform 1 0 81024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_845
timestamp 1679581782
transform 1 0 81696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_852
timestamp 1679581782
transform 1 0 82368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_859
timestamp 1679581782
transform 1 0 83040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_866
timestamp 1679581782
transform 1 0 83712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_873
timestamp 1679581782
transform 1 0 84384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_880
timestamp 1679581782
transform 1 0 85056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_887
timestamp 1679581782
transform 1 0 85728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_894
timestamp 1679581782
transform 1 0 86400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_901
timestamp 1679581782
transform 1 0 87072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_908
timestamp 1679581782
transform 1 0 87744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_915
timestamp 1679581782
transform 1 0 88416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_922
timestamp 1679581782
transform 1 0 89088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_929
timestamp 1679581782
transform 1 0 89760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_936
timestamp 1679581782
transform 1 0 90432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_943
timestamp 1679581782
transform 1 0 91104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_950
timestamp 1679581782
transform 1 0 91776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_957
timestamp 1679581782
transform 1 0 92448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_964
timestamp 1679581782
transform 1 0 93120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_971
timestamp 1679581782
transform 1 0 93792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_978
timestamp 1679581782
transform 1 0 94464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_985
timestamp 1679581782
transform 1 0 95136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_992
timestamp 1679581782
transform 1 0 95808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_999
timestamp 1679581782
transform 1 0 96480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1006
timestamp 1679581782
transform 1 0 97152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1013
timestamp 1679581782
transform 1 0 97824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1020
timestamp 1679581782
transform 1 0 98496 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_1027
timestamp 1677580104
transform 1 0 99168 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_7
timestamp 1677580104
transform 1 0 1248 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_9
timestamp 1677579658
transform 1 0 1440 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_14
timestamp 1679577901
transform 1 0 1920 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_60
timestamp 1677579658
transform 1 0 6336 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_92
timestamp 1679577901
transform 1 0 9408 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_111
timestamp 1677579658
transform 1 0 11232 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_122
timestamp 1677579658
transform 1 0 12288 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_171
timestamp 1677580104
transform 1 0 16992 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_173
timestamp 1677579658
transform 1 0 17184 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_210
timestamp 1679577901
transform 1 0 20736 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_214
timestamp 1677579658
transform 1 0 21120 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_225
timestamp 1679581782
transform 1 0 22176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_232
timestamp 1679577901
transform 1 0 22848 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_236
timestamp 1677580104
transform 1 0 23232 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_259
timestamp 1677580104
transform 1 0 25440 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_320
timestamp 1677580104
transform 1 0 31296 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_322
timestamp 1677579658
transform 1 0 31488 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_341
timestamp 1677579658
transform 1 0 33312 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_369
timestamp 1677579658
transform 1 0 36000 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_411
timestamp 1679581782
transform 1 0 40032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_418
timestamp 1679581782
transform 1 0 40704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_425
timestamp 1679581782
transform 1 0 41376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_432
timestamp 1679581782
transform 1 0 42048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_439
timestamp 1679581782
transform 1 0 42720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_446
timestamp 1679581782
transform 1 0 43392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_453
timestamp 1679581782
transform 1 0 44064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_460
timestamp 1679581782
transform 1 0 44736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_467
timestamp 1679581782
transform 1 0 45408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_474
timestamp 1679581782
transform 1 0 46080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_481
timestamp 1679581782
transform 1 0 46752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_488
timestamp 1679581782
transform 1 0 47424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_495
timestamp 1679581782
transform 1 0 48096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_502
timestamp 1679581782
transform 1 0 48768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_509
timestamp 1679581782
transform 1 0 49440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_516
timestamp 1679581782
transform 1 0 50112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_523
timestamp 1679581782
transform 1 0 50784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_530
timestamp 1679581782
transform 1 0 51456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_537
timestamp 1679581782
transform 1 0 52128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_544
timestamp 1679581782
transform 1 0 52800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_551
timestamp 1679581782
transform 1 0 53472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_558
timestamp 1679581782
transform 1 0 54144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_565
timestamp 1679581782
transform 1 0 54816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_572
timestamp 1679581782
transform 1 0 55488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_579
timestamp 1679581782
transform 1 0 56160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_586
timestamp 1679581782
transform 1 0 56832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_593
timestamp 1679581782
transform 1 0 57504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_600
timestamp 1679581782
transform 1 0 58176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_607
timestamp 1679581782
transform 1 0 58848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_614
timestamp 1679581782
transform 1 0 59520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_621
timestamp 1679581782
transform 1 0 60192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_628
timestamp 1679581782
transform 1 0 60864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_635
timestamp 1679581782
transform 1 0 61536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_642
timestamp 1679581782
transform 1 0 62208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_649
timestamp 1679581782
transform 1 0 62880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_656
timestamp 1679581782
transform 1 0 63552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_663
timestamp 1679581782
transform 1 0 64224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_670
timestamp 1679581782
transform 1 0 64896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_677
timestamp 1679581782
transform 1 0 65568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_684
timestamp 1679581782
transform 1 0 66240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_691
timestamp 1679581782
transform 1 0 66912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_698
timestamp 1679581782
transform 1 0 67584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_705
timestamp 1679581782
transform 1 0 68256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_712
timestamp 1679581782
transform 1 0 68928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_719
timestamp 1679581782
transform 1 0 69600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_726
timestamp 1679581782
transform 1 0 70272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_733
timestamp 1679581782
transform 1 0 70944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_740
timestamp 1679581782
transform 1 0 71616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_747
timestamp 1679581782
transform 1 0 72288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_754
timestamp 1679581782
transform 1 0 72960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_761
timestamp 1679581782
transform 1 0 73632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_768
timestamp 1679581782
transform 1 0 74304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_775
timestamp 1679581782
transform 1 0 74976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_782
timestamp 1679581782
transform 1 0 75648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_789
timestamp 1679581782
transform 1 0 76320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_796
timestamp 1679581782
transform 1 0 76992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_803
timestamp 1679581782
transform 1 0 77664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_810
timestamp 1679581782
transform 1 0 78336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_817
timestamp 1679581782
transform 1 0 79008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_824
timestamp 1679581782
transform 1 0 79680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_831
timestamp 1679581782
transform 1 0 80352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_838
timestamp 1679581782
transform 1 0 81024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_845
timestamp 1679581782
transform 1 0 81696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_852
timestamp 1679581782
transform 1 0 82368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_859
timestamp 1679581782
transform 1 0 83040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_866
timestamp 1679581782
transform 1 0 83712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_873
timestamp 1679581782
transform 1 0 84384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_880
timestamp 1679581782
transform 1 0 85056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_887
timestamp 1679581782
transform 1 0 85728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_894
timestamp 1679581782
transform 1 0 86400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_901
timestamp 1679581782
transform 1 0 87072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_908
timestamp 1679581782
transform 1 0 87744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_915
timestamp 1679581782
transform 1 0 88416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_922
timestamp 1679581782
transform 1 0 89088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_929
timestamp 1679581782
transform 1 0 89760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_936
timestamp 1679581782
transform 1 0 90432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_943
timestamp 1679581782
transform 1 0 91104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_950
timestamp 1679581782
transform 1 0 91776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_957
timestamp 1679581782
transform 1 0 92448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_964
timestamp 1679581782
transform 1 0 93120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_971
timestamp 1679581782
transform 1 0 93792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_978
timestamp 1679581782
transform 1 0 94464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_985
timestamp 1679581782
transform 1 0 95136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_992
timestamp 1679581782
transform 1 0 95808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_999
timestamp 1679581782
transform 1 0 96480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1006
timestamp 1679581782
transform 1 0 97152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1013
timestamp 1679581782
transform 1 0 97824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1020
timestamp 1679581782
transform 1 0 98496 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_1027
timestamp 1677580104
transform 1 0 99168 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_43_0
timestamp 1679577901
transform 1 0 576 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_4
timestamp 1677580104
transform 1 0 960 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_48
timestamp 1677580104
transform 1 0 5184 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_80
timestamp 1679581782
transform 1 0 8256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_87
timestamp 1679577901
transform 1 0 8928 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_138
timestamp 1677580104
transform 1 0 13824 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_158
timestamp 1677580104
transform 1 0 15744 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_160
timestamp 1677579658
transform 1 0 15936 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_182
timestamp 1677579658
transform 1 0 18048 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_43_228
timestamp 1679577901
transform 1 0 22464 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_269
timestamp 1677580104
transform 1 0 26400 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_43_281
timestamp 1679577901
transform 1 0 27552 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_285
timestamp 1677579658
transform 1 0 27936 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_307
timestamp 1679581782
transform 1 0 30048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_398
timestamp 1679581782
transform 1 0 38784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_405
timestamp 1679581782
transform 1 0 39456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_412
timestamp 1679581782
transform 1 0 40128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_419
timestamp 1679581782
transform 1 0 40800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_426
timestamp 1679581782
transform 1 0 41472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_433
timestamp 1679581782
transform 1 0 42144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_440
timestamp 1679581782
transform 1 0 42816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_447
timestamp 1679581782
transform 1 0 43488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_454
timestamp 1679581782
transform 1 0 44160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_461
timestamp 1679581782
transform 1 0 44832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_468
timestamp 1679581782
transform 1 0 45504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_475
timestamp 1679581782
transform 1 0 46176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_482
timestamp 1679581782
transform 1 0 46848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_489
timestamp 1679581782
transform 1 0 47520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_496
timestamp 1679581782
transform 1 0 48192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_503
timestamp 1679581782
transform 1 0 48864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_510
timestamp 1679581782
transform 1 0 49536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_517
timestamp 1679581782
transform 1 0 50208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_524
timestamp 1679581782
transform 1 0 50880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_531
timestamp 1679581782
transform 1 0 51552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_538
timestamp 1679581782
transform 1 0 52224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_545
timestamp 1679581782
transform 1 0 52896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_552
timestamp 1679581782
transform 1 0 53568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_559
timestamp 1679581782
transform 1 0 54240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_566
timestamp 1679581782
transform 1 0 54912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_573
timestamp 1679581782
transform 1 0 55584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_580
timestamp 1679581782
transform 1 0 56256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_587
timestamp 1679581782
transform 1 0 56928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_594
timestamp 1679581782
transform 1 0 57600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_601
timestamp 1679581782
transform 1 0 58272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_608
timestamp 1679581782
transform 1 0 58944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_615
timestamp 1679581782
transform 1 0 59616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_622
timestamp 1679581782
transform 1 0 60288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_629
timestamp 1679581782
transform 1 0 60960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_636
timestamp 1679581782
transform 1 0 61632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_643
timestamp 1679581782
transform 1 0 62304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_650
timestamp 1679581782
transform 1 0 62976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_657
timestamp 1679581782
transform 1 0 63648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_664
timestamp 1679581782
transform 1 0 64320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_671
timestamp 1679581782
transform 1 0 64992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_678
timestamp 1679581782
transform 1 0 65664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_685
timestamp 1679581782
transform 1 0 66336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_692
timestamp 1679581782
transform 1 0 67008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_699
timestamp 1679581782
transform 1 0 67680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_706
timestamp 1679581782
transform 1 0 68352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_713
timestamp 1679581782
transform 1 0 69024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_720
timestamp 1679581782
transform 1 0 69696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_727
timestamp 1679581782
transform 1 0 70368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_734
timestamp 1679581782
transform 1 0 71040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_741
timestamp 1679581782
transform 1 0 71712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_748
timestamp 1679581782
transform 1 0 72384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_755
timestamp 1679581782
transform 1 0 73056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_762
timestamp 1679581782
transform 1 0 73728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_769
timestamp 1679581782
transform 1 0 74400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_776
timestamp 1679581782
transform 1 0 75072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_783
timestamp 1679581782
transform 1 0 75744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_790
timestamp 1679581782
transform 1 0 76416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_797
timestamp 1679581782
transform 1 0 77088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_804
timestamp 1679581782
transform 1 0 77760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_811
timestamp 1679581782
transform 1 0 78432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_818
timestamp 1679581782
transform 1 0 79104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_825
timestamp 1679581782
transform 1 0 79776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_832
timestamp 1679581782
transform 1 0 80448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_839
timestamp 1679581782
transform 1 0 81120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_846
timestamp 1679581782
transform 1 0 81792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_853
timestamp 1679581782
transform 1 0 82464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_860
timestamp 1679581782
transform 1 0 83136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_867
timestamp 1679581782
transform 1 0 83808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_874
timestamp 1679581782
transform 1 0 84480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_881
timestamp 1679581782
transform 1 0 85152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_888
timestamp 1679581782
transform 1 0 85824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_895
timestamp 1679581782
transform 1 0 86496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_902
timestamp 1679581782
transform 1 0 87168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_909
timestamp 1679581782
transform 1 0 87840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_916
timestamp 1679581782
transform 1 0 88512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_923
timestamp 1679581782
transform 1 0 89184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_930
timestamp 1679581782
transform 1 0 89856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_937
timestamp 1679581782
transform 1 0 90528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_944
timestamp 1679581782
transform 1 0 91200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_951
timestamp 1679581782
transform 1 0 91872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_958
timestamp 1679581782
transform 1 0 92544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_965
timestamp 1679581782
transform 1 0 93216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_972
timestamp 1679581782
transform 1 0 93888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_979
timestamp 1679581782
transform 1 0 94560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_986
timestamp 1679581782
transform 1 0 95232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_993
timestamp 1679581782
transform 1 0 95904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1000
timestamp 1679581782
transform 1 0 96576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1007
timestamp 1679581782
transform 1 0 97248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1014
timestamp 1679581782
transform 1 0 97920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1021
timestamp 1679581782
transform 1 0 98592 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_1028
timestamp 1677579658
transform 1 0 99264 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_0
timestamp 1679577901
transform 1 0 576 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_4
timestamp 1677579658
transform 1 0 960 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_36
timestamp 1679577901
transform 1 0 4032 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_101
timestamp 1677579658
transform 1 0 10272 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_181
timestamp 1677579658
transform 1 0 17952 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_205
timestamp 1677580104
transform 1 0 20256 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_256
timestamp 1677580104
transform 1 0 25152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_258
timestamp 1677579658
transform 1 0 25344 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_325
timestamp 1679577901
transform 1 0 31776 0 1 34020
box -48 -56 432 834
use sg13g2_decap_4  FILLER_44_356
timestamp 1679577901
transform 1 0 34752 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_360
timestamp 1677579658
transform 1 0 35136 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_383
timestamp 1679577901
transform 1 0 37344 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_387
timestamp 1677580104
transform 1 0 37728 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_393
timestamp 1679581782
transform 1 0 38304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_400
timestamp 1679581782
transform 1 0 38976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_407
timestamp 1679581782
transform 1 0 39648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_414
timestamp 1679581782
transform 1 0 40320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_421
timestamp 1679581782
transform 1 0 40992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_428
timestamp 1679581782
transform 1 0 41664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_435
timestamp 1679581782
transform 1 0 42336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_442
timestamp 1679581782
transform 1 0 43008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_449
timestamp 1679581782
transform 1 0 43680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_456
timestamp 1679581782
transform 1 0 44352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_463
timestamp 1679581782
transform 1 0 45024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_470
timestamp 1679581782
transform 1 0 45696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_477
timestamp 1679581782
transform 1 0 46368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_484
timestamp 1679581782
transform 1 0 47040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_491
timestamp 1679581782
transform 1 0 47712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_498
timestamp 1679581782
transform 1 0 48384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_505
timestamp 1679581782
transform 1 0 49056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_512
timestamp 1679581782
transform 1 0 49728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_519
timestamp 1679581782
transform 1 0 50400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_526
timestamp 1679581782
transform 1 0 51072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_533
timestamp 1679581782
transform 1 0 51744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_540
timestamp 1679581782
transform 1 0 52416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_547
timestamp 1679581782
transform 1 0 53088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_554
timestamp 1679581782
transform 1 0 53760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_561
timestamp 1679581782
transform 1 0 54432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_568
timestamp 1679581782
transform 1 0 55104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_575
timestamp 1679581782
transform 1 0 55776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_582
timestamp 1679581782
transform 1 0 56448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_589
timestamp 1679581782
transform 1 0 57120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_596
timestamp 1679581782
transform 1 0 57792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_603
timestamp 1679581782
transform 1 0 58464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_610
timestamp 1679581782
transform 1 0 59136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_617
timestamp 1679581782
transform 1 0 59808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_624
timestamp 1679581782
transform 1 0 60480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_631
timestamp 1679581782
transform 1 0 61152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_638
timestamp 1679581782
transform 1 0 61824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_645
timestamp 1679581782
transform 1 0 62496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_652
timestamp 1679581782
transform 1 0 63168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_659
timestamp 1679581782
transform 1 0 63840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_666
timestamp 1679581782
transform 1 0 64512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_673
timestamp 1679581782
transform 1 0 65184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_680
timestamp 1679581782
transform 1 0 65856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_687
timestamp 1679581782
transform 1 0 66528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_694
timestamp 1679581782
transform 1 0 67200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_701
timestamp 1679581782
transform 1 0 67872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_708
timestamp 1679581782
transform 1 0 68544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_715
timestamp 1679581782
transform 1 0 69216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_722
timestamp 1679581782
transform 1 0 69888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_729
timestamp 1679581782
transform 1 0 70560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_736
timestamp 1679581782
transform 1 0 71232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_743
timestamp 1679581782
transform 1 0 71904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_750
timestamp 1679581782
transform 1 0 72576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_757
timestamp 1679581782
transform 1 0 73248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_764
timestamp 1679581782
transform 1 0 73920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_771
timestamp 1679581782
transform 1 0 74592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_778
timestamp 1679581782
transform 1 0 75264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_785
timestamp 1679581782
transform 1 0 75936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_792
timestamp 1679581782
transform 1 0 76608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_799
timestamp 1679581782
transform 1 0 77280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_806
timestamp 1679581782
transform 1 0 77952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_813
timestamp 1679581782
transform 1 0 78624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_820
timestamp 1679581782
transform 1 0 79296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_827
timestamp 1679581782
transform 1 0 79968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_834
timestamp 1679581782
transform 1 0 80640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_841
timestamp 1679581782
transform 1 0 81312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_848
timestamp 1679581782
transform 1 0 81984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_855
timestamp 1679581782
transform 1 0 82656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_862
timestamp 1679581782
transform 1 0 83328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_869
timestamp 1679581782
transform 1 0 84000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_876
timestamp 1679581782
transform 1 0 84672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_883
timestamp 1679581782
transform 1 0 85344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_890
timestamp 1679581782
transform 1 0 86016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_897
timestamp 1679581782
transform 1 0 86688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_904
timestamp 1679581782
transform 1 0 87360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_911
timestamp 1679581782
transform 1 0 88032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_918
timestamp 1679581782
transform 1 0 88704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_925
timestamp 1679581782
transform 1 0 89376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_932
timestamp 1679581782
transform 1 0 90048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_939
timestamp 1679581782
transform 1 0 90720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_946
timestamp 1679581782
transform 1 0 91392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_953
timestamp 1679581782
transform 1 0 92064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_960
timestamp 1679581782
transform 1 0 92736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_967
timestamp 1679581782
transform 1 0 93408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_974
timestamp 1679581782
transform 1 0 94080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_981
timestamp 1679581782
transform 1 0 94752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_988
timestamp 1679581782
transform 1 0 95424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_995
timestamp 1679581782
transform 1 0 96096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1002
timestamp 1679581782
transform 1 0 96768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1009
timestamp 1679581782
transform 1 0 97440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1016
timestamp 1679581782
transform 1 0 98112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_1023
timestamp 1679577901
transform 1 0 98784 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_1027
timestamp 1677580104
transform 1 0 99168 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_18
timestamp 1679581782
transform 1 0 2304 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_25
timestamp 1677580104
transform 1 0 2976 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_125
timestamp 1679577901
transform 1 0 12576 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_138
timestamp 1677580104
transform 1 0 13824 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_149
timestamp 1677580104
transform 1 0 14880 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_164
timestamp 1677580104
transform 1 0 16320 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_212
timestamp 1677579658
transform 1 0 20928 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_226
timestamp 1679581782
transform 1 0 22272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_233
timestamp 1679577901
transform 1 0 22944 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_246
timestamp 1679581782
transform 1 0 24192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_253
timestamp 1679581782
transform 1 0 24864 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_260
timestamp 1677580104
transform 1 0 25536 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_275
timestamp 1679581782
transform 1 0 26976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_282
timestamp 1679581782
transform 1 0 27648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_289
timestamp 1679581782
transform 1 0 28320 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_296
timestamp 1677579658
transform 1 0 28992 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_310
timestamp 1679581782
transform 1 0 30336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_317
timestamp 1679577901
transform 1 0 31008 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_4  FILLER_45_330
timestamp 1679577901
transform 1 0 32256 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_338
timestamp 1679581782
transform 1 0 33024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_345
timestamp 1679581782
transform 1 0 33696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_352
timestamp 1679581782
transform 1 0 34368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_359
timestamp 1679581782
transform 1 0 35040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_366
timestamp 1679581782
transform 1 0 35712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_373
timestamp 1679581782
transform 1 0 36384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_380
timestamp 1679581782
transform 1 0 37056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_387
timestamp 1679581782
transform 1 0 37728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_394
timestamp 1679581782
transform 1 0 38400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_401
timestamp 1679581782
transform 1 0 39072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_408
timestamp 1679581782
transform 1 0 39744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_415
timestamp 1679581782
transform 1 0 40416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_422
timestamp 1679581782
transform 1 0 41088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_429
timestamp 1679581782
transform 1 0 41760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_436
timestamp 1679581782
transform 1 0 42432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_443
timestamp 1679581782
transform 1 0 43104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_450
timestamp 1679581782
transform 1 0 43776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_457
timestamp 1679581782
transform 1 0 44448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_464
timestamp 1679581782
transform 1 0 45120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_471
timestamp 1679581782
transform 1 0 45792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_478
timestamp 1679581782
transform 1 0 46464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_485
timestamp 1679581782
transform 1 0 47136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_492
timestamp 1679581782
transform 1 0 47808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_499
timestamp 1679581782
transform 1 0 48480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_506
timestamp 1679581782
transform 1 0 49152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_513
timestamp 1679581782
transform 1 0 49824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_520
timestamp 1679581782
transform 1 0 50496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_527
timestamp 1679581782
transform 1 0 51168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_534
timestamp 1679581782
transform 1 0 51840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_541
timestamp 1679581782
transform 1 0 52512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_548
timestamp 1679581782
transform 1 0 53184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_555
timestamp 1679581782
transform 1 0 53856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_562
timestamp 1679581782
transform 1 0 54528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_569
timestamp 1679581782
transform 1 0 55200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_576
timestamp 1679581782
transform 1 0 55872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_583
timestamp 1679581782
transform 1 0 56544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_590
timestamp 1679581782
transform 1 0 57216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_597
timestamp 1679581782
transform 1 0 57888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_604
timestamp 1679581782
transform 1 0 58560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_611
timestamp 1679581782
transform 1 0 59232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_618
timestamp 1679581782
transform 1 0 59904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_625
timestamp 1679581782
transform 1 0 60576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_632
timestamp 1679581782
transform 1 0 61248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_639
timestamp 1679581782
transform 1 0 61920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_646
timestamp 1679581782
transform 1 0 62592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_653
timestamp 1679581782
transform 1 0 63264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_660
timestamp 1679581782
transform 1 0 63936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_667
timestamp 1679581782
transform 1 0 64608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_674
timestamp 1679581782
transform 1 0 65280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_681
timestamp 1679581782
transform 1 0 65952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_688
timestamp 1679581782
transform 1 0 66624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_695
timestamp 1679581782
transform 1 0 67296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_702
timestamp 1679581782
transform 1 0 67968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_709
timestamp 1679581782
transform 1 0 68640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_716
timestamp 1679581782
transform 1 0 69312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_723
timestamp 1679581782
transform 1 0 69984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_730
timestamp 1679581782
transform 1 0 70656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_737
timestamp 1679581782
transform 1 0 71328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_744
timestamp 1679581782
transform 1 0 72000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_751
timestamp 1679581782
transform 1 0 72672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_758
timestamp 1679581782
transform 1 0 73344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_765
timestamp 1679581782
transform 1 0 74016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_772
timestamp 1679581782
transform 1 0 74688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_779
timestamp 1679581782
transform 1 0 75360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_786
timestamp 1679581782
transform 1 0 76032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_793
timestamp 1679581782
transform 1 0 76704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_800
timestamp 1679581782
transform 1 0 77376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_807
timestamp 1679581782
transform 1 0 78048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_814
timestamp 1679581782
transform 1 0 78720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_821
timestamp 1679581782
transform 1 0 79392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_828
timestamp 1679581782
transform 1 0 80064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_835
timestamp 1679581782
transform 1 0 80736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_842
timestamp 1679581782
transform 1 0 81408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_849
timestamp 1679581782
transform 1 0 82080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_856
timestamp 1679581782
transform 1 0 82752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_863
timestamp 1679581782
transform 1 0 83424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_870
timestamp 1679581782
transform 1 0 84096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_877
timestamp 1679581782
transform 1 0 84768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_884
timestamp 1679581782
transform 1 0 85440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_891
timestamp 1679581782
transform 1 0 86112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_898
timestamp 1679581782
transform 1 0 86784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_905
timestamp 1679581782
transform 1 0 87456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_912
timestamp 1679581782
transform 1 0 88128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_919
timestamp 1679581782
transform 1 0 88800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_926
timestamp 1679581782
transform 1 0 89472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_933
timestamp 1679581782
transform 1 0 90144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_940
timestamp 1679581782
transform 1 0 90816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_947
timestamp 1679581782
transform 1 0 91488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_954
timestamp 1679581782
transform 1 0 92160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_961
timestamp 1679581782
transform 1 0 92832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_968
timestamp 1679581782
transform 1 0 93504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_975
timestamp 1679581782
transform 1 0 94176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_982
timestamp 1679581782
transform 1 0 94848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_989
timestamp 1679581782
transform 1 0 95520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_996
timestamp 1679581782
transform 1 0 96192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1003
timestamp 1679581782
transform 1 0 96864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1010
timestamp 1679581782
transform 1 0 97536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1017
timestamp 1679581782
transform 1 0 98208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_1024
timestamp 1679577901
transform 1 0 98880 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_1028
timestamp 1677579658
transform 1 0 99264 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_28
timestamp 1679577901
transform 1 0 3264 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_32
timestamp 1677580104
transform 1 0 3648 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_61
timestamp 1677579658
transform 1 0 6432 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_76
timestamp 1677579658
transform 1 0 7872 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_111
timestamp 1677580104
transform 1 0 11232 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_155
timestamp 1677579658
transform 1 0 15456 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_183
timestamp 1677579658
transform 1 0 18144 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_197
timestamp 1679581782
transform 1 0 19488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_204
timestamp 1679581782
transform 1 0 20160 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_211
timestamp 1677580104
transform 1 0 20832 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_216
timestamp 1679581782
transform 1 0 21312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_223
timestamp 1679581782
transform 1 0 21984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_230
timestamp 1679581782
transform 1 0 22656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_237
timestamp 1679581782
transform 1 0 23328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_244
timestamp 1679581782
transform 1 0 24000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_251
timestamp 1679581782
transform 1 0 24672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_258
timestamp 1679581782
transform 1 0 25344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_265
timestamp 1679581782
transform 1 0 26016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_272
timestamp 1679581782
transform 1 0 26688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_279
timestamp 1679581782
transform 1 0 27360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_286
timestamp 1679581782
transform 1 0 28032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_293
timestamp 1679581782
transform 1 0 28704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_300
timestamp 1679581782
transform 1 0 29376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_307
timestamp 1679581782
transform 1 0 30048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_314
timestamp 1679581782
transform 1 0 30720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_321
timestamp 1679581782
transform 1 0 31392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_328
timestamp 1679581782
transform 1 0 32064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_335
timestamp 1679581782
transform 1 0 32736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_342
timestamp 1679581782
transform 1 0 33408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_349
timestamp 1679581782
transform 1 0 34080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_356
timestamp 1679581782
transform 1 0 34752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_363
timestamp 1679581782
transform 1 0 35424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_370
timestamp 1679581782
transform 1 0 36096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_377
timestamp 1679581782
transform 1 0 36768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_384
timestamp 1679581782
transform 1 0 37440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_391
timestamp 1679581782
transform 1 0 38112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_398
timestamp 1679581782
transform 1 0 38784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_405
timestamp 1679581782
transform 1 0 39456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_412
timestamp 1679581782
transform 1 0 40128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_419
timestamp 1679581782
transform 1 0 40800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_426
timestamp 1679581782
transform 1 0 41472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_433
timestamp 1679581782
transform 1 0 42144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_440
timestamp 1679581782
transform 1 0 42816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_447
timestamp 1679581782
transform 1 0 43488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_454
timestamp 1679581782
transform 1 0 44160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_461
timestamp 1679581782
transform 1 0 44832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_468
timestamp 1679581782
transform 1 0 45504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_475
timestamp 1679581782
transform 1 0 46176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_482
timestamp 1679581782
transform 1 0 46848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_489
timestamp 1679581782
transform 1 0 47520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_496
timestamp 1679581782
transform 1 0 48192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_503
timestamp 1679581782
transform 1 0 48864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_510
timestamp 1679581782
transform 1 0 49536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_517
timestamp 1679581782
transform 1 0 50208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_524
timestamp 1679581782
transform 1 0 50880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_531
timestamp 1679581782
transform 1 0 51552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_538
timestamp 1679581782
transform 1 0 52224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_545
timestamp 1679581782
transform 1 0 52896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_552
timestamp 1679581782
transform 1 0 53568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_559
timestamp 1679581782
transform 1 0 54240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_566
timestamp 1679581782
transform 1 0 54912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_573
timestamp 1679581782
transform 1 0 55584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_580
timestamp 1679581782
transform 1 0 56256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_587
timestamp 1679581782
transform 1 0 56928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_594
timestamp 1679581782
transform 1 0 57600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_601
timestamp 1679581782
transform 1 0 58272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_608
timestamp 1679581782
transform 1 0 58944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_615
timestamp 1679581782
transform 1 0 59616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_622
timestamp 1679581782
transform 1 0 60288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_629
timestamp 1679581782
transform 1 0 60960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_636
timestamp 1679581782
transform 1 0 61632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_643
timestamp 1679581782
transform 1 0 62304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_650
timestamp 1679581782
transform 1 0 62976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_657
timestamp 1679581782
transform 1 0 63648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_664
timestamp 1679581782
transform 1 0 64320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_671
timestamp 1679581782
transform 1 0 64992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_678
timestamp 1679581782
transform 1 0 65664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_685
timestamp 1679581782
transform 1 0 66336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_692
timestamp 1679581782
transform 1 0 67008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_699
timestamp 1679581782
transform 1 0 67680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_706
timestamp 1679581782
transform 1 0 68352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_713
timestamp 1679581782
transform 1 0 69024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_720
timestamp 1679581782
transform 1 0 69696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_727
timestamp 1679581782
transform 1 0 70368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_734
timestamp 1679581782
transform 1 0 71040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_741
timestamp 1679581782
transform 1 0 71712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_748
timestamp 1679581782
transform 1 0 72384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_755
timestamp 1679581782
transform 1 0 73056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_762
timestamp 1679581782
transform 1 0 73728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_769
timestamp 1679581782
transform 1 0 74400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_776
timestamp 1679581782
transform 1 0 75072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_783
timestamp 1679581782
transform 1 0 75744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_790
timestamp 1679581782
transform 1 0 76416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_797
timestamp 1679581782
transform 1 0 77088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_804
timestamp 1679581782
transform 1 0 77760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_811
timestamp 1679581782
transform 1 0 78432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_818
timestamp 1679581782
transform 1 0 79104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_825
timestamp 1679581782
transform 1 0 79776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_832
timestamp 1679581782
transform 1 0 80448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_839
timestamp 1679581782
transform 1 0 81120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_846
timestamp 1679581782
transform 1 0 81792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_853
timestamp 1679581782
transform 1 0 82464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_860
timestamp 1679581782
transform 1 0 83136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_867
timestamp 1679581782
transform 1 0 83808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_874
timestamp 1679581782
transform 1 0 84480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_881
timestamp 1679581782
transform 1 0 85152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_888
timestamp 1679581782
transform 1 0 85824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_895
timestamp 1679581782
transform 1 0 86496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_902
timestamp 1679581782
transform 1 0 87168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_909
timestamp 1679581782
transform 1 0 87840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_916
timestamp 1679581782
transform 1 0 88512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_923
timestamp 1679581782
transform 1 0 89184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_930
timestamp 1679581782
transform 1 0 89856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_937
timestamp 1679581782
transform 1 0 90528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_944
timestamp 1679581782
transform 1 0 91200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_951
timestamp 1679581782
transform 1 0 91872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_958
timestamp 1679581782
transform 1 0 92544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_965
timestamp 1679581782
transform 1 0 93216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_972
timestamp 1679581782
transform 1 0 93888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_979
timestamp 1679581782
transform 1 0 94560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_986
timestamp 1679581782
transform 1 0 95232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_993
timestamp 1679581782
transform 1 0 95904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1000
timestamp 1679581782
transform 1 0 96576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1007
timestamp 1679581782
transform 1 0 97248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1014
timestamp 1679581782
transform 1 0 97920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1021
timestamp 1679581782
transform 1 0 98592 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_1028
timestamp 1677579658
transform 1 0 99264 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_35
timestamp 1677580104
transform 1 0 3936 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_37
timestamp 1677579658
transform 1 0 4128 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_46
timestamp 1679581782
transform 1 0 4992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_53
timestamp 1679581782
transform 1 0 5664 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_60
timestamp 1677579658
transform 1 0 6336 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_95
timestamp 1677580104
transform 1 0 9696 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_106
timestamp 1677580104
transform 1 0 10752 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_108
timestamp 1677579658
transform 1 0 10944 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_114
timestamp 1677580104
transform 1 0 11520 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_129
timestamp 1679581782
transform 1 0 12960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_136
timestamp 1679581782
transform 1 0 13632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_143
timestamp 1679577901
transform 1 0 14304 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_147
timestamp 1677579658
transform 1 0 14688 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_151
timestamp 1677580104
transform 1 0 15072 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_179
timestamp 1679581782
transform 1 0 17760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_186
timestamp 1679581782
transform 1 0 18432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_193
timestamp 1679581782
transform 1 0 19104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_200
timestamp 1679581782
transform 1 0 19776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_207
timestamp 1679581782
transform 1 0 20448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_214
timestamp 1679581782
transform 1 0 21120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_221
timestamp 1679581782
transform 1 0 21792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_228
timestamp 1679581782
transform 1 0 22464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_235
timestamp 1679581782
transform 1 0 23136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_242
timestamp 1679581782
transform 1 0 23808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_249
timestamp 1679581782
transform 1 0 24480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_256
timestamp 1679581782
transform 1 0 25152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_263
timestamp 1679581782
transform 1 0 25824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_270
timestamp 1679581782
transform 1 0 26496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_277
timestamp 1679581782
transform 1 0 27168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_284
timestamp 1679581782
transform 1 0 27840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_291
timestamp 1679581782
transform 1 0 28512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_298
timestamp 1679581782
transform 1 0 29184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_305
timestamp 1679581782
transform 1 0 29856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_312
timestamp 1679581782
transform 1 0 30528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_319
timestamp 1679581782
transform 1 0 31200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_326
timestamp 1679581782
transform 1 0 31872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_333
timestamp 1679581782
transform 1 0 32544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_340
timestamp 1679581782
transform 1 0 33216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_347
timestamp 1679581782
transform 1 0 33888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_354
timestamp 1679581782
transform 1 0 34560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_361
timestamp 1679581782
transform 1 0 35232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_368
timestamp 1679581782
transform 1 0 35904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_375
timestamp 1679581782
transform 1 0 36576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_382
timestamp 1679581782
transform 1 0 37248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_389
timestamp 1679581782
transform 1 0 37920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_396
timestamp 1679581782
transform 1 0 38592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_403
timestamp 1679581782
transform 1 0 39264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_410
timestamp 1679581782
transform 1 0 39936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_417
timestamp 1679581782
transform 1 0 40608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_424
timestamp 1679581782
transform 1 0 41280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_431
timestamp 1679581782
transform 1 0 41952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_438
timestamp 1679581782
transform 1 0 42624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_445
timestamp 1679581782
transform 1 0 43296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_452
timestamp 1679581782
transform 1 0 43968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_459
timestamp 1679581782
transform 1 0 44640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_466
timestamp 1679581782
transform 1 0 45312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_473
timestamp 1679581782
transform 1 0 45984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_480
timestamp 1679581782
transform 1 0 46656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_487
timestamp 1679581782
transform 1 0 47328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_494
timestamp 1679581782
transform 1 0 48000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_501
timestamp 1679581782
transform 1 0 48672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_508
timestamp 1679581782
transform 1 0 49344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_515
timestamp 1679581782
transform 1 0 50016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_522
timestamp 1679581782
transform 1 0 50688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_529
timestamp 1679581782
transform 1 0 51360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_536
timestamp 1679581782
transform 1 0 52032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_543
timestamp 1679581782
transform 1 0 52704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_550
timestamp 1679581782
transform 1 0 53376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_557
timestamp 1679581782
transform 1 0 54048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_564
timestamp 1679581782
transform 1 0 54720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_571
timestamp 1679581782
transform 1 0 55392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_578
timestamp 1679581782
transform 1 0 56064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_585
timestamp 1679581782
transform 1 0 56736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_592
timestamp 1679581782
transform 1 0 57408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_599
timestamp 1679581782
transform 1 0 58080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_606
timestamp 1679581782
transform 1 0 58752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_613
timestamp 1679581782
transform 1 0 59424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_620
timestamp 1679581782
transform 1 0 60096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_627
timestamp 1679581782
transform 1 0 60768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_634
timestamp 1679581782
transform 1 0 61440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_641
timestamp 1679581782
transform 1 0 62112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_648
timestamp 1679581782
transform 1 0 62784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_655
timestamp 1679581782
transform 1 0 63456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_662
timestamp 1679581782
transform 1 0 64128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_669
timestamp 1679581782
transform 1 0 64800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_676
timestamp 1679581782
transform 1 0 65472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_683
timestamp 1679581782
transform 1 0 66144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_690
timestamp 1679581782
transform 1 0 66816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_697
timestamp 1679581782
transform 1 0 67488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_704
timestamp 1679581782
transform 1 0 68160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_711
timestamp 1679581782
transform 1 0 68832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_718
timestamp 1679581782
transform 1 0 69504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_725
timestamp 1679581782
transform 1 0 70176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_732
timestamp 1679581782
transform 1 0 70848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_739
timestamp 1679581782
transform 1 0 71520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_746
timestamp 1679581782
transform 1 0 72192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_753
timestamp 1679581782
transform 1 0 72864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_760
timestamp 1679581782
transform 1 0 73536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_767
timestamp 1679581782
transform 1 0 74208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_774
timestamp 1679581782
transform 1 0 74880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_781
timestamp 1679581782
transform 1 0 75552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_788
timestamp 1679581782
transform 1 0 76224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_795
timestamp 1679581782
transform 1 0 76896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_802
timestamp 1679581782
transform 1 0 77568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_809
timestamp 1679581782
transform 1 0 78240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_816
timestamp 1679581782
transform 1 0 78912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_823
timestamp 1679581782
transform 1 0 79584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_830
timestamp 1679581782
transform 1 0 80256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_837
timestamp 1679581782
transform 1 0 80928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_844
timestamp 1679581782
transform 1 0 81600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_851
timestamp 1679581782
transform 1 0 82272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_858
timestamp 1679581782
transform 1 0 82944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_865
timestamp 1679581782
transform 1 0 83616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_872
timestamp 1679581782
transform 1 0 84288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_879
timestamp 1679581782
transform 1 0 84960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_886
timestamp 1679581782
transform 1 0 85632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_893
timestamp 1679581782
transform 1 0 86304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_900
timestamp 1679581782
transform 1 0 86976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_907
timestamp 1679581782
transform 1 0 87648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_914
timestamp 1679581782
transform 1 0 88320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_921
timestamp 1679581782
transform 1 0 88992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_928
timestamp 1679581782
transform 1 0 89664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_935
timestamp 1679581782
transform 1 0 90336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_942
timestamp 1679581782
transform 1 0 91008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_949
timestamp 1679581782
transform 1 0 91680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_956
timestamp 1679581782
transform 1 0 92352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_963
timestamp 1679581782
transform 1 0 93024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_970
timestamp 1679581782
transform 1 0 93696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_977
timestamp 1679581782
transform 1 0 94368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_984
timestamp 1679581782
transform 1 0 95040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_991
timestamp 1679581782
transform 1 0 95712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_998
timestamp 1679581782
transform 1 0 96384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1005
timestamp 1679581782
transform 1 0 97056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1012
timestamp 1679581782
transform 1 0 97728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1019
timestamp 1679581782
transform 1 0 98400 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_1026
timestamp 1677580104
transform 1 0 99072 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_1028
timestamp 1677579658
transform 1 0 99264 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_63
timestamp 1677580104
transform 1 0 6624 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_65
timestamp 1677579658
transform 1 0 6816 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_69
timestamp 1677580104
transform 1 0 7200 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_101
timestamp 1677579658
transform 1 0 10272 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_129
timestamp 1679581782
transform 1 0 12960 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_136
timestamp 1677580104
transform 1 0 13632 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_138
timestamp 1677579658
transform 1 0 13824 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_148
timestamp 1679581782
transform 1 0 14784 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_155
timestamp 1677580104
transform 1 0 15456 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_166
timestamp 1679581782
transform 1 0 16512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_173
timestamp 1679581782
transform 1 0 17184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_180
timestamp 1679581782
transform 1 0 17856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_187
timestamp 1679581782
transform 1 0 18528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_194
timestamp 1679581782
transform 1 0 19200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_201
timestamp 1679581782
transform 1 0 19872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_208
timestamp 1679581782
transform 1 0 20544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_215
timestamp 1679581782
transform 1 0 21216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_222
timestamp 1679581782
transform 1 0 21888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_229
timestamp 1679581782
transform 1 0 22560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_236
timestamp 1679581782
transform 1 0 23232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_243
timestamp 1679581782
transform 1 0 23904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_250
timestamp 1679581782
transform 1 0 24576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_257
timestamp 1679581782
transform 1 0 25248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_264
timestamp 1679581782
transform 1 0 25920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_271
timestamp 1679581782
transform 1 0 26592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_278
timestamp 1679581782
transform 1 0 27264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_285
timestamp 1679581782
transform 1 0 27936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_292
timestamp 1679581782
transform 1 0 28608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_299
timestamp 1679581782
transform 1 0 29280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_306
timestamp 1679581782
transform 1 0 29952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_313
timestamp 1679581782
transform 1 0 30624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_320
timestamp 1679581782
transform 1 0 31296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_327
timestamp 1679581782
transform 1 0 31968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_334
timestamp 1679581782
transform 1 0 32640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_341
timestamp 1679581782
transform 1 0 33312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_348
timestamp 1679581782
transform 1 0 33984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_355
timestamp 1679581782
transform 1 0 34656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_362
timestamp 1679581782
transform 1 0 35328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_369
timestamp 1679581782
transform 1 0 36000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_376
timestamp 1679581782
transform 1 0 36672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_383
timestamp 1679581782
transform 1 0 37344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_390
timestamp 1679581782
transform 1 0 38016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_397
timestamp 1679581782
transform 1 0 38688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_404
timestamp 1679581782
transform 1 0 39360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_411
timestamp 1679581782
transform 1 0 40032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_418
timestamp 1679581782
transform 1 0 40704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_425
timestamp 1679581782
transform 1 0 41376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_432
timestamp 1679581782
transform 1 0 42048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_439
timestamp 1679581782
transform 1 0 42720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_446
timestamp 1679581782
transform 1 0 43392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_453
timestamp 1679581782
transform 1 0 44064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_460
timestamp 1679581782
transform 1 0 44736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_467
timestamp 1679581782
transform 1 0 45408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_474
timestamp 1679581782
transform 1 0 46080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_481
timestamp 1679581782
transform 1 0 46752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_488
timestamp 1679581782
transform 1 0 47424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_495
timestamp 1679581782
transform 1 0 48096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_502
timestamp 1679581782
transform 1 0 48768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_509
timestamp 1679581782
transform 1 0 49440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_516
timestamp 1679581782
transform 1 0 50112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_523
timestamp 1679581782
transform 1 0 50784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_530
timestamp 1679581782
transform 1 0 51456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_537
timestamp 1679581782
transform 1 0 52128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_544
timestamp 1679581782
transform 1 0 52800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_551
timestamp 1679581782
transform 1 0 53472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_558
timestamp 1679581782
transform 1 0 54144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_565
timestamp 1679581782
transform 1 0 54816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_572
timestamp 1679581782
transform 1 0 55488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_579
timestamp 1679581782
transform 1 0 56160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_586
timestamp 1679581782
transform 1 0 56832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_593
timestamp 1679581782
transform 1 0 57504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_600
timestamp 1679581782
transform 1 0 58176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_607
timestamp 1679581782
transform 1 0 58848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_614
timestamp 1679581782
transform 1 0 59520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_621
timestamp 1679581782
transform 1 0 60192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_628
timestamp 1679581782
transform 1 0 60864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_635
timestamp 1679581782
transform 1 0 61536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_642
timestamp 1679581782
transform 1 0 62208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_649
timestamp 1679581782
transform 1 0 62880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_656
timestamp 1679581782
transform 1 0 63552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_663
timestamp 1679581782
transform 1 0 64224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_670
timestamp 1679581782
transform 1 0 64896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_677
timestamp 1679581782
transform 1 0 65568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_684
timestamp 1679581782
transform 1 0 66240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_691
timestamp 1679581782
transform 1 0 66912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_698
timestamp 1679581782
transform 1 0 67584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_705
timestamp 1679581782
transform 1 0 68256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_712
timestamp 1679581782
transform 1 0 68928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_719
timestamp 1679581782
transform 1 0 69600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_726
timestamp 1679581782
transform 1 0 70272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_733
timestamp 1679581782
transform 1 0 70944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_740
timestamp 1679581782
transform 1 0 71616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_747
timestamp 1679581782
transform 1 0 72288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_754
timestamp 1679581782
transform 1 0 72960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_761
timestamp 1679581782
transform 1 0 73632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_768
timestamp 1679581782
transform 1 0 74304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_775
timestamp 1679581782
transform 1 0 74976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_782
timestamp 1679581782
transform 1 0 75648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_789
timestamp 1679581782
transform 1 0 76320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_796
timestamp 1679581782
transform 1 0 76992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_803
timestamp 1679581782
transform 1 0 77664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_810
timestamp 1679581782
transform 1 0 78336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_817
timestamp 1679581782
transform 1 0 79008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_824
timestamp 1679581782
transform 1 0 79680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_831
timestamp 1679581782
transform 1 0 80352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_838
timestamp 1679581782
transform 1 0 81024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_845
timestamp 1679581782
transform 1 0 81696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_852
timestamp 1679581782
transform 1 0 82368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_859
timestamp 1679581782
transform 1 0 83040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_866
timestamp 1679581782
transform 1 0 83712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_873
timestamp 1679581782
transform 1 0 84384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_880
timestamp 1679581782
transform 1 0 85056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_887
timestamp 1679581782
transform 1 0 85728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_894
timestamp 1679581782
transform 1 0 86400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_901
timestamp 1679581782
transform 1 0 87072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_908
timestamp 1679581782
transform 1 0 87744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_915
timestamp 1679581782
transform 1 0 88416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_922
timestamp 1679581782
transform 1 0 89088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_929
timestamp 1679581782
transform 1 0 89760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_936
timestamp 1679581782
transform 1 0 90432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_943
timestamp 1679581782
transform 1 0 91104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_950
timestamp 1679581782
transform 1 0 91776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_957
timestamp 1679581782
transform 1 0 92448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_964
timestamp 1679581782
transform 1 0 93120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_971
timestamp 1679581782
transform 1 0 93792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_978
timestamp 1679581782
transform 1 0 94464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_985
timestamp 1679581782
transform 1 0 95136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_992
timestamp 1679581782
transform 1 0 95808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_999
timestamp 1679581782
transform 1 0 96480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1006
timestamp 1679581782
transform 1 0 97152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1013
timestamp 1679581782
transform 1 0 97824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1020
timestamp 1679581782
transform 1 0 98496 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_1027
timestamp 1677580104
transform 1 0 99168 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_88
timestamp 1679577901
transform 1 0 9024 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_92
timestamp 1677579658
transform 1 0 9408 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_578
timestamp 1679581782
transform 1 0 56064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_585
timestamp 1679581782
transform 1 0 56736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_592
timestamp 1679581782
transform 1 0 57408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_599
timestamp 1679581782
transform 1 0 58080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_606
timestamp 1679581782
transform 1 0 58752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_613
timestamp 1679581782
transform 1 0 59424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679581782
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_627
timestamp 1679581782
transform 1 0 60768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_634
timestamp 1679581782
transform 1 0 61440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_641
timestamp 1679581782
transform 1 0 62112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_648
timestamp 1679581782
transform 1 0 62784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_655
timestamp 1679581782
transform 1 0 63456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_662
timestamp 1679581782
transform 1 0 64128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_669
timestamp 1679581782
transform 1 0 64800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_676
timestamp 1679581782
transform 1 0 65472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_683
timestamp 1679581782
transform 1 0 66144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_690
timestamp 1679581782
transform 1 0 66816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_697
timestamp 1679581782
transform 1 0 67488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_704
timestamp 1679581782
transform 1 0 68160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_711
timestamp 1679581782
transform 1 0 68832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_718
timestamp 1679581782
transform 1 0 69504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_725
timestamp 1679581782
transform 1 0 70176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_732
timestamp 1679581782
transform 1 0 70848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_739
timestamp 1679581782
transform 1 0 71520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_746
timestamp 1679581782
transform 1 0 72192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_753
timestamp 1679581782
transform 1 0 72864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_760
timestamp 1679581782
transform 1 0 73536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_767
timestamp 1679581782
transform 1 0 74208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_774
timestamp 1679581782
transform 1 0 74880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_781
timestamp 1679581782
transform 1 0 75552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_788
timestamp 1679581782
transform 1 0 76224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_795
timestamp 1679581782
transform 1 0 76896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_802
timestamp 1679581782
transform 1 0 77568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_809
timestamp 1679581782
transform 1 0 78240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_816
timestamp 1679581782
transform 1 0 78912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_823
timestamp 1679581782
transform 1 0 79584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_830
timestamp 1679581782
transform 1 0 80256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_837
timestamp 1679581782
transform 1 0 80928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_844
timestamp 1679581782
transform 1 0 81600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_851
timestamp 1679581782
transform 1 0 82272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_858
timestamp 1679581782
transform 1 0 82944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_865
timestamp 1679581782
transform 1 0 83616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_872
timestamp 1679581782
transform 1 0 84288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_879
timestamp 1679581782
transform 1 0 84960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_886
timestamp 1679581782
transform 1 0 85632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_893
timestamp 1679581782
transform 1 0 86304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_900
timestamp 1679581782
transform 1 0 86976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_907
timestamp 1679581782
transform 1 0 87648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_914
timestamp 1679581782
transform 1 0 88320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_921
timestamp 1679581782
transform 1 0 88992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_928
timestamp 1679581782
transform 1 0 89664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_935
timestamp 1679581782
transform 1 0 90336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_942
timestamp 1679581782
transform 1 0 91008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_949
timestamp 1679581782
transform 1 0 91680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_956
timestamp 1679581782
transform 1 0 92352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_963
timestamp 1679581782
transform 1 0 93024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_970
timestamp 1679581782
transform 1 0 93696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_977
timestamp 1679581782
transform 1 0 94368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_984
timestamp 1679581782
transform 1 0 95040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_991
timestamp 1679581782
transform 1 0 95712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_998
timestamp 1679581782
transform 1 0 96384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1005
timestamp 1679581782
transform 1 0 97056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1012
timestamp 1679581782
transform 1 0 97728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1019
timestamp 1679581782
transform 1 0 98400 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_1026
timestamp 1677580104
transform 1 0 99072 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_1028
timestamp 1677579658
transform 1 0 99264 0 -1 38556
box -48 -56 144 834
use sg13g2_tielo  heichips25_ppwm_3
timestamp 1680000637
transform -1 0 1056 0 -1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_4
timestamp 1680000637
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_5
timestamp 1680000637
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_6
timestamp 1680000637
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_7
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_8
timestamp 1680000637
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_9
timestamp 1680000637
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_10
timestamp 1680000637
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_11
timestamp 1680000637
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_12
timestamp 1680000637
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_13
timestamp 1680000637
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_14
timestamp 1680000637
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_15
timestamp 1680000637
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_16
timestamp 1680000637
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_17
timestamp 1680000637
transform -1 0 960 0 -1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_18
timestamp 1680000637
transform -1 0 1344 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_19
timestamp 1680000637
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_20
timestamp 1680000637
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_21
timestamp 1680000637
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_22
timestamp 1680000637
transform -1 0 1344 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_23
timestamp 1680000637
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_24
timestamp 1680000637
transform -1 0 960 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_ppwm_25
timestamp 1680000637
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677672058
transform -1 0 16320 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677672058
transform 1 0 12864 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677672058
transform -1 0 48960 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677672058
transform 1 0 45984 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677672058
transform 1 0 8928 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677672058
transform -1 0 11520 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677672058
transform -1 0 12192 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677672058
transform 1 0 10944 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677672058
transform -1 0 14784 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677672058
transform -1 0 13056 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677672058
transform -1 0 7776 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677672058
transform -1 0 6720 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677672058
transform -1 0 8928 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677672058
transform -1 0 7584 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677672058
transform -1 0 19584 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677672058
transform 1 0 17856 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677672058
transform 1 0 10368 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677672058
transform -1 0 13248 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677672058
transform -1 0 17952 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677672058
transform 1 0 17760 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677672058
transform -1 0 17088 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677672058
transform -1 0 34464 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677672058
transform -1 0 32544 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677672058
transform -1 0 5664 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677672058
transform 1 0 6816 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677672058
transform -1 0 10752 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677672058
transform 1 0 11712 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677672058
transform -1 0 27648 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677672058
transform -1 0 28224 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677672058
transform -1 0 10656 0 -1 38556
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677672058
transform 1 0 10656 0 -1 38556
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677672058
transform 1 0 17760 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677672058
transform 1 0 17184 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677672058
transform -1 0 18048 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677672058
transform -1 0 18816 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677672058
transform -1 0 10848 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677672058
transform 1 0 10848 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677672058
transform -1 0 10368 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677672058
transform -1 0 12096 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677672058
transform -1 0 12192 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677672058
transform -1 0 11232 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677672058
transform -1 0 25728 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677672058
transform -1 0 27168 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677672058
transform -1 0 47808 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677672058
transform -1 0 48672 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1677672058
transform 1 0 5376 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1677672058
transform -1 0 37728 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1677672058
transform 1 0 36576 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1677672058
transform -1 0 15072 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1677672058
transform -1 0 16608 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1677672058
transform -1 0 14400 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1677672058
transform -1 0 14880 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1677672058
transform 1 0 17472 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1677672058
transform -1 0 19776 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1677672058
transform -1 0 5472 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1677672058
transform -1 0 7680 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1677672058
transform 1 0 14016 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1677672058
transform -1 0 15744 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1677672058
transform 1 0 13824 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1677672058
transform -1 0 9984 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1677672058
transform -1 0 10080 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1677672058
transform 1 0 9120 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1677672058
transform -1 0 11424 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1677672058
transform 1 0 43008 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1677672058
transform 1 0 43104 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1677672058
transform 1 0 6720 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1677672058
transform -1 0 17952 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1677672058
transform 1 0 16224 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1677672058
transform -1 0 21312 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1677672058
transform 1 0 18528 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1677672058
transform -1 0 29760 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1677672058
transform -1 0 30048 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1677672058
transform -1 0 29184 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1677672058
transform -1 0 30336 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1677672058
transform -1 0 24288 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1677672058
transform -1 0 22656 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold77
timestamp 1677672058
transform -1 0 44160 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold78
timestamp 1677672058
transform -1 0 41856 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold79
timestamp 1677672058
transform -1 0 43872 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold80
timestamp 1677672058
transform -1 0 36000 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold81
timestamp 1677672058
transform -1 0 36480 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold82
timestamp 1677672058
transform -1 0 48000 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold83
timestamp 1677672058
transform 1 0 48192 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold84
timestamp 1677672058
transform -1 0 45024 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold85
timestamp 1677672058
transform 1 0 43008 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold86
timestamp 1677672058
transform -1 0 41184 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold87
timestamp 1677672058
transform 1 0 40608 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold88
timestamp 1677672058
transform -1 0 24768 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold89
timestamp 1677672058
transform -1 0 24192 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold90
timestamp 1677672058
transform -1 0 35616 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold91
timestamp 1677672058
transform -1 0 36480 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold92
timestamp 1677672058
transform 1 0 8928 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold93
timestamp 1677672058
transform -1 0 10848 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold94
timestamp 1677672058
transform -1 0 7872 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold95
timestamp 1677672058
transform -1 0 43392 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold96
timestamp 1677672058
transform 1 0 42816 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold97
timestamp 1677672058
transform 1 0 4032 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold98
timestamp 1677672058
transform -1 0 3648 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold99
timestamp 1677672058
transform 1 0 4704 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold100
timestamp 1677672058
transform -1 0 43968 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold101
timestamp 1677672058
transform -1 0 13248 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold102
timestamp 1677672058
transform -1 0 11712 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold103
timestamp 1677672058
transform 1 0 11712 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold104
timestamp 1677672058
transform -1 0 12672 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold105
timestamp 1677672058
transform 1 0 13920 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold106
timestamp 1677672058
transform -1 0 16512 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold107
timestamp 1677672058
transform -1 0 20352 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold108
timestamp 1677672058
transform 1 0 3840 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold109
timestamp 1677672058
transform 1 0 11808 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold110
timestamp 1677672058
transform 1 0 10752 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold111
timestamp 1677672058
transform -1 0 31680 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold112
timestamp 1677672058
transform 1 0 37920 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold113
timestamp 1677672058
transform 1 0 38208 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold114
timestamp 1677672058
transform 1 0 13344 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold115
timestamp 1677672058
transform -1 0 15264 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold116
timestamp 1677672058
transform -1 0 26688 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold117
timestamp 1677672058
transform 1 0 15744 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold118
timestamp 1677672058
transform 1 0 18240 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold119
timestamp 1677672058
transform -1 0 26592 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold120
timestamp 1677672058
transform -1 0 4416 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold121
timestamp 1677672058
transform -1 0 6240 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold122
timestamp 1677672058
transform -1 0 31392 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold123
timestamp 1677672058
transform -1 0 32736 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold124
timestamp 1677672058
transform -1 0 16128 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold125
timestamp 1677672058
transform 1 0 13920 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold126
timestamp 1677672058
transform -1 0 34752 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold127
timestamp 1677672058
transform 1 0 33504 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold128
timestamp 1677672058
transform -1 0 4896 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold129
timestamp 1677672058
transform -1 0 4704 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold130
timestamp 1677672058
transform -1 0 17376 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold131
timestamp 1677672058
transform -1 0 36192 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold132
timestamp 1677672058
transform -1 0 33888 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold133
timestamp 1677672058
transform -1 0 40512 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold134
timestamp 1677672058
transform -1 0 40416 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold135
timestamp 1677672058
transform -1 0 10752 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold136
timestamp 1677672058
transform 1 0 7776 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold137
timestamp 1677672058
transform 1 0 25632 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold138
timestamp 1677672058
transform 1 0 39456 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold139
timestamp 1677672058
transform -1 0 34080 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold140
timestamp 1677672058
transform -1 0 32256 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold141
timestamp 1677672058
transform -1 0 21696 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold142
timestamp 1677672058
transform 1 0 20352 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold143
timestamp 1677672058
transform -1 0 50688 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold144
timestamp 1677672058
transform 1 0 48480 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold145
timestamp 1677672058
transform -1 0 11712 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold146
timestamp 1677672058
transform -1 0 7296 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold147
timestamp 1677672058
transform -1 0 7296 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold148
timestamp 1677672058
transform -1 0 3840 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold149
timestamp 1677672058
transform -1 0 42912 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold150
timestamp 1677672058
transform -1 0 17952 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold151
timestamp 1677672058
transform -1 0 11232 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold152
timestamp 1677672058
transform -1 0 21792 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold153
timestamp 1677672058
transform 1 0 18912 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold154
timestamp 1677672058
transform -1 0 40704 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold155
timestamp 1677672058
transform 1 0 37344 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold156
timestamp 1677672058
transform -1 0 47328 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold157
timestamp 1677672058
transform 1 0 46464 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold158
timestamp 1677672058
transform -1 0 11040 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold159
timestamp 1677672058
transform -1 0 5184 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold160
timestamp 1677672058
transform 1 0 4896 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold161
timestamp 1677672058
transform 1 0 40896 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold162
timestamp 1677672058
transform -1 0 42432 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold163
timestamp 1677672058
transform -1 0 21888 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold164
timestamp 1677672058
transform -1 0 44928 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold165
timestamp 1677672058
transform 1 0 12000 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold166
timestamp 1677672058
transform 1 0 13152 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold167
timestamp 1677672058
transform -1 0 7392 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold168
timestamp 1677672058
transform -1 0 35136 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold169
timestamp 1677672058
transform -1 0 8160 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold170
timestamp 1677672058
transform -1 0 10464 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold171
timestamp 1677672058
transform 1 0 8640 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold172
timestamp 1677672058
transform -1 0 4704 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold173
timestamp 1677672058
transform -1 0 38304 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold174
timestamp 1677672058
transform 1 0 32064 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold175
timestamp 1677672058
transform -1 0 49248 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold176
timestamp 1677672058
transform 1 0 49056 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold177
timestamp 1677672058
transform -1 0 28224 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold178
timestamp 1677672058
transform -1 0 6720 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold179
timestamp 1677672058
transform -1 0 4992 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold180
timestamp 1677672058
transform 1 0 3552 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold181
timestamp 1677672058
transform 1 0 5472 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold182
timestamp 1677672058
transform -1 0 5088 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold183
timestamp 1677672058
transform -1 0 50880 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold184
timestamp 1677672058
transform 1 0 47616 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold185
timestamp 1677672058
transform -1 0 32256 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold186
timestamp 1677672058
transform -1 0 36960 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold187
timestamp 1677672058
transform -1 0 35136 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold188
timestamp 1677672058
transform -1 0 36864 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold189
timestamp 1677672058
transform -1 0 30624 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold190
timestamp 1677672058
transform 1 0 44736 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold191
timestamp 1677672058
transform 1 0 29952 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold192
timestamp 1677672058
transform -1 0 42048 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold193
timestamp 1677672058
transform -1 0 49152 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold194
timestamp 1677672058
transform 1 0 43968 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold195
timestamp 1677672058
transform -1 0 51264 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold196
timestamp 1677672058
transform -1 0 47712 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold197
timestamp 1677672058
transform -1 0 9696 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold198
timestamp 1677672058
transform 1 0 6528 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold199
timestamp 1677672058
transform -1 0 8448 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold200
timestamp 1677672058
transform -1 0 17760 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold201
timestamp 1677672058
transform -1 0 9792 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold202
timestamp 1677672058
transform -1 0 39360 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold203
timestamp 1677672058
transform -1 0 8640 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold204
timestamp 1677672058
transform -1 0 7104 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold205
timestamp 1677672058
transform 1 0 4608 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold206
timestamp 1677672058
transform -1 0 5856 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold207
timestamp 1677672058
transform -1 0 48768 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold208
timestamp 1677672058
transform -1 0 47712 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold209
timestamp 1677672058
transform -1 0 50592 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold210
timestamp 1677672058
transform 1 0 47904 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold211
timestamp 1677672058
transform -1 0 7872 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold212
timestamp 1677672058
transform -1 0 4512 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold213
timestamp 1677672058
transform -1 0 47232 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold214
timestamp 1677672058
transform -1 0 19488 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold215
timestamp 1677672058
transform -1 0 12576 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold216
timestamp 1677672058
transform -1 0 6432 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold217
timestamp 1677672058
transform -1 0 37440 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold218
timestamp 1677672058
transform 1 0 38304 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold219
timestamp 1677672058
transform 1 0 5568 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold220
timestamp 1677672058
transform -1 0 6528 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold221
timestamp 1677672058
transform -1 0 4992 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold222
timestamp 1677672058
transform 1 0 42144 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold223
timestamp 1677672058
transform 1 0 43680 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold224
timestamp 1677672058
transform -1 0 13920 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold225
timestamp 1677672058
transform -1 0 9216 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold226
timestamp 1677672058
transform -1 0 9120 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold227
timestamp 1677672058
transform 1 0 9792 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold228
timestamp 1677672058
transform -1 0 32832 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold229
timestamp 1677672058
transform -1 0 39168 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold230
timestamp 1677672058
transform -1 0 37536 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold231
timestamp 1677672058
transform -1 0 45888 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold232
timestamp 1677672058
transform 1 0 43488 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold233
timestamp 1677672058
transform -1 0 3648 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold234
timestamp 1677672058
transform -1 0 3648 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold235
timestamp 1677672058
transform -1 0 2592 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold236
timestamp 1677672058
transform -1 0 46368 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold237
timestamp 1677672058
transform 1 0 44544 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold238
timestamp 1677672058
transform -1 0 3264 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold239
timestamp 1677672058
transform -1 0 4992 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold240
timestamp 1677672058
transform -1 0 40992 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold241
timestamp 1677672058
transform -1 0 38880 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold242
timestamp 1677672058
transform 1 0 38880 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold243
timestamp 1677672058
transform 1 0 3840 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold244
timestamp 1677672058
transform -1 0 6048 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold245
timestamp 1677672058
transform -1 0 4128 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold246
timestamp 1677672058
transform 1 0 16032 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold247
timestamp 1677672058
transform -1 0 19008 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold248
timestamp 1677672058
transform -1 0 18432 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold249
timestamp 1677672058
transform 1 0 4608 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold250
timestamp 1677672058
transform -1 0 8256 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold251
timestamp 1677672058
transform -1 0 7968 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold252
timestamp 1677672058
transform -1 0 40608 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold253
timestamp 1677672058
transform 1 0 37440 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold254
timestamp 1677672058
transform -1 0 41376 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold255
timestamp 1677672058
transform 1 0 38400 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold256
timestamp 1677672058
transform 1 0 4512 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold257
timestamp 1677672058
transform -1 0 10752 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold258
timestamp 1677672058
transform 1 0 8448 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold259
timestamp 1677672058
transform 1 0 42720 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold260
timestamp 1677672058
transform -1 0 42720 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold261
timestamp 1677672058
transform 1 0 42048 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold262
timestamp 1677672058
transform -1 0 45312 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold263
timestamp 1677672058
transform 1 0 43584 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold264
timestamp 1677672058
transform 1 0 45120 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold265
timestamp 1677672058
transform -1 0 40800 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold266
timestamp 1677672058
transform -1 0 39936 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold267
timestamp 1677672058
transform 1 0 37920 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold268
timestamp 1677672058
transform -1 0 5280 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold269
timestamp 1677672058
transform 1 0 4992 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold270
timestamp 1677672058
transform 1 0 4704 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold271
timestamp 1677672058
transform 1 0 47328 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold272
timestamp 1677672058
transform -1 0 45888 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold273
timestamp 1677672058
transform 1 0 43104 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold274
timestamp 1677672058
transform 1 0 13920 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold275
timestamp 1677672058
transform -1 0 18144 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold276
timestamp 1677672058
transform -1 0 7584 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold277
timestamp 1677672058
transform 1 0 36192 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold278
timestamp 1677672058
transform 1 0 37536 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold279
timestamp 1677672058
transform -1 0 6816 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold280
timestamp 1677672058
transform 1 0 18528 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold281
timestamp 1677672058
transform -1 0 21984 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold282
timestamp 1677672058
transform -1 0 18528 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold283
timestamp 1677672058
transform -1 0 4992 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold284
timestamp 1677672058
transform -1 0 4512 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold285
timestamp 1677672058
transform -1 0 47712 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold286
timestamp 1677672058
transform -1 0 39648 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold287
timestamp 1677672058
transform 1 0 43488 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold288
timestamp 1677672058
transform -1 0 41664 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold289
timestamp 1677672058
transform -1 0 18624 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold290
timestamp 1677672058
transform -1 0 16992 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold291
timestamp 1677672058
transform -1 0 44256 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold292
timestamp 1677672058
transform -1 0 34368 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold293
timestamp 1677672058
transform 1 0 34464 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold294
timestamp 1677672058
transform -1 0 27552 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold295
timestamp 1677672058
transform 1 0 17952 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold296
timestamp 1677672058
transform -1 0 21408 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold297
timestamp 1677672058
transform -1 0 45024 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold298
timestamp 1677672058
transform 1 0 44352 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold299
timestamp 1677672058
transform -1 0 33696 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold300
timestamp 1677672058
transform -1 0 39648 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold301
timestamp 1677672058
transform 1 0 24384 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold302
timestamp 1677672058
transform -1 0 22560 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold303
timestamp 1677672058
transform -1 0 32352 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold304
timestamp 1677672058
transform -1 0 17568 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold305
timestamp 1677672058
transform -1 0 26688 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold306
timestamp 1677672058
transform -1 0 23712 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold307
timestamp 1677672058
transform -1 0 17376 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold308
timestamp 1677672058
transform 1 0 34272 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold309
timestamp 1677672058
transform -1 0 26496 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold310
timestamp 1677672058
transform -1 0 37632 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold311
timestamp 1677672058
transform 1 0 33600 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold312
timestamp 1677672058
transform -1 0 41472 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold313
timestamp 1677672058
transform -1 0 36768 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold314
timestamp 1677672058
transform 1 0 35904 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold315
timestamp 1677672058
transform -1 0 23328 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold316
timestamp 1677672058
transform -1 0 21120 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold317
timestamp 1677672058
transform -1 0 20256 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold318
timestamp 1677672058
transform -1 0 20448 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold319
timestamp 1677672058
transform 1 0 41760 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold320
timestamp 1677672058
transform 1 0 38304 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold321
timestamp 1677672058
transform -1 0 30528 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold322
timestamp 1677672058
transform -1 0 32256 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold323
timestamp 1677672058
transform 1 0 3648 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold324
timestamp 1677672058
transform -1 0 32736 0 -1 17388
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_ex__0564_
timestamp 1676382947
transform 1 0 18624 0 1 8316
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_ex__0565_
timestamp 1676382947
transform 1 0 15744 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_4  u_ppwm_u_ex__0566_
timestamp 1676383058
transform 1 0 27456 0 -1 8316
box -48 -56 624 834
use sg13g2_inv_2  u_ppwm_u_ex__0567_
timestamp 1676382947
transform 1 0 28992 0 1 6804
box -48 -56 432 834
use sg13g2_inv_4  u_ppwm_u_ex__0568_
timestamp 1676383058
transform 1 0 34272 0 -1 6804
box -48 -56 624 834
use sg13g2_inv_2  u_ppwm_u_ex__0569_
timestamp 1676382947
transform -1 0 35232 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__0570_
timestamp 1676382929
transform 1 0 35136 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0571_
timestamp 1676382929
transform -1 0 25152 0 1 8316
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__0572_
timestamp 1676382947
transform 1 0 20736 0 1 6804
box -48 -56 432 834
use sg13g2_inv_2  u_ppwm_u_ex__0573_
timestamp 1676382947
transform 1 0 20256 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_ex__0574_
timestamp 1676382929
transform -1 0 31776 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0575_
timestamp 1676382929
transform 1 0 34080 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0576_
timestamp 1676382929
transform -1 0 36384 0 1 11340
box -48 -56 336 834
use sg13g2_inv_4  u_ppwm_u_ex__0577_
timestamp 1676383058
transform -1 0 37536 0 1 11340
box -48 -56 624 834
use sg13g2_inv_1  u_ppwm_u_ex__0578_
timestamp 1676382929
transform 1 0 15648 0 1 14364
box -48 -56 336 834
use sg13g2_inv_4  u_ppwm_u_ex__0579_
timestamp 1676383058
transform -1 0 32640 0 -1 18900
box -48 -56 624 834
use sg13g2_inv_1  u_ppwm_u_ex__0580_
timestamp 1676382929
transform -1 0 22080 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_ex__0581_
timestamp 1676382947
transform -1 0 29568 0 1 9828
box -48 -56 432 834
use sg13g2_inv_4  u_ppwm_u_ex__0582_
timestamp 1676383058
transform -1 0 27456 0 -1 11340
box -48 -56 624 834
use sg13g2_inv_1  u_ppwm_u_ex__0583_
timestamp 1676382929
transform 1 0 16128 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0584_
timestamp 1676382929
transform -1 0 19872 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0585_
timestamp 1676382929
transform -1 0 25440 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0586_
timestamp 1676382929
transform 1 0 34368 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0587_
timestamp 1676382929
transform -1 0 37536 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0588_
timestamp 1676382929
transform -1 0 29088 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0589_
timestamp 1676382929
transform -1 0 33696 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0590_
timestamp 1676382929
transform -1 0 33120 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_ex__0591_
timestamp 1676382929
transform -1 0 35040 0 -1 12852
box -48 -56 336 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0592_
timestamp 1685175443
transform 1 0 16704 0 1 15876
box -48 -56 538 834
use sg13g2_and2_1  u_ppwm_u_ex__0593_
timestamp 1676901763
transform -1 0 24576 0 1 21924
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__0594_
timestamp 1683988354
transform -1 0 22176 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2_2  u_ppwm_u_ex__0595_
timestamp 1683979924
transform -1 0 22848 0 -1 18900
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_ex__0596_
timestamp 1676639442
transform -1 0 21024 0 1 17388
box -48 -56 528 834
use sg13g2_nor2b_2  u_ppwm_u_ex__0597_
timestamp 1685188981
transform 1 0 19104 0 1 9828
box -54 -56 720 834
use sg13g2_nor2_1  u_ppwm_u_ex__0598_
timestamp 1676627187
transform 1 0 15936 0 1 15876
box -48 -56 432 834
use sg13g2_nand3_1  u_ppwm_u_ex__0599_
timestamp 1683988354
transform 1 0 18624 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__0600_
timestamp 1676557249
transform 1 0 19488 0 -1 18900
box -48 -56 432 834
use sg13g2_nand3_1  u_ppwm_u_ex__0601_
timestamp 1683988354
transform -1 0 19488 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0602_
timestamp 1683973020
transform -1 0 17568 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0603_
timestamp 1683973020
transform -1 0 17664 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0604_
timestamp 1685175443
transform -1 0 17760 0 1 17388
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__0605_
timestamp 1676557249
transform 1 0 15840 0 -1 17388
box -48 -56 432 834
use sg13g2_nand4_1  u_ppwm_u_ex__0606_
timestamp 1685201930
transform 1 0 17952 0 -1 17388
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0607_
timestamp 1683973020
transform -1 0 19584 0 1 17388
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0608_
timestamp 1676567195
transform 1 0 20544 0 -1 18900
box -48 -56 528 834
use sg13g2_and3_1  u_ppwm_u_ex__0609_
timestamp 1676971669
transform -1 0 21696 0 -1 18900
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__0610_
timestamp 1683988354
transform -1 0 22848 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0611_
timestamp 1685175443
transform 1 0 25152 0 1 18900
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__0612_
timestamp 1677577977
transform 1 0 25632 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0613_
timestamp 1676627187
transform -1 0 26688 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0614_
timestamp 1685175443
transform 1 0 22944 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0615_
timestamp 1685175443
transform 1 0 25248 0 -1 21924
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__0616_
timestamp 1677577977
transform -1 0 26112 0 -1 20412
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0617_
timestamp 1683973020
transform 1 0 25632 0 1 18900
box -48 -56 528 834
use sg13g2_and3_1  u_ppwm_u_ex__0618_
timestamp 1676971669
transform -1 0 25344 0 -1 20412
box -48 -56 720 834
use sg13g2_or3_1  u_ppwm_u_ex__0619_
timestamp 1677141922
transform 1 0 24960 0 1 20412
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0620_
timestamp 1685175443
transform 1 0 24768 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0621_
timestamp 1683973020
transform 1 0 25728 0 -1 21924
box -48 -56 528 834
use sg13g2_or2_1  u_ppwm_u_ex__0622_
timestamp 1684236171
transform 1 0 23424 0 1 20412
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0623_
timestamp 1676627187
transform -1 0 24096 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0624_
timestamp 1685175443
transform -1 0 24384 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0625_
timestamp 1683973020
transform -1 0 24672 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__0626_
timestamp 1676557249
transform -1 0 24192 0 -1 20412
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0627_
timestamp 1677516600
transform 1 0 22272 0 -1 20412
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0628_
timestamp 1677516600
transform 1 0 23040 0 -1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0629_
timestamp 1685175443
transform 1 0 23616 0 1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0630_
timestamp 1685175443
transform 1 0 22464 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0631_
timestamp 1676627187
transform 1 0 22464 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0632_
timestamp 1685175443
transform -1 0 23616 0 1 18900
box -48 -56 538 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0633_
timestamp 1677516600
transform 1 0 20160 0 1 20412
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0634_
timestamp 1677516600
transform -1 0 21696 0 -1 20412
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0635_
timestamp 1683973020
transform 1 0 21312 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__0636_
timestamp 1676557249
transform -1 0 21120 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0637_
timestamp 1685175443
transform 1 0 21792 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0638_
timestamp 1683973020
transform -1 0 19584 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0639_
timestamp 1685175443
transform -1 0 21600 0 -1 21924
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0640_
timestamp 1676627187
transform 1 0 19776 0 1 20412
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0641_
timestamp 1676557249
transform 1 0 22656 0 1 8316
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0642_
timestamp 1685173987
transform -1 0 31776 0 -1 9828
box -48 -56 624 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0643_
timestamp 1676567195
transform 1 0 33504 0 1 12852
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0644_
timestamp 1685181386
transform -1 0 34464 0 1 12852
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0645_
timestamp 1685181386
transform 1 0 33792 0 -1 14364
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0646_
timestamp 1685197497
transform 1 0 33984 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0647_
timestamp 1676567195
transform 1 0 34080 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0648_
timestamp 1685175443
transform -1 0 35040 0 1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0649_
timestamp 1685173987
transform -1 0 32448 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0650_
timestamp 1685175443
transform -1 0 34080 0 1 11340
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0651_
timestamp 1676627187
transform -1 0 31008 0 -1 9828
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0652_
timestamp 1685197497
transform -1 0 30720 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__0653_
timestamp 1676557249
transform 1 0 29088 0 1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0654_
timestamp 1685175443
transform -1 0 29952 0 1 8316
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0655_
timestamp 1676567195
transform 1 0 23136 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0656_
timestamp 1685175443
transform -1 0 24480 0 1 8316
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__0657_
timestamp 1677577977
transform 1 0 23136 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0658_
timestamp 1676627187
transform 1 0 23904 0 -1 9828
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0659_
timestamp 1676567195
transform -1 0 24000 0 1 8316
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0660_
timestamp 1676627187
transform 1 0 24480 0 1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0661_
timestamp 1685175443
transform -1 0 30624 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0662_
timestamp 1683973020
transform 1 0 23040 0 1 8316
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_ex__0663_
timestamp 1676985977
transform -1 0 22944 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0664_
timestamp 1685181386
transform 1 0 27072 0 1 6804
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0665_
timestamp 1685181386
transform -1 0 39360 0 -1 12852
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0666_
timestamp 1676567195
transform 1 0 37152 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0667_
timestamp 1676567195
transform 1 0 36480 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0668_
timestamp 1685175443
transform 1 0 36096 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0669_
timestamp 1676567195
transform -1 0 38880 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0670_
timestamp 1683973020
transform 1 0 38112 0 -1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0671_
timestamp 1685173987
transform 1 0 36576 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0672_
timestamp 1685175443
transform -1 0 37440 0 1 9828
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0673_
timestamp 1676639442
transform 1 0 36480 0 1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0674_
timestamp 1676567195
transform -1 0 35616 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0675_
timestamp 1685175443
transform 1 0 34656 0 1 5292
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0676_
timestamp 1676567195
transform 1 0 35904 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0677_
timestamp 1685175443
transform 1 0 35616 0 -1 8316
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0678_
timestamp 1676639442
transform -1 0 37344 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0679_
timestamp 1685181386
transform 1 0 33792 0 -1 6804
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0680_
timestamp 1685197497
transform -1 0 36864 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__0681_
timestamp 1676557249
transform -1 0 27936 0 1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0682_
timestamp 1685175443
transform -1 0 27456 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__0683_
timestamp 1676557249
transform -1 0 25632 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0684_
timestamp 1685175443
transform 1 0 24384 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0685_
timestamp 1676627187
transform -1 0 26688 0 1 6804
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0686_
timestamp 1676567195
transform 1 0 24864 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0687_
timestamp 1685175443
transform -1 0 26592 0 1 8316
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0688_
timestamp 1676639442
transform 1 0 25344 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0689_
timestamp 1676627187
transform 1 0 23808 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__0690_
timestamp 1676901763
transform 1 0 26016 0 1 14364
box -48 -56 528 834
use sg13g2_inv_1  u_ppwm_u_ex__0691_
timestamp 1676382929
transform 1 0 25632 0 1 8316
box -48 -56 336 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0692_
timestamp 1685197497
transform -1 0 26592 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__0693_
timestamp 1676557249
transform 1 0 35232 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0694_
timestamp 1685181386
transform 1 0 35328 0 -1 14364
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0695_
timestamp 1676567195
transform 1 0 34848 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0696_
timestamp 1676567195
transform 1 0 34848 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0697_
timestamp 1685175443
transform 1 0 35424 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0698_
timestamp 1676567195
transform 1 0 35808 0 -1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0699_
timestamp 1683973020
transform 1 0 36288 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0700_
timestamp 1685181386
transform 1 0 34272 0 1 9828
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0701_
timestamp 1685181386
transform 1 0 33792 0 1 9828
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0702_
timestamp 1685197497
transform 1 0 35232 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0703_
timestamp 1685175443
transform -1 0 35808 0 -1 9828
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0704_
timestamp 1685173987
transform 1 0 34848 0 1 6804
box -48 -56 624 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0705_
timestamp 1676567195
transform 1 0 29760 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0706_
timestamp 1685175443
transform -1 0 31008 0 1 6804
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0707_
timestamp 1685173987
transform 1 0 29376 0 1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0708_
timestamp 1685175443
transform -1 0 30240 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__0709_
timestamp 1676557249
transform -1 0 22656 0 -1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0710_
timestamp 1685175443
transform 1 0 23616 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0711_
timestamp 1676627187
transform 1 0 24768 0 1 6804
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0712_
timestamp 1676567195
transform 1 0 22464 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0713_
timestamp 1685175443
transform -1 0 24768 0 1 6804
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0714_
timestamp 1676639442
transform 1 0 22656 0 -1 8316
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__0715_
timestamp 1676901763
transform 1 0 22560 0 1 12852
box -48 -56 528 834
use sg13g2_inv_1  u_ppwm_u_ex__0716_
timestamp 1676382929
transform -1 0 22464 0 1 6804
box -48 -56 336 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0717_
timestamp 1685197497
transform 1 0 23520 0 1 6804
box -48 -56 816 834
use sg13g2_and4_1  u_ppwm_u_ex__0718_
timestamp 1676985977
transform -1 0 21792 0 1 17388
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0719_
timestamp 1676627187
transform -1 0 34752 0 1 6804
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0720_
timestamp 1676567195
transform 1 0 34848 0 1 12852
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0721_
timestamp 1685181386
transform 1 0 36096 0 1 12852
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0722_
timestamp 1685181386
transform -1 0 35712 0 -1 12852
box -54 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0723_
timestamp 1685197497
transform 1 0 35328 0 1 12852
box -48 -56 816 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0724_
timestamp 1676567195
transform -1 0 36480 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0725_
timestamp 1685175443
transform 1 0 34752 0 1 9828
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0726_
timestamp 1685181386
transform 1 0 34080 0 -1 9828
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0727_
timestamp 1685181386
transform 1 0 33504 0 1 8316
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0728_
timestamp 1685181386
transform -1 0 36288 0 -1 9828
box -54 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__0729_
timestamp 1677577977
transform 1 0 34656 0 1 8316
box -48 -56 816 834
use sg13g2_nor4_1  u_ppwm_u_ex__0730_
timestamp 1676643125
transform 1 0 34752 0 -1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0731_
timestamp 1685175443
transform -1 0 35904 0 1 8316
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0732_
timestamp 1676639442
transform 1 0 33984 0 -1 8316
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0733_
timestamp 1685197497
transform -1 0 35232 0 -1 8316
box -48 -56 816 834
use sg13g2_a21o_1  u_ppwm_u_ex__0734_
timestamp 1677175127
transform 1 0 33984 0 1 8316
box -48 -56 720 834
use sg13g2_nand2_1  u_ppwm_u_ex__0735_
timestamp 1676557249
transform -1 0 22176 0 1 8316
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0736_
timestamp 1685173987
transform -1 0 20736 0 1 8316
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0737_
timestamp 1676627187
transform -1 0 20640 0 -1 9828
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0738_
timestamp 1685197497
transform 1 0 20640 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__0739_
timestamp 1676557249
transform -1 0 21792 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0740_
timestamp 1683973020
transform -1 0 21120 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__0741_
timestamp 1676557249
transform 1 0 23424 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_2  u_ppwm_u_ex__0742_
timestamp 1683979924
transform 1 0 31296 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0743_
timestamp 1685175443
transform -1 0 20160 0 1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0744_
timestamp 1685175443
transform 1 0 21312 0 1 8316
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0745_
timestamp 1685181386
transform -1 0 37920 0 -1 12852
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0746_
timestamp 1676567195
transform 1 0 36768 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0747_
timestamp 1676567195
transform 1 0 31392 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0748_
timestamp 1685175443
transform 1 0 32352 0 1 11340
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0749_
timestamp 1676567195
transform -1 0 38400 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0750_
timestamp 1683973020
transform 1 0 36960 0 -1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0751_
timestamp 1685173987
transform 1 0 32448 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0752_
timestamp 1685175443
transform -1 0 33504 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0753_
timestamp 1676627187
transform -1 0 33024 0 1 9828
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0754_
timestamp 1685173987
transform 1 0 31296 0 1 9828
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0755_
timestamp 1676627187
transform -1 0 33408 0 1 9828
box -48 -56 432 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0756_
timestamp 1685197497
transform -1 0 32640 0 1 9828
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0757_
timestamp 1676627187
transform 1 0 28320 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_ex__0758_
timestamp 1676627187
transform 1 0 29568 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__0759_
timestamp 1677577977
transform 1 0 27360 0 -1 9828
box -48 -56 816 834
use sg13g2_nor4_1  u_ppwm_u_ex__0760_
timestamp 1676643125
transform -1 0 28704 0 -1 9828
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_ex__0761_
timestamp 1676639442
transform 1 0 27840 0 1 8316
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0762_
timestamp 1685197497
transform -1 0 27840 0 1 8316
box -48 -56 816 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0763_
timestamp 1685181386
transform -1 0 27360 0 -1 9828
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0764_
timestamp 1676567195
transform 1 0 24288 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0765_
timestamp 1685175443
transform 1 0 24768 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0766_
timestamp 1685181386
transform 1 0 24768 0 1 9828
box -54 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__0767_
timestamp 1676643125
transform 1 0 24672 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0768_
timestamp 1685175443
transform -1 0 25728 0 1 9828
box -48 -56 538 834
use sg13g2_nor4_1  u_ppwm_u_ex__0769_
timestamp 1676643125
transform -1 0 22176 0 -1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0770_
timestamp 1685175443
transform 1 0 20160 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0771_
timestamp 1683973020
transform 1 0 20640 0 1 9828
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0772_
timestamp 1685201930
transform -1 0 19104 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0773_
timestamp 1685175443
transform -1 0 16032 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0774_
timestamp 1683973020
transform -1 0 15648 0 1 14364
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__0775_
timestamp 1676901763
transform 1 0 24096 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_2  u_ppwm_u_ex__0776_
timestamp 1685180049
transform 1 0 24096 0 -1 17388
box -48 -56 624 834
use sg13g2_nor3_2  u_ppwm_u_ex__0777_
timestamp 1685180723
transform 1 0 30048 0 1 9828
box -48 -56 912 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0778_
timestamp 1685173987
transform 1 0 32064 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2b_2  u_ppwm_u_ex__0779_
timestamp 1685188981
transform -1 0 22464 0 1 17388
box -54 -56 720 834
use sg13g2_and2_1  u_ppwm_u_ex__0780_
timestamp 1676901763
transform 1 0 22464 0 -1 17388
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__0781_
timestamp 1676557249
transform 1 0 22080 0 -1 17388
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0782_
timestamp 1676557249
transform 1 0 26688 0 1 14364
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__0783_
timestamp 1677577977
transform -1 0 27936 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_2  u_ppwm_u_ex__0784_
timestamp 1683979924
transform -1 0 26784 0 -1 17388
box -48 -56 624 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0785_
timestamp 1685173987
transform -1 0 27552 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0786_
timestamp 1685175443
transform 1 0 33600 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0787_
timestamp 1683973020
transform -1 0 33504 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_2  u_ppwm_u_ex__0788_
timestamp 1685180049
transform -1 0 21984 0 1 15876
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0789_
timestamp 1676627187
transform -1 0 22560 0 1 12852
box -48 -56 432 834
use sg13g2_nor2b_2  u_ppwm_u_ex__0790_
timestamp 1685188981
transform -1 0 22560 0 -1 14364
box -54 -56 720 834
use sg13g2_or2_1  u_ppwm_u_ex__0791_
timestamp 1684236171
transform -1 0 29952 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0792_
timestamp 1685175443
transform -1 0 29472 0 1 12852
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_ex__0793_
timestamp 1677247768
transform -1 0 26688 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_ex__0794_
timestamp 1676557249
transform 1 0 23904 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0795_
timestamp 1685175443
transform -1 0 23904 0 1 14364
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0796_
timestamp 1676627187
transform -1 0 23616 0 1 12852
box -48 -56 432 834
use sg13g2_nor2b_2  u_ppwm_u_ex__0797_
timestamp 1685188981
transform -1 0 23232 0 -1 14364
box -54 -56 720 834
use sg13g2_mux2_1  u_ppwm_u_ex__0798_
timestamp 1677247768
transform -1 0 29760 0 -1 11340
box -48 -56 1008 834
use sg13g2_inv_1  u_ppwm_u_ex__0799_
timestamp 1676382929
transform -1 0 21888 0 -1 12852
box -48 -56 336 834
use sg13g2_mux2_1  u_ppwm_u_ex__0800_
timestamp 1677247768
transform -1 0 28032 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_ex__0801_
timestamp 1677247768
transform 1 0 18240 0 1 12852
box -48 -56 1008 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0802_
timestamp 1685173987
transform -1 0 21888 0 -1 14364
box -48 -56 624 834
use sg13g2_or3_1  u_ppwm_u_ex__0803_
timestamp 1677141922
transform 1 0 24288 0 1 14364
box -48 -56 720 834
use sg13g2_nor2_1  u_ppwm_u_ex__0804_
timestamp 1676627187
transform 1 0 24576 0 -1 18900
box -48 -56 432 834
use sg13g2_nor3_1  u_ppwm_u_ex__0805_
timestamp 1676639442
transform 1 0 24096 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0806_
timestamp 1685175443
transform 1 0 25536 0 -1 17388
box -48 -56 538 834
use sg13g2_nor2b_2  u_ppwm_u_ex__0807_
timestamp 1685188981
transform 1 0 25440 0 1 15876
box -54 -56 720 834
use sg13g2_and2_1  u_ppwm_u_ex__0808_
timestamp 1676901763
transform 1 0 33504 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0809_
timestamp 1685175443
transform 1 0 33984 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0810_
timestamp 1683973020
transform -1 0 34560 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0811_
timestamp 1677247768
transform -1 0 27168 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_ex__0812_
timestamp 1677247768
transform -1 0 30144 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_ex__0813_
timestamp 1677247768
transform -1 0 22848 0 -1 12852
box -48 -56 1008 834
use sg13g2_inv_1  u_ppwm_u_ex__0814_
timestamp 1676382929
transform -1 0 20544 0 1 12852
box -48 -56 336 834
use sg13g2_mux2_1  u_ppwm_u_ex__0815_
timestamp 1677247768
transform -1 0 26016 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_ex__0816_
timestamp 1676557249
transform -1 0 21696 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0817_
timestamp 1685175443
transform -1 0 20736 0 1 14364
box -48 -56 538 834
use sg13g2_and3_2  u_ppwm_u_ex__0818_
timestamp 1683976310
transform -1 0 21216 0 1 15876
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_ex__0819_
timestamp 1683988354
transform 1 0 20064 0 1 15876
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__0820_
timestamp 1683988354
transform -1 0 20544 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0821_
timestamp 1677247768
transform 1 0 19488 0 -1 14364
box -48 -56 1008 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0822_
timestamp 1685173987
transform 1 0 20736 0 1 14364
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__0823_
timestamp 1676557249
transform 1 0 20928 0 -1 17388
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0824_
timestamp 1676557249
transform 1 0 27840 0 1 15876
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0825_
timestamp 1676557249
transform 1 0 27456 0 1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0826_
timestamp 1677516600
transform 1 0 27840 0 1 14364
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0827_
timestamp 1683973020
transform -1 0 29088 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0828_
timestamp 1685175443
transform 1 0 29088 0 1 14364
box -48 -56 538 834
use sg13g2_nand3_1  u_ppwm_u_ex__0829_
timestamp 1683988354
transform 1 0 30336 0 1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0830_
timestamp 1685173987
transform -1 0 33792 0 -1 14364
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__0831_
timestamp 1676557249
transform 1 0 34560 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0832_
timestamp 1685175443
transform 1 0 31872 0 1 14364
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0833_
timestamp 1676639442
transform 1 0 32256 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0834_
timestamp 1685175443
transform -1 0 38496 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0835_
timestamp 1676627187
transform 1 0 37920 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__0836_
timestamp 1676901763
transform -1 0 17280 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_2  u_ppwm_u_ex__0837_
timestamp 1685180049
transform 1 0 17280 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0838_
timestamp 1676627187
transform 1 0 16512 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2b_2  u_ppwm_u_ex__0839_
timestamp 1685211885
transform 1 0 18048 0 1 14364
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0840_
timestamp 1676627187
transform 1 0 16416 0 1 14364
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0841_
timestamp 1685173987
transform 1 0 18816 0 1 14364
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__0842_
timestamp 1676557249
transform 1 0 18336 0 -1 15876
box -48 -56 432 834
use sg13g2_nor3_1  u_ppwm_u_ex__0843_
timestamp 1676639442
transform -1 0 20160 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0844_
timestamp 1677247768
transform -1 0 19104 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_ex__0845_
timestamp 1676557249
transform -1 0 16704 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0846_
timestamp 1685175443
transform -1 0 17664 0 -1 11340
box -48 -56 538 834
use sg13g2_inv_1  u_ppwm_u_ex__0847_
timestamp 1676382929
transform 1 0 18048 0 -1 14364
box -48 -56 336 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0848_
timestamp 1685197497
transform 1 0 20544 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0849_
timestamp 1685175443
transform -1 0 28608 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0850_
timestamp 1676627187
transform -1 0 29568 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__0851_
timestamp 1677577977
transform 1 0 27648 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0852_
timestamp 1677516600
transform 1 0 26208 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0853_
timestamp 1685175443
transform -1 0 28224 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  u_ppwm_u_ex__0854_
timestamp 1677175127
transform -1 0 28800 0 1 12852
box -48 -56 720 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0855_
timestamp 1685173987
transform 1 0 30336 0 -1 12852
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__0856_
timestamp 1676557249
transform 1 0 27072 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0857_
timestamp 1685175443
transform -1 0 30624 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0858_
timestamp 1683973020
transform 1 0 30528 0 1 12852
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0859_
timestamp 1685201930
transform -1 0 30528 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0860_
timestamp 1685175443
transform 1 0 37248 0 1 12852
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0861_
timestamp 1685181386
transform 1 0 37248 0 -1 14364
box -54 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0862_
timestamp 1677516600
transform 1 0 26880 0 -1 12852
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0863_
timestamp 1683973020
transform -1 0 28704 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0864_
timestamp 1683973020
transform -1 0 29184 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0865_
timestamp 1685175443
transform 1 0 27648 0 1 12852
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0866_
timestamp 1676639442
transform -1 0 20064 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0867_
timestamp 1676627187
transform 1 0 19200 0 -1 15876
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0868_
timestamp 1685175443
transform 1 0 20544 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0869_
timestamp 1676627187
transform -1 0 18624 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0870_
timestamp 1683973020
transform -1 0 18144 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0871_
timestamp 1677247768
transform 1 0 16896 0 -1 12852
box -48 -56 1008 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0872_
timestamp 1685173987
transform 1 0 21984 0 1 14364
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__0873_
timestamp 1677175127
transform -1 0 22368 0 -1 15876
box -48 -56 720 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0874_
timestamp 1685173987
transform 1 0 30912 0 -1 12852
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0875_
timestamp 1676627187
transform -1 0 31392 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0876_
timestamp 1683973020
transform -1 0 30048 0 1 14364
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0877_
timestamp 1685201930
transform -1 0 28896 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0878_
timestamp 1685175443
transform 1 0 28896 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0879_
timestamp 1676627187
transform -1 0 30624 0 1 18900
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0880_
timestamp 1676557249
transform 1 0 19968 0 -1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0881_
timestamp 1677516600
transform -1 0 21312 0 1 3780
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0882_
timestamp 1676627187
transform 1 0 28224 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0883_
timestamp 1683973020
transform 1 0 28800 0 1 11340
box -48 -56 528 834
use sg13g2_a21oi_2  u_ppwm_u_ex__0884_
timestamp 1685174172
transform 1 0 27456 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0885_
timestamp 1685175443
transform 1 0 23424 0 -1 3780
box -48 -56 538 834
use sg13g2_a21o_1  u_ppwm_u_ex__0886_
timestamp 1677175127
transform -1 0 24672 0 1 3780
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0887_
timestamp 1685175443
transform -1 0 19200 0 -1 15876
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0888_
timestamp 1676567195
transform -1 0 18816 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0889_
timestamp 1685175443
transform -1 0 19296 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0890_
timestamp 1676627187
transform 1 0 19200 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_ex__0891_
timestamp 1676627187
transform -1 0 17472 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0892_
timestamp 1683973020
transform 1 0 17184 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0893_
timestamp 1677247768
transform 1 0 16896 0 1 11340
box -48 -56 1008 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0894_
timestamp 1685197497
transform 1 0 20160 0 1 11340
box -48 -56 816 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0895_
timestamp 1685173987
transform -1 0 32544 0 -1 6804
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0896_
timestamp 1676627187
transform -1 0 33600 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0897_
timestamp 1683973020
transform -1 0 33024 0 -1 5292
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0898_
timestamp 1685201930
transform -1 0 24672 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0899_
timestamp 1685175443
transform -1 0 25536 0 1 3780
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0900_
timestamp 1685181386
transform 1 0 24672 0 -1 5292
box -54 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0901_
timestamp 1685175443
transform -1 0 20832 0 -1 5292
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__0902_
timestamp 1677577977
transform 1 0 19200 0 -1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0903_
timestamp 1683973020
transform -1 0 20544 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0904_
timestamp 1685175443
transform 1 0 20256 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0905_
timestamp 1683973020
transform -1 0 21024 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0906_
timestamp 1685175443
transform 1 0 21024 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0907_
timestamp 1683973020
transform 1 0 21120 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0908_
timestamp 1676627187
transform -1 0 15840 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0909_
timestamp 1683973020
transform 1 0 16704 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_ex__0910_
timestamp 1677247768
transform 1 0 15936 0 1 11340
box -48 -56 1008 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0911_
timestamp 1685197497
transform 1 0 21024 0 1 11340
box -48 -56 816 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0912_
timestamp 1685173987
transform 1 0 29952 0 1 6804
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0913_
timestamp 1676627187
transform -1 0 29760 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0914_
timestamp 1683973020
transform -1 0 26688 0 1 5292
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0915_
timestamp 1685201930
transform -1 0 21888 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0916_
timestamp 1685175443
transform 1 0 20736 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0917_
timestamp 1685181386
transform -1 0 22080 0 -1 2268
box -54 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0918_
timestamp 1676627187
transform 1 0 16224 0 -1 2268
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__0919_
timestamp 1676901763
transform 1 0 15744 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__0920_
timestamp 1676627187
transform -1 0 17568 0 1 756
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0921_
timestamp 1685175443
transform 1 0 16224 0 -1 3780
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__0922_
timestamp 1676567195
transform -1 0 20064 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0923_
timestamp 1685175443
transform -1 0 17856 0 -1 2268
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__0924_
timestamp 1677577977
transform 1 0 17472 0 1 2268
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__0925_
timestamp 1676557249
transform -1 0 21888 0 1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0926_
timestamp 1685173987
transform 1 0 19584 0 1 12852
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0927_
timestamp 1683973020
transform -1 0 20352 0 -1 12852
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__0928_
timestamp 1676901763
transform 1 0 16704 0 -1 11340
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0929_
timestamp 1685197497
transform 1 0 20352 0 -1 12852
box -48 -56 816 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0930_
timestamp 1685173987
transform -1 0 27744 0 -1 6804
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0931_
timestamp 1676627187
transform 1 0 24288 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0932_
timestamp 1683973020
transform -1 0 24096 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__0933_
timestamp 1683988354
transform -1 0 23520 0 -1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0934_
timestamp 1683973020
transform -1 0 23040 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0935_
timestamp 1685175443
transform 1 0 21216 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0936_
timestamp 1676627187
transform -1 0 22752 0 -1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0937_
timestamp 1683973020
transform 1 0 16224 0 1 2268
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0938_
timestamp 1677516600
transform 1 0 16608 0 -1 2268
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0939_
timestamp 1683973020
transform -1 0 18336 0 -1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0940_
timestamp 1685175443
transform 1 0 18240 0 1 2268
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0941_
timestamp 1685173987
transform 1 0 19104 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0942_
timestamp 1685175443
transform -1 0 20160 0 1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0943_
timestamp 1685173987
transform 1 0 20448 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0944_
timestamp 1685175443
transform 1 0 20832 0 1 8316
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0945_
timestamp 1685173987
transform 1 0 22944 0 1 6804
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__0946_
timestamp 1677175127
transform 1 0 21120 0 1 6804
box -48 -56 720 834
use sg13g2_and3_1  u_ppwm_u_ex__0947_
timestamp 1676971669
transform -1 0 21120 0 1 5292
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0948_
timestamp 1685175443
transform -1 0 19584 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0949_
timestamp 1683973020
transform 1 0 19200 0 1 756
box -48 -56 528 834
use sg13g2_or4_1  u_ppwm_u_ex__0950_
timestamp 1677154604
transform -1 0 17472 0 1 2268
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0951_
timestamp 1685175443
transform 1 0 15744 0 1 2268
box -48 -56 538 834
use sg13g2_and2_1  u_ppwm_u_ex__0952_
timestamp 1676901763
transform 1 0 16704 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0953_
timestamp 1685175443
transform -1 0 18144 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0954_
timestamp 1676627187
transform -1 0 20736 0 1 6804
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__0955_
timestamp 1677577977
transform -1 0 19776 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0956_
timestamp 1683973020
transform 1 0 17472 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0957_
timestamp 1685175443
transform -1 0 19008 0 1 3780
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0958_
timestamp 1685173987
transform 1 0 17856 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0959_
timestamp 1685175443
transform 1 0 18432 0 -1 12852
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0960_
timestamp 1685173987
transform 1 0 18720 0 1 11340
box -48 -56 624 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0961_
timestamp 1685173987
transform 1 0 23616 0 -1 6804
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_ex__0962_
timestamp 1676627187
transform -1 0 24576 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0963_
timestamp 1683973020
transform 1 0 22944 0 1 5292
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_ex__0964_
timestamp 1685201930
transform -1 0 19008 0 1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0965_
timestamp 1685175443
transform 1 0 12864 0 1 5292
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0966_
timestamp 1685181386
transform -1 0 14016 0 -1 6804
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0967_
timestamp 1683973020
transform -1 0 19200 0 -1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0968_
timestamp 1677516600
transform -1 0 18240 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0969_
timestamp 1683973020
transform -1 0 19104 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0970_
timestamp 1685175443
transform -1 0 16992 0 1 5292
box -48 -56 538 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0971_
timestamp 1685173987
transform 1 0 17568 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0972_
timestamp 1685175443
transform -1 0 18528 0 1 11340
box -48 -56 538 834
use sg13g2_nor3_1  u_ppwm_u_ex__0973_
timestamp 1676639442
transform 1 0 22656 0 1 9828
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__0974_
timestamp 1685197497
transform 1 0 23136 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0975_
timestamp 1685175443
transform -1 0 22464 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0976_
timestamp 1683973020
transform 1 0 17664 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0977_
timestamp 1685175443
transform 1 0 16992 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0978_
timestamp 1683973020
transform 1 0 17472 0 1 8316
box -48 -56 528 834
use sg13g2_nor2_2  u_ppwm_u_ex__0979_
timestamp 1683979924
transform 1 0 31104 0 -1 8316
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__0980_
timestamp 1676557249
transform 1 0 32736 0 1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0981_
timestamp 1685173987
transform -1 0 33600 0 1 14364
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__0982_
timestamp 1677175127
transform 1 0 32352 0 1 14364
box -48 -56 720 834
use sg13g2_nor2_1  u_ppwm_u_ex__0983_
timestamp 1676627187
transform 1 0 24672 0 -1 17388
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0984_
timestamp 1685173987
transform -1 0 25152 0 1 17388
box -48 -56 624 834
use sg13g2_nor2b_1  u_ppwm_u_ex__0985_
timestamp 1685181386
transform -1 0 25536 0 -1 17388
box -54 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__0986_
timestamp 1676901763
transform 1 0 27840 0 -1 18900
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__0987_
timestamp 1677577977
transform -1 0 28704 0 1 18900
box -48 -56 816 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0988_
timestamp 1685173987
transform -1 0 28032 0 -1 17388
box -48 -56 624 834
use sg13g2_nand4_1  u_ppwm_u_ex__0989_
timestamp 1685201930
transform 1 0 32256 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__0990_
timestamp 1685175443
transform -1 0 33312 0 -1 18900
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__0991_
timestamp 1676627187
transform 1 0 32064 0 1 18900
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_ex__0992_
timestamp 1676901763
transform 1 0 28992 0 -1 20412
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__0993_
timestamp 1677577977
transform 1 0 28704 0 1 18900
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__0994_
timestamp 1677516600
transform 1 0 29472 0 1 18900
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_ex__0995_
timestamp 1676627187
transform -1 0 30624 0 -1 18900
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0996_
timestamp 1676557249
transform -1 0 31392 0 1 15876
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_ex__0997_
timestamp 1676557249
transform 1 0 31680 0 -1 14364
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__0998_
timestamp 1685173987
transform 1 0 32640 0 -1 14364
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_ex__0999_
timestamp 1683973020
transform 1 0 31392 0 1 14364
box -48 -56 528 834
use sg13g2_nor4_1  u_ppwm_u_ex__1000_
timestamp 1676643125
transform 1 0 31296 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1001_
timestamp 1685175443
transform 1 0 33024 0 1 17388
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_ex__1002_
timestamp 1676627187
transform -1 0 34368 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1003_
timestamp 1683973020
transform 1 0 29280 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__1004_
timestamp 1676557249
transform 1 0 29760 0 -1 18900
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__1005_
timestamp 1677516600
transform 1 0 28320 0 1 17388
box -48 -56 816 834
use sg13g2_or2_1  u_ppwm_u_ex__1006_
timestamp 1684236171
transform 1 0 29184 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1007_
timestamp 1683973020
transform -1 0 29760 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__1008_
timestamp 1676557249
transform 1 0 32256 0 -1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1009_
timestamp 1685173987
transform -1 0 32544 0 1 12852
box -48 -56 624 834
use sg13g2_nand2_1  u_ppwm_u_ex__1010_
timestamp 1676557249
transform -1 0 31872 0 1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1011_
timestamp 1685173987
transform -1 0 30048 0 -1 17388
box -48 -56 624 834
use sg13g2_nand4_1  u_ppwm_u_ex__1012_
timestamp 1685201930
transform 1 0 29568 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1013_
timestamp 1685175443
transform 1 0 37056 0 1 15876
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__1014_
timestamp 1685181386
transform 1 0 36576 0 1 15876
box -54 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__1015_
timestamp 1677516600
transform -1 0 29088 0 -1 18900
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1016_
timestamp 1683973020
transform 1 0 28992 0 -1 17388
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_ex__1017_
timestamp 1683988354
transform 1 0 29664 0 1 17388
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__1018_
timestamp 1676627187
transform -1 0 31296 0 1 17388
box -48 -56 432 834
use sg13g2_nor3_1  u_ppwm_u_ex__1019_
timestamp 1676639442
transform 1 0 31872 0 1 11340
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__1020_
timestamp 1685197497
transform 1 0 31488 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1021_
timestamp 1685175443
transform -1 0 31872 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1022_
timestamp 1683973020
transform 1 0 30432 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1023_
timestamp 1685175443
transform -1 0 31296 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1024_
timestamp 1683973020
transform -1 0 30816 0 -1 17388
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__1025_
timestamp 1676627187
transform -1 0 28512 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__1026_
timestamp 1677577977
transform -1 0 29664 0 1 3780
box -48 -56 816 834
use sg13g2_or2_1  u_ppwm_u_ex__1027_
timestamp 1684236171
transform 1 0 27840 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1028_
timestamp 1685175443
transform 1 0 28032 0 -1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1029_
timestamp 1685175443
transform -1 0 28992 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1030_
timestamp 1683973020
transform 1 0 28128 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1031_
timestamp 1685175443
transform 1 0 29568 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__1032_
timestamp 1676557249
transform -1 0 33216 0 1 5292
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1033_
timestamp 1685173987
transform -1 0 32736 0 1 6804
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__1034_
timestamp 1677175127
transform 1 0 31488 0 1 5292
box -48 -56 720 834
use sg13g2_nand4_1  u_ppwm_u_ex__1035_
timestamp 1685201930
transform -1 0 31296 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1036_
timestamp 1685175443
transform 1 0 31200 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__1037_
timestamp 1685181386
transform 1 0 31680 0 -1 3780
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1038_
timestamp 1683973020
transform 1 0 29088 0 -1 5292
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_ex__1039_
timestamp 1677577977
transform 1 0 28032 0 1 2268
box -48 -56 816 834
use sg13g2_xnor2_1  u_ppwm_u_ex__1040_
timestamp 1677516600
transform 1 0 28608 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1041_
timestamp 1683973020
transform 1 0 28608 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1042_
timestamp 1685175443
transform 1 0 29568 0 1 5292
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__1043_
timestamp 1676557249
transform -1 0 31584 0 -1 6804
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1044_
timestamp 1685173987
transform 1 0 31776 0 -1 8316
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__1045_
timestamp 1677175127
transform 1 0 31296 0 1 6804
box -48 -56 720 834
use sg13g2_nand4_1  u_ppwm_u_ex__1046_
timestamp 1685201930
transform -1 0 30720 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1047_
timestamp 1685175443
transform -1 0 31776 0 1 3780
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__1048_
timestamp 1685181386
transform 1 0 31008 0 1 5292
box -54 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_ex__1049_
timestamp 1676627187
transform -1 0 28896 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_ex__1050_
timestamp 1677577977
transform -1 0 28032 0 1 2268
box -48 -56 816 834
use sg13g2_inv_1  u_ppwm_u_ex__1051_
timestamp 1676382929
transform -1 0 27264 0 1 2268
box -48 -56 336 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1052_
timestamp 1683973020
transform 1 0 28896 0 -1 6804
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_ex__1053_
timestamp 1676901763
transform 1 0 28512 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__1054_
timestamp 1676557249
transform -1 0 29952 0 -1 3780
box -48 -56 432 834
use sg13g2_a21o_1  u_ppwm_u_ex__1055_
timestamp 1677175127
transform 1 0 28224 0 1 3780
box -48 -56 720 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1056_
timestamp 1683973020
transform 1 0 27552 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1057_
timestamp 1685175443
transform 1 0 28032 0 -1 3780
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__1058_
timestamp 1676557249
transform 1 0 31584 0 -1 6804
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1059_
timestamp 1685173987
transform 1 0 32736 0 1 6804
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__1060_
timestamp 1677175127
transform 1 0 32160 0 1 5292
box -48 -56 720 834
use sg13g2_nand4_1  u_ppwm_u_ex__1061_
timestamp 1685201930
transform -1 0 29568 0 -1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1062_
timestamp 1685175443
transform -1 0 30048 0 1 2268
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__1063_
timestamp 1685181386
transform 1 0 29088 0 1 2268
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1064_
timestamp 1683973020
transform -1 0 28224 0 1 3780
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_ex__1065_
timestamp 1677516600
transform -1 0 27264 0 1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1066_
timestamp 1683973020
transform -1 0 26496 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1067_
timestamp 1685175443
transform -1 0 26496 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__1068_
timestamp 1676557249
transform -1 0 24288 0 1 5292
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1069_
timestamp 1685173987
transform 1 0 23040 0 -1 6804
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1070_
timestamp 1683973020
transform -1 0 23904 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_ex__1071_
timestamp 1676557249
transform -1 0 21600 0 1 5292
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_ex__1072_
timestamp 1676627187
transform -1 0 23040 0 -1 5292
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1073_
timestamp 1685175443
transform -1 0 24384 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1074_
timestamp 1683973020
transform 1 0 25536 0 1 3780
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_ex__1075_
timestamp 1676639442
transform 1 0 27264 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1076_
timestamp 1685175443
transform 1 0 26496 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_ex__1077_
timestamp 1676567195
transform -1 0 27456 0 -1 5292
box -48 -56 528 834
use sg13g2_a21oi_2  u_ppwm_u_ex__1078_
timestamp 1685174172
transform -1 0 28224 0 -1 5292
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_ex__1079_
timestamp 1676557249
transform 1 0 15840 0 -1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_ex__1080_
timestamp 1677516600
transform -1 0 18240 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1081_
timestamp 1683973020
transform -1 0 18048 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1082_
timestamp 1685175443
transform 1 0 17184 0 -1 3780
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_ex__1083_
timestamp 1676557249
transform -1 0 25056 0 1 5292
box -48 -56 432 834
use sg13g2_a22oi_1  u_ppwm_u_ex__1084_
timestamp 1685173987
transform 1 0 22464 0 -1 6804
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_ex__1085_
timestamp 1677175127
transform 1 0 21984 0 1 5292
box -48 -56 720 834
use sg13g2_nand4_1  u_ppwm_u_ex__1086_
timestamp 1685201930
transform 1 0 17856 0 -1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1087_
timestamp 1685175443
transform -1 0 19488 0 -1 5292
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_ex__1088_
timestamp 1685181386
transform 1 0 18048 0 1 3780
box -54 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1089_
timestamp 1685175443
transform -1 0 17376 0 1 3780
box -48 -56 538 834
use sg13g2_xor2_1  u_ppwm_u_ex__1090_
timestamp 1677577977
transform -1 0 17760 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1091_
timestamp 1683973020
transform -1 0 16512 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1092_
timestamp 1685175443
transform 1 0 19200 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1093_
timestamp 1683973020
transform -1 0 24000 0 -1 11340
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_ex__1094_
timestamp 1685197497
transform 1 0 23904 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1095_
timestamp 1685175443
transform -1 0 24480 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1096_
timestamp 1683973020
transform -1 0 19872 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_ex__1097_
timestamp 1685175443
transform 1 0 19680 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_ex__1098_
timestamp 1683973020
transform 1 0 16992 0 1 5292
box -48 -56 528 834
use sg13g2_tiehi  u_ppwm_u_ex__1099__52
timestamp 1680000651
transform -1 0 27552 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1099_
timestamp 1746535128
transform 1 0 26688 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1100__51
timestamp 1680000651
transform -1 0 27072 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1100_
timestamp 1746535184
transform 1 0 25728 0 -1 23436
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1101_
timestamp 1746535184
transform 1 0 22848 0 -1 23436
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1101__49
timestamp 1680000651
transform -1 0 23712 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__1102__47
timestamp 1680000651
transform 1 0 19488 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1102_
timestamp 1746535128
transform 1 0 19872 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1103__45
timestamp 1680000651
transform -1 0 14880 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1103_
timestamp 1746535128
transform 1 0 13824 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1104__43
timestamp 1680000651
transform 1 0 14880 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1104_
timestamp 1746535184
transform -1 0 15744 0 -1 15876
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1105__41
timestamp 1680000651
transform -1 0 36288 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1105_
timestamp 1746535184
transform 1 0 35328 0 -1 15876
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1106__39
timestamp 1680000651
transform -1 0 40032 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1106_
timestamp 1746535128
transform 1 0 39168 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1107__37
timestamp 1680000651
transform -1 0 39840 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1107_
timestamp 1746535184
transform 1 0 38976 0 1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1108_
timestamp 1746535184
transform 1 0 29472 0 -1 20412
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1108__35
timestamp 1680000651
transform -1 0 30336 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__1109__33
timestamp 1680000651
transform -1 0 32640 0 -1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1109_
timestamp 1746535128
transform 1 0 31776 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1110__31
timestamp 1680000651
transform -1 0 22560 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1110_
timestamp 1746535128
transform 1 0 21696 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1111__29
timestamp 1680000651
transform -1 0 23712 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1111_
timestamp 1746535128
transform 1 0 22848 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1112__27
timestamp 1680000651
transform 1 0 18528 0 -1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1112_
timestamp 1746535184
transform 1 0 18912 0 -1 2268
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1113__50
timestamp 1680000651
transform -1 0 14400 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1113_
timestamp 1746535184
transform 1 0 13344 0 1 5292
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1114__46
timestamp 1680000651
transform -1 0 14400 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1114_
timestamp 1746535128
transform 1 0 13536 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1115__42
timestamp 1680000651
transform -1 0 33312 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1115_
timestamp 1746535184
transform 1 0 32448 0 1 18900
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1116__38
timestamp 1680000651
transform -1 0 35520 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1116_
timestamp 1746535184
transform 1 0 34464 0 -1 18900
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1117_
timestamp 1746535128
transform 1 0 37248 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1117__34
timestamp 1680000651
transform 1 0 37536 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1118_
timestamp 1746535184
transform 1 0 33216 0 -1 17388
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1118__30
timestamp 1680000651
transform -1 0 34080 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1119_
timestamp 1746535128
transform 1 0 33216 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1119__26
timestamp 1680000651
transform -1 0 34080 0 -1 3780
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__1120__44
timestamp 1680000651
transform -1 0 32736 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1120_
timestamp 1746535184
transform 1 0 31488 0 -1 2268
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1121__36
timestamp 1680000651
transform -1 0 29952 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1121_
timestamp 1746535184
transform 1 0 28800 0 -1 2268
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1122_
timestamp 1746535184
transform 1 0 25536 0 -1 2268
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1122__28
timestamp 1680000651
transform -1 0 26400 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1123_
timestamp 1746535184
transform -1 0 16704 0 1 3780
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1123__40
timestamp 1680000651
transform 1 0 14784 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_ex__1124_
timestamp 1746535184
transform 1 0 14304 0 1 6804
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_ex__1124__53
timestamp 1680000651
transform -1 0 15168 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1125_
timestamp 1746535128
transform -1 0 17280 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1125__54
timestamp 1680000651
transform 1 0 16224 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1126_
timestamp 1746535128
transform 1 0 14688 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_ex__1126__32
timestamp 1680000651
transform 1 0 14976 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_ex__1127__48
timestamp 1680000651
transform 1 0 16704 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_ex__1127_
timestamp 1746535128
transform 1 0 16896 0 1 18900
box -48 -56 2640 834
use sg13g2_inv_1  u_ppwm_u_global_counter__053_
timestamp 1676382929
transform -1 0 41280 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__054_
timestamp 1676382929
transform -1 0 44928 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__055_
timestamp 1676382929
transform 1 0 38112 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__056_
timestamp 1676382929
transform 1 0 38496 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__057_
timestamp 1676382929
transform 1 0 37056 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__058_
timestamp 1676382929
transform -1 0 38304 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_global_counter__059_
timestamp 1676382929
transform 1 0 43872 0 -1 11340
box -48 -56 336 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__060_
timestamp 1677577977
transform 1 0 42720 0 1 12852
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__061_
timestamp 1683988354
transform -1 0 42144 0 1 12852
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_global_counter__062_
timestamp 1677175127
transform -1 0 41472 0 1 14364
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__063_
timestamp 1676901763
transform -1 0 42144 0 -1 14364
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__064_
timestamp 1685201930
transform 1 0 41760 0 -1 12852
box -48 -56 624 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__065_
timestamp 1677516600
transform 1 0 40032 0 1 11340
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__066_
timestamp 1676627187
transform 1 0 41664 0 -1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__067_
timestamp 1677516600
transform 1 0 42336 0 -1 12852
box -48 -56 816 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__068_
timestamp 1677577977
transform 1 0 41376 0 1 6804
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__069_
timestamp 1685201930
transform -1 0 41856 0 1 8316
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__070_
timestamp 1676627187
transform 1 0 39744 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__071_
timestamp 1683973020
transform -1 0 43008 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__072_
timestamp 1676627187
transform 1 0 42144 0 1 5292
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__073_
timestamp 1677577977
transform 1 0 43872 0 1 5292
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__074_
timestamp 1685201930
transform 1 0 43104 0 1 6804
box -48 -56 624 834
use sg13g2_nor3_2  u_ppwm_u_global_counter__075_
timestamp 1685180723
transform 1 0 44256 0 -1 9828
box -48 -56 912 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__076_
timestamp 1683973020
transform 1 0 44640 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_global_counter__077_
timestamp 1676627187
transform -1 0 45600 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__078_
timestamp 1677577977
transform -1 0 47136 0 1 6804
box -48 -56 816 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__079_
timestamp 1683988354
transform -1 0 47520 0 1 12852
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_global_counter__080_
timestamp 1677175127
transform 1 0 42816 0 1 9828
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__081_
timestamp 1676901763
transform 1 0 48768 0 -1 11340
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__082_
timestamp 1685201930
transform 1 0 48192 0 -1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  u_ppwm_u_global_counter__083_
timestamp 1677516600
transform 1 0 46080 0 1 11340
box -48 -56 816 834
use sg13g2_nand4_1  u_ppwm_u_global_counter__084_
timestamp 1685201930
transform 1 0 42048 0 -1 11340
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_global_counter__085_
timestamp 1676639442
transform -1 0 43392 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__086_
timestamp 1685173987
transform 1 0 42144 0 1 12852
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__087_
timestamp 1683973020
transform 1 0 37632 0 -1 11340
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__088_
timestamp 1683988354
transform 1 0 38592 0 -1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_global_counter__089_
timestamp 1685181386
transform 1 0 37440 0 1 9828
box -54 -56 528 834
use sg13g2_and3_2  u_ppwm_u_global_counter__090_
timestamp 1683976310
transform -1 0 39840 0 1 11340
box -48 -56 720 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__091_
timestamp 1685173987
transform 1 0 38400 0 -1 9828
box -48 -56 624 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__092_
timestamp 1683973020
transform -1 0 38400 0 -1 8316
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__093_
timestamp 1683988354
transform 1 0 37248 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_global_counter__094_
timestamp 1685181386
transform 1 0 37536 0 1 8316
box -54 -56 528 834
use sg13g2_and3_2  u_ppwm_u_global_counter__095_
timestamp 1683976310
transform -1 0 38400 0 1 6804
box -48 -56 720 834
use sg13g2_and2_1  u_ppwm_u_global_counter__096_
timestamp 1676901763
transform -1 0 37920 0 -1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__097_
timestamp 1683973020
transform 1 0 40608 0 1 5292
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__098_
timestamp 1683988354
transform -1 0 38400 0 1 2268
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__099_
timestamp 1677577977
transform 1 0 38208 0 -1 6804
box -48 -56 816 834
use sg13g2_and2_1  u_ppwm_u_global_counter__100_
timestamp 1676901763
transform 1 0 35232 0 -1 6804
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_global_counter__101_
timestamp 1683988354
transform 1 0 35712 0 -1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  u_ppwm_u_global_counter__102_
timestamp 1685173987
transform 1 0 36864 0 1 5292
box -48 -56 624 834
use sg13g2_and4_1  u_ppwm_u_global_counter__103_
timestamp 1676985977
transform -1 0 38208 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  u_ppwm_u_global_counter__104_
timestamp 1683973020
transform -1 0 37920 0 1 2268
box -48 -56 528 834
use sg13g2_xor2_1  u_ppwm_u_global_counter__105_
timestamp 1677577977
transform 1 0 35808 0 1 3780
box -48 -56 816 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__106_
timestamp 1746535184
transform 1 0 44064 0 -1 14364
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__107_
timestamp 1746535184
transform 1 0 41664 0 1 14364
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_global_counter__108_
timestamp 1746535128
transform 1 0 40800 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__109_
timestamp 1746535184
transform 1 0 43968 0 -1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__110_
timestamp 1746535184
transform -1 0 44544 0 -1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__111_
timestamp 1746535184
transform -1 0 44448 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__112_
timestamp 1746535184
transform -1 0 47232 0 -1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__113_
timestamp 1746535184
transform -1 0 47424 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__114_
timestamp 1746535184
transform 1 0 46560 0 1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__115_
timestamp 1746535184
transform -1 0 49536 0 1 9828
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__116_
timestamp 1746535184
transform 1 0 46848 0 1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__117_
timestamp 1746535184
transform 1 0 44352 0 1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__118_
timestamp 1746535184
transform -1 0 42720 0 1 9828
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__119_
timestamp 1746535184
transform 1 0 38976 0 -1 9828
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__120_
timestamp 1746535184
transform -1 0 41568 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__121_
timestamp 1746535184
transform 1 0 39168 0 -1 6804
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__122_
timestamp 1746535184
transform 1 0 39168 0 -1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__123_
timestamp 1746535184
transform -1 0 37920 0 -1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__124_
timestamp 1746535184
transform 1 0 38304 0 1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_global_counter__125_
timestamp 1746535184
transform -1 0 39744 0 -1 3780
box -48 -56 2736 834
use sg13g2_inv_1  u_ppwm_u_mem__0613_
timestamp 1676382929
transform -1 0 4992 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0614_
timestamp 1676382929
transform 1 0 6048 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0615_
timestamp 1676382929
transform -1 0 4608 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0616_
timestamp 1676382929
transform -1 0 1056 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0617_
timestamp 1676382929
transform 1 0 5376 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0618_
timestamp 1676382929
transform -1 0 9792 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0619_
timestamp 1676382929
transform 1 0 12960 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0620_
timestamp 1676382929
transform -1 0 7680 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0621_
timestamp 1676382929
transform -1 0 5664 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0622_
timestamp 1676382929
transform -1 0 3936 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0623_
timestamp 1676382929
transform -1 0 3264 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0624_
timestamp 1676382929
transform 1 0 4320 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0625_
timestamp 1676382929
transform 1 0 9216 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0626_
timestamp 1676382929
transform 1 0 13056 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0627_
timestamp 1676382929
transform 1 0 14496 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0628_
timestamp 1676382929
transform -1 0 16512 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0629_
timestamp 1676382929
transform -1 0 18816 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0630_
timestamp 1676382929
transform -1 0 20832 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0631_
timestamp 1676382929
transform -1 0 20928 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0632_
timestamp 1676382929
transform -1 0 14976 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0633_
timestamp 1676382929
transform 1 0 11616 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0634_
timestamp 1676382929
transform -1 0 9504 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0635_
timestamp 1676382929
transform -1 0 14592 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0636_
timestamp 1676382929
transform 1 0 16896 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0637_
timestamp 1676382929
transform -1 0 17952 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0638_
timestamp 1676382929
transform -1 0 18816 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0639_
timestamp 1676382929
transform -1 0 14688 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0640_
timestamp 1676382929
transform -1 0 6720 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0641_
timestamp 1676382929
transform -1 0 5952 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0642_
timestamp 1676382929
transform -1 0 2976 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0643_
timestamp 1676382929
transform -1 0 2592 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0644_
timestamp 1676382929
transform 1 0 7584 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0645_
timestamp 1676382929
transform 1 0 9600 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0646_
timestamp 1676382929
transform -1 0 12672 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0647_
timestamp 1676382929
transform -1 0 13440 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0648_
timestamp 1676382929
transform -1 0 7584 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0649_
timestamp 1676382929
transform -1 0 2784 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0650_
timestamp 1676382929
transform -1 0 2880 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0651_
timestamp 1676382929
transform 1 0 6624 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0652_
timestamp 1676382929
transform -1 0 9600 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0653_
timestamp 1676382929
transform -1 0 14496 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0654_
timestamp 1676382929
transform -1 0 16512 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0655_
timestamp 1676382929
transform -1 0 14784 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0656_
timestamp 1676382929
transform -1 0 6528 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0657_
timestamp 1676382929
transform 1 0 6048 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0658_
timestamp 1676382929
transform 1 0 6432 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0659_
timestamp 1676382929
transform 1 0 9504 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0660_
timestamp 1676382929
transform 1 0 14784 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0661_
timestamp 1676382929
transform 1 0 18144 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0662_
timestamp 1676382929
transform -1 0 20064 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0663_
timestamp 1676382929
transform -1 0 6240 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0664_
timestamp 1676382929
transform 1 0 6240 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0665_
timestamp 1676382929
transform -1 0 7200 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0666_
timestamp 1676382929
transform 1 0 9984 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0667_
timestamp 1676382929
transform 1 0 17472 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0668_
timestamp 1676382929
transform 1 0 21024 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0669_
timestamp 1676382929
transform -1 0 23712 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0670_
timestamp 1676382929
transform -1 0 25728 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0671_
timestamp 1676382929
transform 1 0 28032 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0672_
timestamp 1676382929
transform -1 0 31008 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0673_
timestamp 1676382929
transform 1 0 33696 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0674_
timestamp 1676382929
transform 1 0 35616 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0675_
timestamp 1676382929
transform -1 0 37248 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0676_
timestamp 1676382929
transform -1 0 26784 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0677_
timestamp 1676382929
transform 1 0 26304 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0678_
timestamp 1676382929
transform -1 0 28896 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0679_
timestamp 1676382929
transform 1 0 33024 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0680_
timestamp 1676382929
transform -1 0 35328 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0681_
timestamp 1676382929
transform 1 0 39552 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0682_
timestamp 1676382929
transform -1 0 40224 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0683_
timestamp 1676382929
transform -1 0 33024 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0684_
timestamp 1676382929
transform -1 0 29376 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0685_
timestamp 1676382929
transform -1 0 21888 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0686_
timestamp 1676382929
transform 1 0 27648 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0687_
timestamp 1676382929
transform 1 0 29664 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0688_
timestamp 1676382929
transform -1 0 32256 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0689_
timestamp 1676382929
transform -1 0 32448 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0690_
timestamp 1676382929
transform -1 0 26592 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0691_
timestamp 1676382929
transform -1 0 24960 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0692_
timestamp 1676382929
transform 1 0 26592 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0693_
timestamp 1676382929
transform 1 0 32352 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0694_
timestamp 1676382929
transform -1 0 33504 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0695_
timestamp 1676382929
transform -1 0 35520 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0696_
timestamp 1676382929
transform -1 0 34656 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0697_
timestamp 1676382929
transform 1 0 34080 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0698_
timestamp 1676382929
transform 1 0 38496 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0699_
timestamp 1676382929
transform 1 0 40320 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0700_
timestamp 1676382929
transform -1 0 43392 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0701_
timestamp 1676382929
transform -1 0 46272 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0702_
timestamp 1676382929
transform -1 0 45504 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0703_
timestamp 1676382929
transform -1 0 44160 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0704_
timestamp 1676382929
transform -1 0 39456 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0705_
timestamp 1676382929
transform 1 0 39360 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0706_
timestamp 1676382929
transform 1 0 42048 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0707_
timestamp 1676382929
transform 1 0 45600 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0708_
timestamp 1676382929
transform -1 0 48000 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0709_
timestamp 1676382929
transform -1 0 45696 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0710_
timestamp 1676382929
transform -1 0 44064 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0711_
timestamp 1676382929
transform -1 0 40320 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0712_
timestamp 1676382929
transform -1 0 40992 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0713_
timestamp 1676382929
transform -1 0 43968 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0714_
timestamp 1676382929
transform -1 0 46944 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0715_
timestamp 1676382929
transform -1 0 48000 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0716_
timestamp 1676382929
transform -1 0 44352 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0717_
timestamp 1676382929
transform -1 0 39744 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0718_
timestamp 1676382929
transform 1 0 39552 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0719_
timestamp 1676382929
transform -1 0 40224 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0720_
timestamp 1676382929
transform -1 0 43008 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0721_
timestamp 1676382929
transform 1 0 44928 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0722_
timestamp 1676382929
transform -1 0 49248 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0723_
timestamp 1676382929
transform -1 0 49248 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0724_
timestamp 1676382929
transform -1 0 36768 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_mem__0725_
timestamp 1676382947
transform -1 0 6816 0 -1 14364
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_mem__0726_
timestamp 1676382929
transform -1 0 8640 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0727_
timestamp 1676382929
transform -1 0 36384 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_mem__0728_
timestamp 1676382929
transform 1 0 26016 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_4  u_ppwm_u_mem__0729_
timestamp 1676383058
transform -1 0 23040 0 1 24948
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_mem__0730_
timestamp 1676639442
transform 1 0 6432 0 1 17388
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__0731_
timestamp 1676627187
transform -1 0 8160 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0732_
timestamp 1683973020
transform 1 0 7968 0 -1 18900
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_mem__0733_
timestamp 1683988354
transform 1 0 5952 0 -1 14364
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_mem__0734_
timestamp 1683988354
transform 1 0 4512 0 -1 14364
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__0735_
timestamp 1676639442
transform -1 0 6912 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_mem__0736_
timestamp 1676557249
transform -1 0 7296 0 1 18900
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_mem__0737_
timestamp 1676643125
transform 1 0 6336 0 -1 17388
box -48 -56 624 834
use sg13g2_a21o_1  u_ppwm_u_mem__0738_
timestamp 1677175127
transform -1 0 7584 0 -1 17388
box -48 -56 720 834
use sg13g2_nand3_1  u_ppwm_u_mem__0739_
timestamp 1683988354
transform -1 0 6624 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0740_
timestamp 1685175443
transform -1 0 7104 0 -1 18900
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0741_
timestamp 1677247768
transform 1 0 15360 0 -1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0742_
timestamp 1677247768
transform -1 0 22176 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0743_
timestamp 1676557249
transform -1 0 17280 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0744_
timestamp 1683973020
transform -1 0 16416 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0745_
timestamp 1677247768
transform 1 0 10656 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0746_
timestamp 1676557249
transform 1 0 15168 0 -1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0747_
timestamp 1677247768
transform 1 0 13344 0 1 21924
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0748_
timestamp 1683973020
transform -1 0 15360 0 1 24948
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0749_
timestamp 1685197497
transform 1 0 15648 0 -1 26460
box -48 -56 816 834
use sg13g2_mux4_1  u_ppwm_u_mem__0750_
timestamp 1677257233
transform -1 0 40128 0 1 20412
box -48 -56 2064 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0751_
timestamp 1676567195
transform -1 0 24576 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0752_
timestamp 1677247768
transform -1 0 31584 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0753_
timestamp 1677247768
transform -1 0 30912 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0754_
timestamp 1676557249
transform -1 0 29952 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0755_
timestamp 1683973020
transform 1 0 29568 0 -1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0756_
timestamp 1683973020
transform -1 0 30432 0 -1 24948
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0757_
timestamp 1683996397
transform 1 0 23040 0 1 24948
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0758_
timestamp 1677247768
transform 1 0 12096 0 1 21924
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0759_
timestamp 1677247768
transform 1 0 11040 0 -1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0760_
timestamp 1676557249
transform 1 0 14880 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0761_
timestamp 1683973020
transform -1 0 15840 0 -1 24948
box -48 -56 528 834
use sg13g2_mux4_1  u_ppwm_u_mem__0762_
timestamp 1677257233
transform -1 0 18048 0 -1 34020
box -48 -56 2064 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0763_
timestamp 1685175443
transform 1 0 16512 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0764_
timestamp 1683973020
transform -1 0 16512 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_mem__0765_
timestamp 1676557249
transform 1 0 32832 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0766_
timestamp 1685175443
transform 1 0 33312 0 1 23436
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0767_
timestamp 1676557249
transform 1 0 35616 0 1 29484
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0768_
timestamp 1685175443
transform 1 0 37152 0 -1 29484
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0769_
timestamp 1676557249
transform 1 0 40704 0 1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0770_
timestamp 1685175443
transform -1 0 42048 0 1 21924
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0771_
timestamp 1676557249
transform 1 0 38688 0 -1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0772_
timestamp 1685175443
transform -1 0 38208 0 -1 20412
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0773_
timestamp 1677257233
transform -1 0 38496 0 1 23436
box -48 -56 2064 834
use sg13g2_a21o_2  u_ppwm_u_mem__0774_
timestamp 1683996397
transform 1 0 21312 0 -1 24948
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0775_
timestamp 1677247768
transform 1 0 9792 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0776_
timestamp 1676557249
transform 1 0 12480 0 1 24948
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0777_
timestamp 1677247768
transform -1 0 15936 0 -1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0778_
timestamp 1683973020
transform -1 0 15744 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0779_
timestamp 1677247768
transform 1 0 12576 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0780_
timestamp 1676557249
transform 1 0 13440 0 -1 29484
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0781_
timestamp 1677247768
transform -1 0 15456 0 1 35532
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0782_
timestamp 1683973020
transform -1 0 14976 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0783_
timestamp 1685197497
transform 1 0 14112 0 1 26460
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_mem__0784_
timestamp 1676557249
transform -1 0 35904 0 1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0785_
timestamp 1685175443
transform 1 0 35520 0 1 24948
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0786_
timestamp 1676557249
transform -1 0 37344 0 1 34020
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0787_
timestamp 1685175443
transform 1 0 36384 0 -1 32508
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0788_
timestamp 1676557249
transform 1 0 46080 0 1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0789_
timestamp 1685175443
transform -1 0 46656 0 -1 24948
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0790_
timestamp 1676557249
transform 1 0 42912 0 1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0791_
timestamp 1685175443
transform -1 0 43776 0 -1 23436
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0792_
timestamp 1677257233
transform -1 0 38400 0 1 24948
box -48 -56 2064 834
use sg13g2_a21o_2  u_ppwm_u_mem__0793_
timestamp 1683996397
transform 1 0 21696 0 1 24948
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0794_
timestamp 1677247768
transform 1 0 5664 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0795_
timestamp 1676557249
transform 1 0 8256 0 1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0796_
timestamp 1677247768
transform -1 0 18720 0 -1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0797_
timestamp 1683973020
transform 1 0 14496 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0798_
timestamp 1677247768
transform 1 0 9792 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0799_
timestamp 1676557249
transform 1 0 12096 0 -1 32508
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0800_
timestamp 1677247768
transform 1 0 10272 0 1 35532
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0801_
timestamp 1683973020
transform -1 0 13344 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0802_
timestamp 1685197497
transform 1 0 13344 0 1 26460
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0803_
timestamp 1677247768
transform -1 0 31872 0 -1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0804_
timestamp 1677247768
transform 1 0 30912 0 -1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0805_
timestamp 1683973020
transform 1 0 31296 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0806_
timestamp 1685175443
transform 1 0 30432 0 1 26460
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0807_
timestamp 1677257233
transform -1 0 47712 0 1 24948
box -48 -56 2064 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0808_
timestamp 1683973020
transform 1 0 30912 0 1 26460
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_mem__0809_
timestamp 1677175127
transform 1 0 30240 0 -1 26460
box -48 -56 720 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0810_
timestamp 1685175443
transform 1 0 3840 0 -1 24948
box -48 -56 538 834
use sg13g2_a21o_1  u_ppwm_u_mem__0811_
timestamp 1677175127
transform -1 0 6432 0 1 24948
box -48 -56 720 834
use sg13g2_mux2_1  u_ppwm_u_mem__0812_
timestamp 1677247768
transform 1 0 18912 0 -1 26460
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0813_
timestamp 1683973020
transform -1 0 20352 0 -1 26460
box -48 -56 528 834
use sg13g2_mux4_1  u_ppwm_u_mem__0814_
timestamp 1677257233
transform 1 0 6240 0 -1 34020
box -48 -56 2064 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0815_
timestamp 1685175443
transform 1 0 16992 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0816_
timestamp 1683973020
transform 1 0 17472 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0817_
timestamp 1677247768
transform -1 0 42720 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0818_
timestamp 1676557249
transform -1 0 37536 0 -1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0819_
timestamp 1677247768
transform -1 0 44832 0 -1 26460
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0820_
timestamp 1683973020
transform 1 0 28992 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0821_
timestamp 1685175443
transform -1 0 30432 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0822_
timestamp 1683973020
transform 1 0 30432 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0823_
timestamp 1677247768
transform 1 0 26880 0 1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0824_
timestamp 1683973020
transform -1 0 28224 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0825_
timestamp 1676567195
transform -1 0 29760 0 1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0826_
timestamp 1683973020
transform 1 0 28800 0 1 26460
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0827_
timestamp 1683996397
transform 1 0 28032 0 -1 26460
box -48 -56 816 834
use sg13g2_nor2b_1  u_ppwm_u_mem__0828_
timestamp 1685181386
transform -1 0 6240 0 -1 23436
box -54 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0829_
timestamp 1685175443
transform 1 0 5088 0 1 23436
box -48 -56 538 834
use sg13g2_nand2_1  u_ppwm_u_mem__0830_
timestamp 1676557249
transform 1 0 16320 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_mem__0831_
timestamp 1676567195
transform 1 0 16896 0 1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0832_
timestamp 1683973020
transform -1 0 17856 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0833_
timestamp 1685175443
transform 1 0 5376 0 -1 24948
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0834_
timestamp 1677257233
transform 1 0 4224 0 1 30996
box -48 -56 2064 834
use sg13g2_nor2_1  u_ppwm_u_mem__0835_
timestamp 1676627187
transform -1 0 8064 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0836_
timestamp 1685175443
transform 1 0 18048 0 -1 24948
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0837_
timestamp 1677247768
transform 1 0 25344 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0838_
timestamp 1677247768
transform 1 0 26592 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0839_
timestamp 1677247768
transform -1 0 39360 0 1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0840_
timestamp 1677247768
transform -1 0 42528 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux4_1  u_ppwm_u_mem__0841_
timestamp 1677257233
transform 1 0 26784 0 1 26460
box -48 -56 2064 834
use sg13g2_nand2_1  u_ppwm_u_mem__0842_
timestamp 1676557249
transform -1 0 22272 0 -1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0843_
timestamp 1685175443
transform 1 0 20832 0 -1 24948
box -48 -56 538 834
use sg13g2_mux2_1  u_ppwm_u_mem__0844_
timestamp 1677247768
transform 1 0 5472 0 -1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0845_
timestamp 1676557249
transform 1 0 6144 0 1 26460
box -48 -56 432 834
use sg13g2_mux2_1  u_ppwm_u_mem__0846_
timestamp 1677247768
transform 1 0 12960 0 -1 30996
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0847_
timestamp 1683973020
transform 1 0 13536 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  u_ppwm_u_mem__0848_
timestamp 1677247768
transform 1 0 13344 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0849_
timestamp 1677247768
transform 1 0 7680 0 1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  u_ppwm_u_mem__0850_
timestamp 1676557249
transform 1 0 8544 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0851_
timestamp 1683973020
transform -1 0 14496 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_mem__0852_
timestamp 1685197497
transform -1 0 13824 0 1 24948
box -48 -56 816 834
use sg13g2_mux2_1  u_ppwm_u_mem__0853_
timestamp 1677247768
transform 1 0 25440 0 -1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  u_ppwm_u_mem__0854_
timestamp 1677247768
transform 1 0 25440 0 -1 30996
box -48 -56 1008 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0855_
timestamp 1683973020
transform 1 0 25344 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0856_
timestamp 1685175443
transform 1 0 26304 0 -1 26460
box -48 -56 538 834
use sg13g2_mux4_1  u_ppwm_u_mem__0857_
timestamp 1677257233
transform -1 0 40800 0 -1 24948
box -48 -56 2064 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0858_
timestamp 1683973020
transform 1 0 26880 0 -1 24948
box -48 -56 528 834
use sg13g2_a21o_2  u_ppwm_u_mem__0859_
timestamp 1683996397
transform 1 0 26016 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0860_
timestamp 1685175443
transform -1 0 38304 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0861_
timestamp 1683973020
transform 1 0 38208 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0862_
timestamp 1685175443
transform 1 0 46944 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0863_
timestamp 1683973020
transform 1 0 47424 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0864_
timestamp 1685175443
transform 1 0 48000 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0865_
timestamp 1683973020
transform 1 0 48480 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0866_
timestamp 1685175443
transform 1 0 47328 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0867_
timestamp 1683973020
transform 1 0 48672 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0868_
timestamp 1685175443
transform -1 0 43584 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0869_
timestamp 1683973020
transform -1 0 43104 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0870_
timestamp 1685175443
transform -1 0 41568 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0871_
timestamp 1683973020
transform -1 0 40896 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0872_
timestamp 1685175443
transform 1 0 39840 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0873_
timestamp 1683973020
transform -1 0 40608 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0874_
timestamp 1685175443
transform -1 0 39072 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0875_
timestamp 1683973020
transform 1 0 38112 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0876_
timestamp 1685175443
transform 1 0 43776 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0877_
timestamp 1683973020
transform -1 0 43776 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0878_
timestamp 1685175443
transform 1 0 47136 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0879_
timestamp 1683973020
transform -1 0 48192 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0880_
timestamp 1685175443
transform 1 0 50880 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0881_
timestamp 1683973020
transform -1 0 45696 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0882_
timestamp 1685175443
transform -1 0 44928 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0883_
timestamp 1683973020
transform -1 0 44064 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0884_
timestamp 1685175443
transform 1 0 40896 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0885_
timestamp 1683973020
transform -1 0 41856 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0886_
timestamp 1685175443
transform 1 0 41856 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0887_
timestamp 1683973020
transform -1 0 41568 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0888_
timestamp 1685175443
transform 1 0 40224 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0889_
timestamp 1683973020
transform 1 0 40704 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0890_
timestamp 1685175443
transform 1 0 45984 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0891_
timestamp 1683973020
transform -1 0 47616 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0892_
timestamp 1685175443
transform 1 0 46656 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0893_
timestamp 1683973020
transform -1 0 48192 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0894_
timestamp 1685175443
transform -1 0 44448 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0895_
timestamp 1683973020
transform -1 0 43776 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0896_
timestamp 1685175443
transform -1 0 42912 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0897_
timestamp 1683973020
transform -1 0 40896 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0898_
timestamp 1685175443
transform 1 0 38688 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0899_
timestamp 1683973020
transform 1 0 39360 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0900_
timestamp 1685175443
transform 1 0 38880 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0901_
timestamp 1683973020
transform 1 0 39168 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0902_
timestamp 1685175443
transform -1 0 42624 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0903_
timestamp 1683973020
transform -1 0 42144 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0904_
timestamp 1685175443
transform 1 0 44256 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0905_
timestamp 1683973020
transform -1 0 44640 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0906_
timestamp 1685175443
transform -1 0 46080 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0907_
timestamp 1683973020
transform 1 0 45504 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0908_
timestamp 1685175443
transform -1 0 44256 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0909_
timestamp 1683973020
transform -1 0 43296 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0910_
timestamp 1685175443
transform -1 0 41568 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0911_
timestamp 1683973020
transform -1 0 41088 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0912_
timestamp 1685175443
transform -1 0 38208 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0913_
timestamp 1683973020
transform 1 0 38208 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0914_
timestamp 1685175443
transform 1 0 33792 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0915_
timestamp 1683973020
transform -1 0 34752 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0916_
timestamp 1685175443
transform 1 0 32256 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0917_
timestamp 1683973020
transform 1 0 32544 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0918_
timestamp 1685175443
transform 1 0 35136 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0919_
timestamp 1683973020
transform -1 0 35040 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0920_
timestamp 1685175443
transform -1 0 34080 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0921_
timestamp 1683973020
transform -1 0 33504 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0922_
timestamp 1685175443
transform 1 0 32832 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0923_
timestamp 1683973020
transform 1 0 31680 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0924_
timestamp 1685175443
transform 1 0 26400 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0925_
timestamp 1683973020
transform -1 0 27360 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0926_
timestamp 1685175443
transform -1 0 25344 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0927_
timestamp 1683973020
transform 1 0 24960 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0928_
timestamp 1685175443
transform -1 0 25248 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0929_
timestamp 1683973020
transform 1 0 24576 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0930_
timestamp 1685175443
transform -1 0 31872 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0931_
timestamp 1683973020
transform -1 0 31392 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0932_
timestamp 1685175443
transform -1 0 32736 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0933_
timestamp 1683973020
transform -1 0 31392 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0934_
timestamp 1685175443
transform -1 0 32352 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0935_
timestamp 1683973020
transform -1 0 31872 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0936_
timestamp 1685175443
transform -1 0 28512 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0937_
timestamp 1683973020
transform -1 0 27744 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0938_
timestamp 1685175443
transform 1 0 22656 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0939_
timestamp 1683973020
transform -1 0 22368 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0940_
timestamp 1685175443
transform 1 0 22464 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0941_
timestamp 1683973020
transform 1 0 22944 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0942_
timestamp 1685175443
transform -1 0 32640 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0943_
timestamp 1683973020
transform 1 0 30432 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0944_
timestamp 1685175443
transform -1 0 37344 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0945_
timestamp 1683973020
transform 1 0 36864 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0946_
timestamp 1685175443
transform -1 0 39552 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0947_
timestamp 1683973020
transform -1 0 36864 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0948_
timestamp 1685175443
transform 1 0 36480 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0949_
timestamp 1683973020
transform -1 0 34272 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0950_
timestamp 1685175443
transform -1 0 32352 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0951_
timestamp 1683973020
transform -1 0 32064 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0952_
timestamp 1685175443
transform -1 0 30432 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0953_
timestamp 1683973020
transform -1 0 29760 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0954_
timestamp 1685175443
transform 1 0 27168 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0955_
timestamp 1683973020
transform -1 0 26304 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0956_
timestamp 1685175443
transform -1 0 25440 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0957_
timestamp 1683973020
transform 1 0 25152 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0958_
timestamp 1685175443
transform 1 0 34464 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0959_
timestamp 1683973020
transform 1 0 34944 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0960_
timestamp 1685175443
transform 1 0 35904 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0961_
timestamp 1683973020
transform -1 0 36576 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0962_
timestamp 1685175443
transform 1 0 34944 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0963_
timestamp 1683973020
transform 1 0 35424 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0964_
timestamp 1685175443
transform 1 0 31488 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0965_
timestamp 1683973020
transform -1 0 32448 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0966_
timestamp 1685175443
transform -1 0 31488 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0967_
timestamp 1683973020
transform -1 0 29184 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0968_
timestamp 1685175443
transform 1 0 25632 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0969_
timestamp 1683973020
transform 1 0 25920 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0970_
timestamp 1685175443
transform -1 0 24192 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0971_
timestamp 1683973020
transform -1 0 23328 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0972_
timestamp 1685175443
transform 1 0 21504 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0973_
timestamp 1683973020
transform 1 0 21984 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0974_
timestamp 1685175443
transform 1 0 16512 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0975_
timestamp 1683973020
transform 1 0 16992 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0976_
timestamp 1685175443
transform -1 0 11328 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0977_
timestamp 1683973020
transform -1 0 11520 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0978_
timestamp 1685175443
transform -1 0 9312 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0979_
timestamp 1683973020
transform -1 0 7008 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0980_
timestamp 1685175443
transform -1 0 4896 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0981_
timestamp 1683973020
transform -1 0 3648 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0982_
timestamp 1685175443
transform -1 0 5184 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0983_
timestamp 1683973020
transform 1 0 3744 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0984_
timestamp 1685175443
transform 1 0 17760 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0985_
timestamp 1683973020
transform 1 0 18432 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0986_
timestamp 1685175443
transform -1 0 20256 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0987_
timestamp 1683973020
transform -1 0 18912 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0988_
timestamp 1685175443
transform -1 0 17088 0 -1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0989_
timestamp 1683973020
transform -1 0 15744 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0990_
timestamp 1685175443
transform -1 0 10272 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0991_
timestamp 1683973020
transform 1 0 11520 0 -1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0992_
timestamp 1685175443
transform -1 0 9792 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0993_
timestamp 1683973020
transform -1 0 8448 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0994_
timestamp 1685175443
transform 1 0 6240 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0995_
timestamp 1683973020
transform 1 0 6720 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0996_
timestamp 1685175443
transform -1 0 5184 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0997_
timestamp 1683973020
transform 1 0 4224 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__0998_
timestamp 1685175443
transform 1 0 12480 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__0999_
timestamp 1683973020
transform -1 0 11136 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1000_
timestamp 1685175443
transform 1 0 15264 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1001_
timestamp 1683973020
transform 1 0 15744 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1002_
timestamp 1685175443
transform -1 0 16992 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1003_
timestamp 1683973020
transform -1 0 15264 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1004_
timestamp 1685175443
transform -1 0 12288 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1005_
timestamp 1683973020
transform -1 0 10848 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1006_
timestamp 1685175443
transform -1 0 9984 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1007_
timestamp 1683973020
transform -1 0 7680 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1008_
timestamp 1685175443
transform -1 0 5376 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1009_
timestamp 1683973020
transform -1 0 3360 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1010_
timestamp 1685175443
transform -1 0 5472 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1011_
timestamp 1683973020
transform -1 0 4992 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1012_
timestamp 1685175443
transform -1 0 6624 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1013_
timestamp 1683973020
transform 1 0 6048 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1014_
timestamp 1685175443
transform 1 0 12480 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1015_
timestamp 1683973020
transform 1 0 13920 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1016_
timestamp 1685175443
transform -1 0 14880 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1017_
timestamp 1683973020
transform -1 0 13920 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1018_
timestamp 1685175443
transform -1 0 11808 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1019_
timestamp 1683973020
transform -1 0 11232 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1020_
timestamp 1685175443
transform -1 0 8352 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1021_
timestamp 1683973020
transform 1 0 7104 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1022_
timestamp 1685175443
transform 1 0 3648 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1023_
timestamp 1683973020
transform 1 0 5568 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1024_
timestamp 1685175443
transform -1 0 4512 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1025_
timestamp 1683973020
transform -1 0 4224 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1026_
timestamp 1685175443
transform 1 0 4896 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1027_
timestamp 1683973020
transform 1 0 5664 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1028_
timestamp 1685175443
transform 1 0 6720 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1029_
timestamp 1683973020
transform -1 0 8256 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1030_
timestamp 1685175443
transform 1 0 7968 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1031_
timestamp 1683973020
transform 1 0 8448 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1032_
timestamp 1685175443
transform -1 0 19488 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1033_
timestamp 1683973020
transform -1 0 16896 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1034_
timestamp 1685175443
transform -1 0 19200 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1035_
timestamp 1683973020
transform 1 0 17280 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1036_
timestamp 1685175443
transform -1 0 18432 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1037_
timestamp 1683973020
transform -1 0 17952 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1038_
timestamp 1685175443
transform -1 0 16320 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1039_
timestamp 1683973020
transform -1 0 14208 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1040_
timestamp 1685175443
transform 1 0 10464 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1041_
timestamp 1683973020
transform 1 0 11808 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1042_
timestamp 1685175443
transform -1 0 10656 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1043_
timestamp 1683973020
transform 1 0 9216 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1044_
timestamp 1685175443
transform 1 0 9696 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1045_
timestamp 1683973020
transform 1 0 12384 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1046_
timestamp 1685175443
transform -1 0 20064 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1047_
timestamp 1683973020
transform 1 0 19488 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1048_
timestamp 1685175443
transform 1 0 18528 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1049_
timestamp 1683973020
transform 1 0 19008 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1050_
timestamp 1685175443
transform 1 0 17376 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1051_
timestamp 1683973020
transform 1 0 17856 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1052_
timestamp 1685175443
transform -1 0 17856 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1053_
timestamp 1683973020
transform -1 0 17184 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1054_
timestamp 1685175443
transform -1 0 15840 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1055_
timestamp 1683973020
transform -1 0 14976 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1056_
timestamp 1685175443
transform -1 0 11424 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1057_
timestamp 1683973020
transform 1 0 11328 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1058_
timestamp 1685175443
transform -1 0 9984 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1059_
timestamp 1683973020
transform -1 0 9216 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1060_
timestamp 1685175443
transform -1 0 10272 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1061_
timestamp 1683973020
transform -1 0 6336 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1062_
timestamp 1685175443
transform -1 0 4224 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1063_
timestamp 1683973020
transform 1 0 1824 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1064_
timestamp 1685175443
transform 1 0 2304 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1065_
timestamp 1683973020
transform 1 0 4512 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1066_
timestamp 1685175443
transform -1 0 5952 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1067_
timestamp 1683973020
transform 1 0 4992 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1068_
timestamp 1685175443
transform 1 0 6336 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1069_
timestamp 1683973020
transform -1 0 6528 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1070_
timestamp 1685175443
transform -1 0 11712 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1071_
timestamp 1683973020
transform -1 0 10752 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1072_
timestamp 1685175443
transform -1 0 10272 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1073_
timestamp 1683973020
transform -1 0 9120 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1074_
timestamp 1685175443
transform 1 0 6336 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1075_
timestamp 1683973020
transform 1 0 7680 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1076_
timestamp 1685175443
transform -1 0 4800 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1077_
timestamp 1683973020
transform -1 0 3744 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1078_
timestamp 1685175443
transform -1 0 4704 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1079_
timestamp 1683973020
transform 1 0 3936 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1080_
timestamp 1685175443
transform -1 0 5088 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1081_
timestamp 1683973020
transform 1 0 4704 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_mem__1082_
timestamp 1685175443
transform 1 0 5952 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1083_
timestamp 1683973020
transform 1 0 6432 0 1 18900
box -48 -56 528 834
use sg13g2_nand2b_2  u_ppwm_u_mem__1084_
timestamp 1685211885
transform 1 0 6912 0 1 17388
box -48 -56 816 834
use sg13g2_nand2_2  u_ppwm_u_mem__1085_
timestamp 1685180049
transform -1 0 6048 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_mem__1086_
timestamp 1676627187
transform -1 0 5184 0 -1 20412
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1087_
timestamp 1676901763
transform -1 0 3648 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1088_
timestamp 1676639442
transform 1 0 2688 0 -1 18900
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1089_
timestamp 1676627187
transform -1 0 5856 0 1 20412
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1090_
timestamp 1676901763
transform -1 0 4224 0 -1 20412
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1091_
timestamp 1676639442
transform 1 0 1920 0 1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1092_
timestamp 1683973020
transform 1 0 5472 0 1 18900
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_mem__1093_
timestamp 1676985977
transform -1 0 6336 0 1 17388
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_mem__1094_
timestamp 1676639442
transform -1 0 5472 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1095_
timestamp 1676627187
transform 1 0 1056 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_mem__1096_
timestamp 1676901763
transform -1 0 4416 0 -1 14364
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_mem__1097_
timestamp 1676639442
transform -1 0 1920 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1098_
timestamp 1676627187
transform -1 0 9216 0 1 14364
box -48 -56 432 834
use sg13g2_and3_1  u_ppwm_u_mem__1099_
timestamp 1676971669
transform -1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_nor3_1  u_ppwm_u_mem__1100_
timestamp 1676639442
transform 1 0 5472 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_mem__1101_
timestamp 1676627187
transform 1 0 3744 0 -1 15876
box -48 -56 432 834
use sg13g2_and4_1  u_ppwm_u_mem__1102_
timestamp 1676985977
transform 1 0 4992 0 1 14364
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_mem__1103_
timestamp 1676639442
transform 1 0 5088 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1104_
timestamp 1683973020
transform 1 0 6912 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_mem__1105_
timestamp 1683973020
transform -1 0 7872 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_mem__1106_
timestamp 1685181386
transform -1 0 8736 0 1 15876
box -54 -56 528 834
use sg13g2_tiehi  u_ppwm_u_mem__1107__174
timestamp 1680000651
transform -1 0 36384 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1107_
timestamp 1746535128
transform 1 0 35520 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1108__146
timestamp 1680000651
transform 1 0 48768 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1108_
timestamp 1746535128
transform -1 0 50400 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1109__144
timestamp 1680000651
transform 1 0 49344 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1109_
timestamp 1746535128
transform 1 0 49248 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1110_
timestamp 1746535128
transform 1 0 47808 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1110__142
timestamp 1680000651
transform -1 0 49536 0 1 27972
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1111__140
timestamp 1680000651
transform -1 0 45408 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1111_
timestamp 1746535128
transform 1 0 44064 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1112_
timestamp 1746535128
transform 1 0 40224 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1112__138
timestamp 1680000651
transform 1 0 40032 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1113_
timestamp 1746535128
transform -1 0 43008 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1113__136
timestamp 1680000651
transform 1 0 41472 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1114_
timestamp 1746535128
transform 1 0 37824 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1114__134
timestamp 1680000651
transform -1 0 39456 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1115_
timestamp 1746535184
transform -1 0 46848 0 -1 18900
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1115__132
timestamp 1680000651
transform 1 0 44832 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1116__130
timestamp 1680000651
transform -1 0 50016 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1116_
timestamp 1746535128
transform 1 0 49152 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1117__128
timestamp 1680000651
transform -1 0 51744 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1117_
timestamp 1746535128
transform 1 0 49248 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1118_
timestamp 1746535128
transform 1 0 44928 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1118__126
timestamp 1680000651
transform -1 0 45888 0 1 27972
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1119__124
timestamp 1680000651
transform 1 0 43392 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1119_
timestamp 1746535128
transform -1 0 44448 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1120__122
timestamp 1680000651
transform 1 0 40224 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1120_
timestamp 1746535128
transform 1 0 40608 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1121__120
timestamp 1680000651
transform 1 0 39840 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1121_
timestamp 1746535128
transform 1 0 40416 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1122__118
timestamp 1680000651
transform 1 0 47328 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1122_
timestamp 1746535128
transform 1 0 47712 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1123__116
timestamp 1680000651
transform 1 0 50592 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1123_
timestamp 1746535128
transform -1 0 51936 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1124__114
timestamp 1680000651
transform -1 0 46944 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1124_
timestamp 1746535128
transform 1 0 45792 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1125_
timestamp 1746535128
transform 1 0 41376 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1125__112
timestamp 1680000651
transform -1 0 42240 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1126_
timestamp 1746535128
transform 1 0 39456 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1126__110
timestamp 1680000651
transform -1 0 40320 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1127_
timestamp 1746535128
transform 1 0 37248 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1127__108
timestamp 1680000651
transform -1 0 38112 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1128_
timestamp 1746535128
transform -1 0 44736 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1128__106
timestamp 1680000651
transform 1 0 42624 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1129_
timestamp 1746535128
transform -1 0 47712 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1129__104
timestamp 1680000651
transform 1 0 46464 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1130__102
timestamp 1680000651
transform -1 0 45216 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1130_
timestamp 1746535128
transform 1 0 44352 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1131__100
timestamp 1680000651
transform -1 0 44736 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1131_
timestamp 1746535128
transform 1 0 43968 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1132_
timestamp 1746535128
transform 1 0 40320 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1132__98
timestamp 1680000651
transform 1 0 40224 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1133_
timestamp 1746535128
transform 1 0 36864 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1133__96
timestamp 1680000651
transform -1 0 38016 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1134_
timestamp 1746535128
transform 1 0 34848 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1134__94
timestamp 1680000651
transform 1 0 34464 0 -1 23436
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1135__92
timestamp 1680000651
transform 1 0 31872 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1135_
timestamp 1746535128
transform 1 0 32736 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1136_
timestamp 1746535128
transform 1 0 32928 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1136__90
timestamp 1680000651
transform 1 0 32448 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1137__88
timestamp 1680000651
transform 1 0 32640 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1137_
timestamp 1746535128
transform 1 0 34080 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1138_
timestamp 1746535128
transform 1 0 31776 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1138__86
timestamp 1680000651
transform -1 0 33696 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1139_
timestamp 1746535128
transform 1 0 27360 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1139__84
timestamp 1680000651
transform -1 0 28608 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1140__82
timestamp 1680000651
transform 1 0 24480 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1140_
timestamp 1746535128
transform 1 0 24384 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1141_
timestamp 1746535128
transform 1 0 23520 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1141__80
timestamp 1680000651
transform 1 0 23136 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1142_
timestamp 1746535128
transform -1 0 31680 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1142__78
timestamp 1680000651
transform 1 0 29568 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1143__76
timestamp 1680000651
transform 1 0 30528 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1143_
timestamp 1746535128
transform 1 0 31008 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1144__74
timestamp 1680000651
transform -1 0 33120 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1144_
timestamp 1746535128
transform 1 0 31776 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1145__72
timestamp 1680000651
transform -1 0 29184 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1145_
timestamp 1746535128
transform 1 0 27744 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1146_
timestamp 1746535128
transform 1 0 21312 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1146__70
timestamp 1680000651
transform 1 0 21408 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1147_
timestamp 1746535128
transform 1 0 22464 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1147__68
timestamp 1680000651
transform -1 0 23808 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1148_
timestamp 1746535128
transform 1 0 29376 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1148__66
timestamp 1680000651
transform 1 0 28992 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1149__64
timestamp 1680000651
transform 1 0 37824 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1149_
timestamp 1746535128
transform -1 0 39936 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1150_
timestamp 1746535128
transform 1 0 38304 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1150__62
timestamp 1680000651
transform -1 0 39552 0 -1 32508
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1151__60
timestamp 1680000651
transform 1 0 35232 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1151_
timestamp 1746535128
transform 1 0 35328 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1152_
timestamp 1746535128
transform 1 0 32448 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1152__58
timestamp 1680000651
transform -1 0 33312 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1153_
timestamp 1746535128
transform 1 0 28704 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1153__56
timestamp 1680000651
transform 1 0 28320 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1154_
timestamp 1746535128
transform 1 0 26112 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1154__173
timestamp 1680000651
transform -1 0 28032 0 -1 32508
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1155__171
timestamp 1680000651
transform -1 0 24576 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1155_
timestamp 1746535128
transform 1 0 23712 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1156_
timestamp 1746535184
transform -1 0 37056 0 -1 29484
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1156__169
timestamp 1680000651
transform 1 0 35904 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1157_
timestamp 1746535128
transform 1 0 37440 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1157__167
timestamp 1680000651
transform -1 0 38304 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1158__165
timestamp 1680000651
transform 1 0 33984 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1158_
timestamp 1746535128
transform 1 0 34656 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1159__163
timestamp 1680000651
transform -1 0 33024 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1159_
timestamp 1746535128
transform 1 0 32160 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1160_
timestamp 1746535128
transform 1 0 29184 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1160__161
timestamp 1680000651
transform 1 0 29088 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1161__159
timestamp 1680000651
transform -1 0 26976 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1161_
timestamp 1746535128
transform 1 0 25728 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1162_
timestamp 1746535128
transform 1 0 23328 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1162__157
timestamp 1680000651
transform -1 0 25152 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1163_
timestamp 1746535128
transform 1 0 21312 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1163__155
timestamp 1680000651
transform -1 0 22272 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1164__153
timestamp 1680000651
transform -1 0 19488 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1164_
timestamp 1746535128
transform 1 0 18336 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1165_
timestamp 1746535128
transform 1 0 11904 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1165__151
timestamp 1680000651
transform -1 0 12960 0 -1 37044
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1166__149
timestamp 1680000651
transform 1 0 6720 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1166_
timestamp 1746535128
transform 1 0 7104 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1167__147
timestamp 1680000651
transform -1 0 4608 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1167_
timestamp 1746535128
transform 1 0 3840 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1168__143
timestamp 1680000651
transform -1 0 1920 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1168_
timestamp 1746535128
transform 1 0 1056 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1169_
timestamp 1746535184
transform -1 0 21024 0 -1 32508
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1169__139
timestamp 1680000651
transform 1 0 19392 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1170_
timestamp 1746535128
transform 1 0 18912 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1170__135
timestamp 1680000651
transform 1 0 18048 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1171__131
timestamp 1680000651
transform -1 0 17472 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1171_
timestamp 1746535128
transform 1 0 15552 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1172__127
timestamp 1680000651
transform 1 0 12000 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1172_
timestamp 1746535128
transform -1 0 12960 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1173_
timestamp 1746535128
transform 1 0 7392 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1173__123
timestamp 1680000651
transform -1 0 8352 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1174_
timestamp 1746535128
transform 1 0 4128 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1174__119
timestamp 1680000651
transform -1 0 4992 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1175_
timestamp 1746535128
transform 1 0 1440 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1175__115
timestamp 1680000651
transform 1 0 1056 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1176_
timestamp 1746535128
transform -1 0 10080 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1176__111
timestamp 1680000651
transform 1 0 6624 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1177_
timestamp 1746535128
transform -1 0 19008 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1177__107
timestamp 1680000651
transform -1 0 18720 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1178_
timestamp 1746535128
transform 1 0 14496 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1178__103
timestamp 1680000651
transform 1 0 12960 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1179__99
timestamp 1680000651
transform 1 0 9600 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1179_
timestamp 1746535128
transform 1 0 11232 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1180__95
timestamp 1680000651
transform -1 0 8832 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1180_
timestamp 1746535128
transform 1 0 7680 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1181__91
timestamp 1680000651
transform -1 0 2304 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1181_
timestamp 1746535128
transform 1 0 1440 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1182_
timestamp 1746535128
transform 1 0 1248 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1182__87
timestamp 1680000651
transform -1 0 2112 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1183_
timestamp 1746535128
transform 1 0 4800 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1183__83
timestamp 1680000651
transform -1 0 5664 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1184_
timestamp 1746535128
transform -1 0 15936 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1184__79
timestamp 1680000651
transform 1 0 14784 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1185_
timestamp 1746535128
transform 1 0 13920 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1185__75
timestamp 1680000651
transform -1 0 15264 0 -1 32508
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1186__71
timestamp 1680000651
transform 1 0 9120 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1186_
timestamp 1746535128
transform 1 0 9888 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1187__67
timestamp 1680000651
transform 1 0 6432 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1187_
timestamp 1746535128
transform 1 0 6816 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1188_
timestamp 1746535128
transform 1 0 1152 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1188__63
timestamp 1680000651
transform 1 0 1056 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1189__59
timestamp 1680000651
transform 1 0 864 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1189_
timestamp 1746535128
transform 1 0 1248 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1190__55
timestamp 1680000651
transform -1 0 2016 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1190_
timestamp 1746535128
transform 1 0 1152 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1191__170
timestamp 1680000651
transform 1 0 7584 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1191_
timestamp 1746535128
transform -1 0 9792 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1192_
timestamp 1746535128
transform 1 0 8640 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1192__166
timestamp 1680000651
transform -1 0 10176 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1193__162
timestamp 1680000651
transform 1 0 17952 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1193_
timestamp 1746535128
transform 1 0 18048 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1194_
timestamp 1746535128
transform 1 0 15936 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1194__158
timestamp 1680000651
transform -1 0 16800 0 -1 27972
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1195__154
timestamp 1680000651
transform -1 0 19584 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1195_
timestamp 1746535128
transform 1 0 17952 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1196_
timestamp 1746535128
transform 1 0 14208 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1196__150
timestamp 1680000651
transform -1 0 15072 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1197_
timestamp 1746535128
transform -1 0 13344 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1197__145
timestamp 1680000651
transform 1 0 12192 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1198_
timestamp 1746535128
transform 1 0 8736 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1198__137
timestamp 1680000651
transform 1 0 8832 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1199_
timestamp 1746535128
transform -1 0 13056 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1199__129
timestamp 1680000651
transform 1 0 9792 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1200_
timestamp 1746535128
transform 1 0 19776 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1200__121
timestamp 1680000651
transform -1 0 21024 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1201_
timestamp 1746535128
transform -1 0 23040 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1201__113
timestamp 1680000651
transform 1 0 21216 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1202_
timestamp 1746535128
transform 1 0 18336 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1202__105
timestamp 1680000651
transform -1 0 19200 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1203__97
timestamp 1680000651
transform -1 0 17376 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1203_
timestamp 1746535128
transform 1 0 16512 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1204__89
timestamp 1680000651
transform 1 0 14016 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1204_
timestamp 1746535128
transform 1 0 13920 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1205__81
timestamp 1680000651
transform -1 0 13056 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1205_
timestamp 1746535128
transform 1 0 11808 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1206__73
timestamp 1680000651
transform -1 0 9600 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1206_
timestamp 1746535128
transform 1 0 8736 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1207_
timestamp 1746535128
transform 1 0 6816 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1207__65
timestamp 1680000651
transform -1 0 8448 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1208_
timestamp 1746535128
transform 1 0 960 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1208__57
timestamp 1680000651
transform 1 0 1248 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1209_
timestamp 1746535128
transform 1 0 1056 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1209__168
timestamp 1680000651
transform 1 0 1056 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1210_
timestamp 1746535128
transform 1 0 2016 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1210__160
timestamp 1680000651
transform 1 0 1248 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1211__152
timestamp 1680000651
transform 1 0 5664 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1211_
timestamp 1746535128
transform 1 0 6048 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1212_
timestamp 1746535128
transform 1 0 11616 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1212__141
timestamp 1680000651
transform -1 0 12960 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1213_
timestamp 1746535128
transform 1 0 9504 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1213__125
timestamp 1680000651
transform 1 0 9408 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1214_
timestamp 1746535128
transform -1 0 9216 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1214__109
timestamp 1680000651
transform 1 0 8160 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1215_
timestamp 1746535128
transform 1 0 1632 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1215__93
timestamp 1680000651
transform -1 0 2496 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1216_
timestamp 1746535128
transform 1 0 1344 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1216__77
timestamp 1680000651
transform 1 0 1440 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1217__61
timestamp 1680000651
transform 1 0 1632 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1217_
timestamp 1746535128
transform 1 0 1632 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1218__164
timestamp 1680000651
transform 1 0 5184 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1218_
timestamp 1746535128
transform 1 0 5568 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1219__148
timestamp 1680000651
transform -1 0 2688 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1219_
timestamp 1746535128
transform 1 0 1824 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1220_
timestamp 1746535128
transform 1 0 1152 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1220__117
timestamp 1680000651
transform -1 0 2016 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1221__85
timestamp 1680000651
transform 1 0 768 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1221_
timestamp 1746535128
transform 1 0 1248 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1222__172
timestamp 1680000651
transform -1 0 2016 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1222_
timestamp 1746535184
transform 1 0 1056 0 -1 15876
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1223__133
timestamp 1680000651
transform 1 0 5088 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1223_
timestamp 1746535184
transform 1 0 5760 0 1 14364
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1224__69
timestamp 1680000651
transform 1 0 672 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1224_
timestamp 1746535128
transform 1 0 2304 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1225_
timestamp 1746535128
transform 1 0 7872 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1225__175
timestamp 1680000651
transform -1 0 8832 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_mem__1226_
timestamp 1746535128
transform 1 0 8640 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_mem__1226__176
timestamp 1680000651
transform 1 0 8256 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_mem__1227__156
timestamp 1680000651
transform -1 0 11136 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1227_
timestamp 1746535184
transform 1 0 9312 0 -1 17388
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_mem__1228__101
timestamp 1680000651
transform -1 0 12864 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_mem__1228_
timestamp 1746535184
transform 1 0 12000 0 1 17388
box -48 -56 2736 834
use sg13g2_inv_1  u_ppwm_u_pwm__125_
timestamp 1676382929
transform 1 0 9312 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__126_
timestamp 1676382929
transform -1 0 12096 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__127_
timestamp 1676382929
transform -1 0 9888 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__128_
timestamp 1676382929
transform -1 0 8064 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__129_
timestamp 1676382929
transform 1 0 7008 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__130_
timestamp 1676382929
transform 1 0 9984 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_pwm__131_
timestamp 1676382947
transform -1 0 13920 0 1 3780
box -48 -56 432 834
use sg13g2_inv_1  u_ppwm_u_pwm__132_
timestamp 1676382929
transform 1 0 13248 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__133_
timestamp 1676382929
transform 1 0 10656 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__134_
timestamp 1676382929
transform 1 0 12480 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  u_ppwm_u_pwm__135_
timestamp 1676382929
transform -1 0 13152 0 1 11340
box -48 -56 336 834
use sg13g2_inv_2  u_ppwm_u_pwm__136_
timestamp 1676382947
transform 1 0 4128 0 -1 9828
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_pwm__137_
timestamp 1676643125
transform -1 0 8640 0 1 9828
box -48 -56 624 834
use sg13g2_nor2_1  u_ppwm_u_pwm__138_
timestamp 1676627187
transform 1 0 8544 0 -1 6804
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_pwm__139_
timestamp 1676643125
transform 1 0 7392 0 -1 9828
box -48 -56 624 834
use sg13g2_nand3_1  u_ppwm_u_pwm__140_
timestamp 1683988354
transform 1 0 7584 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__141_
timestamp 1685175443
transform -1 0 14496 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__142_
timestamp 1683973020
transform -1 0 12288 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__143_
timestamp 1685175443
transform -1 0 12960 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__144_
timestamp 1683973020
transform -1 0 12768 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__145_
timestamp 1685175443
transform -1 0 11520 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__146_
timestamp 1683973020
transform -1 0 10272 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__147_
timestamp 1685175443
transform -1 0 12000 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__148_
timestamp 1683973020
transform 1 0 11904 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__149_
timestamp 1685175443
transform -1 0 12192 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__150_
timestamp 1683973020
transform 1 0 13056 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__151_
timestamp 1685175443
transform -1 0 10752 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__152_
timestamp 1683973020
transform -1 0 10272 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__153_
timestamp 1685175443
transform -1 0 11712 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__154_
timestamp 1683973020
transform 1 0 7296 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__155_
timestamp 1685175443
transform -1 0 11232 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__156_
timestamp 1683973020
transform -1 0 8352 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__157_
timestamp 1685175443
transform -1 0 12288 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__158_
timestamp 1683973020
transform -1 0 10368 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__159_
timestamp 1685175443
transform -1 0 10848 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__160_
timestamp 1683973020
transform 1 0 11328 0 1 8316
box -48 -56 528 834
use sg13g2_and2_1  u_ppwm_u_pwm__161_
timestamp 1676901763
transform -1 0 6816 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__162_
timestamp 1685175443
transform -1 0 5952 0 1 12852
box -48 -56 538 834
use sg13g2_nor2_1  u_ppwm_u_pwm__163_
timestamp 1676627187
transform 1 0 3168 0 -1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__164_
timestamp 1685175443
transform 1 0 3744 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__165_
timestamp 1683973020
transform 1 0 4128 0 1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__166_
timestamp 1683973020
transform -1 0 4128 0 1 11340
box -48 -56 528 834
use sg13g2_and4_1  u_ppwm_u_pwm__167_
timestamp 1676985977
transform -1 0 6240 0 -1 11340
box -48 -56 816 834
use sg13g2_nor3_1  u_ppwm_u_pwm__168_
timestamp 1676639442
transform 1 0 4512 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  u_ppwm_u_pwm__169_
timestamp 1676627187
transform -1 0 4032 0 1 8316
box -48 -56 432 834
use sg13g2_and2_1  u_ppwm_u_pwm__170_
timestamp 1676901763
transform -1 0 3840 0 -1 11340
box -48 -56 528 834
use sg13g2_nor3_1  u_ppwm_u_pwm__171_
timestamp 1676639442
transform -1 0 2976 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_pwm__172_
timestamp 1677516600
transform -1 0 2784 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_pwm__173_
timestamp 1676627187
transform 1 0 1632 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__174_
timestamp 1683973020
transform -1 0 1728 0 -1 8316
box -48 -56 528 834
use sg13g2_and3_2  u_ppwm_u_pwm__175_
timestamp 1683976310
transform 1 0 3456 0 1 6804
box -48 -56 720 834
use sg13g2_nor3_1  u_ppwm_u_pwm__176_
timestamp 1676639442
transform 1 0 768 0 -1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  u_ppwm_u_pwm__177_
timestamp 1677516600
transform -1 0 3264 0 -1 6804
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_pwm__178_
timestamp 1676627187
transform 1 0 2112 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__179_
timestamp 1683973020
transform -1 0 4992 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3_1  u_ppwm_u_pwm__180_
timestamp 1683988354
transform 1 0 3840 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__181_
timestamp 1676557249
transform 1 0 4992 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_pwm__182_
timestamp 1676627187
transform 1 0 3456 0 1 5292
box -48 -56 432 834
use sg13g2_or2_1  u_ppwm_u_pwm__183_
timestamp 1684236171
transform 1 0 4512 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__184_
timestamp 1676557249
transform 1 0 5760 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__185_
timestamp 1683973020
transform -1 0 5856 0 -1 6804
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_pwm__186_
timestamp 1685201930
transform 1 0 7776 0 -1 8316
box -48 -56 624 834
use sg13g2_xor2_1  u_ppwm_u_pwm__187_
timestamp 1677577977
transform 1 0 4992 0 -1 8316
box -48 -56 816 834
use sg13g2_nor2_1  u_ppwm_u_pwm__188_
timestamp 1676627187
transform -1 0 6240 0 -1 9828
box -48 -56 432 834
use sg13g2_nand3_1  u_ppwm_u_pwm__189_
timestamp 1683988354
transform -1 0 10176 0 -1 9828
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_pwm__190_
timestamp 1685201930
transform 1 0 9120 0 -1 9828
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_pwm__191_
timestamp 1676639442
transform 1 0 6912 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__192_
timestamp 1685181386
transform 1 0 8544 0 -1 11340
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__193_
timestamp 1685181386
transform 1 0 7872 0 1 11340
box -54 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__194_
timestamp 1685181386
transform -1 0 9984 0 1 9828
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__195_
timestamp 1676567195
transform 1 0 9024 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__196_
timestamp 1685175443
transform 1 0 9792 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__197_
timestamp 1685181386
transform 1 0 8352 0 1 11340
box -54 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__198_
timestamp 1676567195
transform 1 0 8832 0 1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__199_
timestamp 1676567195
transform 1 0 8448 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__200_
timestamp 1683973020
transform 1 0 9312 0 1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__201_
timestamp 1685181386
transform 1 0 8064 0 -1 11340
box -54 -56 528 834
use sg13g2_or4_1  u_ppwm_u_pwm__202_
timestamp 1677154604
transform -1 0 9792 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__203_
timestamp 1685175443
transform -1 0 8064 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__204_
timestamp 1676567195
transform -1 0 7584 0 1 5292
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__205_
timestamp 1676567195
transform 1 0 7584 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__206_
timestamp 1676557249
transform 1 0 7008 0 -1 6804
box -48 -56 432 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__207_
timestamp 1676567195
transform 1 0 7392 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  u_ppwm_u_pwm__208_
timestamp 1676567195
transform 1 0 7584 0 1 5292
box -48 -56 528 834
use sg13g2_nand4_1  u_ppwm_u_pwm__209_
timestamp 1685201930
transform 1 0 8064 0 1 5292
box -48 -56 624 834
use sg13g2_nor2b_1  u_ppwm_u_pwm__210_
timestamp 1685181386
transform 1 0 9312 0 1 3780
box -54 -56 528 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__211_
timestamp 1683973020
transform 1 0 9792 0 -1 5292
box -48 -56 528 834
use sg13g2_a21o_1  u_ppwm_u_pwm__212_
timestamp 1677175127
transform 1 0 9120 0 -1 5292
box -48 -56 720 834
use sg13g2_nor2_1  u_ppwm_u_pwm__213_
timestamp 1676627187
transform 1 0 10272 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_pwm__214_
timestamp 1676627187
transform 1 0 9600 0 1 5292
box -48 -56 432 834
use sg13g2_nor4_1  u_ppwm_u_pwm__215_
timestamp 1676643125
transform 1 0 8544 0 -1 5292
box -48 -56 624 834
use sg13g2_nor3_1  u_ppwm_u_pwm__216_
timestamp 1676639442
transform 1 0 8640 0 -1 3780
box -48 -56 528 834
use sg13g2_a221oi_1  u_ppwm_u_pwm__217_
timestamp 1685197497
transform 1 0 8832 0 1 5292
box -48 -56 816 834
use sg13g2_nand2_1  u_ppwm_u_pwm__218_
timestamp 1676557249
transform -1 0 9312 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_pwm__219_
timestamp 1676627187
transform 1 0 8544 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  u_ppwm_u_pwm__220_
timestamp 1683973020
transform 1 0 9312 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  u_ppwm_u_pwm__221_
timestamp 1676557249
transform -1 0 9312 0 1 6804
box -48 -56 432 834
use sg13g2_nor2_1  u_ppwm_u_pwm__222_
timestamp 1676627187
transform 1 0 8160 0 -1 6804
box -48 -56 432 834
use sg13g2_nand2_1  u_ppwm_u_pwm__223_
timestamp 1676557249
transform -1 0 9984 0 1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__224_
timestamp 1685175443
transform 1 0 9408 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  u_ppwm_u_pwm__225_
timestamp 1685175443
transform 1 0 10368 0 1 8316
box -48 -56 538 834
use sg13g2_or3_1  u_ppwm_u_pwm__226_
timestamp 1677141922
transform 1 0 9888 0 -1 8316
box -48 -56 720 834
use sg13g2_and3_1  u_ppwm_u_pwm__227_
timestamp 1676971669
transform 1 0 10560 0 -1 8316
box -48 -56 720 834
use sg13g2_tiehi  u_ppwm_u_pwm__228__190
timestamp 1680000651
transform -1 0 15264 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__228_
timestamp 1746535128
transform -1 0 15456 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__229__187
timestamp 1680000651
transform 1 0 9600 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__229_
timestamp 1746535128
transform -1 0 12288 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__230__185
timestamp 1680000651
transform 1 0 8544 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__230_
timestamp 1746535128
transform -1 0 10656 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__231_
timestamp 1746535128
transform -1 0 13824 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__231__183
timestamp 1680000651
transform 1 0 11136 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__232__181
timestamp 1680000651
transform -1 0 13056 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__232_
timestamp 1746535128
transform 1 0 11616 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__233__179
timestamp 1680000651
transform 1 0 8928 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__233_
timestamp 1746535128
transform -1 0 10752 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__234__177
timestamp 1680000651
transform -1 0 5088 0 -1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__234_
timestamp 1746535128
transform 1 0 4224 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__235_
timestamp 1746535128
transform 1 0 5280 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__235__197
timestamp 1680000651
transform -1 0 6144 0 1 2268
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__236__195
timestamp 1680000651
transform 1 0 9984 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__236_
timestamp 1746535128
transform 1 0 10368 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__237__193
timestamp 1680000651
transform 1 0 9984 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__237_
timestamp 1746535128
transform 1 0 10176 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__238__191
timestamp 1680000651
transform 1 0 3552 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__238_
timestamp 1746535184
transform 1 0 5568 0 -1 12852
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__239__189
timestamp 1680000651
transform -1 0 3744 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__239_
timestamp 1746535184
transform 1 0 2880 0 -1 12852
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__240_
timestamp 1746535184
transform 1 0 4992 0 1 9828
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__240__186
timestamp 1680000651
transform 1 0 3840 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__241_
timestamp 1746535184
transform 1 0 1440 0 1 9828
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__241__182
timestamp 1680000651
transform -1 0 2304 0 -1 11340
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__242__178
timestamp 1680000651
transform 1 0 1248 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__242_
timestamp 1746535184
transform 1 0 960 0 1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__243_
timestamp 1746535184
transform 1 0 768 0 1 6804
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__243__196
timestamp 1680000651
transform -1 0 1632 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__244_
timestamp 1746535184
transform 1 0 1632 0 -1 5292
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__244__192
timestamp 1680000651
transform -1 0 2592 0 1 5292
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__245__188
timestamp 1680000651
transform -1 0 5760 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__245_
timestamp 1746535184
transform 1 0 4320 0 1 5292
box -48 -56 2736 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__246_
timestamp 1746535128
transform 1 0 5856 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__246__180
timestamp 1680000651
transform 1 0 6144 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  u_ppwm_u_pwm__247__194
timestamp 1680000651
transform 1 0 3744 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_2  u_ppwm_u_pwm__247_
timestamp 1746535184
transform 1 0 4032 0 1 8316
box -48 -56 2736 834
use sg13g2_tiehi  u_ppwm_u_pwm__248__184
timestamp 1680000651
transform -1 0 12384 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__248_
timestamp 1746535128
transform 1 0 11136 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  u_ppwm_u_pwm__249__198
timestamp 1680000651
transform -1 0 12480 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  u_ppwm_u_pwm__249_
timestamp 1746535128
transform 1 0 11616 0 -1 8316
box -48 -56 2640 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel via3 78 36708 78 36708 0 clk
rlabel metal2 38016 18942 38016 18942 0 clknet_0_clk
rlabel metal3 7488 9156 7488 9156 0 clknet_4_0_0_clk
rlabel metal3 45600 11004 45600 11004 0 clknet_4_10_0_clk
rlabel metal3 44352 20748 44352 20748 0 clknet_4_11_0_clk
rlabel metal2 29280 24990 29280 24990 0 clknet_4_12_0_clk
rlabel metal2 30432 29106 30432 29106 0 clknet_4_13_0_clk
rlabel metal2 45504 29064 45504 29064 0 clknet_4_14_0_clk
rlabel metal2 37968 32172 37968 32172 0 clknet_4_15_0_clk
rlabel metal3 6864 17052 6864 17052 0 clknet_4_1_0_clk
rlabel metal2 14016 7896 14016 7896 0 clknet_4_2_0_clk
rlabel metal3 14352 14952 14352 14952 0 clknet_4_3_0_clk
rlabel metal2 6720 27552 6720 27552 0 clknet_4_4_0_clk
rlabel metal2 5760 32088 5760 32088 0 clknet_4_5_0_clk
rlabel metal2 15936 28308 15936 28308 0 clknet_4_6_0_clk
rlabel metal2 17568 32256 17568 32256 0 clknet_4_7_0_clk
rlabel metal2 38208 7896 38208 7896 0 clknet_4_8_0_clk
rlabel metal2 37824 19026 37824 19026 0 clknet_4_9_0_clk
rlabel metal2 2304 7896 2304 7896 0 clknet_5_0__leaf_clk
rlabel metal2 5328 32340 5328 32340 0 clknet_5_10__leaf_clk
rlabel metal2 8160 32760 8160 32760 0 clknet_5_11__leaf_clk
rlabel metal2 14544 29820 14544 29820 0 clknet_5_12__leaf_clk
rlabel metal2 19344 29820 19344 29820 0 clknet_5_13__leaf_clk
rlabel metal2 12720 32928 12720 32928 0 clknet_5_14__leaf_clk
rlabel metal2 19536 32172 19536 32172 0 clknet_5_15__leaf_clk
rlabel metal3 28512 1932 28512 1932 0 clknet_5_16__leaf_clk
rlabel metal2 39648 4032 39648 4032 0 clknet_5_17__leaf_clk
rlabel metal3 34800 18564 34800 18564 0 clknet_5_18__leaf_clk
rlabel metal3 39456 17052 39456 17052 0 clknet_5_19__leaf_clk
rlabel metal3 8016 3444 8016 3444 0 clknet_5_1__leaf_clk
rlabel metal2 40512 15456 40512 15456 0 clknet_5_20__leaf_clk
rlabel metal3 46032 11172 46032 11172 0 clknet_5_21__leaf_clk
rlabel metal3 41904 18564 41904 18564 0 clknet_5_22__leaf_clk
rlabel metal2 45504 19320 45504 19320 0 clknet_5_23__leaf_clk
rlabel metal2 30624 29820 30624 29820 0 clknet_5_24__leaf_clk
rlabel metal2 17856 21924 17856 21924 0 clknet_5_25__leaf_clk
rlabel metal3 29280 28308 29280 28308 0 clknet_5_26__leaf_clk
rlabel metal2 33792 34020 33792 34020 0 clknet_5_27__leaf_clk
rlabel metal3 46224 29148 46224 29148 0 clknet_5_28__leaf_clk
rlabel metal2 50496 22680 50496 22680 0 clknet_5_29__leaf_clk
rlabel metal3 5376 14700 5376 14700 0 clknet_5_2__leaf_clk
rlabel metal3 35424 29148 35424 29148 0 clknet_5_30__leaf_clk
rlabel metal2 38784 33264 38784 33264 0 clknet_5_31__leaf_clk
rlabel metal3 7152 20076 7152 20076 0 clknet_5_3__leaf_clk
rlabel metal2 15648 7056 15648 7056 0 clknet_5_4__leaf_clk
rlabel metal3 15936 4116 15936 4116 0 clknet_5_5__leaf_clk
rlabel metal2 14112 13104 14112 13104 0 clknet_5_6__leaf_clk
rlabel metal2 13104 19236 13104 19236 0 clknet_5_7__leaf_clk
rlabel metal2 2400 23856 2400 23856 0 clknet_5_8__leaf_clk
rlabel metal2 7872 25704 7872 25704 0 clknet_5_9__leaf_clk
rlabel metal2 6144 17304 6144 17304 0 net1
rlabel metal3 366 21588 366 21588 0 net10
rlabel metal2 44448 30156 44448 30156 0 net100
rlabel metal2 12528 17724 12528 17724 0 net101
rlabel metal2 44880 23940 44880 23940 0 net102
rlabel metal3 14112 35028 14112 35028 0 net103
rlabel metal2 46752 20748 46752 20748 0 net104
rlabel metal2 18912 23940 18912 23940 0 net105
rlabel metal3 43584 19404 43584 19404 0 net106
rlabel metal2 18480 31500 18480 31500 0 net107
rlabel metal2 37728 22596 37728 22596 0 net108
rlabel metal2 8592 25956 8592 25956 0 net109
rlabel metal3 366 8988 366 8988 0 net11
rlabel metal2 40032 27300 40032 27300 0 net110
rlabel metal3 8208 31500 8208 31500 0 net111
rlabel metal2 41952 31080 41952 31080 0 net112
rlabel metal3 22032 25956 22032 25956 0 net113
rlabel metal3 46464 29988 46464 29988 0 net114
rlabel metal2 1488 31500 1488 31500 0 net115
rlabel metal2 51168 23940 51168 23940 0 net116
rlabel metal2 1728 18060 1728 18060 0 net117
rlabel metal2 47616 22764 47616 22764 0 net118
rlabel metal2 4752 36540 4752 36540 0 net119
rlabel metal3 366 9828 366 9828 0 net12
rlabel metal3 40512 21420 40512 21420 0 net120
rlabel metal2 20736 29484 20736 29484 0 net121
rlabel metal2 40560 23940 40560 23940 0 net122
rlabel metal2 8064 37926 8064 37926 0 net123
rlabel metal2 43680 24276 43680 24276 0 net124
rlabel metal2 9744 23940 9744 23940 0 net125
rlabel metal2 45552 28476 45552 28476 0 net126
rlabel metal2 12288 37926 12288 37926 0 net127
rlabel metal2 51456 26376 51456 26376 0 net128
rlabel metal2 12576 28098 12576 28098 0 net129
rlabel metal3 366 10668 366 10668 0 net13
rlabel metal2 49680 21420 49680 21420 0 net130
rlabel metal3 16608 36540 16608 36540 0 net131
rlabel metal2 46368 18984 46368 18984 0 net132
rlabel metal3 5808 13356 5808 13356 0 net133
rlabel metal2 39168 19152 39168 19152 0 net134
rlabel metal3 18336 34482 18336 34482 0 net135
rlabel metal2 42000 17892 42000 17892 0 net136
rlabel metal2 9120 26544 9120 26544 0 net137
rlabel metal2 40320 25914 40320 25914 0 net138
rlabel metal2 20544 32592 20544 32592 0 net139
rlabel metal3 366 11508 366 11508 0 net14
rlabel metal2 45024 25452 45024 25452 0 net140
rlabel metal3 12384 21420 12384 21420 0 net141
rlabel metal3 48768 28476 48768 28476 0 net142
rlabel metal2 1632 32886 1632 32886 0 net143
rlabel metal2 49632 24276 49632 24276 0 net144
rlabel metal2 12480 25410 12480 25410 0 net145
rlabel metal3 49488 21420 49488 21420 0 net146
rlabel metal2 4320 36204 4320 36204 0 net147
rlabel metal2 2352 19908 2352 19908 0 net148
rlabel metal3 7296 36540 7296 36540 0 net149
rlabel metal3 366 12348 366 12348 0 net15
rlabel metal2 14736 24444 14736 24444 0 net150
rlabel metal2 12624 36540 12624 36540 0 net151
rlabel metal2 5952 22008 5952 22008 0 net152
rlabel metal3 19008 36036 19008 36036 0 net153
rlabel metal2 19248 24444 19248 24444 0 net154
rlabel metal2 21984 34692 21984 34692 0 net155
rlabel metal2 9792 17724 9792 17724 0 net156
rlabel metal2 24864 34272 24864 34272 0 net157
rlabel metal2 16464 27468 16464 27468 0 net158
rlabel metal3 26448 35028 26448 35028 0 net159
rlabel metal3 366 13188 366 13188 0 net16
rlabel metal2 1968 22428 1968 22428 0 net160
rlabel metal2 29376 35070 29376 35070 0 net161
rlabel metal2 18192 31500 18192 31500 0 net162
rlabel metal2 32736 34692 32736 34692 0 net163
rlabel metal2 5472 19866 5472 19866 0 net164
rlabel metal2 34272 31836 34272 31836 0 net165
rlabel metal2 9888 29568 9888 29568 0 net166
rlabel metal2 37968 34524 37968 34524 0 net167
rlabel metal2 1536 23856 1536 23856 0 net168
rlabel metal2 36576 29820 36576 29820 0 net169
rlabel metal3 366 14028 366 14028 0 net17
rlabel metal2 7872 29484 7872 29484 0 net170
rlabel metal2 24288 31668 24288 31668 0 net171
rlabel metal2 1632 14868 1632 14868 0 net172
rlabel metal2 27744 32382 27744 32382 0 net173
rlabel metal2 36096 20034 36096 20034 0 net174
rlabel metal2 8544 15204 8544 15204 0 net175
rlabel metal3 8832 19404 8832 19404 0 net176
rlabel metal2 4800 3696 4800 3696 0 net177
rlabel metal2 1488 8652 1488 8652 0 net178
rlabel metal2 9216 4116 9216 4116 0 net179
rlabel metal3 558 14868 558 14868 0 net18
rlabel metal2 6432 7476 6432 7476 0 net180
rlabel metal2 12768 4284 12768 4284 0 net181
rlabel metal2 1920 10500 1920 10500 0 net182
rlabel metal3 12384 11592 12384 11592 0 net183
rlabel metal2 12096 16548 12096 16548 0 net184
rlabel metal3 9504 13860 9504 13860 0 net185
rlabel metal3 4800 10836 4800 10836 0 net186
rlabel metal2 11904 14448 11904 14448 0 net187
rlabel metal3 5136 5628 5136 5628 0 net188
rlabel metal2 3408 12516 3408 12516 0 net189
rlabel metal3 366 3108 366 3108 0 net19
rlabel metal2 14976 12516 14976 12516 0 net190
rlabel metal3 4992 13860 4992 13860 0 net191
rlabel metal2 2112 5376 2112 5376 0 net192
rlabel metal2 10272 10080 10272 10080 0 net193
rlabel metal2 4128 9324 4128 9324 0 net194
rlabel metal2 10272 7224 10272 7224 0 net195
rlabel metal2 1344 6720 1344 6720 0 net196
rlabel metal2 5856 3108 5856 3108 0 net197
rlabel metal2 12192 8400 12192 8400 0 net198
rlabel metal3 14304 11676 14304 11676 0 net199
rlabel metal2 14208 7728 14208 7728 0 net2
rlabel metal3 366 3948 366 3948 0 net20
rlabel metal3 14496 12600 14496 12600 0 net200
rlabel metal3 44448 8652 44448 8652 0 net201
rlabel metal2 46704 8652 46704 8652 0 net202
rlabel metal3 10224 12516 10224 12516 0 net203
rlabel metal2 10656 13104 10656 13104 0 net204
rlabel metal2 11424 26376 11424 26376 0 net205
rlabel metal3 12480 24696 12480 24696 0 net206
rlabel metal2 13824 4410 13824 4410 0 net207
rlabel metal2 11712 3612 11712 3612 0 net208
rlabel metal2 7056 2604 7056 2604 0 net209
rlabel metal3 366 4788 366 4788 0 net21
rlabel metal2 4320 4410 4320 4410 0 net210
rlabel metal2 8064 4116 8064 4116 0 net211
rlabel metal2 5376 3654 5376 3654 0 net212
rlabel metal2 18768 23604 18768 23604 0 net213
rlabel metal2 18528 23184 18528 23184 0 net214
rlabel metal2 12576 15414 12576 15414 0 net215
rlabel metal2 12336 14028 12336 14028 0 net216
rlabel metal3 16560 17052 16560 17052 0 net217
rlabel metal3 18912 17724 18912 17724 0 net218
rlabel metal2 16320 17430 16320 17430 0 net219
rlabel metal3 558 5628 558 5628 0 net22
rlabel metal2 32544 23730 32544 23730 0 net220
rlabel metal2 31680 22176 31680 22176 0 net221
rlabel metal2 4896 27762 4896 27762 0 net222
rlabel metal3 8352 25284 8352 25284 0 net223
rlabel metal3 9552 36456 9552 36456 0 net224
rlabel metal2 12000 36162 12000 36162 0 net225
rlabel metal3 26016 29232 26016 29232 0 net226
rlabel metal2 27456 30954 27456 30954 0 net227
rlabel metal2 9552 38220 9552 38220 0 net228
rlabel metal3 12144 37968 12144 37968 0 net229
rlabel metal3 366 6468 366 6468 0 net23
rlabel metal2 18720 28182 18720 28182 0 net230
rlabel metal2 18048 29736 18048 29736 0 net231
rlabel metal3 16560 24612 16560 24612 0 net232
rlabel metal2 18048 25578 18048 25578 0 net233
rlabel metal2 9792 34440 9792 34440 0 net234
rlabel metal2 11328 33978 11328 33978 0 net235
rlabel metal3 8880 32172 8880 32172 0 net236
rlabel metal2 9984 31458 9984 31458 0 net237
rlabel metal2 9792 6720 9792 6720 0 net238
rlabel metal2 10464 6762 10464 6762 0 net239
rlabel metal3 366 7308 366 7308 0 net24
rlabel metal2 25248 31290 25248 31290 0 net240
rlabel metal2 26400 32550 26400 32550 0 net241
rlabel metal2 47040 27132 47040 27132 0 net242
rlabel metal2 47904 27930 47904 27930 0 net243
rlabel metal3 5712 33852 5712 33852 0 net244
rlabel metal3 36336 32172 36336 32172 0 net245
rlabel metal2 37440 32760 37440 32760 0 net246
rlabel metal2 13920 9576 13920 9576 0 net247
rlabel metal3 15744 15540 15744 15540 0 net248
rlabel metal2 13632 32592 13632 32592 0 net249
rlabel metal3 366 8148 366 8148 0 net25
rlabel metal2 14064 32844 14064 32844 0 net250
rlabel metal2 18192 35280 18192 35280 0 net251
rlabel metal2 19008 33978 19008 33978 0 net252
rlabel metal2 4320 26124 4320 26124 0 net253
rlabel metal2 6912 24066 6912 24066 0 net254
rlabel metal2 14400 34650 14400 34650 0 net255
rlabel metal2 14880 33852 14880 33852 0 net256
rlabel metal2 14544 24612 14544 24612 0 net257
rlabel metal2 9264 22260 9264 22260 0 net258
rlabel metal2 8976 20160 8976 20160 0 net259
rlabel metal2 33792 2940 33792 2940 0 net26
rlabel metal2 9984 3444 9984 3444 0 net260
rlabel metal2 10656 2898 10656 2898 0 net261
rlabel metal2 43296 30324 43296 30324 0 net262
rlabel metal2 43968 29736 43968 29736 0 net263
rlabel metal3 6096 34944 6096 34944 0 net264
rlabel metal2 16416 32340 16416 32340 0 net265
rlabel metal3 17952 30744 17952 30744 0 net266
rlabel metal2 19968 33516 19968 33516 0 net267
rlabel metal2 20928 32550 20928 32550 0 net268
rlabel metal2 28896 32172 28896 32172 0 net269
rlabel metal3 19104 1764 19104 1764 0 net27
rlabel metal2 29280 33138 29280 33138 0 net270
rlabel metal2 28128 33474 28128 33474 0 net271
rlabel metal2 29376 34356 29376 34356 0 net272
rlabel metal2 22656 29484 22656 29484 0 net273
rlabel metal3 21648 30744 21648 30744 0 net274
rlabel metal3 41904 21588 41904 21588 0 net275
rlabel metal2 40848 23184 40848 23184 0 net276
rlabel metal3 42144 26124 42144 26124 0 net277
rlabel metal2 35232 33390 35232 33390 0 net278
rlabel metal2 35424 33978 35424 33978 0 net279
rlabel metal2 26064 1932 26064 1932 0 net28
rlabel metal2 47232 26544 47232 26544 0 net280
rlabel metal2 48960 26502 48960 26502 0 net281
rlabel metal2 44352 21000 44352 21000 0 net282
rlabel metal2 44640 20370 44640 20370 0 net283
rlabel metal2 39648 19194 39648 19194 0 net284
rlabel metal2 42912 18144 42912 18144 0 net285
rlabel metal2 23616 32928 23616 32928 0 net286
rlabel metal2 23424 34356 23424 34356 0 net287
rlabel metal2 34176 22344 34176 22344 0 net288
rlabel metal3 35328 23184 35328 23184 0 net289
rlabel metal2 23424 1596 23424 1596 0 net29
rlabel metal2 9696 25032 9696 25032 0 net290
rlabel metal2 9600 22554 9600 22554 0 net291
rlabel metal2 7104 35658 7104 35658 0 net292
rlabel metal2 40896 23730 40896 23730 0 net293
rlabel metal2 44352 24948 44352 24948 0 net294
rlabel metal4 4896 21798 4896 21798 0 net295
rlabel metal2 1536 23184 1536 23184 0 net296
rlabel metal2 5472 32424 5472 32424 0 net297
rlabel metal2 39648 19866 39648 19866 0 net298
rlabel metal2 12000 9324 12000 9324 0 net299
rlabel metal3 414 15708 414 15708 0 net3
rlabel metal2 33792 17052 33792 17052 0 net30
rlabel metal3 10608 9576 10608 9576 0 net300
rlabel metal3 12816 20076 12816 20076 0 net301
rlabel metal2 11904 19530 11904 19530 0 net302
rlabel metal2 14880 36960 14880 36960 0 net303
rlabel metal2 15696 35868 15696 35868 0 net304
rlabel metal3 18720 26796 18720 26796 0 net305
rlabel metal2 4608 32718 4608 32718 0 net306
rlabel metal2 13056 22218 13056 22218 0 net307
rlabel metal2 11616 20664 11616 20664 0 net308
rlabel metal2 34656 30492 34656 30492 0 net309
rlabel metal2 22224 4284 22224 4284 0 net31
rlabel metal3 39168 33432 39168 33432 0 net310
rlabel metal3 38688 30828 38688 30828 0 net311
rlabel metal2 14256 20244 14256 20244 0 net312
rlabel metal2 14016 22386 14016 22386 0 net313
rlabel metal2 25056 26922 25056 26922 0 net314
rlabel metal2 17568 36750 17568 36750 0 net315
rlabel metal3 18720 35280 18720 35280 0 net316
rlabel metal2 25632 34650 25632 34650 0 net317
rlabel metal2 2496 24906 2496 24906 0 net318
rlabel metal2 5472 34692 5472 34692 0 net319
rlabel metal2 15216 16884 15216 16884 0 net32
rlabel metal2 29760 28098 29760 28098 0 net320
rlabel metal2 31920 26796 31920 26796 0 net321
rlabel metal2 13344 31416 13344 31416 0 net322
rlabel metal2 15840 30114 15840 30114 0 net323
rlabel metal3 33504 29820 33504 29820 0 net324
rlabel metal2 34224 27720 34224 27720 0 net325
rlabel metal2 4128 27972 4128 27972 0 net326
rlabel metal3 2640 29232 2640 29232 0 net327
rlabel metal2 16512 22260 16512 22260 0 net328
rlabel metal2 35424 23814 35424 23814 0 net329
rlabel metal2 32352 3696 32352 3696 0 net33
rlabel metal3 32976 21672 32976 21672 0 net330
rlabel metal2 39600 23100 39600 23100 0 net331
rlabel metal2 39600 27720 39600 27720 0 net332
rlabel metal2 8592 20076 8592 20076 0 net333
rlabel metal2 8640 17640 8640 17640 0 net334
rlabel metal2 27744 29400 27744 29400 0 net335
rlabel metal2 40416 26712 40416 26712 0 net336
rlabel metal3 32736 24612 32736 24612 0 net337
rlabel metal2 31248 23184 31248 23184 0 net338
rlabel metal2 20832 25284 20832 25284 0 net339
rlabel metal2 37728 16716 37728 16716 0 net34
rlabel metal3 22032 26292 22032 26292 0 net340
rlabel metal2 49152 25200 49152 25200 0 net341
rlabel metal2 49296 24696 49296 24696 0 net342
rlabel metal2 7584 22302 7584 22302 0 net343
rlabel metal2 6096 21672 6096 21672 0 net344
rlabel metal2 6480 30072 6480 30072 0 net345
rlabel metal2 1344 30114 1344 30114 0 net346
rlabel metal2 39264 19992 39264 19992 0 net347
rlabel metal3 15936 31332 15936 31332 0 net348
rlabel metal2 19872 6426 19872 6426 0 net349
rlabel metal2 29952 20118 29952 20118 0 net35
rlabel metal2 29760 15456 29760 15456 0 net350
rlabel metal2 26400 17850 26400 17850 0 net351
rlabel metal2 16416 5082 16416 5082 0 net352
rlabel metal2 17280 4998 17280 4998 0 net353
rlabel metal2 26112 15708 26112 15708 0 net354
rlabel metal2 32544 7308 32544 7308 0 net355
rlabel metal2 19872 8568 19872 8568 0 net356
rlabel metal2 17904 4116 17904 4116 0 net357
rlabel metal3 23874 17724 23874 17724 0 net358
rlabel metal2 30528 13944 30528 13944 0 net359
rlabel metal2 29280 1596 29280 1596 0 net36
rlabel metal2 31968 14616 31968 14616 0 net360
rlabel metal2 24432 14700 24432 14700 0 net361
rlabel metal2 32256 7560 32256 7560 0 net362
rlabel metal2 24864 11844 24864 11844 0 net363
rlabel metal2 25008 13860 25008 13860 0 net364
rlabel metal2 25632 12936 25632 12936 0 net365
rlabel metal2 26112 14238 26112 14238 0 net366
rlabel metal2 26976 12600 26976 12600 0 net367
rlabel metal2 21600 12936 21600 12936 0 net368
rlabel metal2 18720 15918 18720 15918 0 net369
rlabel metal2 39504 13188 39504 13188 0 net37
rlabel metal3 21024 15204 21024 15204 0 net370
rlabel metal2 19488 3444 19488 3444 0 net371
rlabel metal2 20064 4578 20064 4578 0 net372
rlabel metal2 29280 3906 29280 3906 0 net373
rlabel metal2 19968 5796 19968 5796 0 net374
rlabel metal3 22416 13944 22416 13944 0 net375
rlabel metal2 28800 18144 28800 18144 0 net376
rlabel metal2 22656 12768 22656 12768 0 net377
rlabel metal3 17280 11004 17280 11004 0 net378
rlabel metal2 24768 17136 24768 17136 0 net379
rlabel metal2 34992 18564 34992 18564 0 net38
rlabel metal3 22848 20076 22848 20076 0 net380
rlabel metal3 23472 16212 23472 16212 0 net381
rlabel metal2 23712 15204 23712 15204 0 net382
rlabel metal2 23856 15456 23856 15456 0 net383
rlabel metal2 17088 9660 17088 9660 0 net384
rlabel metal2 19104 9702 19104 9702 0 net385
rlabel metal2 26496 13524 26496 13524 0 net386
rlabel metal2 28656 18732 28656 18732 0 net387
rlabel metal2 21984 17766 21984 17766 0 net388
rlabel metal2 11520 4200 11520 4200 0 net389
rlabel metal2 39744 15792 39744 15792 0 net39
rlabel metal3 12000 8652 12000 8652 0 net390
rlabel metal2 11616 4872 11616 4872 0 net391
rlabel metal2 37968 5376 37968 5376 0 net392
rlabel metal2 28080 27636 28080 27636 0 net393
rlabel metal2 15264 25242 15264 25242 0 net394
rlabel metal3 16032 26796 16032 26796 0 net395
rlabel metal2 20064 26670 20064 26670 0 net396
rlabel metal2 47520 25368 47520 25368 0 net397
rlabel metal2 41568 13188 41568 13188 0 net398
rlabel via1 40896 14530 40896 14530 0 net399
rlabel metal3 366 16548 366 16548 0 net4
rlabel metal2 16176 4032 16176 4032 0 net40
rlabel metal3 4224 20076 4224 20076 0 net400
rlabel metal2 6096 20580 6096 20580 0 net401
rlabel metal2 11616 19782 11616 19782 0 net402
rlabel metal2 2400 24360 2400 24360 0 net403
rlabel metal2 7104 26544 7104 26544 0 net404
rlabel metal2 12096 25494 12096 25494 0 net405
rlabel metal2 11664 21588 11664 21588 0 net406
rlabel metal3 13392 23772 13392 23772 0 net407
rlabel metal3 16704 22932 16704 22932 0 net408
rlabel metal2 5280 34462 5280 34462 0 net409
rlabel metal2 35808 16716 35808 16716 0 net41
rlabel metal2 3744 32970 3744 32970 0 net410
rlabel metal2 12192 29862 12192 29862 0 net411
rlabel metal3 10560 35196 10560 35196 0 net412
rlabel metal2 11760 38220 11760 38220 0 net413
rlabel metal2 11712 32886 11712 32886 0 net414
rlabel metal2 17472 32004 17472 32004 0 net415
rlabel metal2 15408 35196 15408 35196 0 net416
rlabel metal3 19392 29022 19392 29022 0 net417
rlabel metal2 20064 29988 20064 29988 0 net418
rlabel metal2 24096 33264 24096 33264 0 net419
rlabel metal2 32976 19236 32976 19236 0 net42
rlabel metal3 18624 34314 18624 34314 0 net420
rlabel metal2 22752 31416 22752 31416 0 net421
rlabel metal2 13056 30660 13056 30660 0 net422
rlabel metal2 39936 19068 39936 19068 0 net423
rlabel metal2 41280 19950 41280 19950 0 net424
rlabel metal2 33120 21252 33120 21252 0 net425
rlabel metal2 31584 28392 31584 28392 0 net426
rlabel metal2 32928 30114 32928 30114 0 net427
rlabel metal2 31392 33600 31392 33600 0 net428
rlabel metal2 34848 32172 34848 32172 0 net429
rlabel metal2 15216 15540 15216 15540 0 net43
rlabel metal2 36288 32928 36288 32928 0 net430
rlabel metal3 34368 32172 34368 32172 0 net431
rlabel metal2 39360 25830 39360 25830 0 net432
rlabel metal2 49056 26418 49056 26418 0 net433
rlabel metal3 47616 23856 47616 23856 0 net434
rlabel metal2 48768 23856 48768 23856 0 net435
rlabel metal2 40800 29904 40800 29904 0 net436
rlabel metal2 47424 28392 47424 28392 0 net437
rlabel metal2 34272 24360 34272 24360 0 net438
rlabel metal2 38448 5544 38448 5544 0 net439
rlabel metal2 31968 2226 31968 2226 0 net44
rlabel metal2 32160 13020 32160 13020 0 net440
rlabel metal2 46368 10500 46368 10500 0 net441
rlabel metal2 46464 8736 46464 8736 0 net442
rlabel metal2 40416 12054 40416 12054 0 net443
rlabel metal2 41088 14448 41088 14448 0 net444
rlabel metal2 40992 14322 40992 14322 0 net445
rlabel metal2 21600 17850 21600 17850 0 net446
rlabel metal2 19008 20412 19008 20412 0 net447
rlabel metal3 18144 10080 18144 10080 0 net448
rlabel metal2 34080 8190 34080 8190 0 net449
rlabel metal2 14448 11004 14448 11004 0 net45
rlabel metal2 28128 16926 28128 16926 0 net450
rlabel metal2 28704 18018 28704 18018 0 net451
rlabel metal2 35808 13272 35808 13272 0 net452
rlabel metal2 28800 19110 28800 19110 0 net453
rlabel metal2 17856 8106 17856 8106 0 net454
rlabel metal2 19728 5628 19728 5628 0 net455
rlabel metal2 15840 3444 15840 3444 0 net456
rlabel metal2 27936 7516 27936 7516 0 net457
rlabel metal3 17808 3444 17808 3444 0 net458
rlabel metal2 31872 8106 31872 8106 0 net459
rlabel metal2 14064 10332 14064 10332 0 net46
rlabel metal2 16416 3948 16416 3948 0 net460
rlabel metal2 32640 6636 32640 6636 0 net461
rlabel metal2 27552 13902 27552 13902 0 net462
rlabel metal2 26592 11634 26592 11634 0 net463
rlabel metal2 38208 12558 38208 12558 0 net464
rlabel metal2 39744 14784 39744 14784 0 net465
rlabel metal2 27840 15498 27840 15498 0 net466
rlabel metal2 18336 24864 18336 24864 0 net467
rlabel metal2 21408 20538 21408 20538 0 net468
rlabel metal2 21984 20034 21984 20034 0 net469
rlabel metal2 20352 22344 20352 22344 0 net47
rlabel metal2 17040 26124 17040 26124 0 net470
rlabel metal2 12768 25547 12768 25547 0 net471
rlabel metal2 16272 33621 16272 33621 0 net472
rlabel metal2 26016 19992 26016 19992 0 net473
rlabel metal2 29904 26628 29904 26628 0 net474
rlabel metal2 31680 20832 31680 20832 0 net475
rlabel metal2 13536 25452 13536 25452 0 net476
rlabel metal2 13344 27552 13344 27552 0 net477
rlabel metal2 15552 30618 15552 30618 0 net478
rlabel metal3 13680 30660 13680 30660 0 net479
rlabel metal3 17184 19908 17184 19908 0 net48
rlabel metal2 16992 23688 16992 23688 0 net480
rlabel metal2 27120 29820 27120 29820 0 net481
rlabel metal2 35712 29862 35712 29862 0 net482
rlabel metal2 30816 24360 30816 24360 0 net483
rlabel via2 39072 24609 39072 24609 0 net484
rlabel metal2 39216 26796 39216 26796 0 net485
rlabel metal2 31296 29148 31296 29148 0 net486
rlabel metal2 28896 24234 28896 24234 0 net487
rlabel metal4 6432 16968 6432 16968 0 net488
rlabel metal2 5664 13062 5664 13062 0 net489
rlabel metal2 23376 23100 23376 23100 0 net49
rlabel metal3 12576 5628 12576 5628 0 net490
rlabel metal2 19200 5040 19200 5040 0 net491
rlabel metal2 18912 8358 18912 8358 0 net492
rlabel metal2 12000 15330 12000 15330 0 net493
rlabel metal3 5952 30660 5952 30660 0 net494
rlabel metal2 8256 29862 8256 29862 0 net495
rlabel metal2 11040 34482 11040 34482 0 net496
rlabel metal2 9696 35280 9696 35280 0 net497
rlabel metal2 16800 35952 16800 35952 0 net498
rlabel metal2 11520 31668 11520 31668 0 net499
rlabel metal3 366 17388 366 17388 0 net5
rlabel metal2 13824 5964 13824 5964 0 net50
rlabel metal2 11904 30240 11904 30240 0 net500
rlabel metal2 17568 22176 17568 22176 0 net501
rlabel metal2 26688 30576 26688 30576 0 net502
rlabel metal3 19488 30660 19488 30660 0 net503
rlabel metal2 15600 21000 15600 21000 0 net504
rlabel metal2 38736 4116 38736 4116 0 net505
rlabel metal3 34320 15540 34320 15540 0 net506
rlabel metal2 41088 8064 41088 8064 0 net507
rlabel metal2 41280 13230 41280 13230 0 net508
rlabel metal2 42624 16170 42624 16170 0 net509
rlabel metal2 26208 23520 26208 23520 0 net51
rlabel metal2 33120 29778 33120 29778 0 net510
rlabel metal2 36768 33558 36768 33558 0 net511
rlabel metal2 35232 30576 35232 30576 0 net512
rlabel metal2 38736 19236 38736 19236 0 net513
rlabel metal2 47232 21672 47232 21672 0 net514
rlabel metal2 41280 29736 41280 29736 0 net515
rlabel metal2 51168 25788 51168 25788 0 net516
rlabel metal3 46128 23856 46128 23856 0 net517
rlabel metal2 42960 17052 42960 17052 0 net518
rlabel metal2 10032 30744 10032 30744 0 net519
rlabel metal2 27264 22008 27264 22008 0 net52
rlabel metal2 20928 27636 20928 27636 0 net520
rlabel metal2 19776 28224 19776 28224 0 net521
rlabel metal2 40128 31290 40128 31290 0 net522
rlabel metal2 39840 30114 39840 30114 0 net523
rlabel metal2 45408 22218 45408 22218 0 net524
rlabel metal2 47616 20370 47616 20370 0 net525
rlabel metal3 11526 26796 11526 26796 0 net526
rlabel metal2 960 24654 960 24654 0 net527
rlabel metal2 5664 23394 5664 23394 0 net528
rlabel metal2 42144 27888 42144 27888 0 net529
rlabel metal2 14832 7140 14832 7140 0 net53
rlabel metal2 41664 30366 41664 30366 0 net530
rlabel metal2 21120 35616 21120 35616 0 net531
rlabel metal2 43968 25284 43968 25284 0 net532
rlabel metal2 13344 10500 13344 10500 0 net533
rlabel metal2 13728 11214 13728 11214 0 net534
rlabel metal2 6048 19572 6048 19572 0 net535
rlabel metal3 34080 33096 34080 33096 0 net536
rlabel metal2 5568 22470 5568 22470 0 net537
rlabel metal3 7392 28140 7392 28140 0 net538
rlabel metal2 9600 27720 9600 27720 0 net539
rlabel metal2 16656 18564 16656 18564 0 net54
rlabel metal2 3888 30828 3888 30828 0 net540
rlabel metal2 37584 31164 37584 31164 0 net541
rlabel metal2 33120 32424 33120 32424 0 net542
rlabel metal3 46368 29316 46368 29316 0 net543
rlabel metal2 49824 25578 49824 25578 0 net544
rlabel metal2 26496 24654 26496 24654 0 net545
rlabel metal2 5952 6258 5952 6258 0 net546
rlabel metal2 3552 6300 3552 6300 0 net547
rlabel metal2 4368 5628 4368 5628 0 net548
rlabel metal2 3840 12432 3840 12432 0 net549
rlabel metal2 1680 28476 1680 28476 0 net55
rlabel metal2 2976 12768 2976 12768 0 net550
rlabel metal2 45600 25578 45600 25578 0 net551
rlabel metal3 48096 24360 48096 24360 0 net552
rlabel metal2 30912 34314 30912 34314 0 net553
rlabel metal2 35472 26796 35472 26796 0 net554
rlabel metal2 33024 25578 33024 25578 0 net555
rlabel metal2 36096 30408 36096 30408 0 net556
rlabel metal2 29472 29694 29472 29694 0 net557
rlabel metal2 45600 30660 45600 30660 0 net558
rlabel metal2 30768 30408 30768 30408 0 net559
rlabel metal2 29184 33180 29184 33180 0 net56
rlabel metal2 41328 21756 41328 21756 0 net560
rlabel metal2 47328 23016 47328 23016 0 net561
rlabel metal3 45744 18564 45744 18564 0 net562
rlabel metal2 50496 26586 50496 26586 0 net563
rlabel metal2 46944 23352 46944 23352 0 net564
rlabel metal2 7584 15792 7584 15792 0 net565
rlabel metal3 7824 16212 7824 16212 0 net566
rlabel metal2 7968 16212 7968 16212 0 net567
rlabel metal2 14592 29190 14592 29190 0 net568
rlabel metal2 8736 29442 8736 29442 0 net569
rlabel metal2 1536 25620 1536 25620 0 net57
rlabel metal2 38592 23352 38592 23352 0 net570
rlabel metal2 5856 28350 5856 28350 0 net571
rlabel metal2 6336 10710 6336 10710 0 net572
rlabel metal3 5088 10668 5088 10668 0 net573
rlabel metal2 5088 9912 5088 9912 0 net574
rlabel metal2 42240 11214 42240 11214 0 net575
rlabel metal2 46944 11970 46944 11970 0 net576
rlabel metal2 49488 23772 49488 23772 0 net577
rlabel metal2 50304 21126 50304 21126 0 net578
rlabel metal2 6768 31332 6768 31332 0 net579
rlabel metal2 33024 33348 33024 33348 0 net58
rlabel metal2 2496 32592 2496 32592 0 net580
rlabel metal2 46320 28308 46320 28308 0 net581
rlabel metal2 14880 29232 14880 29232 0 net582
rlabel metal2 7488 29568 7488 29568 0 net583
rlabel metal3 5280 29232 5280 29232 0 net584
rlabel metal3 36288 4116 36288 4116 0 net585
rlabel metal2 39600 3444 39600 3444 0 net586
rlabel metal2 5184 14952 5184 14952 0 net587
rlabel metal2 5376 15624 5376 15624 0 net588
rlabel metal2 2400 14994 2400 14994 0 net589
rlabel metal3 1440 28980 1440 28980 0 net59
rlabel metal2 41664 7896 41664 7896 0 net590
rlabel metal2 44448 6720 44448 6720 0 net591
rlabel metal2 13152 32550 13152 32550 0 net592
rlabel metal3 8880 7728 8880 7728 0 net593
rlabel metal3 7680 9492 7680 9492 0 net594
rlabel metal2 10560 12642 10560 12642 0 net595
rlabel metal2 29280 29400 29280 29400 0 net596
rlabel metal2 38112 21630 38112 21630 0 net597
rlabel metal2 35616 21084 35616 21084 0 net598
rlabel metal2 41568 9240 41568 9240 0 net599
rlabel metal3 366 18228 366 18228 0 net6
rlabel metal2 35664 34524 35664 34524 0 net60
rlabel metal2 44064 12768 44064 12768 0 net600
rlabel metal3 3264 7728 3264 7728 0 net601
rlabel metal2 1056 8064 1056 8064 0 net602
rlabel metal2 864 7434 864 7434 0 net603
rlabel metal3 45264 5628 45264 5628 0 net604
rlabel metal3 46224 6468 46224 6468 0 net605
rlabel metal2 2496 16002 2496 16002 0 net606
rlabel metal3 2928 16212 2928 16212 0 net607
rlabel metal2 38304 8232 38304 8232 0 net608
rlabel metal2 37920 8568 37920 8568 0 net609
rlabel metal2 1920 21840 1920 21840 0 net61
rlabel metal2 41472 8022 41472 8022 0 net610
rlabel metal3 4800 17640 4800 17640 0 net611
rlabel metal2 5184 14280 5184 14280 0 net612
rlabel metal2 1440 16548 1440 16548 0 net613
rlabel metal2 16896 17640 16896 17640 0 net614
rlabel metal2 17472 18018 17472 18018 0 net615
rlabel metal2 17184 18816 17184 18816 0 net616
rlabel metal3 3840 18732 3840 18732 0 net617
rlabel metal2 7488 15960 7488 15960 0 net618
rlabel metal2 7104 18564 7104 18564 0 net619
rlabel metal2 39264 31920 39264 31920 0 net62
rlabel metal2 38208 5292 38208 5292 0 net620
rlabel metal2 38304 4116 38304 4116 0 net621
rlabel metal2 38592 5964 38592 5964 0 net622
rlabel metal2 39216 6468 39216 6468 0 net623
rlabel metal2 5952 18018 5952 18018 0 net624
rlabel metal2 9888 18102 9888 18102 0 net625
rlabel metal3 9312 17052 9312 17052 0 net626
rlabel metal2 42912 5964 42912 5964 0 net627
rlabel metal2 42336 7392 42336 7392 0 net628
rlabel metal2 44304 7980 44304 7980 0 net629
rlabel metal2 1344 34104 1344 34104 0 net63
rlabel metal2 44736 5964 44736 5964 0 net630
rlabel metal2 44352 9030 44352 9030 0 net631
rlabel metal2 47328 8610 47328 8610 0 net632
rlabel metal2 40032 10458 40032 10458 0 net633
rlabel metal2 38880 10122 38880 10122 0 net634
rlabel metal2 39072 9786 39072 9786 0 net635
rlabel metal3 3696 6468 3696 6468 0 net636
rlabel metal2 5472 6720 5472 6720 0 net637
rlabel metal2 5328 17976 5328 17976 0 net638
rlabel metal2 46656 10206 46656 10206 0 net639
rlabel metal2 39456 29400 39456 29400 0 net64
rlabel metal2 45120 11256 45120 11256 0 net640
rlabel metal2 43872 12894 43872 12894 0 net641
rlabel metal3 14448 16212 14448 16212 0 net642
rlabel metal3 17184 18732 17184 18732 0 net643
rlabel metal2 8640 7770 8640 7770 0 net644
rlabel metal3 28980 5754 28980 5754 0 net645
rlabel metal2 37824 5040 37824 5040 0 net646
rlabel metal3 6192 11676 6192 11676 0 net647
rlabel metal2 19296 10458 19296 10458 0 net648
rlabel metal2 20736 10248 20736 10248 0 net649
rlabel metal3 7728 24444 7728 24444 0 net65
rlabel metal3 16440 10920 16440 10920 0 net650
rlabel metal3 3984 10416 3984 10416 0 net651
rlabel metal2 2400 9156 2400 9156 0 net652
rlabel metal2 46944 13776 46944 13776 0 net653
rlabel metal2 36672 5586 36672 5586 0 net654
rlabel metal2 44304 10416 44304 10416 0 net655
rlabel metal2 40896 11382 40896 11382 0 net656
rlabel metal2 17856 6846 17856 6846 0 net657
rlabel metal2 14400 7434 14400 7434 0 net658
rlabel metal2 41472 8610 41472 8610 0 net659
rlabel metal2 29568 29988 29568 29988 0 net66
rlabel metal2 33552 17640 33552 17640 0 net660
rlabel metal2 35328 15540 35328 15540 0 net661
rlabel metal3 25536 3444 25536 3444 0 net662
rlabel metal2 19392 4872 19392 4872 0 net663
rlabel metal2 19488 2646 19488 2646 0 net664
rlabel metal2 43488 13314 43488 13314 0 net665
rlabel metal2 44928 9744 44928 9744 0 net666
rlabel metal2 32928 3864 32928 3864 0 net667
rlabel metal3 38304 17724 38304 17724 0 net668
rlabel metal2 25344 2898 25344 2898 0 net669
rlabel metal3 7008 33012 7008 33012 0 net67
rlabel metal2 21792 2898 21792 2898 0 net670
rlabel metal2 31440 2604 31440 2604 0 net671
rlabel metal3 16608 6468 16608 6468 0 net672
rlabel metal2 25776 23772 25776 23772 0 net673
rlabel metal2 22848 21588 22848 21588 0 net674
rlabel metal2 16464 10164 16464 10164 0 net675
rlabel metal2 35040 3864 35040 3864 0 net676
rlabel metal2 25920 2898 25920 2898 0 net677
rlabel metal2 36672 19236 36672 19236 0 net678
rlabel metal2 34464 18564 34464 18564 0 net679
rlabel metal2 23184 29820 23184 29820 0 net68
rlabel metal2 38832 13188 38832 13188 0 net680
rlabel metal2 36000 16506 36000 16506 0 net681
rlabel metal3 36432 3444 36432 3444 0 net682
rlabel metal2 21888 21798 21888 21798 0 net683
rlabel metal2 20064 21084 20064 21084 0 net684
rlabel metal2 19728 21756 19728 21756 0 net685
rlabel metal3 19248 19992 19248 19992 0 net686
rlabel metal2 41952 15792 41952 15792 0 net687
rlabel metal2 39168 16128 39168 16128 0 net688
rlabel metal2 29616 23772 29616 23772 0 net689
rlabel metal2 960 15540 960 15540 0 net69
rlabel metal2 30960 13020 30960 13020 0 net690
rlabel metal3 5232 17724 5232 17724 0 net691
rlabel metal2 31968 13188 31968 13188 0 net692
rlabel metal3 366 19068 366 19068 0 net7
rlabel metal2 21744 31500 21744 31500 0 net70
rlabel metal3 9888 32004 9888 32004 0 net71
rlabel metal2 28896 27678 28896 27678 0 net72
rlabel metal2 9264 19404 9264 19404 0 net73
rlabel metal3 32544 27468 32544 27468 0 net74
rlabel metal2 14976 32424 14976 32424 0 net75
rlabel metal2 30816 23478 30816 23478 0 net76
rlabel metal2 1824 23520 1824 23520 0 net77
rlabel metal3 30528 21420 30528 21420 0 net78
rlabel metal3 15264 30492 15264 30492 0 net79
rlabel metal3 366 19908 366 19908 0 net8
rlabel metal3 23712 26964 23712 26964 0 net80
rlabel metal3 12528 19908 12528 19908 0 net81
rlabel metal2 24768 28644 24768 28644 0 net82
rlabel metal2 5424 30492 5424 30492 0 net83
rlabel metal2 28320 31080 28320 31080 0 net84
rlabel metal2 1056 17472 1056 17472 0 net85
rlabel metal2 32256 29568 32256 29568 0 net86
rlabel metal2 1824 30156 1824 30156 0 net87
rlabel metal2 32928 28140 32928 28140 0 net88
rlabel metal2 14352 22932 14352 22932 0 net89
rlabel metal3 366 20748 366 20748 0 net9
rlabel metal2 32736 24948 32736 24948 0 net90
rlabel metal2 2016 34692 2016 34692 0 net91
rlabel metal3 32688 21420 32688 21420 0 net92
rlabel metal2 2208 26544 2208 26544 0 net93
rlabel metal3 35040 22932 35040 22932 0 net94
rlabel metal2 8544 35868 8544 35868 0 net95
rlabel metal2 37680 28476 37680 28476 0 net96
rlabel metal2 17088 21252 17088 21252 0 net97
rlabel metal2 40512 29778 40512 29778 0 net98
rlabel metal2 11712 33600 11712 33600 0 net99
rlabel metal3 174 37548 174 37548 0 rst_n
rlabel metal2 46656 14364 46656 14364 0 u_ppwm/global_counter\[0\]
rlabel metal2 48672 12390 48672 12390 0 u_ppwm/global_counter\[10\]
rlabel metal2 39264 12390 39264 12390 0 u_ppwm/global_counter\[11\]
rlabel metal3 40464 11004 40464 11004 0 u_ppwm/global_counter\[12\]
rlabel metal2 38208 9828 38208 9828 0 u_ppwm/global_counter\[13\]
rlabel metal2 38976 8148 38976 8148 0 u_ppwm/global_counter\[14\]
rlabel metal2 41280 6804 41280 6804 0 u_ppwm/global_counter\[15\]
rlabel metal2 39552 5754 39552 5754 0 u_ppwm/global_counter\[16\]
rlabel metal2 29856 7014 29856 7014 0 u_ppwm/global_counter\[17\]
rlabel metal2 40512 5544 40512 5544 0 u_ppwm/global_counter\[18\]
rlabel metal2 37296 4116 37296 4116 0 u_ppwm/global_counter\[19\]
rlabel metal2 44928 10878 44928 10878 0 u_ppwm/global_counter\[1\]
rlabel metal2 43536 10164 43536 10164 0 u_ppwm/global_counter\[2\]
rlabel metal2 45792 11760 45792 11760 0 u_ppwm/global_counter\[3\]
rlabel metal3 42144 6384 42144 6384 0 u_ppwm/global_counter\[4\]
rlabel metal3 42384 7980 42384 7980 0 u_ppwm/global_counter\[5\]
rlabel metal4 44736 6510 44736 6510 0 u_ppwm/global_counter\[6\]
rlabel metal2 45216 8610 45216 8610 0 u_ppwm/global_counter\[7\]
rlabel metal2 48912 9492 48912 9492 0 u_ppwm/global_counter\[8\]
rlabel metal2 47424 10710 47424 10710 0 u_ppwm/global_counter\[9\]
rlabel metal2 22656 19320 22656 19320 0 u_ppwm/instr\[0\]
rlabel metal2 20736 18606 20736 18606 0 u_ppwm/instr\[1\]
rlabel metal2 22224 19236 22224 19236 0 u_ppwm/instr\[2\]
rlabel metal2 30336 25578 30336 25578 0 u_ppwm/instr\[3\]
rlabel metal2 28560 20076 28560 20076 0 u_ppwm/instr\[4\]
rlabel metal3 21744 24612 21744 24612 0 u_ppwm/instr\[5\]
rlabel metal2 27552 18858 27552 18858 0 u_ppwm/instr\[6\]
rlabel metal2 11808 17430 11808 17430 0 u_ppwm/mem_write_done
rlabel metal2 29232 21756 29232 21756 0 u_ppwm/pc\[0\]
rlabel metal2 28224 23436 28224 23436 0 u_ppwm/pc\[1\]
rlabel metal2 26112 24696 26112 24696 0 u_ppwm/pc\[2\]
rlabel metal2 22368 22806 22368 22806 0 u_ppwm/pc\[3\]
rlabel metal3 13824 16380 13824 16380 0 u_ppwm/period_start
rlabel metal2 14976 14994 14976 14994 0 u_ppwm/polarity
rlabel metal2 37824 15120 37824 15120 0 u_ppwm/pwm_value\[0\]
rlabel metal2 41760 16212 41760 16212 0 u_ppwm/pwm_value\[1\]
rlabel metal2 41472 13062 41472 13062 0 u_ppwm/pwm_value\[2\]
rlabel metal2 32160 16254 32160 16254 0 u_ppwm/pwm_value\[3\]
rlabel metal3 34080 4368 34080 4368 0 u_ppwm/pwm_value\[4\]
rlabel metal2 24480 3150 24480 3150 0 u_ppwm/pwm_value\[5\]
rlabel metal2 25344 1470 25344 1470 0 u_ppwm/pwm_value\[6\]
rlabel metal2 15792 2604 15792 2604 0 u_ppwm/pwm_value\[7\]
rlabel metal3 16656 5880 16656 5880 0 u_ppwm/pwm_value\[8\]
rlabel metal3 16656 9660 16656 9660 0 u_ppwm/pwm_value\[9\]
rlabel metal2 17376 18102 17376 18102 0 u_ppwm/u_ex/_0000_
rlabel metal2 16992 17304 16992 17304 0 u_ppwm/u_ex/_0001_
rlabel metal2 18048 18732 18048 18732 0 u_ppwm/u_ex/_0002_
rlabel metal2 26592 21756 26592 21756 0 u_ppwm/u_ex/_0003_
rlabel metal2 25920 22428 25920 22428 0 u_ppwm/u_ex/_0004_
rlabel metal2 22656 22428 22656 22428 0 u_ppwm/u_ex/_0005_
rlabel metal2 19968 21168 19968 21168 0 u_ppwm/u_ex/_0006_
rlabel metal3 18432 10710 18432 10710 0 u_ppwm/u_ex/_0007_
rlabel metal2 15456 14868 15456 14868 0 u_ppwm/u_ex/_0008_
rlabel metal2 34512 14952 34512 14952 0 u_ppwm/u_ex/_0009_
rlabel metal2 38400 16296 38400 16296 0 u_ppwm/u_ex/_0010_
rlabel metal2 39072 13482 39072 13482 0 u_ppwm/u_ex/_0011_
rlabel metal2 30336 19530 30336 19530 0 u_ppwm/u_ex/_0012_
rlabel metal2 31872 4326 31872 4326 0 u_ppwm/u_ex/_0013_
rlabel metal3 22128 2100 22128 2100 0 u_ppwm/u_ex/_0014_
rlabel metal3 22752 2016 22752 2016 0 u_ppwm/u_ex/_0015_
rlabel metal2 19248 924 19248 924 0 u_ppwm/u_ex/_0016_
rlabel metal2 13440 5922 13440 5922 0 u_ppwm/u_ex/_0017_
rlabel metal2 17664 8946 17664 8946 0 u_ppwm/u_ex/_0018_
rlabel metal2 32544 19320 32544 19320 0 u_ppwm/u_ex/_0019_
rlabel metal2 34176 17304 34176 17304 0 u_ppwm/u_ex/_0020_
rlabel metal2 37056 16464 37056 16464 0 u_ppwm/u_ex/_0021_
rlabel metal2 33312 16968 33312 16968 0 u_ppwm/u_ex/_0022_
rlabel metal2 33312 2730 33312 2730 0 u_ppwm/u_ex/_0023_
rlabel metal2 31632 1932 31632 1932 0 u_ppwm/u_ex/_0024_
rlabel metal3 29088 2562 29088 2562 0 u_ppwm/u_ex/_0025_
rlabel metal2 25680 3948 25680 3948 0 u_ppwm/u_ex/_0026_
rlabel metal2 16608 4158 16608 4158 0 u_ppwm/u_ex/_0027_
rlabel metal2 17040 5880 17040 5880 0 u_ppwm/u_ex/_0028_
rlabel metal2 36192 11424 36192 11424 0 u_ppwm/u_ex/_0029_
rlabel metal2 32448 11592 32448 11592 0 u_ppwm/u_ex/_0030_
rlabel metal2 15360 14658 15360 14658 0 u_ppwm/u_ex/_0031_
rlabel metal3 18432 17304 18432 17304 0 u_ppwm/u_ex/_0032_
rlabel metal2 21888 17472 21888 17472 0 u_ppwm/u_ex/_0033_
rlabel metal2 29280 12180 29280 12180 0 u_ppwm/u_ex/_0034_
rlabel metal3 25584 12600 25584 12600 0 u_ppwm/u_ex/_0035_
rlabel metal3 16512 14700 16512 14700 0 u_ppwm/u_ex/_0036_
rlabel metal2 17376 16842 17376 16842 0 u_ppwm/u_ex/_0037_
rlabel metal2 24576 7938 24576 7938 0 u_ppwm/u_ex/_0038_
rlabel metal2 34848 5796 34848 5796 0 u_ppwm/u_ex/_0039_
rlabel metal2 37392 9660 37392 9660 0 u_ppwm/u_ex/_0040_
rlabel metal2 28896 8316 28896 8316 0 u_ppwm/u_ex/_0041_
rlabel metal2 31776 10248 31776 10248 0 u_ppwm/u_ex/_0042_
rlabel metal3 32544 11676 32544 11676 0 u_ppwm/u_ex/_0043_
rlabel metal2 34733 12516 34733 12516 0 u_ppwm/u_ex/_0044_
rlabel metal2 17184 20244 17184 20244 0 u_ppwm/u_ex/_0045_
rlabel metal2 23616 21113 23616 21113 0 u_ppwm/u_ex/_0046_
rlabel metal2 20832 18732 20832 18732 0 u_ppwm/u_ex/_0047_
rlabel metal2 22656 18795 22656 18795 0 u_ppwm/u_ex/_0048_
rlabel metal2 19008 17766 19008 17766 0 u_ppwm/u_ex/_0049_
rlabel metal2 19392 10290 19392 10290 0 u_ppwm/u_ex/_0050_
rlabel metal2 16416 16338 16416 16338 0 u_ppwm/u_ex/_0051_
rlabel metal2 19392 18270 19392 18270 0 u_ppwm/u_ex/_0052_
rlabel metal2 17568 17808 17568 17808 0 u_ppwm/u_ex/_0053_
rlabel metal2 17184 19656 17184 19656 0 u_ppwm/u_ex/_0054_
rlabel metal2 17568 16590 17568 16590 0 u_ppwm/u_ex/_0055_
rlabel metal2 16032 17178 16032 17178 0 u_ppwm/u_ex/_0056_
rlabel metal2 18432 17430 18432 17430 0 u_ppwm/u_ex/_0057_
rlabel metal3 22032 18564 22032 18564 0 u_ppwm/u_ex/_0058_
rlabel metal2 21120 18816 21120 18816 0 u_ppwm/u_ex/_0059_
rlabel metal3 21744 19068 21744 19068 0 u_ppwm/u_ex/_0060_
rlabel metal2 25536 18984 25536 18984 0 u_ppwm/u_ex/_0061_
rlabel metal2 26208 21126 26208 21126 0 u_ppwm/u_ex/_0062_
rlabel metal2 24288 20958 24288 20958 0 u_ppwm/u_ex/_0063_
rlabel metal2 26016 21504 26016 21504 0 u_ppwm/u_ex/_0064_
rlabel metal2 25632 19236 25632 19236 0 u_ppwm/u_ex/_0065_
rlabel metal3 25488 19488 25488 19488 0 u_ppwm/u_ex/_0066_
rlabel metal2 24576 20118 24576 20118 0 u_ppwm/u_ex/_0067_
rlabel metal2 25824 21000 25824 21000 0 u_ppwm/u_ex/_0068_
rlabel metal3 25488 21588 25488 21588 0 u_ppwm/u_ex/_0069_
rlabel metal2 24096 20832 24096 20832 0 u_ppwm/u_ex/_0070_
rlabel metal2 24192 21084 24192 21084 0 u_ppwm/u_ex/_0071_
rlabel metal2 23904 19614 23904 19614 0 u_ppwm/u_ex/_0072_
rlabel metal2 23520 19656 23520 19656 0 u_ppwm/u_ex/_0073_
rlabel metal2 23328 19404 23328 19404 0 u_ppwm/u_ex/_0074_
rlabel metal2 23328 20034 23328 20034 0 u_ppwm/u_ex/_0075_
rlabel metal2 23808 19614 23808 19614 0 u_ppwm/u_ex/_0076_
rlabel metal2 24096 19236 24096 19236 0 u_ppwm/u_ex/_0077_
rlabel metal2 22848 20916 22848 20916 0 u_ppwm/u_ex/_0078_
rlabel metal2 23232 19278 23232 19278 0 u_ppwm/u_ex/_0079_
rlabel metal2 21024 20580 21024 20580 0 u_ppwm/u_ex/_0080_
rlabel metal3 19776 19950 19776 19950 0 u_ppwm/u_ex/_0081_
rlabel metal2 21888 20706 21888 20706 0 u_ppwm/u_ex/_0082_
rlabel metal3 21456 20412 21456 20412 0 u_ppwm/u_ex/_0083_
rlabel metal3 20832 20076 20832 20076 0 u_ppwm/u_ex/_0084_
rlabel metal2 19536 19824 19536 19824 0 u_ppwm/u_ex/_0085_
rlabel metal2 21120 21588 21120 21588 0 u_ppwm/u_ex/_0086_
rlabel metal2 23904 9492 23904 9492 0 u_ppwm/u_ex/_0087_
rlabel metal3 30912 8652 30912 8652 0 u_ppwm/u_ex/_0088_
rlabel metal2 34368 12768 34368 12768 0 u_ppwm/u_ex/_0089_
rlabel metal2 34176 12768 34176 12768 0 u_ppwm/u_ex/_0090_
rlabel metal2 34080 12768 34080 12768 0 u_ppwm/u_ex/_0091_
rlabel metal2 33984 11970 33984 11970 0 u_ppwm/u_ex/_0092_
rlabel metal2 34464 11634 34464 11634 0 u_ppwm/u_ex/_0093_
rlabel metal3 34272 11508 34272 11508 0 u_ppwm/u_ex/_0094_
rlabel metal3 32976 10836 32976 10836 0 u_ppwm/u_ex/_0095_
rlabel metal3 33456 11508 33456 11508 0 u_ppwm/u_ex/_0096_
rlabel metal2 30624 8694 30624 8694 0 u_ppwm/u_ex/_0097_
rlabel metal2 30432 8652 30432 8652 0 u_ppwm/u_ex/_0098_
rlabel metal2 29664 8736 29664 8736 0 u_ppwm/u_ex/_0099_
rlabel metal3 29568 8736 29568 8736 0 u_ppwm/u_ex/_0100_
rlabel metal3 23856 8148 23856 8148 0 u_ppwm/u_ex/_0101_
rlabel metal3 24000 8652 24000 8652 0 u_ppwm/u_ex/_0102_
rlabel metal3 24384 9492 24384 9492 0 u_ppwm/u_ex/_0103_
rlabel metal3 23664 9240 23664 9240 0 u_ppwm/u_ex/_0104_
rlabel metal2 24768 8736 24768 8736 0 u_ppwm/u_ex/_0105_
rlabel metal4 30336 8652 30336 8652 0 u_ppwm/u_ex/_0106_
rlabel metal3 22560 9534 22560 9534 0 u_ppwm/u_ex/_0107_
rlabel metal2 23232 8694 23232 8694 0 u_ppwm/u_ex/_0108_
rlabel metal2 22176 9492 22176 9492 0 u_ppwm/u_ex/_0109_
rlabel metal2 27360 7602 27360 7602 0 u_ppwm/u_ex/_0110_
rlabel metal2 38208 11634 38208 11634 0 u_ppwm/u_ex/_0111_
rlabel metal2 37536 11088 37536 11088 0 u_ppwm/u_ex/_0112_
rlabel metal2 36384 10668 36384 10668 0 u_ppwm/u_ex/_0113_
rlabel metal2 37344 10290 37344 10290 0 u_ppwm/u_ex/_0114_
rlabel metal2 38496 11844 38496 11844 0 u_ppwm/u_ex/_0115_
rlabel metal2 37248 10458 37248 10458 0 u_ppwm/u_ex/_0116_
rlabel metal2 37152 10332 37152 10332 0 u_ppwm/u_ex/_0117_
rlabel metal2 36672 8484 36672 8484 0 u_ppwm/u_ex/_0118_
rlabel metal2 37248 8988 37248 8988 0 u_ppwm/u_ex/_0119_
rlabel metal2 35232 5544 35232 5544 0 u_ppwm/u_ex/_0120_
rlabel metal2 36384 7560 36384 7560 0 u_ppwm/u_ex/_0121_
rlabel metal2 36232 8064 36232 8064 0 u_ppwm/u_ex/_0122_
rlabel metal3 36480 7980 36480 7980 0 u_ppwm/u_ex/_0123_
rlabel metal2 36480 7896 36480 7896 0 u_ppwm/u_ex/_0124_
rlabel metal2 34080 6762 34080 6762 0 u_ppwm/u_ex/_0125_
rlabel metal3 36384 8106 36384 8106 0 u_ppwm/u_ex/_0126_
rlabel metal2 27696 7392 27696 7392 0 u_ppwm/u_ex/_0127_
rlabel metal3 26736 7980 26736 7980 0 u_ppwm/u_ex/_0128_
rlabel metal2 24672 8106 24672 8106 0 u_ppwm/u_ex/_0129_
rlabel metal3 25104 7980 25104 7980 0 u_ppwm/u_ex/_0130_
rlabel metal2 26016 7392 26016 7392 0 u_ppwm/u_ex/_0131_
rlabel via1 26013 7980 26013 7980 0 u_ppwm/u_ex/_0132_
rlabel metal2 25728 8106 25728 8106 0 u_ppwm/u_ex/_0133_
rlabel metal2 26208 7896 26208 7896 0 u_ppwm/u_ex/_0134_
rlabel metal3 25440 14700 25440 14700 0 u_ppwm/u_ex/_0135_
rlabel metal2 26496 14280 26496 14280 0 u_ppwm/u_ex/_0136_
rlabel metal2 26496 8232 26496 8232 0 u_ppwm/u_ex/_0137_
rlabel metal3 25344 9282 25344 9282 0 u_ppwm/u_ex/_0138_
rlabel metal3 35232 7224 35232 7224 0 u_ppwm/u_ex/_0139_
rlabel metal2 36336 14028 36336 14028 0 u_ppwm/u_ex/_0140_
rlabel metal2 36576 13944 36576 13944 0 u_ppwm/u_ex/_0141_
rlabel metal2 35712 11088 35712 11088 0 u_ppwm/u_ex/_0142_
rlabel metal2 35712 9702 35712 9702 0 u_ppwm/u_ex/_0143_
rlabel metal3 36432 14028 36432 14028 0 u_ppwm/u_ex/_0144_
rlabel metal2 36336 12516 36336 12516 0 u_ppwm/u_ex/_0145_
rlabel metal3 34992 10164 34992 10164 0 u_ppwm/u_ex/_0146_
rlabel metal2 35328 10122 35328 10122 0 u_ppwm/u_ex/_0147_
rlabel metal2 35520 9744 35520 9744 0 u_ppwm/u_ex/_0148_
rlabel metal2 35232 7392 35232 7392 0 u_ppwm/u_ex/_0149_
rlabel metal2 30144 7812 30144 7812 0 u_ppwm/u_ex/_0150_
rlabel metal2 30144 6678 30144 6678 0 u_ppwm/u_ex/_0151_
rlabel metal2 30624 7560 30624 7560 0 u_ppwm/u_ex/_0152_
rlabel metal2 29952 7812 29952 7812 0 u_ppwm/u_ex/_0153_
rlabel metal4 29856 7560 29856 7560 0 u_ppwm/u_ex/_0154_
rlabel metal3 23184 7980 23184 7980 0 u_ppwm/u_ex/_0155_
rlabel metal2 24000 7896 24000 7896 0 u_ppwm/u_ex/_0156_
rlabel metal2 25104 7392 25104 7392 0 u_ppwm/u_ex/_0157_
rlabel metal2 24101 7056 24101 7056 0 u_ppwm/u_ex/_0158_
rlabel metal2 24384 7686 24384 7686 0 u_ppwm/u_ex/_0159_
rlabel metal2 23904 7476 23904 7476 0 u_ppwm/u_ex/_0160_
rlabel metal2 24672 13146 24672 13146 0 u_ppwm/u_ex/_0161_
rlabel metal3 22944 7140 22944 7140 0 u_ppwm/u_ex/_0162_
rlabel metal2 21888 9240 21888 9240 0 u_ppwm/u_ex/_0163_
rlabel metal3 20736 17892 20736 17892 0 u_ppwm/u_ex/_0164_
rlabel metal2 34464 7812 34464 7812 0 u_ppwm/u_ex/_0165_
rlabel metal3 35472 13188 35472 13188 0 u_ppwm/u_ex/_0166_
rlabel metal2 35520 13146 35520 13146 0 u_ppwm/u_ex/_0167_
rlabel metal2 35424 12936 35424 12936 0 u_ppwm/u_ex/_0168_
rlabel metal3 35952 13020 35952 13020 0 u_ppwm/u_ex/_0169_
rlabel metal2 36096 10164 36096 10164 0 u_ppwm/u_ex/_0170_
rlabel metal2 35712 8988 35712 8988 0 u_ppwm/u_ex/_0171_
rlabel metal2 34848 9408 34848 9408 0 u_ppwm/u_ex/_0172_
rlabel metal3 34368 8736 34368 8736 0 u_ppwm/u_ex/_0173_
rlabel metal2 35040 9366 35040 9366 0 u_ppwm/u_ex/_0174_
rlabel metal2 35184 8484 35184 8484 0 u_ppwm/u_ex/_0175_
rlabel metal3 35424 8652 35424 8652 0 u_ppwm/u_ex/_0176_
rlabel metal3 34992 8484 34992 8484 0 u_ppwm/u_ex/_0177_
rlabel metal2 35136 7896 35136 7896 0 u_ppwm/u_ex/_0178_
rlabel metal2 34992 8148 34992 8148 0 u_ppwm/u_ex/_0179_
rlabel metal4 21408 9156 21408 9156 0 u_ppwm/u_ex/_0180_
rlabel metal2 21984 8862 21984 8862 0 u_ppwm/u_ex/_0181_
rlabel metal2 20064 8526 20064 8526 0 u_ppwm/u_ex/_0182_
rlabel metal2 19968 8736 19968 8736 0 u_ppwm/u_ex/_0183_
rlabel metal2 21696 8064 21696 8064 0 u_ppwm/u_ex/_0184_
rlabel metal2 21600 8274 21600 8274 0 u_ppwm/u_ex/_0185_
rlabel metal2 21312 8652 21312 8652 0 u_ppwm/u_ex/_0186_
rlabel metal3 23808 11676 23808 11676 0 u_ppwm/u_ex/_0187_
rlabel metal2 31968 8148 31968 8148 0 u_ppwm/u_ex/_0188_
rlabel metal3 20640 8652 20640 8652 0 u_ppwm/u_ex/_0189_
rlabel metal2 21744 8568 21744 8568 0 u_ppwm/u_ex/_0190_
rlabel metal2 37056 12474 37056 12474 0 u_ppwm/u_ex/_0191_
rlabel metal2 37200 12516 37200 12516 0 u_ppwm/u_ex/_0192_
rlabel metal2 32640 11508 32640 11508 0 u_ppwm/u_ex/_0193_
rlabel metal3 33072 11592 33072 11592 0 u_ppwm/u_ex/_0194_
rlabel metal2 38016 12600 38016 12600 0 u_ppwm/u_ex/_0195_
rlabel metal3 35184 11760 35184 11760 0 u_ppwm/u_ex/_0196_
rlabel metal3 32976 11004 32976 11004 0 u_ppwm/u_ex/_0197_
rlabel metal2 32256 10374 32256 10374 0 u_ppwm/u_ex/_0198_
rlabel metal3 32256 10248 32256 10248 0 u_ppwm/u_ex/_0199_
rlabel metal3 32016 10164 32016 10164 0 u_ppwm/u_ex/_0200_
rlabel metal2 32544 10248 32544 10248 0 u_ppwm/u_ex/_0201_
rlabel via2 32067 9492 32067 9492 0 u_ppwm/u_ex/_0202_
rlabel metal2 28512 9156 28512 9156 0 u_ppwm/u_ex/_0203_
rlabel metal2 28416 9744 28416 9744 0 u_ppwm/u_ex/_0204_
rlabel metal2 28320 9366 28320 9366 0 u_ppwm/u_ex/_0205_
rlabel metal2 26976 9450 26976 9450 0 u_ppwm/u_ex/_0206_
rlabel metal3 27888 8652 27888 8652 0 u_ppwm/u_ex/_0207_
rlabel metal2 27264 9240 27264 9240 0 u_ppwm/u_ex/_0208_
rlabel metal2 27072 9912 27072 9912 0 u_ppwm/u_ex/_0209_
rlabel metal2 24672 9450 24672 9450 0 u_ppwm/u_ex/_0210_
rlabel metal3 25344 9660 25344 9660 0 u_ppwm/u_ex/_0211_
rlabel metal2 25056 10542 25056 10542 0 u_ppwm/u_ex/_0212_
rlabel metal2 25440 10458 25440 10458 0 u_ppwm/u_ex/_0213_
rlabel metal3 23141 10080 23141 10080 0 u_ppwm/u_ex/_0214_
rlabel metal3 21504 9660 21504 9660 0 u_ppwm/u_ex/_0215_
rlabel metal3 21216 10164 21216 10164 0 u_ppwm/u_ex/_0216_
rlabel metal2 15264 14952 15264 14952 0 u_ppwm/u_ex/_0217_
rlabel metal2 15600 14196 15600 14196 0 u_ppwm/u_ex/_0218_
rlabel metal2 26592 17010 26592 17010 0 u_ppwm/u_ex/_0219_
rlabel metal3 24768 15540 24768 15540 0 u_ppwm/u_ex/_0220_
rlabel metal2 30912 13146 30912 13146 0 u_ppwm/u_ex/_0221_
rlabel metal3 33072 13860 33072 13860 0 u_ppwm/u_ex/_0222_
rlabel metal2 22656 17010 22656 17010 0 u_ppwm/u_ex/_0223_
rlabel metal2 22896 16716 22896 16716 0 u_ppwm/u_ex/_0224_
rlabel metal2 22272 17430 22272 17430 0 u_ppwm/u_ex/_0225_
rlabel metal2 28800 14742 28800 14742 0 u_ppwm/u_ex/_0226_
rlabel metal3 27216 15624 27216 15624 0 u_ppwm/u_ex/_0227_
rlabel metal2 27552 17136 27552 17136 0 u_ppwm/u_ex/_0228_
rlabel metal3 27264 15960 27264 15960 0 u_ppwm/u_ex/_0229_
rlabel metal2 33984 15120 33984 15120 0 u_ppwm/u_ex/_0230_
rlabel metal2 34272 14994 34272 14994 0 u_ppwm/u_ex/_0231_
rlabel metal2 21984 15960 21984 15960 0 u_ppwm/u_ex/_0232_
rlabel metal2 22416 14196 22416 14196 0 u_ppwm/u_ex/_0233_
rlabel metal2 20640 11718 20640 11718 0 u_ppwm/u_ex/_0234_
rlabel metal2 29184 13104 29184 13104 0 u_ppwm/u_ex/_0235_
rlabel metal2 23712 14028 23712 14028 0 u_ppwm/u_ex/_0236_
rlabel metal2 24000 14574 24000 14574 0 u_ppwm/u_ex/_0237_
rlabel metal3 23856 14700 23856 14700 0 u_ppwm/u_ex/_0238_
rlabel metal3 22464 14028 22464 14028 0 u_ppwm/u_ex/_0239_
rlabel metal2 23136 14490 23136 14490 0 u_ppwm/u_ex/_0240_
rlabel metal2 21696 14028 21696 14028 0 u_ppwm/u_ex/_0241_
rlabel metal2 22368 12348 22368 12348 0 u_ppwm/u_ex/_0242_
rlabel metal2 21600 12516 21600 12516 0 u_ppwm/u_ex/_0243_
rlabel metal3 21408 14994 21408 14994 0 u_ppwm/u_ex/_0244_
rlabel metal2 21125 13944 21125 13944 0 u_ppwm/u_ex/_0245_
rlabel metal3 22770 13860 22770 13860 0 u_ppwm/u_ex/_0246_
rlabel metal3 25200 16044 25200 16044 0 u_ppwm/u_ex/_0247_
rlabel metal2 24672 17850 24672 17850 0 u_ppwm/u_ex/_0248_
rlabel metal2 25728 17724 25728 17724 0 u_ppwm/u_ex/_0249_
rlabel metal2 25920 16632 25920 16632 0 u_ppwm/u_ex/_0250_
rlabel metal2 26880 15792 26880 15792 0 u_ppwm/u_ex/_0251_
rlabel metal2 34176 14910 34176 14910 0 u_ppwm/u_ex/_0252_
rlabel metal2 34416 14700 34416 14700 0 u_ppwm/u_ex/_0253_
rlabel metal2 22272 12432 22272 12432 0 u_ppwm/u_ex/_0254_
rlabel metal2 17472 10920 17472 10920 0 u_ppwm/u_ex/_0255_
rlabel metal2 21216 14658 21216 14658 0 u_ppwm/u_ex/_0256_
rlabel metal3 20256 13020 20256 13020 0 u_ppwm/u_ex/_0257_
rlabel metal2 21600 14784 21600 14784 0 u_ppwm/u_ex/_0258_
rlabel metal3 20976 14700 20976 14700 0 u_ppwm/u_ex/_0259_
rlabel metal2 20640 15456 20640 15456 0 u_ppwm/u_ex/_0260_
rlabel metal2 20496 15540 20496 15540 0 u_ppwm/u_ex/_0261_
rlabel metal2 20352 16044 20352 16044 0 u_ppwm/u_ex/_0262_
rlabel metal2 21216 16380 21216 16380 0 u_ppwm/u_ex/_0263_
rlabel metal2 20352 13734 20352 13734 0 u_ppwm/u_ex/_0264_
rlabel metal2 21024 15960 21024 15960 0 u_ppwm/u_ex/_0265_
rlabel metal3 22530 16800 22530 16800 0 u_ppwm/u_ex/_0266_
rlabel metal3 30816 16212 30816 16212 0 u_ppwm/u_ex/_0267_
rlabel metal3 27984 14028 27984 14028 0 u_ppwm/u_ex/_0268_
rlabel metal2 28464 14532 28464 14532 0 u_ppwm/u_ex/_0269_
rlabel metal2 28938 14532 28938 14532 0 u_ppwm/u_ex/_0270_
rlabel metal2 29472 14910 29472 14910 0 u_ppwm/u_ex/_0271_
rlabel metal3 31632 15540 31632 15540 0 u_ppwm/u_ex/_0272_
rlabel metal2 33504 13902 33504 13902 0 u_ppwm/u_ex/_0273_
rlabel metal3 33456 14700 33456 14700 0 u_ppwm/u_ex/_0274_
rlabel metal2 32448 14700 32448 14700 0 u_ppwm/u_ex/_0275_
rlabel metal2 38016 15792 38016 15792 0 u_ppwm/u_ex/_0276_
rlabel metal2 38160 15708 38160 15708 0 u_ppwm/u_ex/_0277_
rlabel metal2 20640 12970 20640 12970 0 u_ppwm/u_ex/_0278_
rlabel metal2 17568 13440 17568 13440 0 u_ppwm/u_ex/_0279_
rlabel metal2 17664 13230 17664 13230 0 u_ppwm/u_ex/_0280_
rlabel metal2 21216 13440 21216 13440 0 u_ppwm/u_ex/_0281_
rlabel metal2 19008 14826 19008 14826 0 u_ppwm/u_ex/_0282_
rlabel metal2 19872 14742 19872 14742 0 u_ppwm/u_ex/_0283_
rlabel metal3 18912 15540 18912 15540 0 u_ppwm/u_ex/_0284_
rlabel metal2 20640 14280 20640 14280 0 u_ppwm/u_ex/_0285_
rlabel metal3 17520 10416 17520 10416 0 u_ppwm/u_ex/_0286_
rlabel metal3 16944 9576 16944 9576 0 u_ppwm/u_ex/_0287_
rlabel metal2 17232 11172 17232 11172 0 u_ppwm/u_ex/_0288_
rlabel metal2 18624 12642 18624 12642 0 u_ppwm/u_ex/_0289_
rlabel metal4 21120 14028 21120 14028 0 u_ppwm/u_ex/_0290_
rlabel metal2 28128 12474 28128 12474 0 u_ppwm/u_ex/_0291_
rlabel metal2 28608 12474 28608 12474 0 u_ppwm/u_ex/_0292_
rlabel metal2 28272 12516 28272 12516 0 u_ppwm/u_ex/_0293_
rlabel metal2 28320 11718 28320 11718 0 u_ppwm/u_ex/_0294_
rlabel metal2 27840 12726 27840 12726 0 u_ppwm/u_ex/_0295_
rlabel metal2 28704 13272 28704 13272 0 u_ppwm/u_ex/_0296_
rlabel metal3 30576 14028 30576 14028 0 u_ppwm/u_ex/_0297_
rlabel metal3 27264 15162 27264 15162 0 u_ppwm/u_ex/_0298_
rlabel metal4 30624 13440 30624 13440 0 u_ppwm/u_ex/_0299_
rlabel metal2 30432 13230 30432 13230 0 u_ppwm/u_ex/_0300_
rlabel metal3 33744 13440 33744 13440 0 u_ppwm/u_ex/_0301_
rlabel metal2 37680 13188 37680 13188 0 u_ppwm/u_ex/_0302_
rlabel metal2 27552 12936 27552 12936 0 u_ppwm/u_ex/_0303_
rlabel metal2 28512 12936 28512 12936 0 u_ppwm/u_ex/_0304_
rlabel metal2 27744 12768 27744 12768 0 u_ppwm/u_ex/_0305_
rlabel metal2 28032 14028 28032 14028 0 u_ppwm/u_ex/_0306_
rlabel metal2 19536 15540 19536 15540 0 u_ppwm/u_ex/_0307_
rlabel metal2 20832 15456 20832 15456 0 u_ppwm/u_ex/_0308_
rlabel metal3 21408 15540 21408 15540 0 u_ppwm/u_ex/_0309_
rlabel metal2 18240 8904 18240 8904 0 u_ppwm/u_ex/_0310_
rlabel metal2 18192 10164 18192 10164 0 u_ppwm/u_ex/_0311_
rlabel metal2 21661 11725 21661 11725 0 u_ppwm/u_ex/_0312_
rlabel metal3 21984 15456 21984 15456 0 u_ppwm/u_ex/_0313_
rlabel metal3 22272 15246 22272 15246 0 u_ppwm/u_ex/_0314_
rlabel metal2 31152 14700 31152 14700 0 u_ppwm/u_ex/_0315_
rlabel metal2 29952 14784 29952 14784 0 u_ppwm/u_ex/_0316_
rlabel metal3 28800 14910 28800 14910 0 u_ppwm/u_ex/_0317_
rlabel metal2 29184 15456 29184 15456 0 u_ppwm/u_ex/_0318_
rlabel metal3 29712 15708 29712 15708 0 u_ppwm/u_ex/_0319_
rlabel metal2 20544 4914 20544 4914 0 u_ppwm/u_ex/_0320_
rlabel metal2 19968 3150 19968 3150 0 u_ppwm/u_ex/_0321_
rlabel metal3 27984 11508 27984 11508 0 u_ppwm/u_ex/_0322_
rlabel metal2 28992 11256 28992 11256 0 u_ppwm/u_ex/_0323_
rlabel metal2 18048 3486 18048 3486 0 u_ppwm/u_ex/_0324_
rlabel metal3 24048 3612 24048 3612 0 u_ppwm/u_ex/_0325_
rlabel metal2 24384 4704 24384 4704 0 u_ppwm/u_ex/_0326_
rlabel metal2 19296 13818 19296 13818 0 u_ppwm/u_ex/_0327_
rlabel metal3 18720 14196 18720 14196 0 u_ppwm/u_ex/_0328_
rlabel metal2 19488 13314 19488 13314 0 u_ppwm/u_ex/_0329_
rlabel metal2 20256 11844 20256 11844 0 u_ppwm/u_ex/_0330_
rlabel metal2 17184 9198 17184 9198 0 u_ppwm/u_ex/_0331_
rlabel metal3 16992 9240 16992 9240 0 u_ppwm/u_ex/_0332_
rlabel metal2 20544 11809 20544 11809 0 u_ppwm/u_ex/_0333_
rlabel metal2 30912 4956 30912 4956 0 u_ppwm/u_ex/_0334_
rlabel metal2 33264 5628 33264 5628 0 u_ppwm/u_ex/_0335_
rlabel metal2 33024 4956 33024 4956 0 u_ppwm/u_ex/_0336_
rlabel metal4 24672 4872 24672 4872 0 u_ppwm/u_ex/_0337_
rlabel metal2 24768 4872 24768 4872 0 u_ppwm/u_ex/_0338_
rlabel metal2 25152 4536 25152 4536 0 u_ppwm/u_ex/_0339_
rlabel metal2 20352 3570 20352 3570 0 u_ppwm/u_ex/_0340_
rlabel metal2 19824 2604 19824 2604 0 u_ppwm/u_ex/_0341_
rlabel metal2 20496 2856 20496 2856 0 u_ppwm/u_ex/_0342_
rlabel metal2 20640 3696 20640 3696 0 u_ppwm/u_ex/_0343_
rlabel metal2 21360 13188 21360 13188 0 u_ppwm/u_ex/_0344_
rlabel metal2 21216 12768 21216 12768 0 u_ppwm/u_ex/_0345_
rlabel metal2 21120 11970 21120 11970 0 u_ppwm/u_ex/_0346_
rlabel metal2 15648 9114 15648 9114 0 u_ppwm/u_ex/_0347_
rlabel metal2 16896 10332 16896 10332 0 u_ppwm/u_ex/_0348_
rlabel metal2 21408 11760 21408 11760 0 u_ppwm/u_ex/_0349_
rlabel metal2 30336 4998 30336 4998 0 u_ppwm/u_ex/_0350_
rlabel metal2 29472 6636 29472 6636 0 u_ppwm/u_ex/_0351_
rlabel metal2 26592 6006 26592 6006 0 u_ppwm/u_ex/_0352_
rlabel metal2 26496 5208 26496 5208 0 u_ppwm/u_ex/_0353_
rlabel metal2 21840 4704 21840 4704 0 u_ppwm/u_ex/_0354_
rlabel metal3 21408 3444 21408 3444 0 u_ppwm/u_ex/_0355_
rlabel metal3 16992 1680 16992 1680 0 u_ppwm/u_ex/_0356_
rlabel metal2 17088 2562 17088 2562 0 u_ppwm/u_ex/_0357_
rlabel metal3 17616 2436 17616 2436 0 u_ppwm/u_ex/_0358_
rlabel metal2 16752 3612 16752 3612 0 u_ppwm/u_ex/_0359_
rlabel metal3 18672 2604 18672 2604 0 u_ppwm/u_ex/_0360_
rlabel metal2 17856 2688 17856 2688 0 u_ppwm/u_ex/_0361_
rlabel metal2 18048 2646 18048 2646 0 u_ppwm/u_ex/_0362_
rlabel metal2 21696 12894 21696 12894 0 u_ppwm/u_ex/_0363_
rlabel metal2 19968 12768 19968 12768 0 u_ppwm/u_ex/_0364_
rlabel metal2 20400 12516 20400 12516 0 u_ppwm/u_ex/_0365_
rlabel metal2 20736 12306 20736 12306 0 u_ppwm/u_ex/_0366_
rlabel metal3 21744 12264 21744 12264 0 u_ppwm/u_ex/_0367_
rlabel metal2 24576 5964 24576 5964 0 u_ppwm/u_ex/_0368_
rlabel metal2 24096 4956 24096 4956 0 u_ppwm/u_ex/_0369_
rlabel metal2 23424 4998 23424 4998 0 u_ppwm/u_ex/_0370_
rlabel metal2 22992 3444 22992 3444 0 u_ppwm/u_ex/_0371_
rlabel metal2 22656 2226 22656 2226 0 u_ppwm/u_ex/_0372_
rlabel metal3 22032 1932 22032 1932 0 u_ppwm/u_ex/_0373_
rlabel metal2 18336 2730 18336 2730 0 u_ppwm/u_ex/_0374_
rlabel metal2 17376 2562 17376 2562 0 u_ppwm/u_ex/_0375_
rlabel metal2 18384 1764 18384 1764 0 u_ppwm/u_ex/_0376_
rlabel metal2 19488 1596 19488 1596 0 u_ppwm/u_ex/_0377_
rlabel via1 19872 11683 19872 11683 0 u_ppwm/u_ex/_0378_
rlabel metal2 20688 11508 20688 11508 0 u_ppwm/u_ex/_0379_
rlabel metal2 21312 6552 21312 6552 0 u_ppwm/u_ex/_0380_
rlabel metal2 21600 7434 21600 7434 0 u_ppwm/u_ex/_0381_
rlabel metal2 21696 7138 21696 7138 0 u_ppwm/u_ex/_0382_
rlabel metal2 20736 6468 20736 6468 0 u_ppwm/u_ex/_0383_
rlabel metal3 20160 1092 20160 1092 0 u_ppwm/u_ex/_0384_
rlabel metal2 19248 1092 19248 1092 0 u_ppwm/u_ex/_0385_
rlabel metal3 17376 2856 17376 2856 0 u_ppwm/u_ex/_0386_
rlabel metal3 16512 2604 16512 2604 0 u_ppwm/u_ex/_0387_
rlabel metal2 17856 3486 17856 3486 0 u_ppwm/u_ex/_0388_
rlabel metal2 18960 4116 18960 4116 0 u_ppwm/u_ex/_0389_
rlabel metal2 20544 6720 20544 6720 0 u_ppwm/u_ex/_0390_
rlabel metal2 19200 5712 19200 5712 0 u_ppwm/u_ex/_0391_
rlabel metal2 18720 4074 18720 4074 0 u_ppwm/u_ex/_0392_
rlabel metal2 18624 4242 18624 4242 0 u_ppwm/u_ex/_0393_
rlabel metal2 18720 12390 18720 12390 0 u_ppwm/u_ex/_0394_
rlabel metal2 18912 12138 18912 12138 0 u_ppwm/u_ex/_0395_
rlabel metal2 18816 5964 18816 5964 0 u_ppwm/u_ex/_0396_
rlabel metal3 24096 6468 24096 6468 0 u_ppwm/u_ex/_0397_
rlabel metal2 23040 5922 23040 5922 0 u_ppwm/u_ex/_0398_
rlabel metal2 18912 5544 18912 5544 0 u_ppwm/u_ex/_0399_
rlabel metal3 16368 5460 16368 5460 0 u_ppwm/u_ex/_0400_
rlabel metal2 13440 6468 13440 6468 0 u_ppwm/u_ex/_0401_
rlabel metal2 18816 7056 18816 7056 0 u_ppwm/u_ex/_0402_
rlabel metal3 17184 5628 17184 5628 0 u_ppwm/u_ex/_0403_
rlabel metal3 17856 5796 17856 5796 0 u_ppwm/u_ex/_0404_
rlabel metal3 17136 7476 17136 7476 0 u_ppwm/u_ex/_0405_
rlabel metal2 18048 11676 18048 11676 0 u_ppwm/u_ex/_0406_
rlabel metal3 18768 11004 18768 11004 0 u_ppwm/u_ex/_0407_
rlabel metal2 23232 10248 23232 10248 0 u_ppwm/u_ex/_0408_
rlabel metal3 22848 10164 22848 10164 0 u_ppwm/u_ex/_0409_
rlabel metal3 17760 10206 17760 10206 0 u_ppwm/u_ex/_0410_
rlabel metal2 17904 8652 17904 8652 0 u_ppwm/u_ex/_0411_
rlabel metal2 17424 8148 17424 8148 0 u_ppwm/u_ex/_0412_
rlabel metal2 31488 7140 31488 7140 0 u_ppwm/u_ex/_0413_
rlabel metal2 32928 13524 32928 13524 0 u_ppwm/u_ex/_0414_
rlabel via2 32928 14530 32928 14530 0 u_ppwm/u_ex/_0415_
rlabel metal2 32544 15918 32544 15918 0 u_ppwm/u_ex/_0416_
rlabel metal2 24912 17220 24912 17220 0 u_ppwm/u_ex/_0417_
rlabel metal2 25152 17472 25152 17472 0 u_ppwm/u_ex/_0418_
rlabel metal2 25248 17472 25248 17472 0 u_ppwm/u_ex/_0419_
rlabel metal2 29568 18606 29568 18606 0 u_ppwm/u_ex/_0420_
rlabel metal2 27840 18018 27840 18018 0 u_ppwm/u_ex/_0421_
rlabel metal2 27744 16674 27744 16674 0 u_ppwm/u_ex/_0422_
rlabel metal3 32832 16380 32832 16380 0 u_ppwm/u_ex/_0423_
rlabel metal3 32640 18732 32640 18732 0 u_ppwm/u_ex/_0424_
rlabel metal2 29376 19194 29376 19194 0 u_ppwm/u_ex/_0425_
rlabel metal2 29712 18564 29712 18564 0 u_ppwm/u_ex/_0426_
rlabel metal2 30336 18816 30336 18816 0 u_ppwm/u_ex/_0427_
rlabel metal2 31488 17094 31488 17094 0 u_ppwm/u_ex/_0428_
rlabel metal3 31392 16380 31392 16380 0 u_ppwm/u_ex/_0429_
rlabel metal2 31776 13776 31776 13776 0 u_ppwm/u_ex/_0430_
rlabel metal2 31776 14532 31776 14532 0 u_ppwm/u_ex/_0431_
rlabel metal2 31440 14952 31440 14952 0 u_ppwm/u_ex/_0432_
rlabel metal3 33024 16212 33024 16212 0 u_ppwm/u_ex/_0433_
rlabel metal2 34080 16926 34080 16926 0 u_ppwm/u_ex/_0434_
rlabel metal2 28896 17136 28896 17136 0 u_ppwm/u_ex/_0435_
rlabel metal2 30000 17724 30000 17724 0 u_ppwm/u_ex/_0436_
rlabel metal2 29424 17892 29424 17892 0 u_ppwm/u_ex/_0437_
rlabel metal2 29856 17640 29856 17640 0 u_ppwm/u_ex/_0438_
rlabel metal2 29616 16464 29616 16464 0 u_ppwm/u_ex/_0439_
rlabel metal2 32448 12642 32448 12642 0 u_ppwm/u_ex/_0440_
rlabel metal3 32016 13188 32016 13188 0 u_ppwm/u_ex/_0441_
rlabel metal2 31680 13482 31680 13482 0 u_ppwm/u_ex/_0442_
rlabel metal2 29664 15792 29664 15792 0 u_ppwm/u_ex/_0443_
rlabel metal3 30096 15372 30096 15372 0 u_ppwm/u_ex/_0444_
rlabel metal3 37200 16044 37200 16044 0 u_ppwm/u_ex/_0445_
rlabel metal3 28272 17892 28272 17892 0 u_ppwm/u_ex/_0446_
rlabel metal2 29040 16884 29040 16884 0 u_ppwm/u_ex/_0447_
rlabel metal2 30720 17808 30720 17808 0 u_ppwm/u_ex/_0448_
rlabel metal2 30816 17808 30816 17808 0 u_ppwm/u_ex/_0449_
rlabel metal2 32064 11970 32064 11970 0 u_ppwm/u_ex/_0450_
rlabel metal2 31872 13146 31872 13146 0 u_ppwm/u_ex/_0451_
rlabel metal2 31488 15708 31488 15708 0 u_ppwm/u_ex/_0452_
rlabel metal2 30432 17304 30432 17304 0 u_ppwm/u_ex/_0453_
rlabel metal2 30816 17052 30816 17052 0 u_ppwm/u_ex/_0454_
rlabel metal2 29184 5040 29184 5040 0 u_ppwm/u_ex/_0455_
rlabel metal2 29376 4914 29376 4914 0 u_ppwm/u_ex/_0456_
rlabel metal2 28800 17304 28800 17304 0 u_ppwm/u_ex/_0457_
rlabel metal3 28560 17052 28560 17052 0 u_ppwm/u_ex/_0458_
rlabel metal2 28752 16044 28752 16044 0 u_ppwm/u_ex/_0459_
rlabel via2 29855 5040 29855 5040 0 u_ppwm/u_ex/_0460_
rlabel metal3 30528 4956 30528 4956 0 u_ppwm/u_ex/_0461_
rlabel metal3 32496 5628 32496 5628 0 u_ppwm/u_ex/_0462_
rlabel metal2 32064 5752 32064 5752 0 u_ppwm/u_ex/_0463_
rlabel metal2 31200 5376 31200 5376 0 u_ppwm/u_ex/_0464_
rlabel metal2 31776 3612 31776 3612 0 u_ppwm/u_ex/_0465_
rlabel metal3 31824 3444 31824 3444 0 u_ppwm/u_ex/_0466_
rlabel metal2 29376 5124 29376 5124 0 u_ppwm/u_ex/_0467_
rlabel metal3 29856 3486 29856 3486 0 u_ppwm/u_ex/_0468_
rlabel metal3 29136 5460 29136 5460 0 u_ppwm/u_ex/_0469_
rlabel metal2 29856 5418 29856 5418 0 u_ppwm/u_ex/_0470_
rlabel metal2 30528 4998 30528 4998 0 u_ppwm/u_ex/_0471_
rlabel metal3 31584 6552 31584 6552 0 u_ppwm/u_ex/_0472_
rlabel metal2 31872 7180 31872 7180 0 u_ppwm/u_ex/_0473_
rlabel metal2 30624 5460 30624 5460 0 u_ppwm/u_ex/_0474_
rlabel metal2 30240 5376 30240 5376 0 u_ppwm/u_ex/_0475_
rlabel metal2 31392 4872 31392 4872 0 u_ppwm/u_ex/_0476_
rlabel metal3 28272 4116 28272 4116 0 u_ppwm/u_ex/_0477_
rlabel metal2 27312 2520 27312 2520 0 u_ppwm/u_ex/_0478_
rlabel metal2 27216 2856 27216 2856 0 u_ppwm/u_ex/_0479_
rlabel metal2 29088 5502 29088 5502 0 u_ppwm/u_ex/_0480_
rlabel metal2 28848 3612 28848 3612 0 u_ppwm/u_ex/_0481_
rlabel metal2 29760 3738 29760 3738 0 u_ppwm/u_ex/_0482_
rlabel metal2 27840 4200 27840 4200 0 u_ppwm/u_ex/_0483_
rlabel metal2 28320 3150 28320 3150 0 u_ppwm/u_ex/_0484_
rlabel metal3 28896 3444 28896 3444 0 u_ppwm/u_ex/_0485_
rlabel metal2 32640 5796 32640 5796 0 u_ppwm/u_ex/_0486_
rlabel metal2 32736 5878 32736 5878 0 u_ppwm/u_ex/_0487_
rlabel metal2 29472 3948 29472 3948 0 u_ppwm/u_ex/_0488_
rlabel metal2 29184 2898 29184 2898 0 u_ppwm/u_ex/_0489_
rlabel metal2 29568 2604 29568 2604 0 u_ppwm/u_ex/_0490_
rlabel metal2 26208 4074 26208 4074 0 u_ppwm/u_ex/_0491_
rlabel metal2 26688 4200 26688 4200 0 u_ppwm/u_ex/_0492_
rlabel metal2 26304 4368 26304 4368 0 u_ppwm/u_ex/_0493_
rlabel metal2 25824 4536 25824 4536 0 u_ppwm/u_ex/_0494_
rlabel metal3 23856 5628 23856 5628 0 u_ppwm/u_ex/_0495_
rlabel metal2 23520 5796 23520 5796 0 u_ppwm/u_ex/_0496_
rlabel metal2 22992 4956 22992 4956 0 u_ppwm/u_ex/_0497_
rlabel metal2 22752 5376 22752 5376 0 u_ppwm/u_ex/_0498_
rlabel metal2 25920 4158 25920 4158 0 u_ppwm/u_ex/_0499_
rlabel metal2 24000 3864 24000 3864 0 u_ppwm/u_ex/_0500_
rlabel metal2 27648 4368 27648 4368 0 u_ppwm/u_ex/_0501_
rlabel metal3 27072 4956 27072 4956 0 u_ppwm/u_ex/_0502_
rlabel metal2 27504 4956 27504 4956 0 u_ppwm/u_ex/_0503_
rlabel metal2 17760 4242 17760 4242 0 u_ppwm/u_ex/_0504_
rlabel metal2 17088 4578 17088 4578 0 u_ppwm/u_ex/_0505_
rlabel metal2 17664 4620 17664 4620 0 u_ppwm/u_ex/_0506_
rlabel metal2 17472 3696 17472 3696 0 u_ppwm/u_ex/_0507_
rlabel metal2 17568 3696 17568 3696 0 u_ppwm/u_ex/_0508_
rlabel metal2 22464 5670 22464 5670 0 u_ppwm/u_ex/_0509_
rlabel metal2 22560 5836 22560 5836 0 u_ppwm/u_ex/_0510_
rlabel metal2 17952 6342 17952 6342 0 u_ppwm/u_ex/_0511_
rlabel metal2 18144 5166 18144 5166 0 u_ppwm/u_ex/_0512_
rlabel metal2 18432 4158 18432 4158 0 u_ppwm/u_ex/_0513_
rlabel metal2 16224 5502 16224 5502 0 u_ppwm/u_ex/_0514_
rlabel metal2 17184 6930 17184 6930 0 u_ppwm/u_ex/_0515_
rlabel metal3 17904 6636 17904 6636 0 u_ppwm/u_ex/_0516_
rlabel metal3 18432 6132 18432 6132 0 u_ppwm/u_ex/_0517_
rlabel metal2 23952 10164 23952 10164 0 u_ppwm/u_ex/_0518_
rlabel metal2 24288 10710 24288 10710 0 u_ppwm/u_ex/_0519_
rlabel metal3 21936 11004 21936 11004 0 u_ppwm/u_ex/_0520_
rlabel metal3 18384 5964 18384 5964 0 u_ppwm/u_ex/_0521_
rlabel metal3 20064 5754 20064 5754 0 u_ppwm/u_ex/_0522_
rlabel metal3 17904 8484 17904 8484 0 u_ppwm/u_ex/_0523_
rlabel metal2 17472 9156 17472 9156 0 u_ppwm/u_ex/_0524_
rlabel metal3 17856 8778 17856 8778 0 u_ppwm/u_ex/_0525_
rlabel metal2 34656 7182 34656 7182 0 u_ppwm/u_ex/_0526_
rlabel metal2 30912 6804 30912 6804 0 u_ppwm/u_ex/_0527_
rlabel metal3 35376 6468 35376 6468 0 u_ppwm/u_ex/_0528_
rlabel metal2 35424 11508 35424 11508 0 u_ppwm/u_ex/_0529_
rlabel metal2 24864 9450 24864 9450 0 u_ppwm/u_ex/_0530_
rlabel metal2 26592 7518 26592 7518 0 u_ppwm/u_ex/_0531_
rlabel metal2 21024 7896 21024 7896 0 u_ppwm/u_ex/_0532_
rlabel metal2 31584 8862 31584 8862 0 u_ppwm/u_ex/_0533_
rlabel metal2 35712 7770 35712 7770 0 u_ppwm/u_ex/_0534_
rlabel metal2 18624 11088 18624 11088 0 u_ppwm/u_ex/cmp_flag_q
rlabel metal3 26976 18732 26976 18732 0 u_ppwm/u_ex/reg_value_q\[0\]
rlabel metal2 37056 18648 37056 18648 0 u_ppwm/u_ex/reg_value_q\[1\]
rlabel metal2 39552 17346 39552 17346 0 u_ppwm/u_ex/reg_value_q\[2\]
rlabel metal2 36672 17010 36672 17010 0 u_ppwm/u_ex/reg_value_q\[3\]
rlabel metal2 35712 4326 35712 4326 0 u_ppwm/u_ex/reg_value_q\[4\]
rlabel metal4 28992 5124 28992 5124 0 u_ppwm/u_ex/reg_value_q\[5\]
rlabel metal2 31248 1932 31248 1932 0 u_ppwm/u_ex/reg_value_q\[6\]
rlabel metal2 20832 7938 20832 7938 0 u_ppwm/u_ex/reg_value_q\[7\]
rlabel metal2 16080 5376 16080 5376 0 u_ppwm/u_ex/reg_value_q\[8\]
rlabel metal2 16896 7182 16896 7182 0 u_ppwm/u_ex/reg_value_q\[9\]
rlabel metal2 14784 18984 14784 18984 0 u_ppwm/u_ex/state_q\[0\]
rlabel metal2 17808 17052 17808 17052 0 u_ppwm/u_ex/state_q\[1\]
rlabel metal2 20352 19572 20352 19572 0 u_ppwm/u_ex/state_q\[2\]
rlabel metal2 43296 13566 43296 13566 0 u_ppwm/u_global_counter/_000_
rlabel metal2 41760 14448 41760 14448 0 u_ppwm/u_global_counter/_001_
rlabel metal2 41568 11256 41568 11256 0 u_ppwm/u_global_counter/_002_
rlabel metal3 43248 12348 43248 12348 0 u_ppwm/u_global_counter/_003_
rlabel metal2 41952 7098 41952 7098 0 u_ppwm/u_global_counter/_004_
rlabel metal2 42432 5460 42432 5460 0 u_ppwm/u_global_counter/_005_
rlabel metal2 44496 5544 44496 5544 0 u_ppwm/u_global_counter/_006_
rlabel metal2 45216 9912 45216 9912 0 u_ppwm/u_global_counter/_007_
rlabel metal2 46560 8274 46560 8274 0 u_ppwm/u_global_counter/_008_
rlabel metal2 49440 10458 49440 10458 0 u_ppwm/u_global_counter/_009_
rlabel metal2 46752 12138 46752 12138 0 u_ppwm/u_global_counter/_010_
rlabel metal3 42816 13356 42816 13356 0 u_ppwm/u_global_counter/_011_
rlabel metal3 41580 10206 41580 10206 0 u_ppwm/u_global_counter/_012_
rlabel metal3 38352 9324 38352 9324 0 u_ppwm/u_global_counter/_013_
rlabel metal2 38976 8736 38976 8736 0 u_ppwm/u_global_counter/_014_
rlabel metal2 40800 5628 40800 5628 0 u_ppwm/u_global_counter/_015_
rlabel metal3 39024 4956 39024 4956 0 u_ppwm/u_global_counter/_016_
rlabel metal3 37392 5628 37392 5628 0 u_ppwm/u_global_counter/_017_
rlabel metal2 37728 3318 37728 3318 0 u_ppwm/u_global_counter/_018_
rlabel metal2 36384 4494 36384 4494 0 u_ppwm/u_global_counter/_019_
rlabel metal2 41088 9366 41088 9366 0 u_ppwm/u_global_counter/_020_
rlabel metal3 43488 11928 43488 11928 0 u_ppwm/u_global_counter/_021_
rlabel metal2 38400 9492 38400 9492 0 u_ppwm/u_global_counter/_022_
rlabel metal3 39792 5628 39792 5628 0 u_ppwm/u_global_counter/_023_
rlabel metal2 36960 5754 36960 5754 0 u_ppwm/u_global_counter/_024_
rlabel metal2 38112 4242 38112 4242 0 u_ppwm/u_global_counter/_025_
rlabel metal3 44256 9492 44256 9492 0 u_ppwm/u_global_counter/_026_
rlabel metal2 40512 11634 40512 11634 0 u_ppwm/u_global_counter/_027_
rlabel metal2 41376 14448 41376 14448 0 u_ppwm/u_global_counter/_028_
rlabel metal3 42384 12348 42384 12348 0 u_ppwm/u_global_counter/_029_
rlabel metal3 42240 5628 42240 5628 0 u_ppwm/u_global_counter/_030_
rlabel metal2 41376 8946 41376 8946 0 u_ppwm/u_global_counter/_031_
rlabel metal2 39936 7266 39936 7266 0 u_ppwm/u_global_counter/_032_
rlabel metal2 42720 7476 42720 7476 0 u_ppwm/u_global_counter/_033_
rlabel metal2 43104 9786 43104 9786 0 u_ppwm/u_global_counter/_034_
rlabel metal3 48000 11004 48000 11004 0 u_ppwm/u_global_counter/_035_
rlabel metal3 44256 5544 44256 5544 0 u_ppwm/u_global_counter/_036_
rlabel metal3 47712 11676 47712 11676 0 u_ppwm/u_global_counter/_037_
rlabel metal2 48960 10710 48960 10710 0 u_ppwm/u_global_counter/_038_
rlabel metal2 45792 10920 45792 10920 0 u_ppwm/u_global_counter/_039_
rlabel metal3 42720 9492 42720 9492 0 u_ppwm/u_global_counter/_040_
rlabel metal2 38784 8106 38784 8106 0 u_ppwm/u_global_counter/_041_
rlabel metal2 37824 10626 37824 10626 0 u_ppwm/u_global_counter/_042_
rlabel metal2 38784 10710 38784 10710 0 u_ppwm/u_global_counter/_043_
rlabel metal3 38928 9408 38928 9408 0 u_ppwm/u_global_counter/_044_
rlabel metal2 38352 7812 38352 7812 0 u_ppwm/u_global_counter/_045_
rlabel metal2 40992 6300 40992 6300 0 u_ppwm/u_global_counter/_046_
rlabel metal2 37872 5292 37872 5292 0 u_ppwm/u_global_counter/_047_
rlabel metal3 39648 6468 39648 6468 0 u_ppwm/u_global_counter/_048_
rlabel metal2 37440 3570 37440 3570 0 u_ppwm/u_global_counter/_049_
rlabel metal2 37056 5586 37056 5586 0 u_ppwm/u_global_counter/_050_
rlabel metal2 37152 2604 37152 2604 0 u_ppwm/u_global_counter/_051_
rlabel metal2 37824 3318 37824 3318 0 u_ppwm/u_global_counter/_052_
rlabel metal2 5568 26418 5568 26418 0 u_ppwm/u_mem/_0000_
rlabel metal3 4464 23268 4464 23268 0 u_ppwm/u_mem/_0001_
rlabel metal3 4992 23100 4992 23100 0 u_ppwm/u_mem/_0002_
rlabel metal2 8256 21210 8256 21210 0 u_ppwm/u_mem/_0003_
rlabel metal2 7872 18018 7872 18018 0 u_ppwm/u_mem/_0004_
rlabel metal2 8544 16968 8544 16968 0 u_ppwm/u_mem/_0005_
rlabel metal2 12096 17808 12096 17808 0 u_ppwm/u_mem/_0006_
rlabel metal3 37536 20076 37536 20076 0 u_ppwm/u_mem/_0007_
rlabel metal2 48000 21630 48000 21630 0 u_ppwm/u_mem/_0008_
rlabel metal2 48672 25032 48672 25032 0 u_ppwm/u_mem/_0009_
rlabel metal2 48576 28392 48576 28392 0 u_ppwm/u_mem/_0010_
rlabel metal3 43584 27048 43584 27048 0 u_ppwm/u_mem/_0011_
rlabel metal3 40560 25284 40560 25284 0 u_ppwm/u_mem/_0012_
rlabel metal2 40704 17808 40704 17808 0 u_ppwm/u_mem/_0013_
rlabel metal2 37920 19152 37920 19152 0 u_ppwm/u_mem/_0014_
rlabel metal2 44064 19110 44064 19110 0 u_ppwm/u_mem/_0015_
rlabel metal3 48624 22176 48624 22176 0 u_ppwm/u_mem/_0016_
rlabel metal2 48288 26208 48288 26208 0 u_ppwm/u_mem/_0017_
rlabel metal2 45024 26418 45024 26418 0 u_ppwm/u_mem/_0018_
rlabel metal2 41664 25032 41664 25032 0 u_ppwm/u_mem/_0019_
rlabel metal2 41472 23142 41472 23142 0 u_ppwm/u_mem/_0020_
rlabel metal2 40512 21042 40512 21042 0 u_ppwm/u_mem/_0021_
rlabel metal2 47712 24528 47712 24528 0 u_ppwm/u_mem/_0022_
rlabel metal2 49152 26040 49152 26040 0 u_ppwm/u_mem/_0023_
rlabel metal3 44736 28224 44736 28224 0 u_ppwm/u_mem/_0024_
rlabel metal2 42336 29526 42336 29526 0 u_ppwm/u_mem/_0025_
rlabel metal3 39888 27048 39888 27048 0 u_ppwm/u_mem/_0026_
rlabel metal2 37344 21966 37344 21966 0 u_ppwm/u_mem/_0027_
rlabel metal3 42528 20244 42528 20244 0 u_ppwm/u_mem/_0028_
rlabel metal2 46560 21084 46560 21084 0 u_ppwm/u_mem/_0029_
rlabel metal2 45696 22428 45696 22428 0 u_ppwm/u_mem/_0030_
rlabel metal2 43200 29190 43200 29190 0 u_ppwm/u_mem/_0031_
rlabel metal2 40416 29442 40416 29442 0 u_ppwm/u_mem/_0032_
rlabel metal2 36960 27048 36960 27048 0 u_ppwm/u_mem/_0033_
rlabel metal2 36384 23730 36384 23730 0 u_ppwm/u_mem/_0034_
rlabel metal2 33792 22218 33792 22218 0 u_ppwm/u_mem/_0035_
rlabel metal2 35040 26376 35040 26376 0 u_ppwm/u_mem/_0036_
rlabel metal2 33600 28392 33600 28392 0 u_ppwm/u_mem/_0037_
rlabel metal2 31824 29232 31824 29232 0 u_ppwm/u_mem/_0038_
rlabel metal2 27312 30492 27312 30492 0 u_ppwm/u_mem/_0039_
rlabel metal2 25008 27468 25008 27468 0 u_ppwm/u_mem/_0040_
rlabel metal2 24768 25368 24768 25368 0 u_ppwm/u_mem/_0041_
rlabel metal2 31344 21420 31344 21420 0 u_ppwm/u_mem/_0042_
rlabel metal2 32160 23856 32160 23856 0 u_ppwm/u_mem/_0043_
rlabel metal2 32640 27888 32640 27888 0 u_ppwm/u_mem/_0044_
rlabel metal2 27840 28182 27840 28182 0 u_ppwm/u_mem/_0045_
rlabel metal2 22272 30702 22272 30702 0 u_ppwm/u_mem/_0046_
rlabel metal3 22848 29316 22848 29316 0 u_ppwm/u_mem/_0047_
rlabel metal2 30528 31626 30528 31626 0 u_ppwm/u_mem/_0048_
rlabel metal2 37056 29778 37056 29778 0 u_ppwm/u_mem/_0049_
rlabel metal2 38304 30702 38304 30702 0 u_ppwm/u_mem/_0050_
rlabel metal2 34176 33726 34176 33726 0 u_ppwm/u_mem/_0051_
rlabel metal2 32208 33096 32208 33096 0 u_ppwm/u_mem/_0052_
rlabel metal2 29904 33684 29904 33684 0 u_ppwm/u_mem/_0053_
rlabel metal2 27072 32088 27072 32088 0 u_ppwm/u_mem/_0054_
rlabel metal3 24624 29736 24624 29736 0 u_ppwm/u_mem/_0055_
rlabel metal2 36960 29400 36960 29400 0 u_ppwm/u_mem/_0056_
rlabel metal2 36672 32928 36672 32928 0 u_ppwm/u_mem/_0057_
rlabel metal2 35616 31038 35616 31038 0 u_ppwm/u_mem/_0058_
rlabel metal2 32256 34062 32256 34062 0 u_ppwm/u_mem/_0059_
rlabel metal3 29616 33852 29616 33852 0 u_ppwm/u_mem/_0060_
rlabel metal2 25968 33852 25968 33852 0 u_ppwm/u_mem/_0061_
rlabel metal2 23136 34524 23136 34524 0 u_ppwm/u_mem/_0062_
rlabel metal2 22176 34062 22176 34062 0 u_ppwm/u_mem/_0063_
rlabel metal2 17184 35574 17184 35574 0 u_ppwm/u_mem/_0064_
rlabel metal3 11616 36540 11616 36540 0 u_ppwm/u_mem/_0065_
rlabel metal2 7056 36120 7056 36120 0 u_ppwm/u_mem/_0066_
rlabel metal2 3456 35532 3456 35532 0 u_ppwm/u_mem/_0067_
rlabel metal2 1152 32844 1152 32844 0 u_ppwm/u_mem/_0068_
rlabel metal2 18672 32844 18672 32844 0 u_ppwm/u_mem/_0069_
rlabel metal2 19680 34440 19680 34440 0 u_ppwm/u_mem/_0070_
rlabel metal3 15984 36876 15984 36876 0 u_ppwm/u_mem/_0071_
rlabel metal2 10752 38136 10752 38136 0 u_ppwm/u_mem/_0072_
rlabel metal2 8352 36708 8352 36708 0 u_ppwm/u_mem/_0073_
rlabel metal3 5520 34608 5520 34608 0 u_ppwm/u_mem/_0074_
rlabel metal2 1536 31206 1536 31206 0 u_ppwm/u_mem/_0075_
rlabel metal2 10944 31500 10944 31500 0 u_ppwm/u_mem/_0076_
rlabel metal2 16320 31290 16320 31290 0 u_ppwm/u_mem/_0077_
rlabel metal3 15408 31584 15408 31584 0 u_ppwm/u_mem/_0078_
rlabel metal2 10944 34440 10944 34440 0 u_ppwm/u_mem/_0079_
rlabel metal2 7776 34230 7776 34230 0 u_ppwm/u_mem/_0080_
rlabel metal2 1728 33684 1728 33684 0 u_ppwm/u_mem/_0081_
rlabel metal2 4896 30156 4896 30156 0 u_ppwm/u_mem/_0082_
rlabel metal2 6288 29820 6288 29820 0 u_ppwm/u_mem/_0083_
rlabel metal2 14016 30828 14016 30828 0 u_ppwm/u_mem/_0084_
rlabel metal2 13728 31794 13728 31794 0 u_ppwm/u_mem/_0085_
rlabel metal2 11808 32508 11808 32508 0 u_ppwm/u_mem/_0086_
rlabel metal2 7248 32340 7248 32340 0 u_ppwm/u_mem/_0087_
rlabel metal2 1248 33516 1248 33516 0 u_ppwm/u_mem/_0088_
rlabel metal2 4608 29064 4608 29064 0 u_ppwm/u_mem/_0089_
rlabel metal2 1248 27258 1248 27258 0 u_ppwm/u_mem/_0090_
rlabel metal2 8064 26670 8064 26670 0 u_ppwm/u_mem/_0091_
rlabel metal2 9696 29778 9696 29778 0 u_ppwm/u_mem/_0092_
rlabel metal2 16704 29652 16704 29652 0 u_ppwm/u_mem/_0093_
rlabel metal3 16752 27720 16752 27720 0 u_ppwm/u_mem/_0094_
rlabel metal3 18288 25536 18288 25536 0 u_ppwm/u_mem/_0095_
rlabel metal2 14304 23856 14304 23856 0 u_ppwm/u_mem/_0096_
rlabel metal2 11040 25368 11040 25368 0 u_ppwm/u_mem/_0097_
rlabel metal2 8832 26670 8832 26670 0 u_ppwm/u_mem/_0098_
rlabel metal2 12480 27636 12480 27636 0 u_ppwm/u_mem/_0099_
rlabel metal3 19296 28308 19296 28308 0 u_ppwm/u_mem/_0100_
rlabel metal2 20448 26376 20448 26376 0 u_ppwm/u_mem/_0101_
rlabel metal2 18000 23268 18000 23268 0 u_ppwm/u_mem/_0102_
rlabel metal2 16656 21672 16656 21672 0 u_ppwm/u_mem/_0103_
rlabel metal2 14880 22806 14880 22806 0 u_ppwm/u_mem/_0104_
rlabel metal2 11424 19782 11424 19782 0 u_ppwm/u_mem/_0105_
rlabel metal2 9984 20706 9984 20706 0 u_ppwm/u_mem/_0106_
rlabel metal2 7584 24654 7584 24654 0 u_ppwm/u_mem/_0107_
rlabel metal3 1536 24780 1536 24780 0 u_ppwm/u_mem/_0108_
rlabel metal3 2928 23688 2928 23688 0 u_ppwm/u_mem/_0109_
rlabel metal2 2112 21504 2112 21504 0 u_ppwm/u_mem/_0110_
rlabel metal2 6432 22806 6432 22806 0 u_ppwm/u_mem/_0111_
rlabel metal2 10848 20832 10848 20832 0 u_ppwm/u_mem/_0112_
rlabel metal2 10752 23016 10752 23016 0 u_ppwm/u_mem/_0113_
rlabel metal2 6912 26040 6912 26040 0 u_ppwm/u_mem/_0114_
rlabel metal2 1728 26418 1728 26418 0 u_ppwm/u_mem/_0115_
rlabel metal2 4032 23982 4032 23982 0 u_ppwm/u_mem/_0116_
rlabel metal3 3312 22176 3312 22176 0 u_ppwm/u_mem/_0117_
rlabel metal2 6528 19782 6528 19782 0 u_ppwm/u_mem/_0118_
rlabel metal2 1920 18942 1920 18942 0 u_ppwm/u_mem/_0119_
rlabel metal3 1680 16380 1680 16380 0 u_ppwm/u_mem/_0120_
rlabel metal2 5040 13860 5040 13860 0 u_ppwm/u_mem/_0121_
rlabel metal3 1440 15540 1440 15540 0 u_ppwm/u_mem/_0122_
rlabel metal2 5760 14196 5760 14196 0 u_ppwm/u_mem/_0123_
rlabel metal2 4896 15498 4896 15498 0 u_ppwm/u_mem/_0124_
rlabel metal2 8352 16758 8352 16758 0 u_ppwm/u_mem/_0125_
rlabel metal2 4800 21378 4800 21378 0 u_ppwm/u_mem/_0126_
rlabel metal2 6432 17724 6432 17724 0 u_ppwm/u_mem/_0127_
rlabel metal2 4320 21000 4320 21000 0 u_ppwm/u_mem/_0128_
rlabel metal2 864 25578 864 25578 0 u_ppwm/u_mem/_0129_
rlabel metal2 8064 26334 8064 26334 0 u_ppwm/u_mem/_0130_
rlabel metal2 8736 23520 8736 23520 0 u_ppwm/u_mem/_0131_
rlabel metal2 10368 21042 10368 21042 0 u_ppwm/u_mem/_0132_
rlabel metal3 6816 22260 6816 22260 0 u_ppwm/u_mem/_0133_
rlabel metal2 5376 21630 5376 21630 0 u_ppwm/u_mem/_0134_
rlabel metal3 4320 23772 4320 23772 0 u_ppwm/u_mem/_0135_
rlabel metal2 2208 25242 2208 25242 0 u_ppwm/u_mem/_0136_
rlabel metal2 5952 24864 5952 24864 0 u_ppwm/u_mem/_0137_
rlabel metal2 8832 21420 8832 21420 0 u_ppwm/u_mem/_0138_
rlabel metal2 11712 20034 11712 20034 0 u_ppwm/u_mem/_0139_
rlabel metal2 14640 21000 14640 21000 0 u_ppwm/u_mem/_0140_
rlabel metal2 16320 22806 16320 22806 0 u_ppwm/u_mem/_0141_
rlabel metal2 18240 23394 18240 23394 0 u_ppwm/u_mem/_0142_
rlabel metal2 19392 26880 19392 26880 0 u_ppwm/u_mem/_0143_
rlabel metal2 19921 29064 19921 29064 0 u_ppwm/u_mem/_0144_
rlabel metal2 12768 27258 12768 27258 0 u_ppwm/u_mem/_0145_
rlabel metal2 9648 26712 9648 26712 0 u_ppwm/u_mem/_0146_
rlabel metal3 12192 25326 12192 25326 0 u_ppwm/u_mem/_0147_
rlabel metal2 13824 24066 13824 24066 0 u_ppwm/u_mem/_0148_
rlabel metal2 17088 25032 17088 25032 0 u_ppwm/u_mem/_0149_
rlabel metal2 17712 27048 17712 27048 0 u_ppwm/u_mem/_0150_
rlabel metal3 17664 29064 17664 29064 0 u_ppwm/u_mem/_0151_
rlabel metal2 14448 28896 14448 28896 0 u_ppwm/u_mem/_0152_
rlabel metal3 7200 26796 7200 26796 0 u_ppwm/u_mem/_0153_
rlabel metal2 6048 27132 6048 27132 0 u_ppwm/u_mem/_0154_
rlabel metal3 3312 27048 3312 27048 0 u_ppwm/u_mem/_0155_
rlabel metal2 2448 33180 2448 33180 0 u_ppwm/u_mem/_0156_
rlabel metal2 7488 32844 7488 32844 0 u_ppwm/u_mem/_0157_
rlabel metal3 10320 31500 10320 31500 0 u_ppwm/u_mem/_0158_
rlabel metal2 13536 31374 13536 31374 0 u_ppwm/u_mem/_0159_
rlabel metal3 13776 31332 13776 31332 0 u_ppwm/u_mem/_0160_
rlabel metal2 7008 28644 7008 28644 0 u_ppwm/u_mem/_0161_
rlabel metal3 3648 29820 3648 29820 0 u_ppwm/u_mem/_0162_
rlabel metal3 2832 32844 2832 32844 0 u_ppwm/u_mem/_0163_
rlabel metal2 6816 32634 6816 32634 0 u_ppwm/u_mem/_0164_
rlabel metal2 9408 34104 9408 34104 0 u_ppwm/u_mem/_0165_
rlabel metal2 14880 31920 14880 31920 0 u_ppwm/u_mem/_0166_
rlabel metal2 16128 31626 16128 31626 0 u_ppwm/u_mem/_0167_
rlabel metal2 14592 30954 14592 30954 0 u_ppwm/u_mem/_0168_
rlabel metal2 6336 31542 6336 31542 0 u_ppwm/u_mem/_0169_
rlabel metal2 6240 33726 6240 33726 0 u_ppwm/u_mem/_0170_
rlabel metal2 8064 36246 8064 36246 0 u_ppwm/u_mem/_0171_
rlabel metal2 11904 38304 11904 38304 0 u_ppwm/u_mem/_0172_
rlabel metal3 15168 36708 15168 36708 0 u_ppwm/u_mem/_0173_
rlabel metal2 18336 34104 18336 34104 0 u_ppwm/u_mem/_0174_
rlabel metal3 19344 33096 19344 33096 0 u_ppwm/u_mem/_0175_
rlabel metal2 6144 32004 6144 32004 0 u_ppwm/u_mem/_0176_
rlabel metal2 6432 32928 6432 32928 0 u_ppwm/u_mem/_0177_
rlabel metal2 6624 36078 6624 36078 0 u_ppwm/u_mem/_0178_
rlabel metal2 11136 36834 11136 36834 0 u_ppwm/u_mem/_0179_
rlabel metal2 17376 35826 17376 35826 0 u_ppwm/u_mem/_0180_
rlabel metal2 22368 34692 22368 34692 0 u_ppwm/u_mem/_0181_
rlabel metal2 23232 33096 23232 33096 0 u_ppwm/u_mem/_0182_
rlabel metal3 25920 33684 25920 33684 0 u_ppwm/u_mem/_0183_
rlabel metal2 28512 33684 28512 33684 0 u_ppwm/u_mem/_0184_
rlabel metal3 31440 33852 31440 33852 0 u_ppwm/u_mem/_0185_
rlabel metal3 34848 30660 34848 30660 0 u_ppwm/u_mem/_0186_
rlabel metal3 36000 32340 36000 32340 0 u_ppwm/u_mem/_0187_
rlabel metal2 35328 29400 35328 29400 0 u_ppwm/u_mem/_0188_
rlabel metal3 26064 29316 26064 29316 0 u_ppwm/u_mem/_0189_
rlabel metal2 26496 31626 26496 31626 0 u_ppwm/u_mem/_0190_
rlabel metal2 29376 31626 29376 31626 0 u_ppwm/u_mem/_0191_
rlabel metal2 33216 32592 33216 32592 0 u_ppwm/u_mem/_0192_
rlabel metal3 34512 32844 34512 32844 0 u_ppwm/u_mem/_0193_
rlabel metal2 36480 32130 36480 32130 0 u_ppwm/u_mem/_0194_
rlabel metal2 37248 29770 37248 29770 0 u_ppwm/u_mem/_0195_
rlabel metal3 31824 32172 31824 32172 0 u_ppwm/u_mem/_0196_
rlabel metal3 29082 29064 29082 29064 0 u_ppwm/u_mem/_0197_
rlabel metal2 21984 29736 21984 29736 0 u_ppwm/u_mem/_0198_
rlabel metal3 27600 29064 27600 29064 0 u_ppwm/u_mem/_0199_
rlabel metal3 30576 27720 30576 27720 0 u_ppwm/u_mem/_0200_
rlabel metal2 31008 24066 31008 24066 0 u_ppwm/u_mem/_0201_
rlabel metal2 32256 21294 32256 21294 0 u_ppwm/u_mem/_0202_
rlabel metal2 26400 25032 26400 25032 0 u_ppwm/u_mem/_0203_
rlabel metal3 25056 27636 25056 27636 0 u_ppwm/u_mem/_0204_
rlabel metal2 26832 30072 26832 30072 0 u_ppwm/u_mem/_0205_
rlabel metal2 32448 29316 32448 29316 0 u_ppwm/u_mem/_0206_
rlabel metal3 32352 27384 32352 27384 0 u_ppwm/u_mem/_0207_
rlabel metal2 35472 26628 35472 26628 0 u_ppwm/u_mem/_0208_
rlabel metal2 32928 22302 32928 22302 0 u_ppwm/u_mem/_0209_
rlabel metal2 34272 23142 34272 23142 0 u_ppwm/u_mem/_0210_
rlabel metal2 38688 24696 38688 24696 0 u_ppwm/u_mem/_0211_
rlabel metal3 40512 29820 40512 29820 0 u_ppwm/u_mem/_0212_
rlabel metal2 43056 31164 43056 31164 0 u_ppwm/u_mem/_0213_
rlabel metal2 46176 26754 46176 26754 0 u_ppwm/u_mem/_0214_
rlabel metal3 44784 21588 44784 21588 0 u_ppwm/u_mem/_0215_
rlabel metal3 42864 20328 42864 20328 0 u_ppwm/u_mem/_0216_
rlabel metal2 39264 20202 39264 20202 0 u_ppwm/u_mem/_0217_
rlabel metal2 40512 24486 40512 24486 0 u_ppwm/u_mem/_0218_
rlabel metal3 41376 27720 41376 27720 0 u_ppwm/u_mem/_0219_
rlabel metal3 44592 30408 44592 30408 0 u_ppwm/u_mem/_0220_
rlabel metal2 47808 27888 47808 27888 0 u_ppwm/u_mem/_0221_
rlabel metal2 46560 24864 46560 24864 0 u_ppwm/u_mem/_0222_
rlabel metal2 41952 22344 41952 22344 0 u_ppwm/u_mem/_0223_
rlabel metal2 41184 22218 41184 22218 0 u_ppwm/u_mem/_0224_
rlabel metal2 40800 24318 40800 24318 0 u_ppwm/u_mem/_0225_
rlabel metal2 43728 25536 43728 25536 0 u_ppwm/u_mem/_0226_
rlabel metal2 45312 27090 45312 27090 0 u_ppwm/u_mem/_0227_
rlabel metal2 47760 22260 47760 22260 0 u_ppwm/u_mem/_0228_
rlabel metal2 43392 22386 43392 22386 0 u_ppwm/u_mem/_0229_
rlabel metal3 39024 19236 39024 19236 0 u_ppwm/u_mem/_0230_
rlabel metal2 40032 17724 40032 17724 0 u_ppwm/u_mem/_0231_
rlabel metal2 40128 24696 40128 24696 0 u_ppwm/u_mem/_0232_
rlabel metal2 42768 26292 42768 26292 0 u_ppwm/u_mem/_0233_
rlabel metal2 49056 28056 49056 28056 0 u_ppwm/u_mem/_0234_
rlabel metal2 48864 25074 48864 25074 0 u_ppwm/u_mem/_0235_
rlabel metal2 47808 21672 47808 21672 0 u_ppwm/u_mem/_0236_
rlabel metal3 38352 20076 38352 20076 0 u_ppwm/u_mem/_0237_
rlabel metal2 6672 17724 6672 17724 0 u_ppwm/u_mem/_0238_
rlabel metal2 8256 19194 8256 19194 0 u_ppwm/u_mem/_0239_
rlabel metal2 36192 25830 36192 25830 0 u_ppwm/u_mem/_0240_
rlabel metal3 25056 24612 25056 24612 0 u_ppwm/u_mem/_0241_
rlabel metal2 15744 26082 15744 26082 0 u_ppwm/u_mem/_0242_
rlabel metal2 6624 18228 6624 18228 0 u_ppwm/u_mem/_0243_
rlabel metal2 8352 18060 8352 18060 0 u_ppwm/u_mem/_0244_
rlabel metal2 6624 15498 6624 15498 0 u_ppwm/u_mem/_0245_
rlabel metal2 6528 14742 6528 14742 0 u_ppwm/u_mem/_0246_
rlabel metal2 7728 18564 7728 18564 0 u_ppwm/u_mem/_0247_
rlabel metal2 6912 18018 6912 18018 0 u_ppwm/u_mem/_0248_
rlabel metal2 7200 17010 7200 17010 0 u_ppwm/u_mem/_0249_
rlabel metal2 6816 18480 6816 18480 0 u_ppwm/u_mem/_0250_
rlabel metal2 16128 27552 16128 27552 0 u_ppwm/u_mem/_0251_
rlabel metal5 19248 26796 19248 26796 0 u_ppwm/u_mem/_0252_
rlabel metal2 16128 26208 16128 26208 0 u_ppwm/u_mem/_0253_
rlabel via1 16226 26124 16226 26124 0 u_ppwm/u_mem/_0254_
rlabel metal2 15264 26082 15264 26082 0 u_ppwm/u_mem/_0255_
rlabel metal3 15696 26124 15696 26124 0 u_ppwm/u_mem/_0256_
rlabel metal2 14976 24570 14976 24570 0 u_ppwm/u_mem/_0257_
rlabel metal2 15456 25536 15456 25536 0 u_ppwm/u_mem/_0258_
rlabel metal2 15744 25620 15744 25620 0 u_ppwm/u_mem/_0259_
rlabel metal2 24576 22176 24576 22176 0 u_ppwm/u_mem/_0260_
rlabel via2 23616 25286 23616 25286 0 u_ppwm/u_mem/_0261_
rlabel metal2 30000 26124 30000 26124 0 u_ppwm/u_mem/_0262_
rlabel metal2 29856 23772 29856 23772 0 u_ppwm/u_mem/_0263_
rlabel metal2 30144 24492 30144 24492 0 u_ppwm/u_mem/_0264_
rlabel metal2 30048 24696 30048 24696 0 u_ppwm/u_mem/_0265_
rlabel metal2 30384 24444 30384 24444 0 u_ppwm/u_mem/_0266_
rlabel metal2 15408 24612 15408 24612 0 u_ppwm/u_mem/_0267_
rlabel metal3 13440 26796 13440 26796 0 u_ppwm/u_mem/_0268_
rlabel metal2 16224 25368 16224 25368 0 u_ppwm/u_mem/_0269_
rlabel metal3 16032 24444 16032 24444 0 u_ppwm/u_mem/_0270_
rlabel metal3 16752 32760 16752 32760 0 u_ppwm/u_mem/_0271_
rlabel metal2 16656 25284 16656 25284 0 u_ppwm/u_mem/_0272_
rlabel metal2 21792 25032 21792 25032 0 u_ppwm/u_mem/_0273_
rlabel metal2 33600 23898 33600 23898 0 u_ppwm/u_mem/_0274_
rlabel metal3 35952 23772 35952 23772 0 u_ppwm/u_mem/_0275_
rlabel metal2 37440 29190 37440 29190 0 u_ppwm/u_mem/_0276_
rlabel metal3 37728 29148 37728 29148 0 u_ppwm/u_mem/_0277_
rlabel metal3 41328 22260 41328 22260 0 u_ppwm/u_mem/_0278_
rlabel metal2 37248 23352 37248 23352 0 u_ppwm/u_mem/_0279_
rlabel metal2 37920 20034 37920 20034 0 u_ppwm/u_mem/_0280_
rlabel metal2 37632 22596 37632 22596 0 u_ppwm/u_mem/_0281_
rlabel metal2 36576 24066 36576 24066 0 u_ppwm/u_mem/_0282_
rlabel metal3 12288 25242 12288 25242 0 u_ppwm/u_mem/_0283_
rlabel metal3 12816 25368 12816 25368 0 u_ppwm/u_mem/_0284_
rlabel metal2 15360 27090 15360 27090 0 u_ppwm/u_mem/_0285_
rlabel metal2 14747 26754 14747 26754 0 u_ppwm/u_mem/_0286_
rlabel metal2 13440 29148 13440 29148 0 u_ppwm/u_mem/_0287_
rlabel metal2 14496 27006 14496 27006 0 u_ppwm/u_mem/_0288_
rlabel metal2 14160 30996 14160 30996 0 u_ppwm/u_mem/_0289_
rlabel metal4 14784 26460 14784 26460 0 u_ppwm/u_mem/_0290_
rlabel metal3 17856 25662 17856 25662 0 u_ppwm/u_mem/_0291_
rlabel metal2 35808 25452 35808 25452 0 u_ppwm/u_mem/_0292_
rlabel metal3 37008 25284 37008 25284 0 u_ppwm/u_mem/_0293_
rlabel metal3 36912 32508 36912 32508 0 u_ppwm/u_mem/_0294_
rlabel metal2 36816 32172 36816 32172 0 u_ppwm/u_mem/_0295_
rlabel metal2 46320 24024 46320 24024 0 u_ppwm/u_mem/_0296_
rlabel metal2 37152 25410 37152 25410 0 u_ppwm/u_mem/_0297_
rlabel metal2 43104 22596 43104 22596 0 u_ppwm/u_mem/_0298_
rlabel metal2 43392 24318 43392 24318 0 u_ppwm/u_mem/_0299_
rlabel metal3 32640 25410 32640 25410 0 u_ppwm/u_mem/_0300_
rlabel metal2 8352 26712 8352 26712 0 u_ppwm/u_mem/_0301_
rlabel metal2 13824 26922 13824 26922 0 u_ppwm/u_mem/_0302_
rlabel metal2 14880 27510 14880 27510 0 u_ppwm/u_mem/_0303_
rlabel metal2 13981 26929 13981 26929 0 u_ppwm/u_mem/_0304_
rlabel metal2 12288 32592 12288 32592 0 u_ppwm/u_mem/_0305_
rlabel metal3 13392 30156 13392 30156 0 u_ppwm/u_mem/_0306_
rlabel metal2 12864 33642 12864 33642 0 u_ppwm/u_mem/_0307_
rlabel metal2 13536 26880 13536 26880 0 u_ppwm/u_mem/_0308_
rlabel metal4 13824 26376 13824 26376 0 u_ppwm/u_mem/_0309_
rlabel metal2 30624 27090 30624 27090 0 u_ppwm/u_mem/_0310_
rlabel metal2 31728 26124 31728 26124 0 u_ppwm/u_mem/_0311_
rlabel metal3 31104 26796 31104 26796 0 u_ppwm/u_mem/_0312_
rlabel metal2 30720 26376 30720 26376 0 u_ppwm/u_mem/_0313_
rlabel metal4 31296 25830 31296 25830 0 u_ppwm/u_mem/_0314_
rlabel metal2 30816 26405 30816 26405 0 u_ppwm/u_mem/_0315_
rlabel metal2 4224 25032 4224 25032 0 u_ppwm/u_mem/_0316_
rlabel metal3 13536 25578 13536 25578 0 u_ppwm/u_mem/_0317_
rlabel metal2 19968 26040 19968 26040 0 u_ppwm/u_mem/_0318_
rlabel metal2 17856 26166 17856 26166 0 u_ppwm/u_mem/_0319_
rlabel metal2 17184 26250 17184 26250 0 u_ppwm/u_mem/_0320_
rlabel metal2 17472 26124 17472 26124 0 u_ppwm/u_mem/_0321_
rlabel metal4 17664 26040 17664 26040 0 u_ppwm/u_mem/_0322_
rlabel metal2 37440 26208 37440 26208 0 u_ppwm/u_mem/_0323_
rlabel metal2 37344 26376 37344 26376 0 u_ppwm/u_mem/_0324_
rlabel metal2 29376 26040 29376 26040 0 u_ppwm/u_mem/_0325_
rlabel metal2 29184 26544 29184 26544 0 u_ppwm/u_mem/_0326_
rlabel metal3 30288 27636 30288 27636 0 u_ppwm/u_mem/_0327_
rlabel metal2 29664 27090 29664 27090 0 u_ppwm/u_mem/_0328_
rlabel metal2 27840 29988 27840 29988 0 u_ppwm/u_mem/_0329_
rlabel metal3 28128 26838 28128 26838 0 u_ppwm/u_mem/_0330_
rlabel metal2 28608 26373 28608 26373 0 u_ppwm/u_mem/_0331_
rlabel metal2 28992 26796 28992 26796 0 u_ppwm/u_mem/_0332_
rlabel metal2 5904 23268 5904 23268 0 u_ppwm/u_mem/_0333_
rlabel metal2 5520 23772 5520 23772 0 u_ppwm/u_mem/_0334_
rlabel metal2 16512 23478 16512 23478 0 u_ppwm/u_mem/_0335_
rlabel metal2 17472 23688 17472 23688 0 u_ppwm/u_mem/_0336_
rlabel metal2 17904 24024 17904 24024 0 u_ppwm/u_mem/_0337_
rlabel metal2 18240 24696 18240 24696 0 u_ppwm/u_mem/_0338_
rlabel metal3 6912 31164 6912 31164 0 u_ppwm/u_mem/_0339_
rlabel metal2 7872 24402 7872 24402 0 u_ppwm/u_mem/_0340_
rlabel metal3 19728 24612 19728 24612 0 u_ppwm/u_mem/_0341_
rlabel metal2 27072 26838 27072 26838 0 u_ppwm/u_mem/_0342_
rlabel metal2 27456 30324 27456 30324 0 u_ppwm/u_mem/_0343_
rlabel metal3 28032 26754 28032 26754 0 u_ppwm/u_mem/_0344_
rlabel metal2 27552 26586 27552 26586 0 u_ppwm/u_mem/_0345_
rlabel metal2 22176 26292 22176 26292 0 u_ppwm/u_mem/_0346_
rlabel metal2 21120 25242 21120 25242 0 u_ppwm/u_mem/_0347_
rlabel metal2 6240 27090 6240 27090 0 u_ppwm/u_mem/_0348_
rlabel metal2 13152 25830 13152 25830 0 u_ppwm/u_mem/_0349_
rlabel metal3 13872 30408 13872 30408 0 u_ppwm/u_mem/_0350_
rlabel metal2 13243 25368 13243 25368 0 u_ppwm/u_mem/_0351_
rlabel metal2 14112 25284 14112 25284 0 u_ppwm/u_mem/_0352_
rlabel metal2 8592 24612 8592 24612 0 u_ppwm/u_mem/_0353_
rlabel metal2 13440 25116 13440 25116 0 u_ppwm/u_mem/_0354_
rlabel metal3 14016 25284 14016 25284 0 u_ppwm/u_mem/_0355_
rlabel metal4 13728 25368 13728 25368 0 u_ppwm/u_mem/_0356_
rlabel metal2 26496 26754 26496 26754 0 u_ppwm/u_mem/_0357_
rlabel metal2 26208 30408 26208 30408 0 u_ppwm/u_mem/_0358_
rlabel metal2 26592 26376 26592 26376 0 u_ppwm/u_mem/_0359_
rlabel metal2 26592 25469 26592 25469 0 u_ppwm/u_mem/_0360_
rlabel metal3 28980 24654 28980 24654 0 u_ppwm/u_mem/_0361_
rlabel metal2 26928 24780 26928 24780 0 u_ppwm/u_mem/_0362_
rlabel metal2 38112 20916 38112 20916 0 u_ppwm/u_mem/_0363_
rlabel metal2 47424 21588 47424 21588 0 u_ppwm/u_mem/_0364_
rlabel metal2 48576 24864 48576 24864 0 u_ppwm/u_mem/_0365_
rlabel metal3 48240 28308 48240 28308 0 u_ppwm/u_mem/_0366_
rlabel metal2 43104 26796 43104 26796 0 u_ppwm/u_mem/_0367_
rlabel metal2 40992 26124 40992 26124 0 u_ppwm/u_mem/_0368_
rlabel metal2 40464 17724 40464 17724 0 u_ppwm/u_mem/_0369_
rlabel metal2 38448 19068 38448 19068 0 u_ppwm/u_mem/_0370_
rlabel metal3 43920 22260 43920 22260 0 u_ppwm/u_mem/_0371_
rlabel metal2 48096 22512 48096 22512 0 u_ppwm/u_mem/_0372_
rlabel metal2 51264 26418 51264 26418 0 u_ppwm/u_mem/_0373_
rlabel metal2 44544 25872 44544 25872 0 u_ppwm/u_mem/_0374_
rlabel metal3 41520 24612 41520 24612 0 u_ppwm/u_mem/_0375_
rlabel metal2 41520 22260 41520 22260 0 u_ppwm/u_mem/_0376_
rlabel metal2 40704 21588 40704 21588 0 u_ppwm/u_mem/_0377_
rlabel metal2 47040 22806 47040 22806 0 u_ppwm/u_mem/_0378_
rlabel metal2 47040 24990 47040 24990 0 u_ppwm/u_mem/_0379_
rlabel metal2 43872 29148 43872 29148 0 u_ppwm/u_mem/_0380_
rlabel metal2 42528 29316 42528 29316 0 u_ppwm/u_mem/_0381_
rlabel metal2 39072 26376 39072 26376 0 u_ppwm/u_mem/_0382_
rlabel metal2 39264 22344 39264 22344 0 u_ppwm/u_mem/_0383_
rlabel metal3 42096 19236 42096 19236 0 u_ppwm/u_mem/_0384_
rlabel metal2 44592 21588 44592 21588 0 u_ppwm/u_mem/_0385_
rlabel metal2 45600 22596 45600 22596 0 u_ppwm/u_mem/_0386_
rlabel metal3 43536 28308 43536 28308 0 u_ppwm/u_mem/_0387_
rlabel metal2 41088 29820 41088 29820 0 u_ppwm/u_mem/_0388_
rlabel metal2 38304 26166 38304 26166 0 u_ppwm/u_mem/_0389_
rlabel metal2 34176 23856 34176 23856 0 u_ppwm/u_mem/_0390_
rlabel metal2 32640 22008 32640 22008 0 u_ppwm/u_mem/_0391_
rlabel metal2 35520 26376 35520 26376 0 u_ppwm/u_mem/_0392_
rlabel metal2 33600 27804 33600 27804 0 u_ppwm/u_mem/_0393_
rlabel metal2 33216 30240 33216 30240 0 u_ppwm/u_mem/_0394_
rlabel metal2 27264 30702 27264 30702 0 u_ppwm/u_mem/_0395_
rlabel metal2 24960 29064 24960 29064 0 u_ppwm/u_mem/_0396_
rlabel metal2 24672 25956 24672 25956 0 u_ppwm/u_mem/_0397_
rlabel metal2 31392 21588 31392 21588 0 u_ppwm/u_mem/_0398_
rlabel metal3 31824 23772 31824 23772 0 u_ppwm/u_mem/_0399_
rlabel metal2 31872 28308 31872 28308 0 u_ppwm/u_mem/_0400_
rlabel metal3 27888 29148 27888 29148 0 u_ppwm/u_mem/_0401_
rlabel metal2 22320 29820 22320 29820 0 u_ppwm/u_mem/_0402_
rlabel metal2 22944 29148 22944 29148 0 u_ppwm/u_mem/_0403_
rlabel metal2 32256 31164 32256 31164 0 u_ppwm/u_mem/_0404_
rlabel metal2 36960 30240 36960 30240 0 u_ppwm/u_mem/_0405_
rlabel metal3 37968 30660 37968 30660 0 u_ppwm/u_mem/_0406_
rlabel metal2 34176 32886 34176 32886 0 u_ppwm/u_mem/_0407_
rlabel metal2 31968 32592 31968 32592 0 u_ppwm/u_mem/_0408_
rlabel metal2 29664 31374 29664 31374 0 u_ppwm/u_mem/_0409_
rlabel metal3 26880 32172 26880 32172 0 u_ppwm/u_mem/_0410_
rlabel metal2 25248 30072 25248 30072 0 u_ppwm/u_mem/_0411_
rlabel metal2 34992 29820 34992 29820 0 u_ppwm/u_mem/_0412_
rlabel metal2 36384 32340 36384 32340 0 u_ppwm/u_mem/_0413_
rlabel metal2 35424 30660 35424 30660 0 u_ppwm/u_mem/_0414_
rlabel metal2 32352 33600 32352 33600 0 u_ppwm/u_mem/_0415_
rlabel metal3 30096 33684 30096 33684 0 u_ppwm/u_mem/_0416_
rlabel metal2 26064 32844 26064 32844 0 u_ppwm/u_mem/_0417_
rlabel metal2 23808 33054 23808 33054 0 u_ppwm/u_mem/_0418_
rlabel metal2 21984 33684 21984 33684 0 u_ppwm/u_mem/_0419_
rlabel metal2 17088 35238 17088 35238 0 u_ppwm/u_mem/_0420_
rlabel metal2 11520 35994 11520 35994 0 u_ppwm/u_mem/_0421_
rlabel metal3 7920 35784 7920 35784 0 u_ppwm/u_mem/_0422_
rlabel metal3 4032 34356 4032 34356 0 u_ppwm/u_mem/_0423_
rlabel metal3 4320 33684 4320 33684 0 u_ppwm/u_mem/_0424_
rlabel metal2 18144 32886 18144 32886 0 u_ppwm/u_mem/_0425_
rlabel metal3 19344 34356 19344 34356 0 u_ppwm/u_mem/_0426_
rlabel metal3 16176 36708 16176 36708 0 u_ppwm/u_mem/_0427_
rlabel metal2 11568 38220 11568 38220 0 u_ppwm/u_mem/_0428_
rlabel metal3 8880 35868 8880 35868 0 u_ppwm/u_mem/_0429_
rlabel metal2 6720 34356 6720 34356 0 u_ppwm/u_mem/_0430_
rlabel metal2 4512 30828 4512 30828 0 u_ppwm/u_mem/_0431_
rlabel metal2 11040 30912 11040 30912 0 u_ppwm/u_mem/_0432_
rlabel metal2 15744 31332 15744 31332 0 u_ppwm/u_mem/_0433_
rlabel metal2 15120 31332 15120 31332 0 u_ppwm/u_mem/_0434_
rlabel metal2 11904 33432 11904 33432 0 u_ppwm/u_mem/_0435_
rlabel metal3 7584 34398 7584 34398 0 u_ppwm/u_mem/_0436_
rlabel metal3 4224 32844 4224 32844 0 u_ppwm/u_mem/_0437_
rlabel metal2 4992 29820 4992 29820 0 u_ppwm/u_mem/_0438_
rlabel metal2 6096 29820 6096 29820 0 u_ppwm/u_mem/_0439_
rlabel metal3 13392 30828 13392 30828 0 u_ppwm/u_mem/_0440_
rlabel metal2 13824 31752 13824 31752 0 u_ppwm/u_mem/_0441_
rlabel metal2 11280 32844 11280 32844 0 u_ppwm/u_mem/_0442_
rlabel metal3 7584 32172 7584 32172 0 u_ppwm/u_mem/_0443_
rlabel metal2 5616 32844 5616 32844 0 u_ppwm/u_mem/_0444_
rlabel metal2 4128 29316 4128 29316 0 u_ppwm/u_mem/_0445_
rlabel metal2 5760 27342 5760 27342 0 u_ppwm/u_mem/_0446_
rlabel metal2 8160 27216 8160 27216 0 u_ppwm/u_mem/_0447_
rlabel metal3 8448 29820 8448 29820 0 u_ppwm/u_mem/_0448_
rlabel metal3 17952 29148 17952 29148 0 u_ppwm/u_mem/_0449_
rlabel metal2 17376 27552 17376 27552 0 u_ppwm/u_mem/_0450_
rlabel metal2 17904 25284 17904 25284 0 u_ppwm/u_mem/_0451_
rlabel metal2 14064 23772 14064 23772 0 u_ppwm/u_mem/_0452_
rlabel metal3 11376 25284 11376 25284 0 u_ppwm/u_mem/_0453_
rlabel metal3 9792 26796 9792 26796 0 u_ppwm/u_mem/_0454_
rlabel metal2 12480 26712 12480 26712 0 u_ppwm/u_mem/_0455_
rlabel metal2 19584 29232 19584 29232 0 u_ppwm/u_mem/_0456_
rlabel metal2 18912 26586 18912 26586 0 u_ppwm/u_mem/_0457_
rlabel metal2 17856 23100 17856 23100 0 u_ppwm/u_mem/_0458_
rlabel metal2 17424 22260 17424 22260 0 u_ppwm/u_mem/_0459_
rlabel metal2 14928 22260 14928 22260 0 u_ppwm/u_mem/_0460_
rlabel metal2 11520 19656 11520 19656 0 u_ppwm/u_mem/_0461_
rlabel metal2 9120 21168 9120 21168 0 u_ppwm/u_mem/_0462_
rlabel metal2 6240 24864 6240 24864 0 u_ppwm/u_mem/_0463_
rlabel metal2 1920 25662 1920 25662 0 u_ppwm/u_mem/_0464_
rlabel metal2 4608 24192 4608 24192 0 u_ppwm/u_mem/_0465_
rlabel metal2 5136 21588 5136 21588 0 u_ppwm/u_mem/_0466_
rlabel metal2 6720 21504 6720 21504 0 u_ppwm/u_mem/_0467_
rlabel metal3 10992 20748 10992 20748 0 u_ppwm/u_mem/_0468_
rlabel metal2 9024 23184 9024 23184 0 u_ppwm/u_mem/_0469_
rlabel metal2 6672 24780 6672 24780 0 u_ppwm/u_mem/_0470_
rlabel metal3 4032 26796 4032 26796 0 u_ppwm/u_mem/_0471_
rlabel metal3 4176 22260 4176 22260 0 u_ppwm/u_mem/_0472_
rlabel metal2 4704 21126 4704 21126 0 u_ppwm/u_mem/_0473_
rlabel metal2 6432 19236 6432 19236 0 u_ppwm/u_mem/_0474_
rlabel metal2 7488 17598 7488 17598 0 u_ppwm/u_mem/_0475_
rlabel metal2 2016 17388 2016 17388 0 u_ppwm/u_mem/_0476_
rlabel metal2 2976 19194 2976 19194 0 u_ppwm/u_mem/_0477_
rlabel metal2 4032 20034 4032 20034 0 u_ppwm/u_mem/_0478_
rlabel metal2 2208 16254 2208 16254 0 u_ppwm/u_mem/_0479_
rlabel metal2 2304 17640 2304 17640 0 u_ppwm/u_mem/_0480_
rlabel metal2 5760 17052 5760 17052 0 u_ppwm/u_mem/_0481_
rlabel metal2 1344 15162 1344 15162 0 u_ppwm/u_mem/_0482_
rlabel metal3 4896 16170 4896 16170 0 u_ppwm/u_mem/_0483_
rlabel metal2 1632 15456 1632 15456 0 u_ppwm/u_mem/_0484_
rlabel metal3 5760 14070 5760 14070 0 u_ppwm/u_mem/_0485_
rlabel metal2 5088 16002 5088 16002 0 u_ppwm/u_mem/_0486_
rlabel metal2 3936 15834 3936 15834 0 u_ppwm/u_mem/_0487_
rlabel metal2 5472 15288 5472 15288 0 u_ppwm/u_mem/_0488_
rlabel metal3 6864 15708 6864 15708 0 u_ppwm/u_mem/_0489_
rlabel metal3 8160 15708 8160 15708 0 u_ppwm/u_mem/_0490_
rlabel metal2 4704 19278 4704 19278 0 u_ppwm/u_mem/bit_count\[0\]
rlabel metal3 4224 17808 4224 17808 0 u_ppwm/u_mem/bit_count\[1\]
rlabel metal2 3744 17472 3744 17472 0 u_ppwm/u_mem/bit_count\[2\]
rlabel metal2 3552 15120 3552 15120 0 u_ppwm/u_mem/bit_count\[3\]
rlabel metal3 6768 14868 6768 14868 0 u_ppwm/u_mem/bit_count\[4\]
rlabel metal2 4800 15036 4800 15036 0 u_ppwm/u_mem/bit_count\[5\]
rlabel metal3 9984 15708 9984 15708 0 u_ppwm/u_mem/bit_count\[6\]
rlabel metal2 39072 21168 39072 21168 0 u_ppwm/u_mem/memory\[0\]
rlabel metal2 10272 24780 10272 24780 0 u_ppwm/u_mem/memory\[100\]
rlabel metal2 5376 25830 5376 25830 0 u_ppwm/u_mem/memory\[101\]
rlabel metal2 3792 24612 3792 24612 0 u_ppwm/u_mem/memory\[102\]
rlabel metal2 4992 22890 4992 22890 0 u_ppwm/u_mem/memory\[103\]
rlabel metal3 7584 21504 7584 21504 0 u_ppwm/u_mem/memory\[104\]
rlabel metal2 13920 21588 13920 21588 0 u_ppwm/u_mem/memory\[105\]
rlabel metal2 11904 23436 11904 23436 0 u_ppwm/u_mem/memory\[106\]
rlabel metal2 9024 24654 9024 24654 0 u_ppwm/u_mem/memory\[107\]
rlabel metal3 51456 27048 51456 27048 0 u_ppwm/u_mem/memory\[10\]
rlabel metal2 47424 26250 47424 26250 0 u_ppwm/u_mem/memory\[11\]
rlabel metal3 41952 26250 41952 26250 0 u_ppwm/u_mem/memory\[12\]
rlabel metal3 42672 23772 42672 23772 0 u_ppwm/u_mem/memory\[13\]
rlabel metal3 41136 21000 41136 21000 0 u_ppwm/u_mem/memory\[14\]
rlabel metal2 47616 23688 47616 23688 0 u_ppwm/u_mem/memory\[15\]
rlabel metal2 50784 25830 50784 25830 0 u_ppwm/u_mem/memory\[16\]
rlabel metal2 49104 29148 49104 29148 0 u_ppwm/u_mem/memory\[17\]
rlabel metal2 42720 29778 42720 29778 0 u_ppwm/u_mem/memory\[18\]
rlabel metal2 40992 27888 40992 27888 0 u_ppwm/u_mem/memory\[19\]
rlabel metal3 39168 19950 39168 19950 0 u_ppwm/u_mem/memory\[1\]
rlabel metal2 39744 22596 39744 22596 0 u_ppwm/u_mem/memory\[20\]
rlabel metal3 40560 20580 40560 20580 0 u_ppwm/u_mem/memory\[21\]
rlabel metal2 44928 20958 44928 20958 0 u_ppwm/u_mem/memory\[22\]
rlabel metal2 47184 22260 47184 22260 0 u_ppwm/u_mem/memory\[23\]
rlabel metal2 46512 29652 46512 29652 0 u_ppwm/u_mem/memory\[24\]
rlabel metal3 42480 29064 42480 29064 0 u_ppwm/u_mem/memory\[25\]
rlabel metal2 39360 27972 39360 27972 0 u_ppwm/u_mem/memory\[26\]
rlabel metal2 37344 23310 37344 23310 0 u_ppwm/u_mem/memory\[27\]
rlabel metal2 35520 23436 35520 23436 0 u_ppwm/u_mem/memory\[28\]
rlabel metal2 35856 24612 35856 24612 0 u_ppwm/u_mem/memory\[29\]
rlabel metal2 50496 23814 50496 23814 0 u_ppwm/u_mem/memory\[2\]
rlabel metal3 35232 27468 35232 27468 0 u_ppwm/u_mem/memory\[30\]
rlabel metal2 34272 29568 34272 29568 0 u_ppwm/u_mem/memory\[31\]
rlabel metal2 29856 30324 29856 30324 0 u_ppwm/u_mem/memory\[32\]
rlabel metal3 26304 29148 26304 29148 0 u_ppwm/u_mem/memory\[33\]
rlabel metal2 26016 26544 26016 26544 0 u_ppwm/u_mem/memory\[34\]
rlabel metal2 30336 23016 30336 23016 0 u_ppwm/u_mem/memory\[35\]
rlabel metal3 33312 23268 33312 23268 0 u_ppwm/u_mem/memory\[36\]
rlabel metal3 33216 27048 33216 27048 0 u_ppwm/u_mem/memory\[37\]
rlabel metal2 31296 28350 31296 28350 0 u_ppwm/u_mem/memory\[38\]
rlabel metal2 23808 30324 23808 30324 0 u_ppwm/u_mem/memory\[39\]
rlabel metal2 50304 27636 50304 27636 0 u_ppwm/u_mem/memory\[3\]
rlabel metal3 25440 29652 25440 29652 0 u_ppwm/u_mem/memory\[40\]
rlabel metal2 32736 29652 32736 29652 0 u_ppwm/u_mem/memory\[41\]
rlabel metal2 36768 29568 36768 29568 0 u_ppwm/u_mem/memory\[42\]
rlabel metal3 40080 31164 40080 31164 0 u_ppwm/u_mem/memory\[43\]
rlabel metal2 37824 34104 37824 34104 0 u_ppwm/u_mem/memory\[44\]
rlabel metal2 34944 33390 34944 33390 0 u_ppwm/u_mem/memory\[45\]
rlabel metal3 31632 32928 31632 32928 0 u_ppwm/u_mem/memory\[46\]
rlabel metal2 29664 32550 29664 32550 0 u_ppwm/u_mem/memory\[47\]
rlabel metal2 26016 31584 26016 31584 0 u_ppwm/u_mem/memory\[48\]
rlabel metal2 34464 29232 34464 29232 0 u_ppwm/u_mem/memory\[49\]
rlabel metal2 47712 27006 47712 27006 0 u_ppwm/u_mem/memory\[4\]
rlabel via2 38208 32004 38208 32004 0 u_ppwm/u_mem/memory\[50\]
rlabel metal2 37344 34524 37344 34524 0 u_ppwm/u_mem/memory\[51\]
rlabel metal2 35040 33516 35040 33516 0 u_ppwm/u_mem/memory\[52\]
rlabel metal3 31920 34608 31920 34608 0 u_ppwm/u_mem/memory\[53\]
rlabel metal2 29088 34188 29088 34188 0 u_ppwm/u_mem/memory\[54\]
rlabel metal3 26160 33600 26160 33600 0 u_ppwm/u_mem/memory\[55\]
rlabel metal2 23760 34188 23760 34188 0 u_ppwm/u_mem/memory\[56\]
rlabel metal2 17760 34314 17760 34314 0 u_ppwm/u_mem/memory\[57\]
rlabel metal2 14976 35784 14976 35784 0 u_ppwm/u_mem/memory\[58\]
rlabel metal2 10656 36666 10656 36666 0 u_ppwm/u_mem/memory\[59\]
rlabel metal2 42720 25662 42720 25662 0 u_ppwm/u_mem/memory\[5\]
rlabel metal3 6576 35700 6576 35700 0 u_ppwm/u_mem/memory\[60\]
rlabel metal3 4032 31920 4032 31920 0 u_ppwm/u_mem/memory\[61\]
rlabel metal2 13824 32634 13824 32634 0 u_ppwm/u_mem/memory\[62\]
rlabel metal2 21360 33852 21360 33852 0 u_ppwm/u_mem/memory\[63\]
rlabel metal2 17568 35238 17568 35238 0 u_ppwm/u_mem/memory\[64\]
rlabel metal2 14016 37296 14016 37296 0 u_ppwm/u_mem/memory\[65\]
rlabel metal2 9888 37002 9888 37002 0 u_ppwm/u_mem/memory\[66\]
rlabel metal3 7200 35112 7200 35112 0 u_ppwm/u_mem/memory\[67\]
rlabel metal2 4896 31374 4896 31374 0 u_ppwm/u_mem/memory\[68\]
rlabel metal2 12672 31206 12672 31206 0 u_ppwm/u_mem/memory\[69\]
rlabel metal2 40512 18984 40512 18984 0 u_ppwm/u_mem/memory\[6\]
rlabel metal3 17184 30828 17184 30828 0 u_ppwm/u_mem/memory\[70\]
rlabel metal2 17280 33222 17280 33222 0 u_ppwm/u_mem/memory\[71\]
rlabel metal3 13920 33852 13920 33852 0 u_ppwm/u_mem/memory\[72\]
rlabel metal2 10176 34650 10176 34650 0 u_ppwm/u_mem/memory\[73\]
rlabel metal2 5472 33852 5472 33852 0 u_ppwm/u_mem/memory\[74\]
rlabel metal2 4608 30366 4608 30366 0 u_ppwm/u_mem/memory\[75\]
rlabel metal3 6480 29064 6480 29064 0 u_ppwm/u_mem/memory\[76\]
rlabel metal2 13440 30156 13440 30156 0 u_ppwm/u_mem/memory\[77\]
rlabel metal3 15360 32172 15360 32172 0 u_ppwm/u_mem/memory\[78\]
rlabel metal2 12384 31542 12384 31542 0 u_ppwm/u_mem/memory\[79\]
rlabel metal3 40704 18312 40704 18312 0 u_ppwm/u_mem/memory\[7\]
rlabel metal2 10368 32886 10368 32886 0 u_ppwm/u_mem/memory\[80\]
rlabel metal2 6096 34356 6096 34356 0 u_ppwm/u_mem/memory\[81\]
rlabel metal2 4320 29778 4320 29778 0 u_ppwm/u_mem/memory\[82\]
rlabel metal2 4800 27930 4800 27930 0 u_ppwm/u_mem/memory\[83\]
rlabel metal2 8544 27846 8544 27846 0 u_ppwm/u_mem/memory\[84\]
rlabel metal2 11520 28266 11520 28266 0 u_ppwm/u_mem/memory\[85\]
rlabel metal2 17664 29274 17664 29274 0 u_ppwm/u_mem/memory\[86\]
rlabel metal2 17856 29064 17856 29064 0 u_ppwm/u_mem/memory\[87\]
rlabel metal3 18816 26124 18816 26124 0 u_ppwm/u_mem/memory\[88\]
rlabel metal2 17088 23982 17088 23982 0 u_ppwm/u_mem/memory\[89\]
rlabel metal2 38976 19782 38976 19782 0 u_ppwm/u_mem/memory\[8\]
rlabel metal2 13920 25200 13920 25200 0 u_ppwm/u_mem/memory\[90\]
rlabel metal2 11232 26502 11232 26502 0 u_ppwm/u_mem/memory\[91\]
rlabel metal2 10944 27678 10944 27678 0 u_ppwm/u_mem/memory\[92\]
rlabel metal2 19440 29148 19440 29148 0 u_ppwm/u_mem/memory\[93\]
rlabel metal2 18720 26922 18720 26922 0 u_ppwm/u_mem/memory\[94\]
rlabel metal2 17568 23236 17568 23236 0 u_ppwm/u_mem/memory\[95\]
rlabel metal2 19008 22764 19008 22764 0 u_ppwm/u_mem/memory\[96\]
rlabel metal2 15648 23184 15648 23184 0 u_ppwm/u_mem/memory\[97\]
rlabel metal2 13440 19950 13440 19950 0 u_ppwm/u_mem/memory\[98\]
rlabel metal2 11808 21924 11808 21924 0 u_ppwm/u_mem/memory\[99\]
rlabel metal2 49056 22176 49056 22176 0 u_ppwm/u_mem/memory\[9\]
rlabel metal2 11136 18270 11136 18270 0 u_ppwm/u_mem/state_q\[0\]
rlabel metal2 21552 19824 21552 19824 0 u_ppwm/u_mem/state_q\[2\]
rlabel metal2 12960 12558 12960 12558 0 u_ppwm/u_pwm/_000_
rlabel metal2 12576 13440 12576 13440 0 u_ppwm/u_pwm/_001_
rlabel metal2 11424 13020 11424 13020 0 u_ppwm/u_pwm/_002_
rlabel metal3 12672 11508 12672 11508 0 u_ppwm/u_pwm/_003_
rlabel metal2 12960 4200 12960 4200 0 u_ppwm/u_pwm/_004_
rlabel metal2 11328 3528 11328 3528 0 u_ppwm/u_pwm/_005_
rlabel metal2 7392 3906 7392 3906 0 u_ppwm/u_pwm/_006_
rlabel metal2 8160 3780 8160 3780 0 u_ppwm/u_pwm/_007_
rlabel metal3 10656 6636 10656 6636 0 u_ppwm/u_pwm/_008_
rlabel metal2 11424 9492 11424 9492 0 u_ppwm/u_pwm/_009_
rlabel metal2 5664 12558 5664 12558 0 u_ppwm/u_pwm/_010_
rlabel metal2 4560 11508 4560 11508 0 u_ppwm/u_pwm/_011_
rlabel metal2 5760 9408 5760 9408 0 u_ppwm/u_pwm/_012_
rlabel metal2 1536 10500 1536 10500 0 u_ppwm/u_pwm/_013_
rlabel metal2 1056 8946 1056 8946 0 u_ppwm/u_pwm/_014_
rlabel metal2 2496 7896 2496 7896 0 u_ppwm/u_pwm/_015_
rlabel metal2 1728 5628 1728 5628 0 u_ppwm/u_pwm/_016_
rlabel metal2 3648 6090 3648 6090 0 u_ppwm/u_pwm/_017_
rlabel metal2 5808 6300 5808 6300 0 u_ppwm/u_pwm/_018_
rlabel metal2 4128 8736 4128 8736 0 u_ppwm/u_pwm/_019_
rlabel metal3 8448 11928 8448 11928 0 u_ppwm/u_pwm/_020_
rlabel metal3 11424 8064 11424 8064 0 u_ppwm/u_pwm/_021_
rlabel metal3 3216 8820 3216 8820 0 u_ppwm/u_pwm/_022_
rlabel metal2 1344 8442 1344 8442 0 u_ppwm/u_pwm/_023_
rlabel metal2 1920 9450 1920 9450 0 u_ppwm/u_pwm/_024_
rlabel metal2 1584 8148 1584 8148 0 u_ppwm/u_pwm/_025_
rlabel metal2 1248 7644 1248 7644 0 u_ppwm/u_pwm/_026_
rlabel metal2 2400 6426 2400 6426 0 u_ppwm/u_pwm/_027_
rlabel metal2 4800 5082 4800 5082 0 u_ppwm/u_pwm/_028_
rlabel metal3 4656 5460 4656 5460 0 u_ppwm/u_pwm/_029_
rlabel metal3 4464 5040 4464 5040 0 u_ppwm/u_pwm/_030_
rlabel metal3 5136 7980 5136 7980 0 u_ppwm/u_pwm/_031_
rlabel metal2 5808 6468 5808 6468 0 u_ppwm/u_pwm/_032_
rlabel metal2 8304 8148 8304 8148 0 u_ppwm/u_pwm/_033_
rlabel metal2 5712 8148 5712 8148 0 u_ppwm/u_pwm/_034_
rlabel metal2 7200 9576 7200 9576 0 u_ppwm/u_pwm/_035_
rlabel metal2 7296 9408 7296 9408 0 u_ppwm/u_pwm/_036_
rlabel metal2 9168 11004 9168 11004 0 u_ppwm/u_pwm/_037_
rlabel metal3 8832 11424 8832 11424 0 u_ppwm/u_pwm/_038_
rlabel metal2 9552 10416 9552 10416 0 u_ppwm/u_pwm/_039_
rlabel metal2 10080 10878 10080 10878 0 u_ppwm/u_pwm/_040_
rlabel metal2 7776 11046 7776 11046 0 u_ppwm/u_pwm/_041_
rlabel metal3 9024 11676 9024 11676 0 u_ppwm/u_pwm/_042_
rlabel metal2 9216 11424 9216 11424 0 u_ppwm/u_pwm/_043_
rlabel metal2 9696 11718 9696 11718 0 u_ppwm/u_pwm/_044_
rlabel metal3 8736 11508 8736 11508 0 u_ppwm/u_pwm/_045_
rlabel metal2 9696 10920 9696 10920 0 u_ppwm/u_pwm/_046_
rlabel metal2 7872 11088 7872 11088 0 u_ppwm/u_pwm/_047_
rlabel metal2 9024 5712 9024 5712 0 u_ppwm/u_pwm/_048_
rlabel metal3 7824 5460 7824 5460 0 u_ppwm/u_pwm/_049_
rlabel metal2 8352 5964 8352 5964 0 u_ppwm/u_pwm/_050_
rlabel metal2 9312 5922 9312 5922 0 u_ppwm/u_pwm/_051_
rlabel metal2 8256 5880 8256 5880 0 u_ppwm/u_pwm/_052_
rlabel metal3 8786 5628 8786 5628 0 u_ppwm/u_pwm/_053_
rlabel metal2 8592 4956 8592 4956 0 u_ppwm/u_pwm/_054_
rlabel metal2 9504 4578 9504 4578 0 u_ppwm/u_pwm/_055_
rlabel metal2 8928 3402 8928 3402 0 u_ppwm/u_pwm/_056_
rlabel metal3 8976 4956 8976 4956 0 u_ppwm/u_pwm/_057_
rlabel metal3 9648 4872 9648 4872 0 u_ppwm/u_pwm/_058_
rlabel metal2 9072 3444 9072 3444 0 u_ppwm/u_pwm/_059_
rlabel metal2 8784 5124 8784 5124 0 u_ppwm/u_pwm/_060_
rlabel metal2 8928 5586 8928 5586 0 u_ppwm/u_pwm/_061_
rlabel metal2 8256 6384 8256 6384 0 u_ppwm/u_pwm/_062_
rlabel metal2 9024 7266 9024 7266 0 u_ppwm/u_pwm/_063_
rlabel metal3 9504 7140 9504 7140 0 u_ppwm/u_pwm/_064_
rlabel metal2 9216 7182 9216 7182 0 u_ppwm/u_pwm/_065_
rlabel metal3 8784 6468 8784 6468 0 u_ppwm/u_pwm/_066_
rlabel metal2 10176 7392 10176 7392 0 u_ppwm/u_pwm/_067_
rlabel metal2 9696 8106 9696 8106 0 u_ppwm/u_pwm/_068_
rlabel metal3 10272 7980 10272 7980 0 u_ppwm/u_pwm/_069_
rlabel metal2 10800 7980 10800 7980 0 u_ppwm/u_pwm/_070_
rlabel metal2 10944 7896 10944 7896 0 u_ppwm/u_pwm/_071_
rlabel metal2 5568 6636 5568 6636 0 u_ppwm/u_pwm/_072_
rlabel metal2 11616 8610 11616 8610 0 u_ppwm/u_pwm/_073_
rlabel metal3 9456 6300 9456 6300 0 u_ppwm/u_pwm/_074_
rlabel metal2 8064 3696 8064 3696 0 u_ppwm/u_pwm/_075_
rlabel metal3 7392 2604 7392 2604 0 u_ppwm/u_pwm/_076_
rlabel metal2 9984 4872 9984 4872 0 u_ppwm/u_pwm/_077_
rlabel metal3 13488 4116 13488 4116 0 u_ppwm/u_pwm/_078_
rlabel metal3 12816 10164 12816 10164 0 u_ppwm/u_pwm/_079_
rlabel metal3 10416 11676 10416 11676 0 u_ppwm/u_pwm/_080_
rlabel metal2 12480 13524 12480 13524 0 u_ppwm/u_pwm/_081_
rlabel metal2 12912 11928 12912 11928 0 u_ppwm/u_pwm/_082_
rlabel metal2 864 7938 864 7938 0 u_ppwm/u_pwm/_083_
rlabel metal2 7968 9324 7968 9324 0 u_ppwm/u_pwm/_084_
rlabel metal2 8688 6300 8688 6300 0 u_ppwm/u_pwm/_085_
rlabel metal2 7680 8736 7680 8736 0 u_ppwm/u_pwm/_086_
rlabel metal2 8256 8568 8256 8568 0 u_ppwm/u_pwm/_087_
rlabel metal2 14112 11760 14112 11760 0 u_ppwm/u_pwm/_088_
rlabel metal2 12672 13860 12672 13860 0 u_ppwm/u_pwm/_089_
rlabel metal2 10176 11718 10176 11718 0 u_ppwm/u_pwm/_090_
rlabel metal2 11808 11844 11808 11844 0 u_ppwm/u_pwm/_091_
rlabel metal3 12480 4116 12480 4116 0 u_ppwm/u_pwm/_092_
rlabel metal2 10272 4116 10272 4116 0 u_ppwm/u_pwm/_093_
rlabel metal2 11424 3318 11424 3318 0 u_ppwm/u_pwm/_094_
rlabel metal2 8256 3486 8256 3486 0 u_ppwm/u_pwm/_095_
rlabel metal2 11904 6048 11904 6048 0 u_ppwm/u_pwm/_096_
rlabel metal2 10752 9282 10752 9282 0 u_ppwm/u_pwm/_097_
rlabel metal2 4512 11802 4512 11802 0 u_ppwm/u_pwm/_098_
rlabel metal3 4608 13188 4608 13188 0 u_ppwm/u_pwm/_099_
rlabel metal2 4272 11676 4272 11676 0 u_ppwm/u_pwm/_100_
rlabel metal2 4704 11760 4704 11760 0 u_ppwm/u_pwm/_101_
rlabel metal2 3648 11088 3648 11088 0 u_ppwm/u_pwm/_102_
rlabel metal3 14592 13356 14592 13356 0 u_ppwm/u_pwm/cmp_value\[0\]
rlabel metal3 10128 14196 10128 14196 0 u_ppwm/u_pwm/cmp_value\[1\]
rlabel metal3 8592 12516 8592 12516 0 u_ppwm/u_pwm/cmp_value\[2\]
rlabel metal2 12144 11676 12144 11676 0 u_ppwm/u_pwm/cmp_value\[3\]
rlabel metal3 14400 3612 14400 3612 0 u_ppwm/u_pwm/cmp_value\[4\]
rlabel metal2 9216 3150 9216 3150 0 u_ppwm/u_pwm/cmp_value\[5\]
rlabel metal2 7632 4956 7632 4956 0 u_ppwm/u_pwm/cmp_value\[6\]
rlabel metal2 8784 4116 8784 4116 0 u_ppwm/u_pwm/cmp_value\[7\]
rlabel metal2 12864 6888 12864 6888 0 u_ppwm/u_pwm/cmp_value\[8\]
rlabel metal2 12672 9912 12672 9912 0 u_ppwm/u_pwm/cmp_value\[9\]
rlabel metal2 8064 12852 8064 12852 0 u_ppwm/u_pwm/counter\[0\]
rlabel metal2 5568 12096 5568 12096 0 u_ppwm/u_pwm/counter\[1\]
rlabel metal3 7248 10416 7248 10416 0 u_ppwm/u_pwm/counter\[2\]
rlabel metal2 7776 11676 7776 11676 0 u_ppwm/u_pwm/counter\[3\]
rlabel metal2 1440 8022 1440 8022 0 u_ppwm/u_pwm/counter\[4\]
rlabel metal2 9696 5502 9696 5502 0 u_ppwm/u_pwm/counter\[5\]
rlabel metal2 7488 6552 7488 6552 0 u_ppwm/u_pwm/counter\[6\]
rlabel metal2 6624 6384 6624 6384 0 u_ppwm/u_pwm/counter\[7\]
rlabel metal2 9120 7770 9120 7770 0 u_ppwm/u_pwm/counter\[8\]
rlabel metal3 8352 8148 8352 8148 0 u_ppwm/u_pwm/counter\[9\]
rlabel metal3 366 22428 366 22428 0 ui_in[0]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
