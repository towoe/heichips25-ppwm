* NGSPICE file created from heichips25_ppwm.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

.subckt heichips25_ppwm VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_28_907 VPWR VGND sg13g2_decap_8
XFILLER_36_951 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__627_ hold306/A net325 u_ppwm_u_ex__636_/A VPWR VGND sg13g2_and2_1
XFILLER_23_623 VPWR VGND sg13g2_decap_8
XFILLER_35_1009 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__558_ u_ppwm_u_ex__560_/C u_ppwm_u_ex__558_/B u_ppwm_u_ex__558_/C u_ppwm_u_ex__558_/Y
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_ex__489_ net631 VPWR u_ppwm_u_ex__489_/Y VGND u_ppwm_u_ex__487_/Y u_ppwm_u_ex__488_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__1163__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_2_527 VPWR VGND sg13g2_decap_8
XFILLER_19_929 VPWR VGND sg13g2_decap_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_26_461 VPWR VGND sg13g2_decap_8
XFILLER_42_965 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_8
XFILLER_41_486 VPWR VGND sg13g2_fill_1
XFILLER_6_811 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__182_ net626 u_ppwm_u_pwm__182_/C net580 u_ppwm_u_pwm__185_/B VPWR VGND
+ sg13g2_nand3_1
XFILLER_6_888 VPWR VGND sg13g2_decap_8
XFILLER_5_332 VPWR VGND sg13g2_decap_8
XFILLER_1_582 VPWR VGND sg13g2_decap_8
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_37_715 VPWR VGND sg13g2_decap_8
XFILLER_18_940 VPWR VGND sg13g2_decap_8
XFILLER_33_932 VPWR VGND sg13g2_decap_8
XFILLER_17_494 VPWR VGND sg13g2_decap_8
XFILLER_32_420 VPWR VGND sg13g2_fill_2
XFILLER_20_615 VPWR VGND sg13g2_decap_8
XFILLER_34_1020 VPWR VGND sg13g2_decap_8
XFILLER_8_181 VPWR VGND sg13g2_decap_8
XFILLER_9_682 VPWR VGND sg13g2_decap_8
XFILLER_28_704 VPWR VGND sg13g2_decap_8
XFILLER_24_965 VPWR VGND sg13g2_decap_8
XFILLER_23_497 VPWR VGND sg13g2_decap_8
XFILLER_7_608 VPWR VGND sg13g2_decap_8
XFILLER_11_659 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_3_803 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_2_324 VPWR VGND sg13g2_decap_8
Xhold170 hold170/A VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold192 hold192/A VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold181 hold181/A VPWR VGND net524 sg13g2_dlygate4sd3_1
XFILLER_19_726 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_15_921 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_42_762 VPWR VGND sg13g2_decap_8
XFILLER_41_250 VPWR VGND sg13g2_fill_2
XFILLER_14_464 VPWR VGND sg13g2_decap_8
XFILLER_15_998 VPWR VGND sg13g2_decap_8
XFILLER_30_902 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0992_ net430 VPWR u_ppwm_u_mem__0992_/Y VGND net349 hold106/A sg13g2_o21ai_1
XFILLER_30_979 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__234_ net195 VGND VPWR net265 hold67/A clknet_5_5__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__165_ u_ppwm_u_pwm__165_/A u_ppwm_u_pwm__165_/B u_ppwm_u_pwm__236_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_685 VPWR VGND sg13g2_decap_8
XFILLER_2_891 VPWR VGND sg13g2_decap_8
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_37_589 VPWR VGND sg13g2_decap_8
XFILLER_21_913 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
XFILLER_20_489 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1121__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_0_806 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_11 VPWR VGND uio_out[0] sg13g2_tielo
Xheichips25_ppwm_22 VPWR VGND uo_out[4] sg13g2_tielo
XFILLER_16_707 VPWR VGND sg13g2_decap_8
XFILLER_28_578 VPWR VGND sg13g2_decap_8
XFILLER_43_537 VPWR VGND sg13g2_decap_8
XFILLER_24_762 VPWR VGND sg13g2_decap_8
XFILLER_8_917 VPWR VGND sg13g2_decap_8
XFILLER_7_405 VPWR VGND sg13g2_decap_8
XFILLER_11_456 VPWR VGND sg13g2_decap_8
XFILLER_12_957 VPWR VGND sg13g2_decap_8
XFILLER_3_600 VPWR VGND sg13g2_decap_8
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
XFILLER_2_121 VPWR VGND sg13g2_decap_4
XFILLER_3_677 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_fill_2
XFILLER_19_523 VPWR VGND sg13g2_decap_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1191_ net169 VGND VPWR net486 hold231/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_537 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_9_22 VPWR VGND sg13g2_fill_1
XFILLER_15_795 VPWR VGND sg13g2_decap_8
XFILLER_9_66 VPWR VGND sg13g2_decap_4
XFILLER_14_294 VPWR VGND sg13g2_fill_1
XFILLER_30_776 VPWR VGND sg13g2_decap_8
XFILLER_31_1012 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0975_ VGND VPWR net350 u_ppwm_u_mem__0667_/Y u_ppwm_u_mem__1164_/D
+ u_ppwm_u_mem__0974_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__217_ VPWR VGND u_ppwm_u_pwm__203_/X u_ppwm_u_pwm__216_/X u_ppwm_u_pwm__215_/Y
+ u_ppwm_u_pwm__211_/Y u_ppwm_u_pwm__217_/Y u_ppwm_u_pwm__215_/C sg13g2_a221oi_1
XFILLER_7_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__148_ VGND VPWR u_ppwm_u_pwm__136_/Y net328 hold220/A u_ppwm_u_pwm__147_/Y
+ sg13g2_a21oi_1
XFILLER_6_482 VPWR VGND sg13g2_decap_8
XFILLER_38_865 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__097_ VGND VPWR u_ppwm_u_global_counter__056_/Y u_ppwm_u_global_counter__093_/Y
+ hold235/A u_ppwm_u_global_counter__099_/B sg13g2_a21oi_1
XFILLER_25_548 VPWR VGND sg13g2_decap_8
XFILLER_37_397 VPWR VGND sg13g2_fill_1
XFILLER_21_710 VPWR VGND sg13g2_decap_8
XFILLER_20_220 VPWR VGND sg13g2_fill_1
XFILLER_21_787 VPWR VGND sg13g2_decap_8
XFILLER_4_419 VPWR VGND sg13g2_decap_8
XFILLER_0_603 VPWR VGND sg13g2_decap_8
XFILLER_18_20 VPWR VGND sg13g2_decap_4
XFILLER_29_843 VPWR VGND sg13g2_decap_8
XFILLER_44_802 VPWR VGND sg13g2_decap_8
XFILLER_16_504 VPWR VGND sg13g2_decap_8
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_12_754 VPWR VGND sg13g2_decap_8
XFILLER_34_85 VPWR VGND sg13g2_decap_4
XFILLER_8_714 VPWR VGND sg13g2_decap_8
XFILLER_11_286 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0760_ u_ppwm_u_mem__0760_/Y net334 u_ppwm_u_mem__0760_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0691_ VPWR u_ppwm_u_mem__0691_/Y net606 VGND sg13g2_inv_1
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_3_474 VPWR VGND sg13g2_decap_8
XFILLER_39_618 VPWR VGND sg13g2_decap_8
XFILLER_47_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1174_ net118 VGND VPWR net209 hold46/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__660_ net319 VPWR u_ppwm_u_ex__660_/Y VGND net394 net396 sg13g2_o21ai_1
XFILLER_35_813 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__591_ u_ppwm_u_ex__591_/A u_ppwm_u_ex__593_/B u_ppwm_u_ex__591_/C u_ppwm_u_ex__591_/D
+ u_ppwm_u_ex__591_/X VPWR VGND sg13g2_and4_1
XFILLER_15_592 VPWR VGND sg13g2_decap_8
XFILLER_30_573 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0958_ net449 VPWR u_ppwm_u_mem__0958_/Y VGND net368 hold172/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0889_ VGND VPWR net360 u_ppwm_u_mem__0710_/Y hold247/A u_ppwm_u_mem__0888_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1204__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_38_662 VPWR VGND sg13g2_decap_8
XFILLER_26_846 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__789_ u_ppwm_u_ex__789_/Y net379 net322 VPWR VGND sg13g2_nand2_1
XFILLER_13_518 VPWR VGND sg13g2_decap_8
XFILLER_21_584 VPWR VGND sg13g2_decap_8
XFILLER_5_717 VPWR VGND sg13g2_decap_8
XFILLER_20_65 VPWR VGND sg13g2_fill_1
XFILLER_0_400 VPWR VGND sg13g2_decap_8
XFILLER_1_967 VPWR VGND sg13g2_decap_8
XFILLER_49_938 VPWR VGND sg13g2_decap_8
Xhold41 hold41/A VPWR VGND net238 sg13g2_dlygate4sd3_1
Xhold30 hold30/A VPWR VGND net227 sg13g2_dlygate4sd3_1
XFILLER_0_477 VPWR VGND sg13g2_decap_8
XFILLER_48_459 VPWR VGND sg13g2_decap_8
Xhold63 hold63/A VPWR VGND net260 sg13g2_dlygate4sd3_1
Xhold74 hold74/A VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold52 hold52/A VPWR VGND net249 sg13g2_dlygate4sd3_1
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
XFILLER_29_85 VPWR VGND sg13g2_decap_4
XFILLER_29_640 VPWR VGND sg13g2_decap_8
Xhold85 hold85/A VPWR VGND net282 sg13g2_dlygate4sd3_1
XFILLER_17_802 VPWR VGND sg13g2_decap_8
Xhold96 hold96/A VPWR VGND net293 sg13g2_dlygate4sd3_1
XFILLER_44_676 VPWR VGND sg13g2_decap_8
XFILLER_16_334 VPWR VGND sg13g2_fill_1
XFILLER_17_879 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_fill_1
XFILLER_43_186 VPWR VGND sg13g2_fill_1
XFILLER_31_326 VPWR VGND sg13g2_decap_8
XFILLER_8_511 VPWR VGND sg13g2_decap_8
XFILLER_12_551 VPWR VGND sg13g2_decap_8
XFILLER_8_588 VPWR VGND sg13g2_decap_8
XFILLER_6_34 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0812_ hold61/A hold98/A net412 u_ppwm_u_mem__0812_/X VPWR VGND sg13g2_mux2_1
XFILLER_6_56 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0743_ u_ppwm_u_mem__0743_/Y net334 u_ppwm_u_mem__0743_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0674_ VPWR u_ppwm_u_mem__0674_/Y net237 VGND sg13g2_inv_1
XFILLER_4_783 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__712_ u_ppwm_u_ex__712_/A u_ppwm_u_ex__712_/B hold309/A VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__1226_ net175 VGND VPWR net514 hold170/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_610 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1157_ net166 VGND VPWR net238 hold63/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__643_ u_ppwm_u_ex__644_/B net396 net319 VPWR VGND sg13g2_xnor2_1
XFILLER_23_805 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__574_ u_ppwm_u_ex__574_/Y hold209/A u_ppwm_u_ex__424_/Y hold234/A u_ppwm_u_ex__583_/A
+ VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1088_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1088_/B u_ppwm_u_mem__1090_/B
+ u_ppwm_u_mem__1219_/D VPWR VGND sg13g2_nor3_1
XFILLER_35_687 VPWR VGND sg13g2_decap_8
XFILLER_31_893 VPWR VGND sg13g2_decap_8
XFILLER_2_709 VPWR VGND sg13g2_decap_8
XFILLER_39_982 VPWR VGND sg13g2_decap_8
XFILLER_25_142 VPWR VGND sg13g2_decap_4
XFILLER_26_643 VPWR VGND sg13g2_decap_8
XFILLER_13_315 VPWR VGND sg13g2_fill_2
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_4
XFILLER_41_668 VPWR VGND sg13g2_decap_8
XFILLER_5_514 VPWR VGND sg13g2_decap_8
XFILLER_1_764 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_decap_8
XFILLER_0_274 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_45_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1011_ VGND VPWR net346 u_ppwm_u_mem__0649_/Y u_ppwm_u_mem__1182_/D
+ u_ppwm_u_mem__1010_/Y sg13g2_a21oi_1
XFILLER_44_473 VPWR VGND sg13g2_decap_8
XFILLER_16_175 VPWR VGND sg13g2_fill_2
XFILLER_17_676 VPWR VGND sg13g2_decap_8
XFILLER_31_145 VPWR VGND sg13g2_fill_2
XFILLER_32_668 VPWR VGND sg13g2_decap_8
XFILLER_13_882 VPWR VGND sg13g2_decap_8
XFILLER_8_341 VPWR VGND sg13g2_fill_2
XFILLER_9_864 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0726_ VPWR u_ppwm_u_mem__0726_/Y net513 VGND sg13g2_inv_1
XFILLER_4_580 VPWR VGND sg13g2_decap_8
Xfanout309 fanout309/A net309 VPWR VGND sg13g2_buf_8
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0657_ VPWR u_ppwm_u_mem__0657_/Y net208 VGND sg13g2_inv_1
XFILLER_39_256 VPWR VGND sg13g2_fill_2
XFILLER_36_930 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1209_ net167 VGND VPWR u_ppwm_u_mem__1209_/D hold128/A clknet_5_13__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_23_602 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__626_ fanout315/A u_ppwm_u_ex__637_/A VPWR VGND net317 sg13g2_nand2b_2
Xu_ppwm_u_ex__557_ hold185/A net393 u_ppwm_u_ex__558_/C VPWR VGND sg13g2_xor2_1
XFILLER_22_156 VPWR VGND sg13g2_fill_2
XFILLER_23_679 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__488_ u_ppwm_u_ex__488_/Y u_ppwm_u_ex__488_/A u_ppwm_u_ex__488_/B VPWR
+ VGND sg13g2_nand2_1
XFILLER_31_690 VPWR VGND sg13g2_decap_8
XFILLER_2_506 VPWR VGND sg13g2_decap_8
Xhold330 hold330/A VPWR VGND net673 sg13g2_dlygate4sd3_1
XFILLER_19_908 VPWR VGND sg13g2_decap_8
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_18_429 VPWR VGND sg13g2_decap_8
XFILLER_27_952 VPWR VGND sg13g2_decap_8
XFILLER_42_944 VPWR VGND sg13g2_decap_8
XFILLER_14_646 VPWR VGND sg13g2_decap_8
XFILLER_13_145 VPWR VGND sg13g2_fill_1
XFILLER_10_830 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__181_ u_ppwm_u_pwm__242_/D net422 u_ppwm_u_pwm__181_/B u_ppwm_u_pwm__181_/C
+ VPWR VGND sg13g2_and3_1
XFILLER_6_867 VPWR VGND sg13g2_decap_8
XFILLER_5_388 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_4
XFILLER_1_561 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_36_215 VPWR VGND sg13g2_decap_8
XFILLER_17_473 VPWR VGND sg13g2_decap_8
XFILLER_18_996 VPWR VGND sg13g2_decap_8
XFILLER_33_911 VPWR VGND sg13g2_decap_8
XFILLER_32_454 VPWR VGND sg13g2_fill_1
XFILLER_33_988 VPWR VGND sg13g2_decap_8
XFILLER_9_661 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0709_ VPWR u_ppwm_u_mem__0709_/Y net591 VGND sg13g2_inv_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
XFILLER_43_719 VPWR VGND sg13g2_decap_8
XFILLER_42_218 VPWR VGND sg13g2_decap_8
XFILLER_24_944 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__609_ VPWR VGND u_ppwm_u_ex__608_/Y u_ppwm_u_ex__595_/Y u_ppwm_u_ex__607_/Y
+ u_ppwm_u_ex__519_/A u_ppwm_u_ex__609_/Y hold118/A sg13g2_a221oi_1
XFILLER_11_638 VPWR VGND sg13g2_decap_8
XFILLER_23_476 VPWR VGND sg13g2_decap_8
XFILLER_6_108 VPWR VGND sg13g2_fill_1
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_fill_1
XFILLER_12_55 VPWR VGND sg13g2_fill_1
XFILLER_3_859 VPWR VGND sg13g2_decap_8
Xhold171 hold171/A VPWR VGND net514 sg13g2_dlygate4sd3_1
Xhold160 hold160/A VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold193 hold193/A VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold182 hold182/A VPWR VGND net525 sg13g2_dlygate4sd3_1
XFILLER_19_705 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_15_900 VPWR VGND sg13g2_decap_8
XFILLER_34_719 VPWR VGND sg13g2_decap_8
XFILLER_42_741 VPWR VGND sg13g2_decap_8
XFILLER_14_443 VPWR VGND sg13g2_decap_8
XFILLER_15_977 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0991_ VGND VPWR net349 u_ppwm_u_mem__0659_/Y u_ppwm_u_mem__1172_/D
+ u_ppwm_u_mem__0990_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__233_ net197 VGND VPWR net250 hold52/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_30_958 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__164_ net422 VPWR u_ppwm_u_pwm__165_/B VGND net625 net630 sg13g2_o21ai_1
XFILLER_6_664 VPWR VGND sg13g2_decap_8
XFILLER_2_870 VPWR VGND sg13g2_decap_8
XFILLER_37_568 VPWR VGND sg13g2_decap_8
XFILLER_18_793 VPWR VGND sg13g2_decap_8
XFILLER_33_785 VPWR VGND sg13g2_decap_8
XFILLER_21_969 VPWR VGND sg13g2_decap_8
XFILLER_20_468 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_23 VPWR VGND uo_out[5] sg13g2_tielo
Xheichips25_ppwm_12 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_28_557 VPWR VGND sg13g2_decap_8
XFILLER_43_516 VPWR VGND sg13g2_decap_8
XFILLER_15_207 VPWR VGND sg13g2_fill_1
XFILLER_24_741 VPWR VGND sg13g2_decap_8
XFILLER_12_936 VPWR VGND sg13g2_decap_8
XFILLER_11_435 VPWR VGND sg13g2_decap_8
XFILLER_3_656 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1176__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_2_177 VPWR VGND sg13g2_decap_4
XFILLER_47_822 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_19_502 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1190_ net54 VGND VPWR u_ppwm_u_mem__1190_/D hold173/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_19_579 VPWR VGND sg13g2_decap_8
XFILLER_15_774 VPWR VGND sg13g2_decap_8
XFILLER_30_755 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0974_ net434 VPWR u_ppwm_u_mem__0974_/Y VGND net355 net214 sg13g2_o21ai_1
Xu_ppwm_u_pwm__216_ u_ppwm_u_pwm__216_/A u_ppwm_u_pwm__216_/B u_ppwm_u_pwm__216_/X
+ VPWR VGND sg13g2_and2_1
XFILLER_7_951 VPWR VGND sg13g2_decap_8
XFILLER_6_461 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__147_ net425 VPWR u_ppwm_u_pwm__147_/Y VGND net396 net329 sg13g2_o21ai_1
XFILLER_9_1025 VPWR VGND sg13g2_decap_4
XFILLER_38_844 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__096_ net331 u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__099_/B
+ VPWR VGND sg13g2_and2_1
XFILLER_25_527 VPWR VGND sg13g2_decap_8
XFILLER_18_590 VPWR VGND sg13g2_decap_8
XFILLER_33_582 VPWR VGND sg13g2_decap_8
XFILLER_20_254 VPWR VGND sg13g2_decap_8
XFILLER_20_265 VPWR VGND sg13g2_fill_1
XFILLER_21_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__231__179 VPWR VGND net179 sg13g2_tiehi
Xu_ppwm_u_mem__1207__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_0_659 VPWR VGND sg13g2_decap_8
XFILLER_29_822 VPWR VGND sg13g2_decap_8
XFILLER_29_899 VPWR VGND sg13g2_decap_8
XFILLER_44_858 VPWR VGND sg13g2_decap_8
XFILLER_12_733 VPWR VGND sg13g2_decap_8
XFILLER_15_1019 VPWR VGND sg13g2_decap_8
XFILLER_11_243 VPWR VGND sg13g2_fill_1
XFILLER_11_254 VPWR VGND sg13g2_fill_2
XFILLER_11_276 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0690_ VPWR u_ppwm_u_mem__0690_/Y net289 VGND sg13g2_inv_1
XFILLER_4_965 VPWR VGND sg13g2_decap_8
XFILLER_3_453 VPWR VGND sg13g2_decap_8
XFILLER_19_310 VPWR VGND sg13g2_fill_1
XFILLER_19_321 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1173_ net122 VGND VPWR net244 hold106/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_47_696 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__590_ u_ppwm_u_ex__591_/D hold333/A hold221/A VPWR VGND sg13g2_nand2b_1
XFILLER_34_313 VPWR VGND sg13g2_fill_2
XFILLER_35_869 VPWR VGND sg13g2_decap_8
XFILLER_43_880 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_30_552 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0957_ VGND VPWR net367 u_ppwm_u_mem__0676_/Y u_ppwm_u_mem__1155_/D
+ u_ppwm_u_mem__0956_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0888_ net447 VPWR u_ppwm_u_mem__0888_/Y VGND net360 net506 sg13g2_o21ai_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_29_107 VPWR VGND sg13g2_fill_2
XFILLER_38_641 VPWR VGND sg13g2_decap_8
XFILLER_26_825 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__079_ net657 u_ppwm_u_global_counter__082_/D net291 u_ppwm_u_global_counter__083_/B
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__788_ VGND VPWR u_ppwm_u_ex__753_/B u_ppwm_u_ex__785_/Y u_ppwm_u_ex__788_/Y
+ u_ppwm_u_ex__787_/Y sg13g2_a21oi_1
XFILLER_38_1019 VPWR VGND sg13g2_decap_8
XFILLER_25_379 VPWR VGND sg13g2_decap_8
XFILLER_34_880 VPWR VGND sg13g2_decap_8
XFILLER_21_563 VPWR VGND sg13g2_decap_8
XFILLER_20_44 VPWR VGND sg13g2_fill_1
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_1_946 VPWR VGND sg13g2_decap_8
Xhold20 hold20/A VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold31 hold31/A VPWR VGND net228 sg13g2_dlygate4sd3_1
XFILLER_0_456 VPWR VGND sg13g2_decap_8
XFILLER_48_438 VPWR VGND sg13g2_decap_8
Xhold64 hold64/A VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold53 hold53/A VPWR VGND net250 sg13g2_dlygate4sd3_1
Xhold42 hold42/A VPWR VGND net239 sg13g2_dlygate4sd3_1
Xhold86 hold86/A VPWR VGND net283 sg13g2_dlygate4sd3_1
Xhold97 hold97/A VPWR VGND net294 sg13g2_dlygate4sd3_1
Xhold75 hold75/A VPWR VGND net272 sg13g2_dlygate4sd3_1
XFILLER_29_696 VPWR VGND sg13g2_decap_8
XFILLER_44_655 VPWR VGND sg13g2_decap_8
XFILLER_17_858 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1131__99 VPWR VGND net99 sg13g2_tiehi
XFILLER_12_530 VPWR VGND sg13g2_decap_8
XFILLER_25_891 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1110__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_8_567 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0811_ net412 u_ppwm_u_mem__0616_/Y u_ppwm_u_mem__0810_/Y u_ppwm_u_mem__0811_/X
+ VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_mem__0742_ hold85/A hold144/A net413 u_ppwm_u_mem__0743_/B VPWR VGND sg13g2_mux2_1
XFILLER_4_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0673_ VPWR u_ppwm_u_mem__0673_/Y net306 VGND sg13g2_inv_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1225_ net174 VGND VPWR net551 hold206/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__711_ net426 VPWR u_ppwm_u_ex__712_/B VGND net651 net310 sg13g2_o21ai_1
XFILLER_19_173 VPWR VGND sg13g2_decap_8
XFILLER_47_493 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1156_ net168 VGND VPWR net261 hold172/A clknet_5_30__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__642_ VGND VPWR u_ppwm_u_ex__636_/A u_ppwm_u_ex__636_/B u_ppwm_u_ex__644_/A
+ u_ppwm_u_ex__634_/X sg13g2_a21oi_1
XFILLER_35_666 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__573_ u_ppwm_u_ex__594_/B u_ppwm_u_ex__573_/C u_ppwm_u_ex__573_/A u_ppwm_u_ex__617_/B
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__1087_ net618 net338 u_ppwm_u_mem__1090_/B VPWR VGND sg13g2_and2_1
XFILLER_31_872 VPWR VGND sg13g2_decap_8
XFILLER_44_1012 VPWR VGND sg13g2_decap_8
XFILLER_45_408 VPWR VGND sg13g2_fill_2
XFILLER_39_961 VPWR VGND sg13g2_decap_8
XFILLER_26_622 VPWR VGND sg13g2_decap_8
XFILLER_38_493 VPWR VGND sg13g2_fill_2
XFILLER_14_828 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_26_699 VPWR VGND sg13g2_decap_8
XFILLER_41_647 VPWR VGND sg13g2_decap_8
XFILLER_22_894 VPWR VGND sg13g2_decap_8
XFILLER_31_32 VPWR VGND sg13g2_decap_4
XFILLER_1_743 VPWR VGND sg13g2_decap_8
XFILLER_49_714 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_45_920 VPWR VGND sg13g2_decap_8
XFILLER_17_655 VPWR VGND sg13g2_decap_8
XFILLER_29_493 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1010_ net430 VPWR u_ppwm_u_mem__1010_/Y VGND net346 net524 sg13g2_o21ai_1
XFILLER_45_997 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_4
XFILLER_32_647 VPWR VGND sg13g2_decap_8
XFILLER_13_861 VPWR VGND sg13g2_decap_8
XFILLER_9_843 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0725_ u_ppwm_u_mem__1094_/A net423 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0656_ VPWR u_ppwm_u_mem__0656_/Y net620 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1208_ net56 VGND VPWR net472 hold236/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1139_ net83 VGND VPWR net273 hold19/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
Xheichips25_ppwm_3 VPWR VGND uio_oe[0] sg13g2_tielo
Xu_ppwm_u_ex__625_ u_ppwm/instr\[0\] net317 fanout316/A VPWR VGND sg13g2_nor2_2
XFILLER_36_986 VPWR VGND sg13g2_decap_8
XFILLER_22_113 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__556_ hold203/A net395 u_ppwm_u_ex__558_/B VPWR VGND sg13g2_nor2b_1
XFILLER_23_658 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__487_ net400 u_ppwm_u_ex__442_/Y u_ppwm_u_ex__487_/Y VPWR VGND sg13g2_nor2b_1
Xhold320 hold320/A VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold331 hold331/A VPWR VGND net674 sg13g2_dlygate4sd3_1
XFILLER_46_728 VPWR VGND sg13g2_decap_8
XFILLER_45_216 VPWR VGND sg13g2_fill_2
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_42_923 VPWR VGND sg13g2_decap_8
XFILLER_14_625 VPWR VGND sg13g2_decap_8
XFILLER_26_98 VPWR VGND sg13g2_fill_2
XFILLER_26_496 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__180_ u_ppwm_u_pwm__181_/C net626 u_ppwm_u_pwm__182_/C VPWR VGND sg13g2_nand2_1
XFILLER_22_691 VPWR VGND sg13g2_decap_8
XFILLER_6_846 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_5_367 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_1_540 VPWR VGND sg13g2_decap_8
XFILLER_49_511 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_17_452 VPWR VGND sg13g2_decap_8
XFILLER_18_975 VPWR VGND sg13g2_decap_8
XFILLER_45_794 VPWR VGND sg13g2_decap_8
XFILLER_32_422 VPWR VGND sg13g2_fill_1
XFILLER_32_433 VPWR VGND sg13g2_fill_1
XFILLER_33_967 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__814__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_9_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0708_ VPWR u_ppwm_u_mem__0708_/Y net483 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0639_ VPWR u_ppwm_u_mem__0639_/Y net231 VGND sg13g2_inv_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
XFILLER_28_739 VPWR VGND sg13g2_decap_8
XFILLER_24_923 VPWR VGND sg13g2_decap_8
XFILLER_36_783 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__608_ u_ppwm_u_ex__608_/Y net380 u_ppwm_u_ex__608_/B VPWR VGND sg13g2_nand2_1
XFILLER_23_455 VPWR VGND sg13g2_decap_8
XFILLER_11_617 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__539_ u_ppwm_u_ex__543_/B net378 hold308/A VPWR VGND sg13g2_xnor2_1
XFILLER_3_838 VPWR VGND sg13g2_decap_8
Xhold150 hold150/A VPWR VGND net493 sg13g2_dlygate4sd3_1
Xhold161 hold161/A VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold172 hold172/A VPWR VGND net515 sg13g2_dlygate4sd3_1
XFILLER_2_359 VPWR VGND sg13g2_decap_8
Xhold194 hold194/A VPWR VGND net537 sg13g2_dlygate4sd3_1
Xhold183 hold183/A VPWR VGND net526 sg13g2_dlygate4sd3_1
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_37_20 VPWR VGND sg13g2_fill_2
XFILLER_42_720 VPWR VGND sg13g2_decap_8
XFILLER_14_422 VPWR VGND sg13g2_decap_8
XFILLER_41_230 VPWR VGND sg13g2_decap_8
XFILLER_15_956 VPWR VGND sg13g2_decap_8
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_293 VPWR VGND sg13g2_fill_2
XFILLER_42_797 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_decap_8
XFILLER_30_937 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0990_ net431 VPWR u_ppwm_u_mem__0990_/Y VGND net351 net270 sg13g2_o21ai_1
Xu_ppwm_u_pwm__232_ net177 VGND VPWR net221 hold23/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__811__28 VPWR VGND net28 sg13g2_tiehi
Xu_ppwm_u_pwm__163_ net625 net630 u_ppwm_u_pwm__165_/A VPWR VGND sg13g2_and2_1
XFILLER_6_643 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_49_385 VPWR VGND sg13g2_decap_8
XFILLER_37_547 VPWR VGND sg13g2_decap_8
XFILLER_18_772 VPWR VGND sg13g2_decap_8
XFILLER_25_709 VPWR VGND sg13g2_decap_8
XFILLER_45_591 VPWR VGND sg13g2_decap_8
XFILLER_17_293 VPWR VGND sg13g2_fill_1
XFILLER_33_764 VPWR VGND sg13g2_decap_8
XFILLER_21_948 VPWR VGND sg13g2_decap_8
XFILLER_20_447 VPWR VGND sg13g2_decap_8
XFILLER_32_296 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1201__112 VPWR VGND net112 sg13g2_tiehi
Xheichips25_ppwm_24 VPWR VGND uo_out[6] sg13g2_tielo
Xheichips25_ppwm_13 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_28_536 VPWR VGND sg13g2_decap_8
XFILLER_24_720 VPWR VGND sg13g2_decap_8
XFILLER_36_580 VPWR VGND sg13g2_decap_8
XFILLER_11_414 VPWR VGND sg13g2_decap_8
XFILLER_12_915 VPWR VGND sg13g2_decap_8
XFILLER_23_274 VPWR VGND sg13g2_fill_2
XFILLER_24_797 VPWR VGND sg13g2_decap_8
XFILLER_23_99 VPWR VGND sg13g2_fill_1
XFILLER_3_635 VPWR VGND sg13g2_decap_8
XFILLER_2_156 VPWR VGND sg13g2_fill_1
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_801 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_19_558 VPWR VGND sg13g2_decap_8
XFILLER_15_753 VPWR VGND sg13g2_decap_8
XFILLER_42_594 VPWR VGND sg13g2_decap_8
XFILLER_30_734 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0973_ VGND VPWR net355 u_ppwm_u_mem__0668_/Y hold18/A u_ppwm_u_mem__0972_/Y
+ sg13g2_a21oi_1
XFILLER_10_480 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__215_ u_ppwm_u_pwm__215_/A u_ppwm_u_pwm__215_/B u_ppwm_u_pwm__215_/C
+ u_ppwm_u_pwm__215_/D u_ppwm_u_pwm__215_/Y VPWR VGND sg13g2_nor4_1
XFILLER_7_930 VPWR VGND sg13g2_decap_8
XFILLER_11_981 VPWR VGND sg13g2_decap_8
XFILLER_6_440 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__146_ VGND VPWR u_ppwm_u_pwm__137_/Y net328 hold22/A u_ppwm_u_pwm__145_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1216__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_9_1004 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1120__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_38_823 VPWR VGND sg13g2_decap_8
XFILLER_49_182 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__095_ u_ppwm_u_global_counter__103_/C net552 net577 u_ppwm_u_global_counter__095_/C
+ VPWR VGND sg13g2_and3_2
XFILLER_25_506 VPWR VGND sg13g2_decap_8
XFILLER_33_561 VPWR VGND sg13g2_decap_8
XFILLER_21_745 VPWR VGND sg13g2_decap_8
XFILLER_0_638 VPWR VGND sg13g2_decap_8
XFILLER_47_108 VPWR VGND sg13g2_decap_8
XFILLER_29_801 VPWR VGND sg13g2_decap_8
XFILLER_29_878 VPWR VGND sg13g2_decap_8
XFILLER_44_837 VPWR VGND sg13g2_decap_8
XFILLER_16_539 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1143__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_43_358 VPWR VGND sg13g2_decap_8
XFILLER_12_712 VPWR VGND sg13g2_decap_8
XFILLER_11_222 VPWR VGND sg13g2_decap_4
XFILLER_24_594 VPWR VGND sg13g2_decap_8
XFILLER_12_789 VPWR VGND sg13g2_decap_8
XFILLER_8_749 VPWR VGND sg13g2_decap_8
XFILLER_4_944 VPWR VGND sg13g2_decap_8
XFILLER_3_432 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__247__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_47_675 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1172_ net126 VGND VPWR u_ppwm_u_mem__1172_/D hold73/A clknet_5_14__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_848 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
XFILLER_22_509 VPWR VGND sg13g2_decap_8
XFILLER_30_531 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0956_ net444 VPWR u_ppwm_u_mem__0956_/Y VGND net367 net247 sg13g2_o21ai_1
Xu_ppwm_u_mem__0887_ VGND VPWR net362 u_ppwm_u_mem__0711_/Y hold164/A u_ppwm_u_mem__0886_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__129_ VPWR u_ppwm_u_pwm__129_/Y net568 VGND sg13g2_inv_1
XFILLER_34_0 VPWR VGND sg13g2_decap_4
XFILLER_38_620 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_804 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_fill_2
XFILLER_37_163 VPWR VGND sg13g2_fill_2
XFILLER_38_697 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__078_ u_ppwm_u_global_counter__082_/D net291 hold95/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__787_ u_ppwm_u_ex__787_/Y u_ppwm_u_ex__787_/A u_ppwm_u_ex__787_/B VPWR
+ VGND sg13g2_nand2_1
XFILLER_25_347 VPWR VGND sg13g2_decap_4
XFILLER_41_829 VPWR VGND sg13g2_decap_8
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_20_12 VPWR VGND sg13g2_decap_8
XFILLER_20_23 VPWR VGND sg13g2_fill_2
XFILLER_20_34 VPWR VGND sg13g2_fill_1
XFILLER_1_925 VPWR VGND sg13g2_decap_8
XFILLER_0_435 VPWR VGND sg13g2_decap_8
XFILLER_48_417 VPWR VGND sg13g2_decap_8
Xhold32 hold32/A VPWR VGND net229 sg13g2_dlygate4sd3_1
Xhold21 hold21/A VPWR VGND net218 sg13g2_dlygate4sd3_1
Xhold10 hold10/A VPWR VGND net207 sg13g2_dlygate4sd3_1
Xhold54 hold54/A VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold65 hold65/A VPWR VGND net262 sg13g2_dlygate4sd3_1
Xhold43 hold43/A VPWR VGND net240 sg13g2_dlygate4sd3_1
Xhold76 hold76/A VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold98 hold98/A VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold87 hold87/A VPWR VGND net284 sg13g2_dlygate4sd3_1
XFILLER_43_100 VPWR VGND sg13g2_fill_2
XFILLER_17_837 VPWR VGND sg13g2_decap_8
XFILLER_29_675 VPWR VGND sg13g2_decap_8
XFILLER_44_634 VPWR VGND sg13g2_decap_8
XFILLER_16_325 VPWR VGND sg13g2_decap_4
XFILLER_28_196 VPWR VGND sg13g2_decap_4
XFILLER_25_870 VPWR VGND sg13g2_decap_8
XFILLER_32_829 VPWR VGND sg13g2_decap_8
XFILLER_40_884 VPWR VGND sg13g2_decap_8
XFILLER_8_546 VPWR VGND sg13g2_decap_8
XFILLER_12_586 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0810_ net404 VPWR u_ppwm_u_mem__0810_/Y VGND hold128/A net411 sg13g2_o21ai_1
Xu_ppwm_u_mem__0741_ hold110/A hold182/A net411 u_ppwm_u_mem__0741_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0672_ VPWR u_ppwm_u_mem__0672_/Y net576 VGND sg13g2_inv_1
XFILLER_4_741 VPWR VGND sg13g2_decap_8
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1224_ net68 VGND VPWR net599 hold254/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__710_ VPWR VGND net316 net309 u_ppwm_u_ex__709_/Y net386 u_ppwm_u_ex__712_/A
+ net311 sg13g2_a221oi_1
XFILLER_48_984 VPWR VGND sg13g2_decap_8
XFILLER_47_472 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__641_ VGND VPWR u_ppwm_u_ex__638_/Y u_ppwm_u_ex__639_/Y u_ppwm_u_ex__808_/D
+ u_ppwm_u_ex__640_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__1155_ net170 VGND VPWR u_ppwm_u_mem__1155_/D hold50/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_645 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__572_ VGND VPWR u_ppwm_u_ex__538_/B hold314/A u_ppwm_u_ex__573_/C net324
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1086_ net618 net338 u_ppwm_u_mem__1088_/B VPWR VGND sg13g2_nor2_1
XFILLER_34_155 VPWR VGND sg13g2_decap_8
XFILLER_34_166 VPWR VGND sg13g2_fill_2
XFILLER_22_328 VPWR VGND sg13g2_fill_2
XFILLER_31_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0939_ VGND VPWR net366 u_ppwm_u_mem__0685_/Y u_ppwm_u_mem__1146_/D
+ u_ppwm_u_mem__0938_/Y sg13g2_a21oi_1
XFILLER_39_940 VPWR VGND sg13g2_decap_8
XFILLER_26_601 VPWR VGND sg13g2_decap_8
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_26_678 VPWR VGND sg13g2_decap_8
XFILLER_41_626 VPWR VGND sg13g2_decap_8
XFILLER_13_317 VPWR VGND sg13g2_fill_1
XFILLER_21_361 VPWR VGND sg13g2_decap_4
XFILLER_22_873 VPWR VGND sg13g2_decap_8
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_5_549 VPWR VGND sg13g2_decap_8
XFILLER_1_722 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_1_799 VPWR VGND sg13g2_decap_8
XFILLER_17_634 VPWR VGND sg13g2_decap_8
XFILLER_45_976 VPWR VGND sg13g2_decap_8
XFILLER_32_626 VPWR VGND sg13g2_decap_8
XFILLER_13_840 VPWR VGND sg13g2_decap_8
XFILLER_40_681 VPWR VGND sg13g2_decap_8
XFILLER_8_321 VPWR VGND sg13g2_fill_1
XFILLER_8_310 VPWR VGND sg13g2_decap_8
XFILLER_9_822 VPWR VGND sg13g2_decap_8
XFILLER_8_343 VPWR VGND sg13g2_fill_1
XFILLER_9_899 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0724_ VPWR u_ppwm_u_mem__0724_/Y net511 VGND sg13g2_inv_1
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0655_ VPWR u_ppwm_u_mem__0655_/Y net453 VGND sg13g2_inv_1
XFILLER_39_258 VPWR VGND sg13g2_fill_1
XFILLER_48_781 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1207_ net64 VGND VPWR u_ppwm_u_mem__1207_/D hold89/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_965 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1138_ net85 VGND VPWR net217 hold174/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
Xheichips25_ppwm_4 VPWR VGND uio_oe[1] sg13g2_tielo
Xu_ppwm_u_ex__624_ fanout317/A u_ppwm/instr\[1\] VPWR VGND u_ppwm/instr\[2\] sg13g2_nand2b_2
XFILLER_35_453 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__555_ hold243/A hold332/A u_ppwm_u_ex__560_/C VPWR VGND sg13g2_nor2b_1
XFILLER_23_637 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1069_ VGND VPWR net338 u_ppwm_u_mem__0620_/Y hold224/A u_ppwm_u_mem__1068_/Y
+ sg13g2_a21oi_1
XFILLER_10_309 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__486_ u_ppwm_u_ex__488_/B u_ppwm_u_ex__486_/B u_ppwm_u_ex__486_/Y VPWR
+ VGND sg13g2_nor2_1
XFILLER_30_191 VPWR VGND sg13g2_fill_1
XFILLER_11_1023 VPWR VGND sg13g2_decap_4
Xhold310 hold310/A VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold332 hold332/A VPWR VGND net675 sg13g2_dlygate4sd3_1
Xhold321 hold321/A VPWR VGND net664 sg13g2_dlygate4sd3_1
XFILLER_46_707 VPWR VGND sg13g2_decap_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_42_902 VPWR VGND sg13g2_decap_8
XFILLER_14_604 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__808__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_26_475 VPWR VGND sg13g2_decap_8
XFILLER_42_979 VPWR VGND sg13g2_decap_8
XFILLER_22_670 VPWR VGND sg13g2_decap_8
XFILLER_6_825 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_5_346 VPWR VGND sg13g2_decap_8
XFILLER_1_596 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_37_729 VPWR VGND sg13g2_decap_8
XFILLER_17_431 VPWR VGND sg13g2_decap_8
XFILLER_18_954 VPWR VGND sg13g2_decap_8
XFILLER_36_239 VPWR VGND sg13g2_decap_8
XFILLER_45_773 VPWR VGND sg13g2_decap_8
XFILLER_33_946 VPWR VGND sg13g2_decap_8
XFILLER_20_629 VPWR VGND sg13g2_decap_8
XFILLER_41_990 VPWR VGND sg13g2_decap_8
XFILLER_9_696 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0707_ VPWR u_ppwm_u_mem__0707_/Y net301 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0638_ VPWR u_ppwm_u_mem__0638_/Y net284 VGND sg13g2_inv_1
XFILLER_28_718 VPWR VGND sg13g2_decap_8
XFILLER_24_902 VPWR VGND sg13g2_decap_8
XFILLER_36_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1130__101 VPWR VGND net101 sg13g2_tiehi
Xu_ppwm_u_ex__607_ u_ppwm_u_ex__606_/Y VPWR u_ppwm_u_ex__607_/Y VGND u_ppwm_u_ex__600_/Y
+ u_ppwm_u_ex__604_/Y sg13g2_o21ai_1
XFILLER_23_434 VPWR VGND sg13g2_decap_8
XFILLER_24_979 VPWR VGND sg13g2_decap_8
XFILLER_10_106 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__538_ net378 u_ppwm_u_ex__538_/B u_ppwm_u_ex__538_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_ex__469_ u_ppwm_u_ex__488_/B u_ppwm_u_ex__469_/B u_ppwm_u_ex__469_/C u_ppwm_u_ex__469_/X
+ VPWR VGND sg13g2_or3_1
XFILLER_32_990 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_3_817 VPWR VGND sg13g2_decap_8
Xhold140 hold140/A VPWR VGND net483 sg13g2_dlygate4sd3_1
XFILLER_2_338 VPWR VGND sg13g2_decap_8
Xhold162 hold162/A VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold151 hold151/A VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold195 hold195/A VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold184 hold184/A VPWR VGND net527 sg13g2_dlygate4sd3_1
Xhold173 hold173/A VPWR VGND net516 sg13g2_dlygate4sd3_1
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_2_1010 VPWR VGND sg13g2_decap_8
XFILLER_15_935 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_42_776 VPWR VGND sg13g2_decap_8
XFILLER_14_478 VPWR VGND sg13g2_decap_8
XFILLER_30_916 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__231_ net179 VGND VPWR net223 hold25/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_622 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__162_ VGND VPWR u_ppwm_u_pwm__129_/Y net330 hold226/A u_ppwm_u_pwm__161_/Y
+ sg13g2_a21oi_1
XFILLER_6_699 VPWR VGND sg13g2_decap_8
XFILLER_1_393 VPWR VGND sg13g2_decap_8
XFILLER_49_364 VPWR VGND sg13g2_decap_8
XFILLER_18_751 VPWR VGND sg13g2_decap_8
XFILLER_45_570 VPWR VGND sg13g2_decap_8
XFILLER_17_250 VPWR VGND sg13g2_decap_8
XFILLER_33_743 VPWR VGND sg13g2_decap_8
XFILLER_21_927 VPWR VGND sg13g2_decap_8
XFILLER_20_426 VPWR VGND sg13g2_decap_8
XFILLER_9_493 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_25 VPWR VGND uo_out[7] sg13g2_tielo
Xheichips25_ppwm_14 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_28_515 VPWR VGND sg13g2_decap_8
XFILLER_23_231 VPWR VGND sg13g2_fill_2
XFILLER_24_776 VPWR VGND sg13g2_decap_8
XFILLER_7_419 VPWR VGND sg13g2_decap_8
XFILLER_23_78 VPWR VGND sg13g2_decap_8
XFILLER_20_993 VPWR VGND sg13g2_decap_8
XFILLER_23_89 VPWR VGND sg13g2_fill_2
XFILLER_3_614 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_24_1000 VPWR VGND sg13g2_decap_8
Xfanout450 net451 net450 VPWR VGND sg13g2_buf_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_19_537 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_15_732 VPWR VGND sg13g2_decap_8
XFILLER_42_573 VPWR VGND sg13g2_decap_8
XFILLER_30_713 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0972_ net434 VPWR u_ppwm_u_mem__0972_/Y VGND net355 hold85/A sg13g2_o21ai_1
XFILLER_11_960 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__214_ hold278/A u_ppwm_u_pwm__214_/B u_ppwm_u_pwm__215_/D VPWR VGND
+ sg13g2_nor2_1
XFILLER_31_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_986 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__145_ net424 VPWR u_ppwm_u_pwm__145_/Y VGND net398 net328 sg13g2_o21ai_1
XFILLER_6_496 VPWR VGND sg13g2_decap_8
XFILLER_38_802 VPWR VGND sg13g2_decap_8
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__094_ net553 u_ppwm_u_global_counter__093_/Y hold211/A VPWR
+ VGND sg13g2_nor2b_1
XFILLER_38_879 VPWR VGND sg13g2_decap_8
XFILLER_33_540 VPWR VGND sg13g2_decap_8
XFILLER_21_724 VPWR VGND sg13g2_decap_8
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_617 VPWR VGND sg13g2_decap_8
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_29_857 VPWR VGND sg13g2_decap_8
XFILLER_16_518 VPWR VGND sg13g2_decap_8
XFILLER_37_890 VPWR VGND sg13g2_decap_8
XFILLER_24_573 VPWR VGND sg13g2_decap_8
XFILLER_8_728 VPWR VGND sg13g2_decap_8
XFILLER_12_768 VPWR VGND sg13g2_decap_8
XFILLER_11_267 VPWR VGND sg13g2_decap_8
XFILLER_20_790 VPWR VGND sg13g2_decap_8
XFILLER_4_923 VPWR VGND sg13g2_decap_8
XFILLER_3_411 VPWR VGND sg13g2_decap_8
XFILLER_3_488 VPWR VGND sg13g2_decap_8
XFILLER_47_654 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1171_ net130 VGND VPWR net271 hold124/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_304 VPWR VGND sg13g2_fill_1
XFILLER_35_827 VPWR VGND sg13g2_decap_8
XFILLER_30_587 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0955_ VGND VPWR net367 u_ppwm_u_mem__0677_/Y hold51/A u_ppwm_u_mem__0954_/Y
+ sg13g2_a21oi_1
XFILLER_7_783 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0886_ net448 VPWR u_ppwm_u_mem__0886_/Y VGND net362 net491 sg13g2_o21ai_1
Xu_ppwm_u_pwm__128_ VPWR u_ppwm_u_pwm__128_/Y hold192/A VGND sg13g2_inv_1
Xu_ppwm_u_pwm__230__181 VPWR VGND net181 sg13g2_tiehi
Xu_ppwm_u_mem__1159__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__786_ net321 VPWR u_ppwm_u_ex__787_/B VGND hold310/A hold296/A sg13g2_o21ai_1
XFILLER_38_676 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__077_ u_ppwm_u_global_counter__082_/D net462 hold120/A VPWR
+ VGND sg13g2_nor2_1
XFILLER_41_808 VPWR VGND sg13g2_decap_8
XFILLER_21_521 VPWR VGND sg13g2_decap_8
XFILLER_33_381 VPWR VGND sg13g2_decap_8
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
XFILLER_21_598 VPWR VGND sg13g2_decap_8
XFILLER_1_904 VPWR VGND sg13g2_decap_8
XFILLER_0_414 VPWR VGND sg13g2_decap_8
Xhold22 hold22/A VPWR VGND net219 sg13g2_dlygate4sd3_1
XFILLER_29_33 VPWR VGND sg13g2_fill_1
Xhold11 hold11/A VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold55 hold55/A VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold44 hold44/A VPWR VGND net241 sg13g2_dlygate4sd3_1
Xhold33 hold33/A VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_654 VPWR VGND sg13g2_decap_8
Xhold66 hold66/A VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold99 hold99/A VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold77 hold77/A VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold88 hold88/A VPWR VGND net285 sg13g2_dlygate4sd3_1
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_613 VPWR VGND sg13g2_decap_8
XFILLER_17_816 VPWR VGND sg13g2_decap_8
XFILLER_32_808 VPWR VGND sg13g2_decap_8
XFILLER_40_863 VPWR VGND sg13g2_decap_8
XFILLER_8_525 VPWR VGND sg13g2_decap_8
XFILLER_12_565 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0740_ u_ppwm_u_mem__0739_/Y VPWR u_ppwm_u_mem__1228_/D VGND net603
+ u_ppwm_u_mem__0737_/D sg13g2_o21ai_1
Xu_ppwm_u_mem__0671_ VPWR u_ppwm_u_mem__0671_/Y net256 VGND sg13g2_inv_1
XFILLER_4_720 VPWR VGND sg13g2_decap_8
XFILLER_10_90 VPWR VGND sg13g2_fill_2
XFILLER_4_797 VPWR VGND sg13g2_decap_8
XFILLER_0_981 VPWR VGND sg13g2_decap_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1223_ net132 VGND VPWR u_ppwm_u_mem__1223_/D hold259/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_47_451 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__640_ net426 VPWR u_ppwm_u_ex__640_/Y VGND net398 fanout310/A sg13g2_o21ai_1
XFILLER_35_624 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1154_ net172 VGND VPWR net248 hold112/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__829__43 VPWR VGND net43 sg13g2_tiehi
Xu_ppwm_u_ex__571_ net327 net325 u_ppwm_u_ex__594_/B VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__1085_ u_ppwm_u_mem__1103_/A net423 u_ppwm_u_mem__1085_/B VPWR VGND
+ sg13g2_nand2_2
XFILLER_23_819 VPWR VGND sg13g2_decap_8
XFILLER_16_882 VPWR VGND sg13g2_decap_8
XFILLER_31_830 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0938_ net444 VPWR u_ppwm_u_mem__0938_/Y VGND net366 net280 sg13g2_o21ai_1
XFILLER_7_580 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0869_ VGND VPWR net362 u_ppwm_u_mem__0720_/Y hold190/A u_ppwm_u_mem__0868_/Y
+ sg13g2_a21oi_1
XFILLER_39_996 VPWR VGND sg13g2_decap_8
XFILLER_26_657 VPWR VGND sg13g2_decap_8
XFILLER_41_605 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__769_ VPWR u_ppwm_u_ex__769_/Y u_ppwm_u_ex__787_/A VGND sg13g2_inv_1
XFILLER_15_46 VPWR VGND sg13g2_fill_1
XFILLER_25_178 VPWR VGND sg13g2_decap_8
XFILLER_22_852 VPWR VGND sg13g2_decap_8
XFILLER_5_528 VPWR VGND sg13g2_decap_8
XFILLER_1_701 VPWR VGND sg13g2_decap_8
XFILLER_0_222 VPWR VGND sg13g2_decap_8
XFILLER_1_778 VPWR VGND sg13g2_decap_8
XFILLER_49_749 VPWR VGND sg13g2_decap_8
XFILLER_0_288 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_17_613 VPWR VGND sg13g2_decap_8
XFILLER_29_451 VPWR VGND sg13g2_fill_2
XFILLER_45_955 VPWR VGND sg13g2_decap_8
XFILLER_32_605 VPWR VGND sg13g2_decap_8
XFILLER_44_487 VPWR VGND sg13g2_decap_8
XFILLER_9_801 VPWR VGND sg13g2_decap_8
XFILLER_40_660 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_13_896 VPWR VGND sg13g2_decap_8
XFILLER_9_878 VPWR VGND sg13g2_decap_8
XFILLER_8_399 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0723_ VPWR u_ppwm_u_mem__0723_/Y net585 VGND sg13g2_inv_1
XFILLER_4_594 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0654_ VPWR u_ppwm_u_mem__0654_/Y net276 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1117__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_48_760 VPWR VGND sg13g2_decap_8
XFILLER_47_270 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1206_ net72 VGND VPWR u_ppwm_u_mem__1206_/D hold15/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_421 VPWR VGND sg13g2_decap_8
XFILLER_35_432 VPWR VGND sg13g2_fill_1
XFILLER_36_944 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1137_ net87 VGND VPWR net518 hold187/A clknet_5_30__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__623_ fanout309/A u_ppwm_u_ex__714_/B VPWR VGND net327 sg13g2_nand2b_2
Xheichips25_ppwm_5 VPWR VGND uio_oe[2] sg13g2_tielo
Xu_ppwm_u_ex__554_ u_ppwm_u_ex__553_/Y VPWR u_ppwm_u_ex__554_/Y VGND net397 u_ppwm_u_ex__440_/Y
+ sg13g2_o21ai_1
XFILLER_23_616 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1068_ net429 VPWR u_ppwm_u_mem__1068_/Y VGND net338 net477 sg13g2_o21ai_1
Xu_ppwm_u_ex__485_ u_ppwm_u_ex__485_/B u_ppwm_u_ex__485_/C u_ppwm_u_ex__485_/A u_ppwm_u_ex__485_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_11_1002 VPWR VGND sg13g2_decap_8
Xhold300 hold300/A VPWR VGND net643 sg13g2_dlygate4sd3_1
Xhold311 hold311/A VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold322 hold322/A VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold333 hold333/A VPWR VGND net676 sg13g2_dlygate4sd3_1
XFILLER_39_793 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_fill_2
XFILLER_42_958 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_6_804 VPWR VGND sg13g2_decap_8
XFILLER_5_325 VPWR VGND sg13g2_decap_8
XFILLER_1_575 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_37_708 VPWR VGND sg13g2_decap_8
XFILLER_18_933 VPWR VGND sg13g2_decap_8
XFILLER_45_752 VPWR VGND sg13g2_decap_8
XFILLER_17_487 VPWR VGND sg13g2_decap_8
XFILLER_33_925 VPWR VGND sg13g2_decap_8
XFILLER_20_608 VPWR VGND sg13g2_decap_8
XFILLER_34_1013 VPWR VGND sg13g2_decap_8
XFILLER_13_693 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1227__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_9_675 VPWR VGND sg13g2_decap_8
XFILLER_5_892 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0706_ VPWR u_ppwm_u_mem__0706_/Y net503 VGND sg13g2_inv_1
XFILLER_4_391 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0637_ VPWR u_ppwm_u_mem__0637_/Y net258 VGND sg13g2_inv_1
XFILLER_27_207 VPWR VGND sg13g2_decap_8
XFILLER_36_741 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__606_ VGND VPWR u_ppwm_u_ex__417_/Y hold243/A u_ppwm_u_ex__606_/Y u_ppwm_u_ex__605_/Y
+ sg13g2_a21oi_1
XFILLER_24_958 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__537_ u_ppwm_u_ex__519_/Y VPWR u_ppwm_u_ex__543_/A VGND u_ppwm_u_ex__520_/Y
+ u_ppwm_u_ex__536_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__468_ u_ppwm_u_ex__468_/A u_ppwm_u_ex__468_/B u_ppwm_u_ex__469_/C VPWR
+ VGND sg13g2_nor2_1
XFILLER_12_25 VPWR VGND sg13g2_decap_8
Xhold141 hold141/A VPWR VGND net484 sg13g2_dlygate4sd3_1
XFILLER_2_317 VPWR VGND sg13g2_decap_8
Xhold130 hold130/A VPWR VGND net473 sg13g2_dlygate4sd3_1
Xhold152 hold152/A VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold174 hold174/A VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold185 hold185/A VPWR VGND net528 sg13g2_dlygate4sd3_1
Xhold163 hold163/A VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold196 hold196/A VPWR VGND net539 sg13g2_dlygate4sd3_1
XFILLER_19_719 VPWR VGND sg13g2_decap_8
XFILLER_37_11 VPWR VGND sg13g2_fill_1
XFILLER_39_590 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_37_99 VPWR VGND sg13g2_decap_8
XFILLER_15_914 VPWR VGND sg13g2_decap_8
XFILLER_42_755 VPWR VGND sg13g2_decap_8
XFILLER_26_295 VPWR VGND sg13g2_fill_1
XFILLER_41_243 VPWR VGND sg13g2_decap_8
XFILLER_14_457 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__230_ net181 VGND VPWR net305 hold107/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__161_ net425 VPWR u_ppwm_u_pwm__161_/Y VGND hold308/A net329 sg13g2_o21ai_1
XFILLER_6_601 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_678 VPWR VGND sg13g2_decap_8
XFILLER_5_177 VPWR VGND sg13g2_fill_1
XFILLER_2_884 VPWR VGND sg13g2_decap_8
XFILLER_1_372 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
XFILLER_18_730 VPWR VGND sg13g2_decap_8
XFILLER_33_722 VPWR VGND sg13g2_decap_8
XFILLER_21_906 VPWR VGND sg13g2_decap_8
XFILLER_33_799 VPWR VGND sg13g2_decap_8
XFILLER_13_490 VPWR VGND sg13g2_decap_8
XFILLER_9_472 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__810__30 VPWR VGND net30 sg13g2_tiehi
Xheichips25_ppwm_15 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_24_755 VPWR VGND sg13g2_decap_8
XFILLER_11_449 VPWR VGND sg13g2_decap_8
XFILLER_20_972 VPWR VGND sg13g2_decap_8
XFILLER_2_125 VPWR VGND sg13g2_fill_2
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 net442 net440 VPWR VGND sg13g2_buf_8
Xfanout451 net452 net451 VPWR VGND sg13g2_buf_8
XFILLER_47_836 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_19_516 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_42_552 VPWR VGND sg13g2_decap_8
XFILLER_15_788 VPWR VGND sg13g2_decap_8
XFILLER_14_287 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0971_ VGND VPWR net356 u_ppwm_u_mem__0669_/Y hold86/A u_ppwm_u_mem__0970_/Y
+ sg13g2_a21oi_1
XFILLER_30_769 VPWR VGND sg13g2_decap_8
XFILLER_31_1005 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__213_ u_ppwm_u_pwm__214_/B hold278/A u_ppwm_u_pwm__212_/Y u_ppwm_u_pwm__215_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_7_965 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__144_ VGND VPWR u_ppwm_u_pwm__138_/Y net328 hold4/A u_ppwm_u_pwm__143_/Y
+ sg13g2_a21oi_1
XFILLER_6_475 VPWR VGND sg13g2_decap_8
XFILLER_2_681 VPWR VGND sg13g2_decap_8
XFILLER_49_140 VPWR VGND sg13g2_decap_8
XFILLER_1_191 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__093_ net331 u_ppwm_u_global_counter__095_/C net552 u_ppwm_u_global_counter__093_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_38_858 VPWR VGND sg13g2_decap_8
XFILLER_21_703 VPWR VGND sg13g2_decap_8
XFILLER_33_596 VPWR VGND sg13g2_decap_8
XFILLER_18_13 VPWR VGND sg13g2_decap_8
XFILLER_29_836 VPWR VGND sg13g2_decap_8
XFILLER_28_379 VPWR VGND sg13g2_fill_1
XFILLER_24_552 VPWR VGND sg13g2_decap_8
XFILLER_12_747 VPWR VGND sg13g2_decap_8
XFILLER_8_707 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_5_1__leaf_clk clkload0/X VPWR VGND sg13g2_buf_1
XFILLER_4_902 VPWR VGND sg13g2_decap_8
XFILLER_4_979 VPWR VGND sg13g2_decap_8
XFILLER_3_467 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_633 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1170_ net134 VGND VPWR net468 hold144/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_806 VPWR VGND sg13g2_decap_8
XFILLER_46_187 VPWR VGND sg13g2_fill_2
XFILLER_43_894 VPWR VGND sg13g2_decap_8
XFILLER_15_585 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0954_ net444 VPWR u_ppwm_u_mem__0954_/Y VGND net366 hold112/A sg13g2_o21ai_1
XFILLER_30_566 VPWR VGND sg13g2_decap_8
XFILLER_7_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0885_ VGND VPWR net359 u_ppwm_u_mem__0712_/Y hold149/A u_ppwm_u_mem__0884_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__127_ VPWR u_ppwm_u_pwm__127_/Y hold268/A VGND sg13g2_inv_1
XFILLER_38_655 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__785_ u_ppwm_u_ex__785_/A u_ppwm_u_ex__785_/B u_ppwm_u_ex__785_/C u_ppwm_u_ex__785_/D
+ u_ppwm_u_ex__785_/Y VPWR VGND sg13g2_nor4_1
XFILLER_26_839 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__076_ VGND VPWR net202 u_ppwm_u_global_counter__073_/B hold119/A
+ net461 sg13g2_a21oi_1
XFILLER_1_93 VPWR VGND sg13g2_fill_1
XFILLER_19_880 VPWR VGND sg13g2_decap_8
XFILLER_21_500 VPWR VGND sg13g2_decap_8
XFILLER_34_894 VPWR VGND sg13g2_decap_8
XFILLER_21_577 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1127__107 VPWR VGND net107 sg13g2_tiehi
Xhold12 hold12/A VPWR VGND net209 sg13g2_dlygate4sd3_1
Xhold23 hold23/A VPWR VGND net220 sg13g2_dlygate4sd3_1
Xhold56 hold56/A VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold45 hold45/A VPWR VGND net242 sg13g2_dlygate4sd3_1
Xhold34 hold34/A VPWR VGND net231 sg13g2_dlygate4sd3_1
Xhold67 hold67/A VPWR VGND net264 sg13g2_dlygate4sd3_1
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
XFILLER_28_132 VPWR VGND sg13g2_fill_2
XFILLER_29_633 VPWR VGND sg13g2_decap_8
Xhold89 hold89/A VPWR VGND net286 sg13g2_dlygate4sd3_1
Xhold78 hold78/A VPWR VGND net275 sg13g2_dlygate4sd3_1
XFILLER_28_143 VPWR VGND sg13g2_fill_1
XFILLER_45_44 VPWR VGND sg13g2_decap_4
XFILLER_16_316 VPWR VGND sg13g2_decap_4
XFILLER_44_669 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_4
XFILLER_40_842 VPWR VGND sg13g2_decap_8
XFILLER_8_504 VPWR VGND sg13g2_decap_8
XFILLER_12_544 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0670_ VPWR u_ppwm_u_mem__0670_/Y net559 VGND sg13g2_inv_1
XFILLER_4_776 VPWR VGND sg13g2_decap_8
XFILLER_0_960 VPWR VGND sg13g2_decap_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
XFILLER_47_430 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1222_ net171 VGND VPWR u_ppwm_u_mem__1222_/D hold281/A clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_mem__1153_ net55 VGND VPWR net456 hold114/A clknet_5_27__leaf_clk sg13g2_dfrbpq_2
XFILLER_35_603 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__570_ u_ppwm_u_ex__569_/Y VPWR u_ppwm_u_ex__573_/A VGND u_ppwm_u_ex__565_/Y
+ u_ppwm_u_ex__568_/Y sg13g2_o21ai_1
XFILLER_16_861 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1084_ u_ppwm_u_mem__1085_/B net513 VPWR VGND net338 sg13g2_nand2b_2
XFILLER_43_691 VPWR VGND sg13g2_decap_8
XFILLER_31_886 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0937_ VGND VPWR net366 u_ppwm_u_mem__0686_/Y hold84/A u_ppwm_u_mem__0936_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0868_ net448 VPWR u_ppwm_u_mem__0868_/Y VGND net362 net527 sg13g2_o21ai_1
Xu_ppwm_u_mem__1189__58 VPWR VGND net58 sg13g2_tiehi
Xu_ppwm_u_mem__1196__149 VPWR VGND net149 sg13g2_tiehi
Xu_ppwm_u_mem__0799_ u_ppwm_u_mem__0799_/Y net405 u_ppwm_u_mem__0799_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_975 VPWR VGND sg13g2_decap_8
XFILLER_26_636 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__059_ VPWR u_ppwm_u_global_counter__075_/A net336 VGND sg13g2_inv_1
Xu_ppwm_u_ex__768_ net321 VPWR u_ppwm_u_ex__787_/A VGND net381 hold293/A sg13g2_o21ai_1
XFILLER_25_135 VPWR VGND sg13g2_decap_8
XFILLER_25_146 VPWR VGND sg13g2_fill_1
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_15_36 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__699_ VGND VPWR u_ppwm_u_ex__664_/B u_ppwm_u_ex__696_/Y u_ppwm_u_ex__699_/Y
+ u_ppwm_u_ex__698_/Y sg13g2_a21oi_1
XFILLER_22_831 VPWR VGND sg13g2_decap_8
XFILLER_34_691 VPWR VGND sg13g2_decap_8
XFILLER_5_507 VPWR VGND sg13g2_decap_8
XFILLER_0_201 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_fill_2
XFILLER_1_757 VPWR VGND sg13g2_decap_8
XFILLER_49_728 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_45_934 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_decap_8
XFILLER_44_466 VPWR VGND sg13g2_decap_8
XFILLER_44_444 VPWR VGND sg13g2_fill_2
XFILLER_17_669 VPWR VGND sg13g2_decap_8
XFILLER_13_875 VPWR VGND sg13g2_decap_8
XFILLER_8_334 VPWR VGND sg13g2_decap_8
XFILLER_9_857 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0722_ VPWR u_ppwm_u_mem__0722_/Y net501 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0653_ VPWR u_ppwm_u_mem__0653_/Y net278 VGND sg13g2_inv_1
XFILLER_4_573 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1205_ net80 VGND VPWR net213 hold65/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_923 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_6 VPWR VGND uio_oe[3] sg13g2_tielo
Xu_ppwm_u_ex__622_ u_ppwm/instr\[2\] net327 u_ppwm_u_ex__622_/C fanout310/A VPWR VGND
+ sg13g2_nor3_2
Xu_ppwm_u_mem__1136_ net89 VGND VPWR net531 hold232/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__553_ u_ppwm_u_ex__553_/Y hold203/A net395 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1067_ VGND VPWR net339 u_ppwm_u_mem__0621_/Y hold135/A u_ppwm_u_mem__1066_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__484_ VGND VPWR u_ppwm_u_ex__485_/A u_ppwm_u_ex__485_/B u_ppwm_u_ex__486_/B
+ u_ppwm_u_ex__485_/C sg13g2_a21oi_1
XFILLER_31_683 VPWR VGND sg13g2_decap_8
Xhold301 hold301/A VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold312 hold312/A VPWR VGND net655 sg13g2_dlygate4sd3_1
Xhold323 hold323/A VPWR VGND net666 sg13g2_dlygate4sd3_1
XFILLER_39_772 VPWR VGND sg13g2_decap_8
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_26_57 VPWR VGND sg13g2_fill_1
XFILLER_38_293 VPWR VGND sg13g2_fill_1
XFILLER_42_937 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
XFILLER_41_458 VPWR VGND sg13g2_fill_1
XFILLER_42_34 VPWR VGND sg13g2_fill_1
XFILLER_9_109 VPWR VGND sg13g2_fill_2
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_21_182 VPWR VGND sg13g2_fill_2
XFILLER_21_193 VPWR VGND sg13g2_fill_2
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_1_554 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_18_912 VPWR VGND sg13g2_decap_8
XFILLER_45_731 VPWR VGND sg13g2_decap_8
XFILLER_33_904 VPWR VGND sg13g2_decap_8
XFILLER_17_466 VPWR VGND sg13g2_decap_8
XFILLER_18_989 VPWR VGND sg13g2_decap_8
XFILLER_32_447 VPWR VGND sg13g2_fill_2
XFILLER_13_672 VPWR VGND sg13g2_decap_8
XFILLER_9_654 VPWR VGND sg13g2_decap_8
XFILLER_5_871 VPWR VGND sg13g2_decap_8
XFILLER_4_370 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0705_ VPWR u_ppwm_u_mem__0705_/Y net537 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0636_ VPWR u_ppwm_u_mem__0636_/Y net245 VGND sg13g2_inv_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__227__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_36_720 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1182__86 VPWR VGND net86 sg13g2_tiehi
Xu_ppwm_u_ex__605_ u_ppwm_u_ex__605_/A u_ppwm_u_ex__604_/A u_ppwm_u_ex__605_/Y VPWR
+ VGND sg13g2_nor2b_1
XFILLER_24_937 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1119_ net123 VGND VPWR net492 hold126/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_797 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__536_ VPWR VGND u_ppwm_u_ex__528_/Y u_ppwm_u_ex__535_/Y u_ppwm_u_ex__534_/Y
+ u_ppwm_u_ex__534_/B u_ppwm_u_ex__536_/Y u_ppwm_u_ex__532_/Y sg13g2_a221oi_1
XFILLER_23_469 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__467_ u_ppwm_u_ex__468_/A u_ppwm_u_ex__468_/B u_ppwm_u_ex__469_/B VPWR
+ VGND sg13g2_and2_1
Xhold120 hold120/A VPWR VGND net463 sg13g2_dlygate4sd3_1
XFILLER_2_307 VPWR VGND sg13g2_fill_1
Xhold153 hold153/A VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold131 hold131/A VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold142 hold142/A VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold175 hold175/A VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold186 hold186/A VPWR VGND net529 sg13g2_dlygate4sd3_1
Xhold164 hold164/A VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold197 hold197/A VPWR VGND net540 sg13g2_dlygate4sd3_1
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_37_45 VPWR VGND sg13g2_fill_1
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_42_734 VPWR VGND sg13g2_decap_8
XFILLER_14_436 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__160_ VGND VPWR u_ppwm_u_pwm__218_/B net330 hold68/A u_ppwm_u_pwm__159_/Y
+ sg13g2_a21oi_1
XFILLER_5_112 VPWR VGND sg13g2_fill_2
XFILLER_6_657 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_2_863 VPWR VGND sg13g2_decap_8
XFILLER_1_351 VPWR VGND sg13g2_decap_8
XFILLER_49_322 VPWR VGND sg13g2_decap_8
XFILLER_49_399 VPWR VGND sg13g2_decap_8
XFILLER_18_786 VPWR VGND sg13g2_decap_8
XFILLER_33_701 VPWR VGND sg13g2_decap_8
XFILLER_32_222 VPWR VGND sg13g2_decap_8
XFILLER_33_778 VPWR VGND sg13g2_decap_8
XFILLER_9_451 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0619_ VPWR u_ppwm_u_mem__0619_/Y net233 VGND sg13g2_inv_1
Xheichips25_ppwm_16 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_43_509 VPWR VGND sg13g2_decap_8
XFILLER_24_734 VPWR VGND sg13g2_decap_8
XFILLER_36_594 VPWR VGND sg13g2_decap_8
XFILLER_12_929 VPWR VGND sg13g2_decap_8
XFILLER_23_233 VPWR VGND sg13g2_fill_1
XFILLER_11_428 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__519_ u_ppwm_u_ex__519_/Y u_ppwm_u_ex__519_/A net388 VPWR VGND sg13g2_nand2_1
XFILLER_23_266 VPWR VGND sg13g2_fill_2
XFILLER_20_951 VPWR VGND sg13g2_decap_8
XFILLER_3_649 VPWR VGND sg13g2_decap_8
Xfanout430 net431 net430 VPWR VGND sg13g2_buf_8
Xfanout441 net442 net441 VPWR VGND sg13g2_buf_8
XFILLER_47_815 VPWR VGND sg13g2_decap_8
Xfanout452 rst_n net452 VPWR VGND sg13g2_buf_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_34_509 VPWR VGND sg13g2_fill_1
XFILLER_42_531 VPWR VGND sg13g2_decap_8
XFILLER_9_27 VPWR VGND sg13g2_decap_4
XFILLER_15_767 VPWR VGND sg13g2_decap_8
XFILLER_30_748 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0970_ net435 VPWR u_ppwm_u_mem__0970_/Y VGND net356 hold216/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__212_ hold25/A hold300/A u_ppwm_u_pwm__212_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_7_944 VPWR VGND sg13g2_decap_8
XFILLER_11_995 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_6_454 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__143_ net424 VPWR u_ppwm_u_pwm__143_/Y VGND hold306/A net328 sg13g2_o21ai_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_2_660 VPWR VGND sg13g2_decap_8
XFILLER_9_1018 VPWR VGND sg13g2_decap_8
XFILLER_37_303 VPWR VGND sg13g2_fill_1
XFILLER_38_837 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__092_ VGND VPWR net331 u_ppwm_u_global_counter__095_/C hold210/A
+ net552 sg13g2_a21oi_1
XFILLER_18_583 VPWR VGND sg13g2_decap_8
XFILLER_33_575 VPWR VGND sg13g2_decap_8
XFILLER_21_759 VPWR VGND sg13g2_decap_8
XFILLER_9_281 VPWR VGND sg13g2_decap_4
XFILLER_29_815 VPWR VGND sg13g2_decap_8
XFILLER_24_531 VPWR VGND sg13g2_decap_8
XFILLER_11_203 VPWR VGND sg13g2_fill_1
XFILLER_12_726 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_5_3__leaf_clk clkload1/X VPWR VGND sg13g2_buf_1
XFILLER_4_958 VPWR VGND sg13g2_decap_8
XFILLER_3_446 VPWR VGND sg13g2_decap_8
XFILLER_47_612 VPWR VGND sg13g2_decap_8
XFILLER_19_314 VPWR VGND sg13g2_decap_8
XFILLER_47_689 VPWR VGND sg13g2_decap_8
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_15_564 VPWR VGND sg13g2_decap_8
XFILLER_30_545 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0953_ VGND VPWR net369 u_ppwm_u_mem__0678_/Y hold113/A u_ppwm_u_mem__0952_/Y
+ sg13g2_a21oi_1
XFILLER_10_280 VPWR VGND sg13g2_decap_8
XFILLER_7_741 VPWR VGND sg13g2_decap_8
XFILLER_11_792 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__126_ VPWR u_ppwm_u_pwm__126_/Y net580 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0884_ net448 VPWR u_ppwm_u_mem__0884_/Y VGND net359 net469 sg13g2_o21ai_1
XFILLER_38_634 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__075_ u_ppwm_u_global_counter__075_/A u_ppwm_u_global_counter__085_/A
+ u_ppwm_u_global_counter__085_/B u_ppwm_u_global_counter__082_/D VPWR VGND sg13g2_nor3_2
Xu_ppwm_u_ex__784_ VGND VPWR u_ppwm_u_ex__781_/Y u_ppwm_u_ex__782_/Y u_ppwm_u_ex__824_/D
+ u_ppwm_u_ex__783_/Y sg13g2_a21oi_1
XFILLER_26_818 VPWR VGND sg13g2_decap_8
XFILLER_34_873 VPWR VGND sg13g2_decap_8
XFILLER_21_556 VPWR VGND sg13g2_decap_8
XFILLER_1_939 VPWR VGND sg13g2_decap_8
XFILLER_0_449 VPWR VGND sg13g2_decap_8
Xhold13 hold13/A VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold46 hold46/A VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold24 hold24/A VPWR VGND net221 sg13g2_dlygate4sd3_1
XFILLER_29_612 VPWR VGND sg13g2_decap_8
Xhold35 hold35/A VPWR VGND net232 sg13g2_dlygate4sd3_1
Xhold79 hold79/A VPWR VGND net276 sg13g2_dlygate4sd3_1
Xhold68 hold68/A VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold57 hold57/A VPWR VGND net254 sg13g2_dlygate4sd3_1
XFILLER_29_689 VPWR VGND sg13g2_decap_8
XFILLER_44_648 VPWR VGND sg13g2_decap_8
XFILLER_40_821 VPWR VGND sg13g2_decap_8
XFILLER_25_884 VPWR VGND sg13g2_decap_8
XFILLER_12_523 VPWR VGND sg13g2_decap_8
XFILLER_40_898 VPWR VGND sg13g2_decap_8
XFILLER_4_755 VPWR VGND sg13g2_decap_8
XFILLER_48_921 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1221_ net84 VGND VPWR net584 hold239/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_998 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1152_ net57 VGND VPWR u_ppwm_u_mem__1152_/D hold100/A clknet_5_30__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_47_486 VPWR VGND sg13g2_decap_8
XFILLER_16_840 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1083_ VGND VPWR u_ppwm_u_mem__0730_/A net339 u_ppwm_u_mem__1218_/D
+ u_ppwm_u_mem__1082_/Y sg13g2_a21oi_1
XFILLER_34_125 VPWR VGND sg13g2_fill_2
XFILLER_35_659 VPWR VGND sg13g2_decap_8
XFILLER_43_670 VPWR VGND sg13g2_decap_8
XFILLER_15_361 VPWR VGND sg13g2_fill_1
XFILLER_37_1023 VPWR VGND sg13g2_decap_4
XFILLER_31_865 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0936_ net446 VPWR u_ppwm_u_mem__0936_/Y VGND net366 hold123/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0867_ VGND VPWR net370 u_ppwm_u_mem__0721_/Y u_ppwm_u_mem__1110_/D
+ u_ppwm_u_mem__0866_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0798_ hold167/A hold165/A net414 u_ppwm_u_mem__0799_/B VPWR VGND sg13g2_mux2_1
XFILLER_44_1005 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_39_954 VPWR VGND sg13g2_decap_8
XFILLER_26_615 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__058_ VPWR u_ppwm_u_global_counter__058_/Y net564 VGND sg13g2_inv_1
Xu_ppwm_u_ex__767_ u_ppwm_u_ex__785_/C net380 net321 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__698_ u_ppwm_u_ex__698_/Y u_ppwm_u_ex__698_/A u_ppwm_u_ex__698_/B VPWR
+ VGND sg13g2_nand2_1
XFILLER_22_810 VPWR VGND sg13g2_decap_8
XFILLER_34_670 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__237__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_22_887 VPWR VGND sg13g2_decap_8
XFILLER_1_736 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_45_913 VPWR VGND sg13g2_decap_8
XFILLER_17_648 VPWR VGND sg13g2_decap_8
XFILLER_16_158 VPWR VGND sg13g2_fill_2
XFILLER_16_169 VPWR VGND sg13g2_fill_1
XFILLER_13_854 VPWR VGND sg13g2_decap_8
XFILLER_25_681 VPWR VGND sg13g2_decap_8
XFILLER_9_836 VPWR VGND sg13g2_decap_8
XFILLER_40_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0721_ VPWR u_ppwm_u_mem__0721_/Y net527 VGND sg13g2_inv_1
XFILLER_4_552 VPWR VGND sg13g2_decap_8
XFILLER_21_91 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0652_ VPWR u_ppwm_u_mem__0652_/Y net510 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1204_ net88 VGND VPWR net263 hold146/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_902 VPWR VGND sg13g2_decap_8
XFILLER_48_795 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__621_ u_ppwm/instr\[2\] u_ppwm_u_ex__622_/C u_ppwm_u_ex__714_/B VPWR
+ VGND sg13g2_nor2_2
XFILLER_47_294 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1135_ net91 VGND VPWR u_ppwm_u_mem__1135_/D hold38/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_979 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__552_ VPWR VGND u_ppwm_u_ex__550_/Y u_ppwm_u_ex__551_/Y u_ppwm_u_ex__549_/Y
+ net397 u_ppwm_u_ex__552_/Y u_ppwm_u_ex__440_/Y sg13g2_a221oi_1
Xu_ppwm_u_mem__1066_ net423 VPWR u_ppwm_u_mem__1066_/Y VGND net339 hold191/A sg13g2_o21ai_1
Xheichips25_ppwm_7 VPWR VGND uio_oe[4] sg13g2_tielo
Xu_ppwm_u_ex__817__37 VPWR VGND net37 sg13g2_tiehi
Xu_ppwm_u_ex__483_ u_ppwm_u_ex__485_/C net400 net320 VPWR VGND sg13g2_xnor2_1
XFILLER_31_662 VPWR VGND sg13g2_decap_8
Xhold302 hold302/A VPWR VGND net645 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0919_ VGND VPWR net365 u_ppwm_u_mem__0695_/Y hold188/A u_ppwm_u_mem__0918_/Y
+ sg13g2_a21oi_1
Xhold313 hold313/A VPWR VGND net656 sg13g2_dlygate4sd3_1
Xhold324 hold324/A VPWR VGND net667 sg13g2_dlygate4sd3_1
XFILLER_39_751 VPWR VGND sg13g2_decap_8
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_38_272 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__819_ net29 VGND VPWR u_ppwm_u_ex__819_/D hold315/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_42_916 VPWR VGND sg13g2_decap_8
XFILLER_14_618 VPWR VGND sg13g2_decap_8
XFILLER_26_489 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_22_684 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_6_839 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_1_533 VPWR VGND sg13g2_decap_8
XFILLER_49_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_45_710 VPWR VGND sg13g2_decap_8
XFILLER_17_445 VPWR VGND sg13g2_decap_8
XFILLER_18_968 VPWR VGND sg13g2_decap_8
XFILLER_45_787 VPWR VGND sg13g2_decap_8
XFILLER_13_651 VPWR VGND sg13g2_decap_8
XFILLER_9_633 VPWR VGND sg13g2_decap_8
XFILLER_5_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0704_ VPWR u_ppwm_u_mem__0704_/Y net479 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0635_ VPWR u_ppwm_u_mem__0635_/Y net210 VGND sg13g2_inv_1
XFILLER_48_592 VPWR VGND sg13g2_decap_8
XFILLER_35_220 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__604_ u_ppwm_u_ex__605_/A u_ppwm_u_ex__604_/C u_ppwm_u_ex__604_/A u_ppwm_u_ex__604_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_24_916 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1118_ net125 VGND VPWR net470 hold121/A clknet_5_23__leaf_clk sg13g2_dfrbpq_2
XFILLER_36_776 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__535_ net380 net390 u_ppwm_u_ex__535_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_23_448 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1049_ VGND VPWR net354 u_ppwm_u_mem__0630_/Y hold99/A u_ppwm_u_mem__1048_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__466_ u_ppwm_u_ex__468_/B net415 fanout327/A VPWR VGND sg13g2_nand2_1
XFILLER_31_492 VPWR VGND sg13g2_fill_1
Xhold110 hold110/A VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold132 hold132/A VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold121 hold121/A VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold143 hold143/A VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold176 hold176/A VPWR VGND net519 sg13g2_dlygate4sd3_1
Xhold154 hold154/A VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold165 hold165/A VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold187 hold187/A VPWR VGND net530 sg13g2_dlygate4sd3_1
Xhold198 hold198/A VPWR VGND net541 sg13g2_dlygate4sd3_1
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_2_1024 VPWR VGND sg13g2_decap_4
XFILLER_26_231 VPWR VGND sg13g2_decap_8
XFILLER_42_713 VPWR VGND sg13g2_decap_8
XFILLER_14_415 VPWR VGND sg13g2_decap_8
XFILLER_15_949 VPWR VGND sg13g2_decap_8
XFILLER_26_286 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_22_481 VPWR VGND sg13g2_decap_8
XFILLER_6_636 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_135 VPWR VGND sg13g2_fill_1
XFILLER_2_842 VPWR VGND sg13g2_decap_8
XFILLER_1_330 VPWR VGND sg13g2_decap_8
XFILLER_49_301 VPWR VGND sg13g2_decap_8
XFILLER_49_378 VPWR VGND sg13g2_decap_8
XFILLER_18_765 VPWR VGND sg13g2_decap_8
XFILLER_45_584 VPWR VGND sg13g2_decap_8
XFILLER_33_757 VPWR VGND sg13g2_decap_8
XFILLER_14_982 VPWR VGND sg13g2_decap_8
XFILLER_9_430 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0618_ VPWR u_ppwm_u_mem__0618_/Y net543 VGND sg13g2_inv_1
Xheichips25_ppwm_17 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_28_529 VPWR VGND sg13g2_decap_8
XFILLER_24_713 VPWR VGND sg13g2_decap_8
XFILLER_36_573 VPWR VGND sg13g2_decap_8
XFILLER_12_908 VPWR VGND sg13g2_decap_8
XFILLER_11_407 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__518_ VGND VPWR u_ppwm_u_ex__508_/Y u_ppwm_u_ex__515_/Y u_ppwm_u_ex__518_/Y
+ u_ppwm_u_ex__517_/Y sg13g2_a21oi_1
XFILLER_20_930 VPWR VGND sg13g2_decap_8
XFILLER_23_48 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__449_ u_ppwm_u_ex__449_/Y net377 u_ppwm_u_ex__448_/Y VPWR VGND sg13g2_nand2b_1
XFILLER_3_628 VPWR VGND sg13g2_decap_8
Xfanout420 net421 net420 VPWR VGND sg13g2_buf_2
Xfanout431 net432 net431 VPWR VGND sg13g2_buf_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_24_1014 VPWR VGND sg13g2_decap_8
Xfanout442 net452 net442 VPWR VGND sg13g2_buf_8
XFILLER_42_510 VPWR VGND sg13g2_decap_8
XFILLER_15_746 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_14_256 VPWR VGND sg13g2_decap_4
XFILLER_42_587 VPWR VGND sg13g2_decap_8
XFILLER_30_727 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__211_ u_ppwm_u_pwm__215_/A u_ppwm_u_pwm__215_/B u_ppwm_u_pwm__211_/Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_7_923 VPWR VGND sg13g2_decap_8
XFILLER_11_974 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_6_433 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__142_ u_ppwm_u_pwm__185_/A u_ppwm_u_pwm__142_/C u_ppwm_u_pwm__219_/A
+ fanout330/A VPWR VGND u_ppwm_u_pwm__142_/D sg13g2_nand4_1
XFILLER_49_175 VPWR VGND sg13g2_decap_8
XFILLER_38_816 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1137__87 VPWR VGND net87 sg13g2_tiehi
Xu_ppwm_u_global_counter__091_ hold273/A u_ppwm_u_global_counter__095_/C net331 u_ppwm_u_global_counter__088_/Y
+ u_ppwm_u_global_counter__055_/Y VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1152__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_18_562 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
XFILLER_33_554 VPWR VGND sg13g2_decap_8
XFILLER_21_738 VPWR VGND sg13g2_decap_8
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
XFILLER_24_510 VPWR VGND sg13g2_decap_8
XFILLER_12_705 VPWR VGND sg13g2_decap_8
XFILLER_24_587 VPWR VGND sg13g2_decap_8
XFILLER_34_69 VPWR VGND sg13g2_fill_2
XFILLER_11_226 VPWR VGND sg13g2_fill_1
Xclkload2 clknet_5_4__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_4_937 VPWR VGND sg13g2_decap_8
XFILLER_3_425 VPWR VGND sg13g2_decap_8
XFILLER_47_668 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_fill_1
XFILLER_28_893 VPWR VGND sg13g2_decap_8
XFILLER_43_852 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_30_524 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0952_ net445 VPWR u_ppwm_u_mem__0952_/Y VGND net369 hold114/A sg13g2_o21ai_1
XFILLER_7_720 VPWR VGND sg13g2_decap_8
XFILLER_11_771 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__125_ u_ppwm_u_pwm__185_/A net604 VPWR VGND sg13g2_inv_2
Xu_ppwm_u_mem__0883_ VGND VPWR net362 u_ppwm_u_mem__0713_/Y hold127/A u_ppwm_u_mem__0882_/Y
+ sg13g2_a21oi_1
XFILLER_7_797 VPWR VGND sg13g2_decap_8
XFILLER_3_992 VPWR VGND sg13g2_decap_8
XFILLER_34_4 VPWR VGND sg13g2_fill_2
XFILLER_38_613 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__074_ hold311/A net202 net268 u_ppwm_u_global_counter__085_/B
+ VPWR VGND net461 sg13g2_nand4_1
Xu_ppwm_u_ex__783_ net441 VPWR u_ppwm_u_ex__783_/Y VGND net653 net308 sg13g2_o21ai_1
XFILLER_37_134 VPWR VGND sg13g2_decap_4
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_25_318 VPWR VGND sg13g2_fill_2
XFILLER_25_329 VPWR VGND sg13g2_fill_1
XFILLER_34_852 VPWR VGND sg13g2_decap_8
XFILLER_33_351 VPWR VGND sg13g2_decap_8
XFILLER_21_535 VPWR VGND sg13g2_decap_8
XFILLER_33_395 VPWR VGND sg13g2_decap_4
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
XFILLER_20_49 VPWR VGND sg13g2_fill_1
XFILLER_1_918 VPWR VGND sg13g2_decap_8
XFILLER_0_428 VPWR VGND sg13g2_decap_8
Xhold14 hold14/A VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold47 hold47/A VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold25 hold25/A VPWR VGND net222 sg13g2_dlygate4sd3_1
Xhold36 hold36/A VPWR VGND net233 sg13g2_dlygate4sd3_1
Xhold69 hold69/A VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold58 hold58/A VPWR VGND net255 sg13g2_dlygate4sd3_1
XFILLER_29_668 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_4
XFILLER_44_627 VPWR VGND sg13g2_decap_8
XFILLER_40_800 VPWR VGND sg13g2_decap_8
XFILLER_12_502 VPWR VGND sg13g2_decap_8
XFILLER_25_863 VPWR VGND sg13g2_decap_8
XFILLER_40_877 VPWR VGND sg13g2_decap_8
XFILLER_12_579 VPWR VGND sg13g2_decap_8
XFILLER_8_539 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_4_734 VPWR VGND sg13g2_decap_8
XFILLER_48_900 VPWR VGND sg13g2_decap_8
XFILLER_0_995 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1220_ net116 VGND VPWR u_ppwm_u_mem__1220_/D hold276/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_47_465 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1151_ net59 VGND VPWR net298 hold205/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_638 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1082_ net423 VPWR u_ppwm_u_mem__1082_/Y VGND net206 net339 sg13g2_o21ai_1
XFILLER_28_690 VPWR VGND sg13g2_decap_8
XFILLER_37_1002 VPWR VGND sg13g2_decap_8
XFILLER_16_896 VPWR VGND sg13g2_decap_8
XFILLER_31_844 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0935_ VGND VPWR net365 u_ppwm_u_mem__0687_/Y u_ppwm_u_mem__1144_/D
+ u_ppwm_u_mem__0934_/Y sg13g2_a21oi_1
XFILLER_7_594 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0866_ net450 VPWR u_ppwm_u_mem__0866_/Y VGND net370 net501 sg13g2_o21ai_1
Xu_ppwm_u_mem__0797_ VGND VPWR net334 u_ppwm_u_mem__0796_/X u_ppwm_u_mem__0797_/Y
+ net333 sg13g2_a21oi_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_933 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__057_ VPWR u_ppwm_u_global_counter__057_/Y net614 VGND sg13g2_inv_1
Xu_ppwm_u_ex__766_ u_ppwm_u_ex__779_/A net380 net321 VPWR VGND sg13g2_nand2_1
XFILLER_41_619 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__697_ net318 VPWR u_ppwm_u_ex__698_/B VGND net387 net389 sg13g2_o21ai_1
XFILLER_33_181 VPWR VGND sg13g2_fill_1
XFILLER_22_866 VPWR VGND sg13g2_decap_8
XFILLER_21_365 VPWR VGND sg13g2_fill_2
XFILLER_1_715 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_decap_8
XFILLER_17_627 VPWR VGND sg13g2_decap_8
XFILLER_45_969 VPWR VGND sg13g2_decap_8
XFILLER_25_660 VPWR VGND sg13g2_decap_8
XFILLER_32_619 VPWR VGND sg13g2_decap_8
XFILLER_13_833 VPWR VGND sg13g2_decap_8
XFILLER_31_118 VPWR VGND sg13g2_fill_2
XFILLER_9_815 VPWR VGND sg13g2_decap_8
XFILLER_40_674 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0720_ VPWR u_ppwm_u_mem__0720_/Y net532 VGND sg13g2_inv_1
XFILLER_4_531 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0651_ VPWR u_ppwm_u_mem__0651_/Y net293 VGND sg13g2_inv_1
XFILLER_0_792 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1156__168 VPWR VGND net168 sg13g2_tiehi
Xu_ppwm_u_mem__1203_ net96 VGND VPWR net490 hold130/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_774 VPWR VGND sg13g2_decap_8
XFILLER_47_251 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__620_ u_ppwm_u_ex__622_/C net377 u_ppwm_u_ex__620_/B VPWR VGND sg13g2_nand2_1
XFILLER_47_284 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1134_ net93 VGND VPWR net236 hold57/A clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_958 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__551_ hold311/A net398 u_ppwm_u_ex__551_/Y VPWR VGND sg13g2_nor2b_1
Xheichips25_ppwm_8 VPWR VGND uio_oe[5] sg13g2_tielo
Xu_ppwm_u_mem__1065_ VGND VPWR net339 u_ppwm_u_mem__0622_/Y u_ppwm_u_mem__1209_/D
+ u_ppwm_u_mem__1064_/Y sg13g2_a21oi_1
XFILLER_35_468 VPWR VGND sg13g2_decap_4
XFILLER_44_991 VPWR VGND sg13g2_decap_8
XFILLER_16_693 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__482_ u_ppwm_u_ex__482_/A u_ppwm_u_ex__482_/B u_ppwm_u_ex__804_/D VPWR
+ VGND sg13g2_nor2_1
XFILLER_31_641 VPWR VGND sg13g2_decap_8
XFILLER_30_184 VPWR VGND sg13g2_decap_8
XFILLER_11_1016 VPWR VGND sg13g2_decap_8
XFILLER_11_1027 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0918_ net449 VPWR u_ppwm_u_mem__0918_/Y VGND net365 hold232/A sg13g2_o21ai_1
XFILLER_7_391 VPWR VGND sg13g2_decap_8
Xhold314 hold314/A VPWR VGND net657 sg13g2_dlygate4sd3_1
Xhold325 hold325/A VPWR VGND net668 sg13g2_dlygate4sd3_1
Xhold303 hold303/A VPWR VGND net646 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0849_ hold134/A hold9/A net410 u_ppwm_u_mem__0850_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__1185__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_27_903 VPWR VGND sg13g2_decap_8
XFILLER_39_730 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__109_ net438 VGND VPWR net547 hold203/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__818_ net33 VGND VPWR net642 hold328/A clknet_5_6__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__749_ net322 VPWR u_ppwm_u_ex__749_/Y VGND fanout383/A hold315/A sg13g2_o21ai_1
XFILLER_26_468 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_fill_2
XFILLER_42_58 VPWR VGND sg13g2_fill_1
XFILLER_21_140 VPWR VGND sg13g2_fill_1
XFILLER_22_663 VPWR VGND sg13g2_decap_8
XFILLER_6_818 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_5_339 VPWR VGND sg13g2_decap_8
XFILLER_1_512 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_589 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_decap_8
XFILLER_18_947 VPWR VGND sg13g2_decap_8
XFILLER_45_766 VPWR VGND sg13g2_decap_8
XFILLER_44_243 VPWR VGND sg13g2_fill_1
XFILLER_44_276 VPWR VGND sg13g2_fill_2
XFILLER_33_939 VPWR VGND sg13g2_decap_8
XFILLER_13_630 VPWR VGND sg13g2_decap_8
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_9_612 VPWR VGND sg13g2_decap_8
XFILLER_34_1027 VPWR VGND sg13g2_fill_2
XFILLER_8_188 VPWR VGND sg13g2_fill_2
XFILLER_9_689 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0703_ VPWR u_ppwm_u_mem__0703_/Y net500 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0634_ VPWR u_ppwm_u_mem__0634_/Y net266 VGND sg13g2_inv_1
XFILLER_48_571 VPWR VGND sg13g2_decap_8
XFILLER_36_755 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__603_ u_ppwm_u_ex__604_/C u_ppwm_u_ex__439_/Y net383 u_ppwm_u_ex__560_/B
+ net382 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1117_ net127 VGND VPWR net465 hold180/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__534_ u_ppwm_u_ex__534_/A u_ppwm_u_ex__534_/B u_ppwm_u_ex__534_/C u_ppwm_u_ex__534_/Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_17_991 VPWR VGND sg13g2_decap_8
XFILLER_23_427 VPWR VGND sg13g2_decap_8
XFILLER_16_490 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1048_ net433 VPWR u_ppwm_u_mem__1048_/Y VGND net354 hold115/A sg13g2_o21ai_1
Xu_ppwm_u_ex__465_ u_ppwm_u_ex__468_/A net407 net326 VPWR VGND sg13g2_xnor2_1
XFILLER_32_983 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
Xhold100 hold100/A VPWR VGND net297 sg13g2_dlygate4sd3_1
Xhold144 hold144/A VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold122 hold122/A VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold133 hold133/A VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold111 hold111/A VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold177 hold177/A VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold166 hold166/A VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold155 hold155/A VPWR VGND net498 sg13g2_dlygate4sd3_1
Xhold199 hold199/A VPWR VGND net542 sg13g2_dlygate4sd3_1
Xhold188 hold188/A VPWR VGND net531 sg13g2_dlygate4sd3_1
XFILLER_2_1003 VPWR VGND sg13g2_decap_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_15_928 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_42_769 VPWR VGND sg13g2_decap_8
XFILLER_30_909 VPWR VGND sg13g2_decap_8
XFILLER_22_460 VPWR VGND sg13g2_decap_8
XFILLER_23_994 VPWR VGND sg13g2_decap_8
XFILLER_6_615 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_5_114 VPWR VGND sg13g2_fill_1
XFILLER_2_821 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1149__63 VPWR VGND net63 sg13g2_tiehi
XFILLER_2_898 VPWR VGND sg13g2_decap_8
XFILLER_1_386 VPWR VGND sg13g2_decap_8
XFILLER_49_357 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1192__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_17_210 VPWR VGND sg13g2_fill_2
XFILLER_18_744 VPWR VGND sg13g2_decap_8
XFILLER_45_563 VPWR VGND sg13g2_decap_8
XFILLER_17_243 VPWR VGND sg13g2_decap_8
XFILLER_33_736 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
XFILLER_41_780 VPWR VGND sg13g2_decap_8
XFILLER_9_486 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0617_ VPWR u_ppwm_u_mem__0617_/Y net558 VGND sg13g2_inv_1
Xheichips25_ppwm_18 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_28_508 VPWR VGND sg13g2_decap_8
XFILLER_36_552 VPWR VGND sg13g2_decap_8
XFILLER_24_769 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__517_ u_ppwm_u_ex__517_/B u_ppwm_u_ex__517_/C net324 u_ppwm_u_ex__517_/Y
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__448_ u_ppwm/instr\[2\] net320 u_ppwm_u_ex__448_/C u_ppwm_u_ex__620_/B
+ u_ppwm_u_ex__448_/Y VPWR VGND sg13g2_nor4_1
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_32_780 VPWR VGND sg13g2_decap_8
XFILLER_20_986 VPWR VGND sg13g2_decap_8
XFILLER_3_607 VPWR VGND sg13g2_decap_8
Xfanout421 net672 net421 VPWR VGND sg13g2_buf_8
Xfanout410 net411 net410 VPWR VGND sg13g2_buf_8
Xfanout432 net436 net432 VPWR VGND sg13g2_buf_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
Xfanout443 net446 net443 VPWR VGND sg13g2_buf_8
XFILLER_14_213 VPWR VGND sg13g2_fill_1
XFILLER_15_725 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_4
XFILLER_42_566 VPWR VGND sg13g2_decap_8
XFILLER_30_706 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__210_ u_ppwm_u_pwm__210_/B u_ppwm_u_pwm__216_/B u_ppwm_u_pwm__210_/A
+ u_ppwm_u_pwm__215_/B VPWR VGND u_ppwm_u_pwm__210_/D sg13g2_nand4_1
XFILLER_23_791 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_7_902 VPWR VGND sg13g2_decap_8
XFILLER_11_953 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_31_1019 VPWR VGND sg13g2_decap_8
XFILLER_6_412 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__141_ hold237/A hold283/A hold300/A hold278/A u_ppwm_u_pwm__142_/D VPWR
+ VGND sg13g2_nor4_1
XFILLER_7_979 VPWR VGND sg13g2_decap_8
XFILLER_6_489 VPWR VGND sg13g2_decap_8
XFILLER_2_695 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__090_ u_ppwm_u_global_counter__095_/C net555 net615 hold318/A
+ VPWR VGND sg13g2_and3_2
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_18_541 VPWR VGND sg13g2_decap_8
XFILLER_33_533 VPWR VGND sg13g2_decap_8
XFILLER_21_717 VPWR VGND sg13g2_decap_8
XFILLER_9_250 VPWR VGND sg13g2_fill_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1215__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_44_809 VPWR VGND sg13g2_decap_8
XFILLER_28_349 VPWR VGND sg13g2_fill_2
XFILLER_36_360 VPWR VGND sg13g2_fill_1
XFILLER_36_371 VPWR VGND sg13g2_fill_2
XFILLER_37_883 VPWR VGND sg13g2_decap_8
XFILLER_24_566 VPWR VGND sg13g2_decap_8
XFILLER_7_209 VPWR VGND sg13g2_fill_2
Xclkload3 clknet_5_7__leaf_clk clkload3/X VPWR VGND sg13g2_buf_1
XFILLER_20_783 VPWR VGND sg13g2_decap_8
XFILLER_4_916 VPWR VGND sg13g2_decap_8
XFILLER_3_404 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1221__84 VPWR VGND net84 sg13g2_tiehi
XFILLER_47_647 VPWR VGND sg13g2_decap_8
XFILLER_19_338 VPWR VGND sg13g2_fill_2
XFILLER_28_872 VPWR VGND sg13g2_decap_8
XFILLER_43_831 VPWR VGND sg13g2_decap_8
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_15_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0951_ VGND VPWR net368 u_ppwm_u_mem__0679_/Y u_ppwm_u_mem__1152_/D
+ u_ppwm_u_mem__0950_/Y sg13g2_a21oi_1
XFILLER_11_750 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0882_ net448 VPWR u_ppwm_u_mem__0882_/Y VGND net362 net464 sg13g2_o21ai_1
XFILLER_7_776 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__124_ u_ppwm_u_pwm__219_/A net594 VPWR VGND sg13g2_inv_2
XFILLER_3_971 VPWR VGND sg13g2_decap_8
XFILLER_2_492 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__073_ u_ppwm_u_global_counter__073_/B net202 hold6/A VPWR
+ VGND sg13g2_xor2_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__782_ VPWR VGND net639 u_ppwm_u_ex__714_/Y fanout312/A net379 u_ppwm_u_ex__782_/Y
+ fanout314/A sg13g2_a221oi_1
XFILLER_38_669 VPWR VGND sg13g2_decap_8
XFILLER_19_894 VPWR VGND sg13g2_decap_8
XFILLER_18_393 VPWR VGND sg13g2_fill_2
XFILLER_34_831 VPWR VGND sg13g2_decap_8
XFILLER_21_514 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1166__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_407 VPWR VGND sg13g2_decap_8
Xhold26 hold26/A VPWR VGND net223 sg13g2_dlygate4sd3_1
Xhold37 hold37/A VPWR VGND net234 sg13g2_dlygate4sd3_1
XFILLER_29_59 VPWR VGND sg13g2_decap_4
Xhold15 hold15/A VPWR VGND net212 sg13g2_dlygate4sd3_1
Xhold59 hold59/A VPWR VGND net256 sg13g2_dlygate4sd3_1
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_fill_1
XFILLER_28_113 VPWR VGND sg13g2_decap_4
Xhold48 hold48/A VPWR VGND net245 sg13g2_dlygate4sd3_1
XFILLER_29_647 VPWR VGND sg13g2_decap_8
XFILLER_44_606 VPWR VGND sg13g2_decap_8
XFILLER_17_809 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_25_842 VPWR VGND sg13g2_decap_8
XFILLER_37_680 VPWR VGND sg13g2_decap_8
XFILLER_40_856 VPWR VGND sg13g2_decap_8
XFILLER_8_518 VPWR VGND sg13g2_decap_8
XFILLER_12_558 VPWR VGND sg13g2_decap_8
XFILLER_20_580 VPWR VGND sg13g2_decap_8
XFILLER_4_713 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_8
XFILLER_10_61 VPWR VGND sg13g2_fill_2
XFILLER_3_267 VPWR VGND sg13g2_fill_2
XFILLER_0_974 VPWR VGND sg13g2_decap_8
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_47_444 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1150_ net61 VGND VPWR u_ppwm_u_mem__1150_/D hold176/A clknet_5_31__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_19_124 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1081_ VGND VPWR u_ppwm_u_mem__0613_/Y net339 hold10/A u_ppwm_u_mem__1080_/Y
+ sg13g2_a21oi_1
XFILLER_35_617 VPWR VGND sg13g2_decap_8
XFILLER_16_875 VPWR VGND sg13g2_decap_8
XFILLER_30_322 VPWR VGND sg13g2_decap_4
XFILLER_31_823 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0934_ net445 VPWR u_ppwm_u_mem__0934_/Y VGND net365 net459 sg13g2_o21ai_1
XFILLER_7_573 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0865_ VGND VPWR net370 u_ppwm_u_mem__0722_/Y hold159/A u_ppwm_u_mem__0864_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0796_ hold87/A hold115/A net413 u_ppwm_u_mem__0796_/X VPWR VGND sg13g2_mux2_1
XFILLER_39_912 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__125_ net441 VGND VPWR net205 hold7/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__765_ VGND VPWR u_ppwm_u_ex__762_/Y u_ppwm_u_ex__763_/Y u_ppwm_u_ex__822_/D
+ u_ppwm_u_ex__764_/Y sg13g2_a21oi_1
XFILLER_39_989 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__056_ VPWR u_ppwm_u_global_counter__056_/Y net577 VGND sg13g2_inv_1
XFILLER_19_691 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__696_ u_ppwm_u_ex__696_/A u_ppwm_u_ex__696_/B u_ppwm_u_ex__696_/C u_ppwm_u_ex__696_/D
+ u_ppwm_u_ex__696_/Y VPWR VGND sg13g2_nor4_1
XFILLER_22_845 VPWR VGND sg13g2_decap_8
XFILLER_0_215 VPWR VGND sg13g2_decap_8
XFILLER_17_606 VPWR VGND sg13g2_decap_8
XFILLER_45_948 VPWR VGND sg13g2_decap_8
XFILLER_16_127 VPWR VGND sg13g2_fill_2
XFILLER_13_812 VPWR VGND sg13g2_decap_8
XFILLER_40_653 VPWR VGND sg13g2_decap_8
XFILLER_12_322 VPWR VGND sg13g2_decap_4
XFILLER_13_889 VPWR VGND sg13g2_decap_8
XFILLER_4_510 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0650_ VPWR u_ppwm_u_mem__0650_/Y net524 VGND sg13g2_inv_1
XFILLER_4_587 VPWR VGND sg13g2_decap_8
XFILLER_0_771 VPWR VGND sg13g2_decap_8
XFILLER_48_753 VPWR VGND sg13g2_decap_8
XFILLER_47_230 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1202_ net104 VGND VPWR net474 hold98/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_274 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1133_ net95 VGND VPWR net255 hold227/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_414 VPWR VGND sg13g2_decap_8
XFILLER_36_937 VPWR VGND sg13g2_decap_8
XFILLER_44_970 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__550_ hold71/A hold306/A u_ppwm_u_ex__550_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_23_609 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_9 VPWR VGND uio_oe[6] sg13g2_tielo
Xu_ppwm_u_mem__1064_ net429 VPWR u_ppwm_u_mem__1064_/Y VGND net339 net471 sg13g2_o21ai_1
XFILLER_16_672 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__481_ net443 VPWR u_ppwm_u_ex__482_/B VGND net631 net402 sg13g2_o21ai_1
XFILLER_31_620 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_697 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__236__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_8_882 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0917_ VGND VPWR net358 u_ppwm_u_mem__0696_/Y u_ppwm_u_mem__1135_/D
+ u_ppwm_u_mem__0916_/Y sg13g2_a21oi_1
Xhold326 hold326/A VPWR VGND net669 sg13g2_dlygate4sd3_1
Xhold315 hold315/A VPWR VGND net658 sg13g2_dlygate4sd3_1
Xhold304 hold304/A VPWR VGND net647 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0848_ hold13/A hold146/A net410 u_ppwm_u_mem__0848_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0779_ hold81/A hold195/A net411 u_ppwm_u_mem__0780_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_ex__817_ net37 VGND VPWR net635 hold298/A clknet_5_18__leaf_clk sg13g2_dfrbpq_2
XFILLER_39_786 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__108_ net438 VGND VPWR net252 hold54/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_26_38 VPWR VGND sg13g2_fill_1
XFILLER_27_959 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__748_ VGND VPWR u_ppwm_u_ex__748_/X u_ppwm_u_ex__748_/B u_ppwm_u_ex__748_/A
+ sg13g2_or2_1
Xu_ppwm_u_ex__679_ net318 VPWR u_ppwm_u_ex__698_/A VGND net391 net392 sg13g2_o21ai_1
XFILLER_35_981 VPWR VGND sg13g2_decap_8
XFILLER_22_642 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_1_568 VPWR VGND sg13g2_decap_8
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_18_926 VPWR VGND sg13g2_decap_8
XFILLER_45_745 VPWR VGND sg13g2_decap_8
XFILLER_33_918 VPWR VGND sg13g2_decap_8
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_34_1006 VPWR VGND sg13g2_decap_8
XFILLER_13_686 VPWR VGND sg13g2_decap_8
XFILLER_9_668 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0702_ VPWR u_ppwm_u_mem__0702_/Y net505 VGND sg13g2_inv_1
XFILLER_5_885 VPWR VGND sg13g2_decap_8
XFILLER_4_384 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0633_ VPWR u_ppwm_u_mem__0633_/Y net498 VGND sg13g2_inv_1
XFILLER_48_550 VPWR VGND sg13g2_decap_8
XFILLER_36_734 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__602_ u_ppwm_u_ex__605_/A hold185/A net382 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1116_ net129 VGND VPWR u_ppwm_u_mem__1116_/D hold44/A clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__533_ u_ppwm_u_ex__532_/Y VPWR u_ppwm_u_ex__534_/C VGND u_ppwm_u_ex__418_/Y
+ net393 sg13g2_o21ai_1
XFILLER_17_970 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1047_ VGND VPWR net354 u_ppwm_u_mem__0631_/Y u_ppwm_u_mem__1200_/D
+ u_ppwm_u_mem__1046_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__464_ u_ppwm_u_ex__463_/Y VPWR u_ppwm_u_ex__464_/Y VGND net407 net415
+ sg13g2_o21ai_1
XFILLER_32_962 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
Xhold101 hold101/A VPWR VGND net298 sg13g2_dlygate4sd3_1
Xhold112 hold112/A VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold134 hold134/A VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold123 hold123/A VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold145 hold145/A VPWR VGND net488 sg13g2_dlygate4sd3_1
Xhold167 hold167/A VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold156 hold156/A VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold178 hold178/A VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold189 hold189/A VPWR VGND net532 sg13g2_dlygate4sd3_1
XFILLER_39_583 VPWR VGND sg13g2_decap_8
XFILLER_15_907 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_42_748 VPWR VGND sg13g2_decap_8
XFILLER_23_973 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__804__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_2_800 VPWR VGND sg13g2_decap_8
XFILLER_2_877 VPWR VGND sg13g2_decap_8
XFILLER_1_365 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_40_1010 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__226__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_18_723 VPWR VGND sg13g2_decap_8
XFILLER_45_542 VPWR VGND sg13g2_decap_8
XFILLER_33_715 VPWR VGND sg13g2_decap_8
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_13_483 VPWR VGND sg13g2_decap_8
XFILLER_9_465 VPWR VGND sg13g2_decap_8
XFILLER_5_682 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0616_ VPWR u_ppwm_u_mem__0616_/Y net592 VGND sg13g2_inv_1
XFILLER_4_96 VPWR VGND sg13g2_decap_4
Xheichips25_ppwm_19 VPWR VGND uo_out[1] sg13g2_tielo
XFILLER_36_531 VPWR VGND sg13g2_decap_8
XFILLER_24_748 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__516_ VGND VPWR u_ppwm_u_ex__511_/B u_ppwm_u_ex__515_/D u_ppwm_u_ex__517_/C
+ u_ppwm_u_ex__509_/Y sg13g2_a21oi_1
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__447_ VGND VPWR u_ppwm_u_ex__620_/B u_ppwm/instr\[1\] u_ppwm/instr\[0\]
+ sg13g2_or2_1
XFILLER_20_965 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout422 net437 net422 VPWR VGND sg13g2_buf_8
Xfanout400 fanout401/A net400 VPWR VGND sg13g2_buf_8
Xfanout411 net414 net411 VPWR VGND sg13g2_buf_8
Xfanout444 net445 net444 VPWR VGND sg13g2_buf_8
Xfanout433 net436 net433 VPWR VGND sg13g2_buf_8
XFILLER_47_829 VPWR VGND sg13g2_decap_8
XFILLER_19_509 VPWR VGND sg13g2_decap_8
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_15_704 VPWR VGND sg13g2_decap_8
XFILLER_42_545 VPWR VGND sg13g2_decap_8
XFILLER_11_932 VPWR VGND sg13g2_decap_8
XFILLER_23_770 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__140_ net337 hold268/A hold192/A hold287/A u_ppwm_u_pwm__142_/C VPWR
+ VGND sg13g2_nor4_1
XFILLER_7_958 VPWR VGND sg13g2_decap_8
XFILLER_6_468 VPWR VGND sg13g2_decap_8
XFILLER_2_674 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_1_184 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_18_520 VPWR VGND sg13g2_decap_8
XFILLER_46_840 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_18_597 VPWR VGND sg13g2_decap_8
XFILLER_33_589 VPWR VGND sg13g2_decap_8
XFILLER_9_240 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1199__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_29_829 VPWR VGND sg13g2_decap_8
XFILLER_37_862 VPWR VGND sg13g2_decap_8
XFILLER_24_545 VPWR VGND sg13g2_decap_8
Xclkload4 clknet_5_12__leaf_clk clkload4/X VPWR VGND sg13g2_buf_1
XFILLER_20_762 VPWR VGND sg13g2_decap_8
XFILLER_47_626 VPWR VGND sg13g2_decap_8
XFILLER_28_851 VPWR VGND sg13g2_decap_8
XFILLER_43_810 VPWR VGND sg13g2_decap_8
XFILLER_15_501 VPWR VGND sg13g2_decap_8
XFILLER_27_361 VPWR VGND sg13g2_decap_4
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0950_ net449 VPWR u_ppwm_u_mem__0950_/Y VGND net374 net297 sg13g2_o21ai_1
XFILLER_30_559 VPWR VGND sg13g2_decap_8
XFILLER_6_210 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0881_ VGND VPWR net370 u_ppwm_u_mem__0714_/Y hold122/A u_ppwm_u_mem__0880_/Y
+ sg13g2_a21oi_1
XFILLER_7_755 VPWR VGND sg13g2_decap_8
XFILLER_3_950 VPWR VGND sg13g2_decap_8
XFILLER_2_471 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__072_ u_ppwm_u_global_counter__073_/B net587 hold245/A VPWR
+ VGND sg13g2_nor2_1
XFILLER_1_42 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__781_ u_ppwm_u_ex__781_/B u_ppwm_u_ex__781_/C fanout316/A u_ppwm_u_ex__781_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_38_648 VPWR VGND sg13g2_decap_8
XFILLER_18_361 VPWR VGND sg13g2_decap_4
XFILLER_19_873 VPWR VGND sg13g2_decap_8
XFILLER_34_810 VPWR VGND sg13g2_decap_8
XFILLER_34_887 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1203__96 VPWR VGND net96 sg13g2_tiehi
Xhold27 hold27/A VPWR VGND net224 sg13g2_dlygate4sd3_1
XFILLER_29_49 VPWR VGND sg13g2_fill_1
Xhold16 hold16/A VPWR VGND net213 sg13g2_dlygate4sd3_1
Xhold38 hold38/A VPWR VGND net235 sg13g2_dlygate4sd3_1
XFILLER_29_626 VPWR VGND sg13g2_decap_8
Xhold49 hold49/A VPWR VGND net246 sg13g2_dlygate4sd3_1
XFILLER_45_48 VPWR VGND sg13g2_fill_1
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_40_835 VPWR VGND sg13g2_decap_8
XFILLER_12_537 VPWR VGND sg13g2_decap_8
XFILLER_25_898 VPWR VGND sg13g2_decap_8
XFILLER_4_769 VPWR VGND sg13g2_decap_8
XFILLER_0_953 VPWR VGND sg13g2_decap_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
XFILLER_47_423 VPWR VGND sg13g2_decap_8
XFILLER_47_412 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1080_ net426 VPWR u_ppwm_u_mem__1080_/Y VGND net345 hold178/A sg13g2_o21ai_1
XFILLER_16_854 VPWR VGND sg13g2_decap_8
XFILLER_31_802 VPWR VGND sg13g2_decap_8
XFILLER_43_684 VPWR VGND sg13g2_decap_8
XFILLER_30_312 VPWR VGND sg13g2_fill_2
XFILLER_31_879 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0933_ VGND VPWR net365 u_ppwm_u_mem__0688_/Y hold117/A u_ppwm_u_mem__0932_/Y
+ sg13g2_a21oi_1
XFILLER_7_552 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0864_ net450 VPWR u_ppwm_u_mem__0864_/Y VGND net370 hold242/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0795_ u_ppwm_u_mem__0795_/Y net404 u_ppwm_u_mem__0795_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_44_1019 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__124_ net440 VGND VPWR net565 hold221/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_968 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__055_ VPWR u_ppwm_u_global_counter__055_/Y net615 VGND sg13g2_inv_1
Xu_ppwm_u_ex__764_ net441 VPWR u_ppwm_u_ex__764_/Y VGND net381 net307 sg13g2_o21ai_1
XFILLER_26_629 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_19_670 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__695_ VGND VPWR u_ppwm_u_ex__692_/Y u_ppwm_u_ex__693_/Y hold331/A u_ppwm_u_ex__694_/Y
+ sg13g2_a21oi_1
XFILLER_22_824 VPWR VGND sg13g2_decap_8
XFILLER_34_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1188__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_45_927 VPWR VGND sg13g2_decap_8
XFILLER_44_459 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_fill_2
XFILLER_25_695 VPWR VGND sg13g2_decap_8
XFILLER_40_632 VPWR VGND sg13g2_decap_8
XFILLER_13_868 VPWR VGND sg13g2_decap_8
XFILLER_4_566 VPWR VGND sg13g2_decap_8
XFILLER_0_750 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1195__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_48_732 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1201_ net112 VGND VPWR net296 hold115/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_916 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1132_ net97 VGND VPWR net571 hold102/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_990 VPWR VGND sg13g2_decap_8
XFILLER_35_437 VPWR VGND sg13g2_fill_2
XFILLER_46_91 VPWR VGND sg13g2_fill_1
XFILLER_16_651 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1063_ VGND VPWR net343 u_ppwm_u_mem__0623_/Y hold129/A u_ppwm_u_mem__1062_/Y
+ sg13g2_a21oi_1
XFILLER_35_459 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__480_ u_ppwm_u_ex__482_/A u_ppwm_u_ex__485_/B u_ppwm_u_ex__479_/Y u_ppwm_u_ex__474_/Y
+ u_ppwm_u_ex__472_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_43_481 VPWR VGND sg13g2_decap_8
XFILLER_15_183 VPWR VGND sg13g2_fill_1
XFILLER_31_676 VPWR VGND sg13g2_decap_8
XFILLER_8_861 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0916_ net446 VPWR u_ppwm_u_mem__0916_/Y VGND net358 net235 sg13g2_o21ai_1
Xhold316 hold316/A VPWR VGND net659 sg13g2_dlygate4sd3_1
Xhold305 hold305/A VPWR VGND net648 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0847_ VGND VPWR net335 u_ppwm_u_mem__0846_/X u_ppwm_u_mem__0847_/Y
+ net403 sg13g2_a21oi_1
Xhold327 hold327/A VPWR VGND net670 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0778_ VGND VPWR net334 u_ppwm_u_mem__0777_/X u_ppwm_u_mem__0778_/Y
+ net333 sg13g2_a21oi_1
XFILLER_30_0 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__816_ net41 VGND VPWR net652 hold308/A clknet_5_6__leaf_clk sg13g2_dfrbpq_2
XFILLER_39_765 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__107_ net438 VGND VPWR net656 hold311/A clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_27_938 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__747_ VGND VPWR u_ppwm_u_ex__744_/Y u_ppwm_u_ex__745_/Y hold316/A u_ppwm_u_ex__746_/Y
+ sg13g2_a21oi_1
XFILLER_35_960 VPWR VGND sg13g2_decap_8
XFILLER_41_429 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__678_ u_ppwm_u_ex__696_/C net389 net318 VPWR VGND sg13g2_xnor2_1
XFILLER_22_621 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_22_698 VPWR VGND sg13g2_decap_8
XFILLER_1_547 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1155__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_18_905 VPWR VGND sg13g2_decap_8
XFILLER_29_231 VPWR VGND sg13g2_fill_2
XFILLER_29_253 VPWR VGND sg13g2_fill_1
XFILLER_45_724 VPWR VGND sg13g2_decap_8
XFILLER_44_212 VPWR VGND sg13g2_decap_4
XFILLER_44_256 VPWR VGND sg13g2_fill_2
XFILLER_17_459 VPWR VGND sg13g2_decap_8
XFILLER_26_993 VPWR VGND sg13g2_decap_8
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_25_492 VPWR VGND sg13g2_decap_8
XFILLER_13_665 VPWR VGND sg13g2_decap_8
XFILLER_9_647 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0701_ VPWR u_ppwm_u_mem__0701_/Y net475 VGND sg13g2_inv_1
XFILLER_5_864 VPWR VGND sg13g2_decap_8
XFILLER_4_363 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0632_ VPWR u_ppwm_u_mem__0632_/Y net274 VGND sg13g2_inv_1
XFILLER_36_713 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__601_ u_ppwm_u_ex__604_/A net381 hold243/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1115_ net131 VGND VPWR net242 hold217/A clknet_5_29__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__532_ u_ppwm_u_ex__532_/Y net381 net391 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1046_ net435 VPWR u_ppwm_u_mem__1046_/Y VGND net353 net274 sg13g2_o21ai_1
Xu_ppwm_u_ex__463_ u_ppwm_u_ex__463_/Y net377 u_ppwm_u_ex__474_/B VPWR VGND sg13g2_nand2_1
XFILLER_32_941 VPWR VGND sg13g2_decap_8
Xhold113 hold113/A VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold124 hold124/A VPWR VGND net467 sg13g2_dlygate4sd3_1
Xhold135 hold135/A VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold102 hold102/A VPWR VGND net299 sg13g2_dlygate4sd3_1
Xhold146 hold146/A VPWR VGND net489 sg13g2_dlygate4sd3_1
Xhold157 hold157/A VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold168 hold168/A VPWR VGND net511 sg13g2_dlygate4sd3_1
Xhold179 hold179/A VPWR VGND net522 sg13g2_dlygate4sd3_1
XFILLER_37_16 VPWR VGND sg13g2_decap_4
XFILLER_39_562 VPWR VGND sg13g2_decap_8
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_26_245 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1181__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_42_727 VPWR VGND sg13g2_decap_8
XFILLER_14_429 VPWR VGND sg13g2_decap_8
XFILLER_41_237 VPWR VGND sg13g2_fill_1
XFILLER_23_952 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_22_495 VPWR VGND sg13g2_decap_8
XFILLER_2_856 VPWR VGND sg13g2_decap_8
XFILLER_1_344 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_18_702 VPWR VGND sg13g2_decap_8
XFILLER_45_521 VPWR VGND sg13g2_decap_8
XFILLER_18_779 VPWR VGND sg13g2_decap_8
XFILLER_45_598 VPWR VGND sg13g2_decap_8
XFILLER_26_790 VPWR VGND sg13g2_decap_8
XFILLER_9_444 VPWR VGND sg13g2_decap_8
XFILLER_13_462 VPWR VGND sg13g2_decap_8
XFILLER_14_996 VPWR VGND sg13g2_decap_8
XFILLER_5_661 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0615_ VPWR u_ppwm_u_mem__0615_/Y net521 VGND sg13g2_inv_1
XFILLER_49_882 VPWR VGND sg13g2_decap_8
XFILLER_24_727 VPWR VGND sg13g2_decap_8
XFILLER_36_587 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__515_ u_ppwm_u_ex__515_/A u_ppwm_u_ex__515_/B u_ppwm_u_ex__515_/C u_ppwm_u_ex__515_/D
+ u_ppwm_u_ex__515_/Y VPWR VGND sg13g2_nor4_1
Xu_ppwm_u_mem__1029_ VGND VPWR net347 u_ppwm_u_mem__0640_/Y hold143/A u_ppwm_u_mem__1028_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__446_ u_ppwm_u_ex__448_/C u_ppwm_u_ex__517_/B net324 VPWR VGND sg13g2_nand2b_1
XFILLER_20_944 VPWR VGND sg13g2_decap_8
Xfanout423 net437 net423 VPWR VGND sg13g2_buf_8
Xfanout401 fanout401/A net401 VPWR VGND sg13g2_buf_1
Xfanout412 net413 net412 VPWR VGND sg13g2_buf_8
Xfanout445 net446 net445 VPWR VGND sg13g2_buf_8
Xfanout434 net435 net434 VPWR VGND sg13g2_buf_8
XFILLER_47_808 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1113__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_42_524 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_11_911 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_7_937 VPWR VGND sg13g2_decap_8
XFILLER_11_988 VPWR VGND sg13g2_decap_8
XFILLER_6_447 VPWR VGND sg13g2_decap_8
XFILLER_2_653 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_fill_2
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_18_576 VPWR VGND sg13g2_decap_8
XFILLER_33_568 VPWR VGND sg13g2_decap_8
XFILLER_14_793 VPWR VGND sg13g2_decap_8
XFILLER_13_281 VPWR VGND sg13g2_decap_8
XFILLER_9_285 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__199_ VPWR VGND u_ppwm_u_pwm__128_/Y u_ppwm_u_pwm__197_/Y hold21/A u_ppwm_u_pwm__127_/Y
+ u_ppwm_u_pwm__199_/Y hold219/A sg13g2_a221oi_1
XFILLER_29_808 VPWR VGND sg13g2_decap_8
XFILLER_37_841 VPWR VGND sg13g2_decap_8
XFILLER_24_524 VPWR VGND sg13g2_decap_8
XFILLER_12_719 VPWR VGND sg13g2_decap_8
XFILLER_20_741 VPWR VGND sg13g2_decap_8
Xclkload5 clknet_5_14__leaf_clk clkload5/X VPWR VGND sg13g2_buf_1
Xu_ppwm_u_ex__429_ VPWR u_ppwm_u_ex__429_/Y net336 VGND sg13g2_inv_1
XFILLER_30_1021 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1206__72 VPWR VGND net72 sg13g2_tiehi
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_439 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_8_1022 VPWR VGND sg13g2_decap_8
XFILLER_47_605 VPWR VGND sg13g2_decap_8
XFILLER_28_830 VPWR VGND sg13g2_decap_8
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_42_365 VPWR VGND sg13g2_decap_4
XFILLER_30_538 VPWR VGND sg13g2_decap_8
XFILLER_7_734 VPWR VGND sg13g2_decap_8
XFILLER_11_785 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0880_ net447 VPWR u_ppwm_u_mem__0880_/Y VGND net371 hold180/A sg13g2_o21ai_1
XFILLER_2_450 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_38_627 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__071_ VGND VPWR net528 u_ppwm_u_global_counter__068_/B hold244/A
+ net586 sg13g2_a21oi_1
XFILLER_19_852 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__780_ u_ppwm_u_ex__779_/B u_ppwm_u_ex__779_/A u_ppwm_u_ex__785_/D u_ppwm_u_ex__781_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_37_148 VPWR VGND sg13g2_fill_2
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_18_395 VPWR VGND sg13g2_fill_1
XFILLER_33_310 VPWR VGND sg13g2_fill_1
XFILLER_33_332 VPWR VGND sg13g2_decap_8
XFILLER_34_866 VPWR VGND sg13g2_decap_8
XFILLER_33_365 VPWR VGND sg13g2_fill_2
XFILLER_14_590 VPWR VGND sg13g2_decap_8
XFILLER_21_549 VPWR VGND sg13g2_decap_8
XFILLER_20_19 VPWR VGND sg13g2_decap_4
Xhold17 hold17/A VPWR VGND net214 sg13g2_dlygate4sd3_1
Xhold28 hold28/A VPWR VGND net225 sg13g2_dlygate4sd3_1
XFILLER_29_605 VPWR VGND sg13g2_decap_8
Xhold39 hold39/A VPWR VGND net236 sg13g2_dlygate4sd3_1
XFILLER_25_800 VPWR VGND sg13g2_decap_8
XFILLER_24_343 VPWR VGND sg13g2_fill_2
XFILLER_25_877 VPWR VGND sg13g2_decap_8
XFILLER_40_814 VPWR VGND sg13g2_decap_8
XFILLER_12_516 VPWR VGND sg13g2_decap_8
XFILLER_4_748 VPWR VGND sg13g2_decap_8
XFILLER_0_932 VPWR VGND sg13g2_decap_8
XFILLER_48_914 VPWR VGND sg13g2_decap_8
XFILLER_47_479 VPWR VGND sg13g2_decap_8
XFILLER_16_833 VPWR VGND sg13g2_decap_8
XFILLER_43_663 VPWR VGND sg13g2_decap_8
XFILLER_37_1016 VPWR VGND sg13g2_decap_8
XFILLER_15_387 VPWR VGND sg13g2_fill_2
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
XFILLER_31_858 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1165__150 VPWR VGND net150 sg13g2_tiehi
Xu_ppwm_u_mem__0932_ net445 VPWR u_ppwm_u_mem__0932_/Y VGND net365 hold151/A sg13g2_o21ai_1
XFILLER_7_531 VPWR VGND sg13g2_decap_8
XFILLER_11_582 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0863_ VGND VPWR net361 u_ppwm_u_mem__0723_/Y u_ppwm_u_mem__1108_/D
+ u_ppwm_u_mem__0862_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0794_ hold236/A hold215/A net410 u_ppwm_u_mem__0795_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_global_counter__123_ net440 VGND VPWR u_ppwm_u_global_counter__123_/D hold271/A
+ clknet_5_20__leaf_clk sg13g2_dfrbpq_2
XFILLER_39_947 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__054_ VPWR u_ppwm_u_global_counter__054_/Y net609 VGND sg13g2_inv_1
Xu_ppwm_u_ex__763_ VPWR VGND net636 u_ppwm_u_ex__714_/Y fanout312/A net380 u_ppwm_u_ex__763_/Y
+ net314 sg13g2_a221oi_1
XFILLER_26_608 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__694_ net426 VPWR u_ppwm_u_ex__694_/Y VGND net387 net310 sg13g2_o21ai_1
XFILLER_22_803 VPWR VGND sg13g2_decap_8
XFILLER_33_140 VPWR VGND sg13g2_fill_2
XFILLER_34_663 VPWR VGND sg13g2_decap_8
XFILLER_21_313 VPWR VGND sg13g2_decap_4
XFILLER_1_729 VPWR VGND sg13g2_decap_8
XFILLER_29_402 VPWR VGND sg13g2_fill_1
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
XFILLER_45_906 VPWR VGND sg13g2_decap_8
XFILLER_38_991 VPWR VGND sg13g2_decap_8
XFILLER_40_611 VPWR VGND sg13g2_decap_8
XFILLER_25_674 VPWR VGND sg13g2_decap_8
XFILLER_13_847 VPWR VGND sg13g2_decap_8
XFILLER_40_688 VPWR VGND sg13g2_decap_8
XFILLER_8_317 VPWR VGND sg13g2_fill_1
XFILLER_9_829 VPWR VGND sg13g2_decap_8
XFILLER_21_51 VPWR VGND sg13g2_fill_1
XFILLER_4_545 VPWR VGND sg13g2_decap_8
XFILLER_21_84 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_fill_1
XFILLER_48_711 VPWR VGND sg13g2_decap_8
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1200_ net120 VGND VPWR u_ppwm_u_mem__1200_/D hold77/A clknet_5_24__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_48_788 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1131_ net99 VGND VPWR net300 hold132/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_298 VPWR VGND sg13g2_fill_2
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_16_630 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1062_ net429 VPWR u_ppwm_u_mem__1062_/Y VGND net342 hold236/A sg13g2_o21ai_1
XFILLER_31_655 VPWR VGND sg13g2_decap_8
XFILLER_8_840 VPWR VGND sg13g2_decap_8
XFILLER_12_880 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0915_ VGND VPWR net358 u_ppwm_u_mem__0697_/Y hold39/A u_ppwm_u_mem__0914_/Y
+ sg13g2_a21oi_1
Xhold317 hold317/A VPWR VGND net660 sg13g2_dlygate4sd3_1
Xhold306 hold306/A VPWR VGND net649 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0846_ hold274/A hold277/A net411 u_ppwm_u_mem__0846_/X VPWR VGND sg13g2_mux2_1
Xhold328 hold328/A VPWR VGND net671 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0777_ hold34/A hold77/A net413 u_ppwm_u_mem__0777_/X VPWR VGND sg13g2_mux2_1
XFILLER_39_744 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__106_ net438 VGND VPWR net269 hold71/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__815_ net45 VGND VPWR u_ppwm_u_ex__815_/D hold333/A clknet_5_7__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_42_909 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__746_ net441 VPWR u_ppwm_u_ex__746_/Y VGND net383 net307 sg13g2_o21ai_1
Xu_ppwm_u_ex__677_ u_ppwm_u_ex__690_/A net389 net318 VPWR VGND sg13g2_nand2_1
XFILLER_22_600 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__816__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_22_677 VPWR VGND sg13g2_decap_8
XFILLER_1_526 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_210 VPWR VGND sg13g2_decap_8
XFILLER_45_703 VPWR VGND sg13g2_decap_8
XFILLER_17_438 VPWR VGND sg13g2_decap_8
XFILLER_26_972 VPWR VGND sg13g2_decap_8
XFILLER_41_920 VPWR VGND sg13g2_decap_8
XFILLER_13_644 VPWR VGND sg13g2_decap_8
XFILLER_25_471 VPWR VGND sg13g2_decap_8
XFILLER_9_626 VPWR VGND sg13g2_decap_8
XFILLER_12_143 VPWR VGND sg13g2_fill_2
XFILLER_41_997 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1123__115 VPWR VGND net115 sg13g2_tiehi
Xu_ppwm_u_mem__0700_ VPWR u_ppwm_u_mem__0700_/Y net299 VGND sg13g2_inv_1
XFILLER_5_843 VPWR VGND sg13g2_decap_8
XFILLER_4_342 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0631_ VPWR u_ppwm_u_mem__0631_/Y net458 VGND sg13g2_inv_1
XFILLER_48_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__600_ VPWR VGND u_ppwm_u_ex__420_/Y u_ppwm_u_ex__599_/Y hold54/A u_ppwm_u_ex__419_/Y
+ u_ppwm_u_ex__600_/Y hold203/A sg13g2_a221oi_1
XFILLER_24_909 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1114_ net133 VGND VPWR net561 hold138/A clknet_5_23__leaf_clk sg13g2_dfrbpq_2
XFILLER_36_769 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__531_ u_ppwm_u_ex__530_/Y VPWR u_ppwm_u_ex__534_/B VGND net381 u_ppwm_u_ex__583_/A
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__1045_ VGND VPWR net353 u_ppwm_u_mem__0632_/Y hold78/A u_ppwm_u_mem__1044_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__462_ u_ppwm_u_ex__474_/B u_ppwm_u_ex__472_/B u_ppwm_u_ex__488_/B VPWR
+ VGND sg13g2_nand2_1
XFILLER_32_920 VPWR VGND sg13g2_decap_8
XFILLER_32_997 VPWR VGND sg13g2_decap_8
Xhold114 hold114/A VPWR VGND net457 sg13g2_dlygate4sd3_1
Xhold125 hold125/A VPWR VGND net468 sg13g2_dlygate4sd3_1
Xhold103 hold103/A VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold147 hold147/A VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold136 hold136/A VPWR VGND net479 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0829_ net404 VPWR u_ppwm_u_mem__0829_/Y VGND hold191/A net412 sg13g2_o21ai_1
Xhold158 hold158/A VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold169 hold169/A VPWR VGND net512 sg13g2_dlygate4sd3_1
XFILLER_39_541 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_42_706 VPWR VGND sg13g2_decap_8
XFILLER_14_408 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__729_ net442 VPWR u_ppwm_u_ex__729_/Y VGND net634 net307 sg13g2_o21ai_1
XFILLER_23_931 VPWR VGND sg13g2_decap_8
XFILLER_22_474 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_6_629 VPWR VGND sg13g2_decap_8
XFILLER_2_835 VPWR VGND sg13g2_decap_8
XFILLER_1_323 VPWR VGND sg13g2_decap_8
XFILLER_45_500 VPWR VGND sg13g2_decap_8
XFILLER_18_758 VPWR VGND sg13g2_decap_8
XFILLER_45_577 VPWR VGND sg13g2_decap_8
XFILLER_17_257 VPWR VGND sg13g2_fill_1
XFILLER_17_268 VPWR VGND sg13g2_decap_4
XFILLER_13_441 VPWR VGND sg13g2_decap_8
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_41_794 VPWR VGND sg13g2_decap_8
XFILLER_9_423 VPWR VGND sg13g2_decap_8
XFILLER_40_260 VPWR VGND sg13g2_fill_2
XFILLER_5_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0614_ VPWR u_ppwm_u_mem__0730_/A net1 VGND sg13g2_inv_1
XFILLER_1_890 VPWR VGND sg13g2_decap_8
XFILLER_49_861 VPWR VGND sg13g2_decap_8
XFILLER_48_382 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__240__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_24_706 VPWR VGND sg13g2_decap_8
XFILLER_36_566 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__514_ net379 hold221/A u_ppwm_u_ex__515_/D VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_mem__1028_ net429 VPWR u_ppwm_u_mem__1028_/Y VGND net347 hold231/A sg13g2_o21ai_1
Xu_ppwm_u_ex__445_ net325 net327 u_ppwm_u_ex__517_/B VPWR VGND sg13g2_nor2b_1
XFILLER_20_923 VPWR VGND sg13g2_decap_8
XFILLER_32_794 VPWR VGND sg13g2_decap_8
XFILLER_31_293 VPWR VGND sg13g2_decap_4
XFILLER_9_990 VPWR VGND sg13g2_decap_8
Xfanout402 net638 net402 VPWR VGND sg13g2_buf_8
Xfanout413 net414 net413 VPWR VGND sg13g2_buf_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
Xfanout424 net427 net424 VPWR VGND sg13g2_buf_8
XFILLER_24_1007 VPWR VGND sg13g2_decap_8
Xfanout446 net452 net446 VPWR VGND sg13g2_buf_8
Xfanout435 net436 net435 VPWR VGND sg13g2_buf_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1146__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_42_503 VPWR VGND sg13g2_decap_8
XFILLER_15_739 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_7_916 VPWR VGND sg13g2_decap_8
XFILLER_11_967 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_6_426 VPWR VGND sg13g2_decap_8
XFILLER_13_96 VPWR VGND sg13g2_fill_2
XFILLER_2_632 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1200__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_38_809 VPWR VGND sg13g2_decap_8
XFILLER_49_168 VPWR VGND sg13g2_decap_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_18_555 VPWR VGND sg13g2_decap_8
XFILLER_33_547 VPWR VGND sg13g2_decap_8
XFILLER_13_260 VPWR VGND sg13g2_fill_1
XFILLER_14_772 VPWR VGND sg13g2_decap_8
XFILLER_41_591 VPWR VGND sg13g2_decap_8
XFILLER_9_264 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_pwm__198_ VGND VPWR u_ppwm_u_pwm__194_/Y u_ppwm_u_pwm__196_/Y u_ppwm_u_pwm__198_/Y
+ u_ppwm_u_pwm__197_/Y sg13g2_a21oi_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_6_993 VPWR VGND sg13g2_decap_8
XFILLER_37_820 VPWR VGND sg13g2_decap_8
XFILLER_24_503 VPWR VGND sg13g2_decap_8
XFILLER_36_385 VPWR VGND sg13g2_decap_4
XFILLER_37_897 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__428_ VPWR u_ppwm_u_ex__637_/B net325 VGND sg13g2_inv_1
XFILLER_20_720 VPWR VGND sg13g2_decap_8
XFILLER_32_591 VPWR VGND sg13g2_decap_8
Xclkload6 clknet_5_21__leaf_clk clkload6/X VPWR VGND sg13g2_buf_1
XFILLER_30_1000 VPWR VGND sg13g2_decap_8
XFILLER_20_797 VPWR VGND sg13g2_decap_8
XFILLER_3_418 VPWR VGND sg13g2_decap_8
XFILLER_8_1001 VPWR VGND sg13g2_decap_8
XFILLER_19_308 VPWR VGND sg13g2_fill_2
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_43_845 VPWR VGND sg13g2_decap_8
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_42_344 VPWR VGND sg13g2_fill_1
XFILLER_30_517 VPWR VGND sg13g2_decap_8
XFILLER_7_713 VPWR VGND sg13g2_decap_8
XFILLER_11_764 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_4
XFILLER_6_245 VPWR VGND sg13g2_fill_1
XFILLER_3_985 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_4
XFILLER_38_606 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__070_ u_ppwm_u_global_counter__070_/A u_ppwm_u_global_counter__085_/A
+ u_ppwm_u_global_counter__073_/B VPWR VGND sg13g2_nor2_1
XFILLER_19_831 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_decap_8
XFILLER_34_845 VPWR VGND sg13g2_decap_8
XFILLER_21_528 VPWR VGND sg13g2_decap_8
XFILLER_33_388 VPWR VGND sg13g2_decap_8
XFILLER_33_399 VPWR VGND sg13g2_fill_2
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_790 VPWR VGND sg13g2_decap_8
Xhold18 hold18/A VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold29 hold29/A VPWR VGND net226 sg13g2_dlygate4sd3_1
Xu_ppwm_u_pwm__246__184 VPWR VGND net184 sg13g2_tiehi
Xu_ppwm_u_mem__1214__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_45_39 VPWR VGND sg13g2_fill_1
XFILLER_37_694 VPWR VGND sg13g2_decap_8
XFILLER_25_856 VPWR VGND sg13g2_decap_8
XFILLER_36_193 VPWR VGND sg13g2_fill_1
XFILLER_20_594 VPWR VGND sg13g2_decap_8
XFILLER_4_727 VPWR VGND sg13g2_decap_8
XFILLER_0_911 VPWR VGND sg13g2_decap_8
XFILLER_0_988 VPWR VGND sg13g2_decap_8
XFILLER_47_458 VPWR VGND sg13g2_decap_8
XFILLER_15_311 VPWR VGND sg13g2_decap_8
XFILLER_16_812 VPWR VGND sg13g2_decap_8
XFILLER_28_683 VPWR VGND sg13g2_decap_8
XFILLER_43_642 VPWR VGND sg13g2_decap_8
XFILLER_16_889 VPWR VGND sg13g2_decap_8
XFILLER_31_837 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0931_ VGND VPWR net364 u_ppwm_u_mem__0689_/Y hold152/A u_ppwm_u_mem__0930_/Y
+ sg13g2_a21oi_1
XFILLER_7_510 VPWR VGND sg13g2_decap_8
XFILLER_11_561 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0862_ net451 VPWR u_ppwm_u_mem__0862_/Y VGND net361 net511 sg13g2_o21ai_1
XFILLER_7_587 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0793_ u_ppwm_u_mem__0792_/X u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0783_/Y
+ u_ppwm/instr\[2\] VPWR VGND sg13g2_a21o_2
XFILLER_3_782 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_39_926 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__122_ net440 VGND VPWR net199 hold1/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__053_ VPWR u_ppwm_u_global_counter__066_/A net546 VGND sg13g2_inv_1
Xu_ppwm_u_ex__762_ u_ppwm_u_ex__762_/B u_ppwm_u_ex__762_/C fanout316/A u_ppwm_u_ex__762_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_20_1021 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__693_ VPWR VGND net389 net309 net311 net386 u_ppwm_u_ex__693_/Y net313
+ sg13g2_a221oi_1
XFILLER_34_642 VPWR VGND sg13g2_decap_8
XFILLER_22_859 VPWR VGND sg13g2_decap_8
XFILLER_30_881 VPWR VGND sg13g2_decap_8
XFILLER_1_708 VPWR VGND sg13g2_decap_8
XFILLER_0_229 VPWR VGND sg13g2_decap_8
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_25_653 VPWR VGND sg13g2_decap_8
XFILLER_37_480 VPWR VGND sg13g2_fill_2
XFILLER_13_826 VPWR VGND sg13g2_decap_8
XFILLER_9_808 VPWR VGND sg13g2_decap_8
XFILLER_40_667 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_4
XFILLER_21_892 VPWR VGND sg13g2_decap_8
XFILLER_4_524 VPWR VGND sg13g2_decap_8
XFILLER_0_785 VPWR VGND sg13g2_decap_8
XFILLER_48_767 VPWR VGND sg13g2_decap_8
XFILLER_47_244 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1130_ net101 VGND VPWR net476 hold162/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1061_ VGND VPWR net340 u_ppwm_u_mem__0624_/Y u_ppwm_u_mem__1207_/D
+ u_ppwm_u_mem__1060_/Y sg13g2_a21oi_1
XFILLER_35_428 VPWR VGND sg13g2_decap_4
XFILLER_35_439 VPWR VGND sg13g2_fill_1
XFILLER_44_984 VPWR VGND sg13g2_decap_8
XFILLER_16_686 VPWR VGND sg13g2_decap_8
XFILLER_31_634 VPWR VGND sg13g2_decap_8
XFILLER_30_155 VPWR VGND sg13g2_fill_1
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_11_380 VPWR VGND sg13g2_fill_2
XFILLER_11_1009 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0914_ net446 VPWR u_ppwm_u_mem__0914_/Y VGND net358 hold57/A sg13g2_o21ai_1
XFILLER_8_896 VPWR VGND sg13g2_decap_8
Xhold307 hold307/A VPWR VGND net650 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0845_ u_ppwm_u_mem__0845_/Y net404 u_ppwm_u_mem__0845_/B VPWR VGND
+ sg13g2_nand2_1
Xhold318 hold318/A VPWR VGND net661 sg13g2_dlygate4sd3_1
Xhold329 hold329/A VPWR VGND net672 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0776_ u_ppwm_u_mem__0776_/Y net404 u_ppwm_u_mem__0776_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_39_723 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__105_ u_ppwm_u_global_counter__105_/B net204 hold8/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__814_ net47 VGND VPWR net674 hold330/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__745_ VPWR VGND net658 u_ppwm_u_ex__714_/Y net312 net382 u_ppwm_u_ex__745_/Y
+ net314 sg13g2_a221oi_1
Xu_ppwm_u_ex__676_ VGND VPWR u_ppwm_u_ex__673_/Y u_ppwm_u_ex__674_/Y u_ppwm_u_ex__812_/D
+ u_ppwm_u_ex__675_/Y sg13g2_a21oi_1
XFILLER_21_100 VPWR VGND sg13g2_fill_2
XFILLER_35_995 VPWR VGND sg13g2_decap_8
XFILLER_22_656 VPWR VGND sg13g2_decap_8
XFILLER_1_505 VPWR VGND sg13g2_decap_8
XFILLER_29_233 VPWR VGND sg13g2_fill_1
XFILLER_17_417 VPWR VGND sg13g2_decap_8
XFILLER_45_759 VPWR VGND sg13g2_decap_8
XFILLER_26_951 VPWR VGND sg13g2_decap_8
XFILLER_29_299 VPWR VGND sg13g2_fill_1
XFILLER_25_450 VPWR VGND sg13g2_decap_8
XFILLER_13_623 VPWR VGND sg13g2_decap_8
XFILLER_16_96 VPWR VGND sg13g2_fill_2
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_9_605 VPWR VGND sg13g2_decap_8
XFILLER_32_73 VPWR VGND sg13g2_fill_2
XFILLER_5_822 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0630_ VPWR u_ppwm_u_mem__0630_/Y net295 VGND sg13g2_inv_1
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_4_398 VPWR VGND sg13g2_decap_8
XFILLER_0_582 VPWR VGND sg13g2_decap_8
XFILLER_48_564 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1113_ net135 VGND VPWR net482 hold257/A clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_748 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__530_ u_ppwm_u_ex__530_/Y net393 net382 VPWR VGND sg13g2_nand2b_1
XFILLER_17_984 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1044_ net433 VPWR u_ppwm_u_mem__1044_/Y VGND net353 hold155/A sg13g2_o21ai_1
XFILLER_44_781 VPWR VGND sg13g2_decap_8
XFILLER_16_483 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__461_ VGND VPWR u_ppwm_u_ex__426_/Y u_ppwm_u_ex__459_/Y u_ppwm_u_ex__802_/D
+ u_ppwm_u_ex__460_/Y sg13g2_a21oi_1
XFILLER_31_431 VPWR VGND sg13g2_fill_1
XFILLER_32_976 VPWR VGND sg13g2_decap_8
Xhold104 hold104/A VPWR VGND net301 sg13g2_dlygate4sd3_1
XFILLER_8_693 VPWR VGND sg13g2_decap_8
Xhold126 hold126/A VPWR VGND net469 sg13g2_dlygate4sd3_1
Xhold115 hold115/A VPWR VGND net458 sg13g2_dlygate4sd3_1
Xhold148 hold148/A VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold137 hold137/A VPWR VGND net480 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0828_ hold178/A net412 u_ppwm_u_mem__0828_/Y VPWR VGND sg13g2_nor2b_1
Xhold159 hold159/A VPWR VGND net502 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0759_ hold142/A hold155/A net412 u_ppwm_u_mem__0760_/B VPWR VGND sg13g2_mux2_1
XFILLER_39_520 VPWR VGND sg13g2_decap_8
XFILLER_39_597 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__728_ VPWR VGND net641 u_ppwm_u_ex__726_/Y net312 net323 u_ppwm_u_ex__728_/Y
+ fanout317/A sg13g2_a221oi_1
XFILLER_23_910 VPWR VGND sg13g2_decap_8
XFILLER_35_792 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__659_ u_ppwm_u_ex__659_/Y u_ppwm_u_ex__659_/B u_ppwm_u_ex__644_/B VPWR
+ VGND sg13g2_nand2b_1
XFILLER_22_453 VPWR VGND sg13g2_decap_8
XFILLER_23_987 VPWR VGND sg13g2_decap_8
XFILLER_6_608 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_814 VPWR VGND sg13g2_decap_8
XFILLER_1_302 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_379 VPWR VGND sg13g2_decap_8
XFILLER_40_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_236 VPWR VGND sg13g2_decap_8
XFILLER_18_737 VPWR VGND sg13g2_decap_8
XFILLER_45_556 VPWR VGND sg13g2_decap_8
XFILLER_33_729 VPWR VGND sg13g2_decap_8
XFILLER_13_420 VPWR VGND sg13g2_decap_8
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_41_773 VPWR VGND sg13g2_decap_8
XFILLER_9_402 VPWR VGND sg13g2_decap_8
XFILLER_13_497 VPWR VGND sg13g2_decap_8
XFILLER_9_479 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__233__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_5_696 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0613_ VPWR u_ppwm_u_mem__0613_/Y net206 VGND sg13g2_inv_1
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_48_361 VPWR VGND sg13g2_decap_8
XFILLER_36_545 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1169__138 VPWR VGND net138 sg13g2_tiehi
Xu_ppwm_u_ex__513_ u_ppwm_u_ex__519_/A hold271/A u_ppwm_u_ex__515_/C VPWR VGND sg13g2_nor2_1
XFILLER_17_781 VPWR VGND sg13g2_decap_8
XFILLER_23_206 VPWR VGND sg13g2_fill_1
XFILLER_16_280 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1027_ VGND VPWR net341 u_ppwm_u_mem__0641_/Y u_ppwm_u_mem__1190_/D
+ u_ppwm_u_mem__1026_/Y sg13g2_a21oi_1
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_902 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__444_ VPWR u_ppwm_u_ex__444_/Y u_ppwm_u_ex__488_/A VGND sg13g2_inv_1
XFILLER_32_773 VPWR VGND sg13g2_decap_8
XFILLER_31_272 VPWR VGND sg13g2_decap_8
XFILLER_20_979 VPWR VGND sg13g2_decap_8
XFILLER_8_490 VPWR VGND sg13g2_decap_8
Xfanout403 hold295/A net403 VPWR VGND sg13g2_buf_8
Xfanout414 net421 net414 VPWR VGND sg13g2_buf_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
Xfanout425 net427 net425 VPWR VGND sg13g2_buf_1
Xfanout436 net437 net436 VPWR VGND sg13g2_buf_8
Xfanout447 net448 net447 VPWR VGND sg13g2_buf_8
XFILLER_39_383 VPWR VGND sg13g2_decap_8
XFILLER_15_718 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_14_206 VPWR VGND sg13g2_decap_8
XFILLER_42_559 VPWR VGND sg13g2_decap_8
XFILLER_23_784 VPWR VGND sg13g2_decap_8
XFILLER_11_946 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_6_405 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_2_611 VPWR VGND sg13g2_decap_8
XFILLER_2_688 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_1_198 VPWR VGND sg13g2_decap_8
XFILLER_18_534 VPWR VGND sg13g2_decap_8
XFILLER_46_854 VPWR VGND sg13g2_decap_8
XFILLER_14_751 VPWR VGND sg13g2_decap_8
XFILLER_41_570 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__197_ net337 hold153/A u_ppwm_u_pwm__197_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_6_972 VPWR VGND sg13g2_decap_8
XFILLER_5_493 VPWR VGND sg13g2_decap_8
XFILLER_36_353 VPWR VGND sg13g2_decap_8
XFILLER_37_876 VPWR VGND sg13g2_decap_8
XFILLER_24_559 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__427_ u_ppwm_u_ex__637_/A u_ppwm/instr\[0\] VPWR VGND sg13g2_inv_2
XFILLER_32_570 VPWR VGND sg13g2_decap_8
XFILLER_20_776 VPWR VGND sg13g2_decap_8
Xclkload7 clknet_5_22__leaf_clk clkload7/X VPWR VGND sg13g2_buf_1
Xu_ppwm_u_mem__1223__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_4_909 VPWR VGND sg13g2_decap_8
XFILLER_27_342 VPWR VGND sg13g2_decap_8
XFILLER_28_865 VPWR VGND sg13g2_decap_8
XFILLER_43_824 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_decap_8
XFILLER_11_743 VPWR VGND sg13g2_decap_8
XFILLER_23_581 VPWR VGND sg13g2_decap_8
XFILLER_7_769 VPWR VGND sg13g2_decap_8
XFILLER_6_279 VPWR VGND sg13g2_decap_4
XFILLER_3_964 VPWR VGND sg13g2_decap_8
XFILLER_2_485 VPWR VGND sg13g2_decap_8
XFILLER_37_106 VPWR VGND sg13g2_fill_1
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_810 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_19_887 VPWR VGND sg13g2_decap_8
XFILLER_34_824 VPWR VGND sg13g2_decap_8
XFILLER_45_183 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1133__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_33_367 VPWR VGND sg13g2_fill_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
Xhold19 hold19/A VPWR VGND net216 sg13g2_dlygate4sd3_1
XFILLER_28_117 VPWR VGND sg13g2_fill_2
XFILLER_25_835 VPWR VGND sg13g2_decap_8
XFILLER_37_673 VPWR VGND sg13g2_decap_8
XFILLER_36_183 VPWR VGND sg13g2_decap_4
XFILLER_24_367 VPWR VGND sg13g2_fill_2
XFILLER_40_849 VPWR VGND sg13g2_decap_8
XFILLER_33_890 VPWR VGND sg13g2_decap_8
XFILLER_20_573 VPWR VGND sg13g2_decap_8
XFILLER_4_706 VPWR VGND sg13g2_decap_8
XFILLER_0_967 VPWR VGND sg13g2_decap_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_47_437 VPWR VGND sg13g2_decap_8
XFILLER_19_117 VPWR VGND sg13g2_decap_8
XFILLER_28_662 VPWR VGND sg13g2_decap_8
XFILLER_43_621 VPWR VGND sg13g2_decap_8
XFILLER_16_868 VPWR VGND sg13g2_decap_8
XFILLER_31_816 VPWR VGND sg13g2_decap_8
XFILLER_43_698 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_fill_1
XFILLER_30_326 VPWR VGND sg13g2_fill_2
XFILLER_11_540 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0930_ net443 VPWR u_ppwm_u_mem__0930_/Y VGND net364 net289 sg13g2_o21ai_1
Xu_ppwm_u_mem__0861_ VGND VPWR net360 u_ppwm_u_mem__0724_/Y hold169/A u_ppwm_u_mem__0860_/Y
+ sg13g2_a21oi_1
XFILLER_7_566 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0792_ net408 u_ppwm_u_mem__0785_/Y u_ppwm_u_mem__0787_/Y u_ppwm_u_mem__0791_/Y
+ u_ppwm_u_mem__0789_/Y fanout333/A u_ppwm_u_mem__0792_/X VPWR VGND sg13g2_mux4_1
XFILLER_3_761 VPWR VGND sg13g2_decap_8
XFILLER_39_905 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__121_ net440 VGND VPWR net578 hold234/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__761_ u_ppwm_u_ex__761_/B u_ppwm_u_ex__785_/B u_ppwm_u_ex__761_/A u_ppwm_u_ex__762_/C
+ VPWR VGND sg13g2_nand3_1
XFILLER_20_1000 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__692_ u_ppwm_u_ex__692_/B u_ppwm_u_ex__692_/C net316 u_ppwm_u_ex__692_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_19_684 VPWR VGND sg13g2_decap_8
XFILLER_34_621 VPWR VGND sg13g2_decap_8
XFILLER_22_838 VPWR VGND sg13g2_decap_8
XFILLER_34_698 VPWR VGND sg13g2_decap_8
XFILLER_30_860 VPWR VGND sg13g2_decap_8
XFILLER_0_208 VPWR VGND sg13g2_decap_8
XFILLER_16_109 VPWR VGND sg13g2_fill_1
XFILLER_25_632 VPWR VGND sg13g2_decap_8
XFILLER_13_805 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_fill_2
XFILLER_40_646 VPWR VGND sg13g2_decap_8
XFILLER_21_871 VPWR VGND sg13g2_decap_8
XFILLER_4_503 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1179__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_0_764 VPWR VGND sg13g2_decap_8
XFILLER_48_746 VPWR VGND sg13g2_decap_8
XFILLER_47_223 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1060_ net428 VPWR u_ppwm_u_mem__1060_/Y VGND net340 net286 sg13g2_o21ai_1
XFILLER_44_963 VPWR VGND sg13g2_decap_8
XFILLER_16_665 VPWR VGND sg13g2_decap_8
XFILLER_43_495 VPWR VGND sg13g2_decap_8
XFILLER_31_613 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0913_ VGND VPWR net359 u_ppwm_u_mem__0698_/Y hold58/A u_ppwm_u_mem__0912_/Y
+ sg13g2_a21oi_1
XFILLER_8_875 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_fill_2
Xhold308 hold308/A VPWR VGND net651 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0844_ hold201/A hold173/A net410 u_ppwm_u_mem__0845_/B VPWR VGND sg13g2_mux2_1
Xhold319 hold319/A VPWR VGND net662 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0775_ hold89/A hold200/A net410 u_ppwm_u_mem__0776_/B VPWR VGND sg13g2_mux2_1
XFILLER_39_702 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__243__188 VPWR VGND net188 sg13g2_tiehi
Xu_ppwm_u_ex__813_ net49 VGND VPWR net669 hold325/A clknet_5_3__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_global_counter__104_ VGND VPWR u_ppwm_u_global_counter__058_/Y u_ppwm_u_global_counter__101_/Y
+ hold222/A u_ppwm_u_global_counter__105_/B sg13g2_a21oi_1
XFILLER_39_779 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__744_ u_ppwm_u_ex__744_/B u_ppwm_u_ex__744_/C net316 u_ppwm_u_ex__744_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_26_429 VPWR VGND sg13g2_decap_4
XFILLER_19_481 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__675_ net425 VPWR u_ppwm_u_ex__675_/Y VGND net391 net310 sg13g2_o21ai_1
Xu_ppwm_u_mem__1189_ net58 VGND VPWR u_ppwm_u_mem__1189_/D hold28/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_974 VPWR VGND sg13g2_decap_8
XFILLER_22_635 VPWR VGND sg13g2_decap_8
XFILLER_18_919 VPWR VGND sg13g2_decap_8
XFILLER_45_738 VPWR VGND sg13g2_decap_8
XFILLER_26_930 VPWR VGND sg13g2_decap_8
XFILLER_13_602 VPWR VGND sg13g2_decap_8
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_12_145 VPWR VGND sg13g2_fill_1
XFILLER_13_679 VPWR VGND sg13g2_decap_8
XFILLER_5_801 VPWR VGND sg13g2_decap_8
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_4_377 VPWR VGND sg13g2_decap_8
XFILLER_0_561 VPWR VGND sg13g2_decap_8
XFILLER_48_543 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1112_ net137 VGND VPWR net601 hold189/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_727 VPWR VGND sg13g2_decap_8
XFILLER_44_760 VPWR VGND sg13g2_decap_8
XFILLER_17_963 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1043_ VGND VPWR net342 u_ppwm_u_mem__0633_/Y hold156/A u_ppwm_u_mem__1042_/Y
+ sg13g2_a21oi_1
XFILLER_35_248 VPWR VGND sg13g2_fill_2
XFILLER_16_462 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__460_ net443 VPWR u_ppwm_u_ex__460_/Y VGND u_ppwm_u_ex__426_/Y u_ppwm_u_ex__459_/Y
+ sg13g2_o21ai_1
XFILLER_32_955 VPWR VGND sg13g2_decap_8
XFILLER_8_672 VPWR VGND sg13g2_decap_8
Xhold105 hold105/A VPWR VGND net302 sg13g2_dlygate4sd3_1
XFILLER_7_193 VPWR VGND sg13g2_fill_2
Xhold116 hold116/A VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold149 hold149/A VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold127 hold127/A VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold138 hold138/A VPWR VGND net481 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0827_ u_ppwm_u_mem__0826_/Y u_ppwm_u_mem__0825_/Y u_ppwm_u_mem__0816_/Y
+ fanout326/A VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_mem__0758_ hold15/A hold36/A net410 u_ppwm_u_mem__0758_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0689_ VPWR u_ppwm_u_mem__0689_/Y net494 VGND sg13g2_inv_1
XFILLER_39_576 VPWR VGND sg13g2_decap_8
XFILLER_27_749 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__727_ VGND VPWR net384 net314 u_ppwm_u_ex__727_/Y u_ppwm_u_ex__714_/Y
+ sg13g2_a21oi_1
XFILLER_26_259 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__658_ VGND VPWR u_ppwm_u_ex__655_/Y u_ppwm_u_ex__656_/Y hold322/A u_ppwm_u_ex__657_/Y
+ sg13g2_a21oi_1
XFILLER_34_270 VPWR VGND sg13g2_decap_4
XFILLER_35_771 VPWR VGND sg13g2_decap_8
XFILLER_22_432 VPWR VGND sg13g2_decap_8
XFILLER_23_966 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__589_ u_ppwm_u_ex__591_/C net388 hold271/A VPWR VGND sg13g2_nand2b_1
XFILLER_1_358 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_40_1003 VPWR VGND sg13g2_decap_8
XFILLER_18_716 VPWR VGND sg13g2_decap_8
XFILLER_45_535 VPWR VGND sg13g2_decap_8
XFILLER_33_708 VPWR VGND sg13g2_decap_8
XFILLER_14_933 VPWR VGND sg13g2_decap_8
XFILLER_41_752 VPWR VGND sg13g2_decap_8
XFILLER_13_476 VPWR VGND sg13g2_decap_8
XFILLER_40_262 VPWR VGND sg13g2_fill_1
XFILLER_9_458 VPWR VGND sg13g2_decap_8
XFILLER_5_675 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_fill_2
XFILLER_48_340 VPWR VGND sg13g2_decap_8
XFILLER_49_896 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__512_ hold221/A net379 u_ppwm_u_ex__515_/B VPWR VGND sg13g2_nor2b_1
XFILLER_17_760 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1026_ net428 VPWR u_ppwm_u_mem__1026_/Y VGND net340 net516 sg13g2_o21ai_1
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_32_752 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__443_ net402 net406 net400 u_ppwm_u_ex__488_/A VPWR VGND net413 sg13g2_nand4_1
XFILLER_31_240 VPWR VGND sg13g2_decap_8
XFILLER_20_958 VPWR VGND sg13g2_decap_8
Xfanout404 net406 net404 VPWR VGND sg13g2_buf_8
Xfanout426 net427 net426 VPWR VGND sg13g2_buf_8
Xfanout437 net452 net437 VPWR VGND sg13g2_buf_8
Xfanout448 net451 net448 VPWR VGND sg13g2_buf_8
Xfanout415 net421 net415 VPWR VGND sg13g2_buf_8
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_42_538 VPWR VGND sg13g2_decap_8
XFILLER_14_218 VPWR VGND sg13g2_fill_2
XFILLER_11_925 VPWR VGND sg13g2_decap_8
XFILLER_23_763 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_22_262 VPWR VGND sg13g2_fill_2
XFILLER_2_667 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_1_177 VPWR VGND sg13g2_decap_8
XFILLER_46_833 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1145__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_18_513 VPWR VGND sg13g2_decap_8
XFILLER_45_398 VPWR VGND sg13g2_fill_2
XFILLER_14_730 VPWR VGND sg13g2_decap_8
XFILLER_9_233 VPWR VGND sg13g2_fill_2
XFILLER_10_991 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__196_ u_ppwm_u_pwm__196_/Y net337 hold153/A VPWR VGND sg13g2_nand2b_1
XFILLER_6_951 VPWR VGND sg13g2_decap_8
XFILLER_5_472 VPWR VGND sg13g2_decap_8
XFILLER_49_693 VPWR VGND sg13g2_decap_8
XFILLER_37_855 VPWR VGND sg13g2_decap_8
XFILLER_24_538 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1009_ VGND VPWR net347 u_ppwm_u_mem__0650_/Y u_ppwm_u_mem__1181_/D
+ u_ppwm_u_mem__1008_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__426_ VPWR u_ppwm_u_ex__426_/Y net415 VGND sg13g2_inv_1
XFILLER_20_755 VPWR VGND sg13g2_decap_8
Xclkload8 clknet_5_25__leaf_clk clkload8/X VPWR VGND sg13g2_buf_1
XFILLER_47_619 VPWR VGND sg13g2_decap_8
XFILLER_43_803 VPWR VGND sg13g2_decap_8
XFILLER_27_321 VPWR VGND sg13g2_decap_8
XFILLER_28_844 VPWR VGND sg13g2_decap_8
XFILLER_23_560 VPWR VGND sg13g2_decap_8
XFILLER_11_722 VPWR VGND sg13g2_decap_8
XFILLER_7_748 VPWR VGND sg13g2_decap_8
XFILLER_11_799 VPWR VGND sg13g2_decap_8
XFILLER_10_287 VPWR VGND sg13g2_decap_4
XFILLER_6_269 VPWR VGND sg13g2_decap_4
XFILLER_40_96 VPWR VGND sg13g2_fill_1
XFILLER_3_943 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_46_630 VPWR VGND sg13g2_decap_8
XFILLER_19_866 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_decap_8
XFILLER_18_376 VPWR VGND sg13g2_decap_4
XFILLER_34_803 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__239__182 VPWR VGND net182 sg13g2_tiehi
Xu_ppwm_u_pwm__179_ VGND VPWR u_ppwm_u_pwm__181_/B u_ppwm_u_pwm__182_/C net626 sg13g2_or2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_29_619 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_49_490 VPWR VGND sg13g2_decap_8
XFILLER_37_652 VPWR VGND sg13g2_decap_8
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_40_828 VPWR VGND sg13g2_decap_8
XFILLER_20_552 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_0_946 VPWR VGND sg13g2_decap_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
XFILLER_19_31 VPWR VGND sg13g2_fill_2
XFILLER_28_641 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_decap_8
XFILLER_16_847 VPWR VGND sg13g2_decap_8
XFILLER_43_677 VPWR VGND sg13g2_decap_8
XFILLER_15_357 VPWR VGND sg13g2_decap_4
XFILLER_30_305 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0860_ net447 VPWR u_ppwm_u_mem__0860_/Y VGND net360 u_ppwm_u_mem__1107_/Q
+ sg13g2_o21ai_1
XFILLER_7_545 VPWR VGND sg13g2_decap_8
XFILLER_11_596 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0791_ u_ppwm_u_mem__0790_/Y VPWR u_ppwm_u_mem__0791_/Y VGND u_ppwm_u_mem__0723_/Y
+ net418 sg13g2_o21ai_1
XFILLER_3_740 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__120_ net440 VGND VPWR net554 hold209/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__760_ u_ppwm_u_ex__761_/B u_ppwm_u_ex__761_/A u_ppwm_u_ex__785_/B u_ppwm_u_ex__762_/B
+ VPWR VGND sg13g2_a21o_1
XFILLER_47_983 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__691_ u_ppwm_u_ex__690_/B u_ppwm_u_ex__690_/A u_ppwm_u_ex__696_/D u_ppwm_u_ex__692_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_19_663 VPWR VGND sg13g2_decap_8
XFILLER_34_600 VPWR VGND sg13g2_decap_8
XFILLER_22_817 VPWR VGND sg13g2_decap_8
XFILLER_34_677 VPWR VGND sg13g2_decap_8
XFILLER_33_187 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0989_ VGND VPWR net351 u_ppwm_u_mem__0660_/Y hold74/A u_ppwm_u_mem__0988_/Y
+ sg13g2_a21oi_1
XFILLER_25_611 VPWR VGND sg13g2_decap_8
XFILLER_37_482 VPWR VGND sg13g2_fill_1
XFILLER_40_625 VPWR VGND sg13g2_decap_8
XFILLER_25_688 VPWR VGND sg13g2_decap_8
XFILLER_21_850 VPWR VGND sg13g2_decap_8
XFILLER_4_559 VPWR VGND sg13g2_decap_8
XFILLER_0_743 VPWR VGND sg13g2_decap_8
XFILLER_48_725 VPWR VGND sg13g2_decap_8
XFILLER_47_202 VPWR VGND sg13g2_decap_8
XFILLER_36_909 VPWR VGND sg13g2_decap_8
XFILLER_47_257 VPWR VGND sg13g2_fill_2
XFILLER_29_983 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_fill_1
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_15_110 VPWR VGND sg13g2_decap_4
XFILLER_16_644 VPWR VGND sg13g2_decap_8
XFILLER_43_474 VPWR VGND sg13g2_decap_8
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_15_176 VPWR VGND sg13g2_decap_8
XFILLER_31_669 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0912_ net443 VPWR u_ppwm_u_mem__0912_/Y VGND net358 hold227/A sg13g2_o21ai_1
XFILLER_8_854 VPWR VGND sg13g2_decap_8
XFILLER_12_894 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0843_ u_ppwm_u_mem__0842_/Y VPWR fanout324/A VGND u_ppwm_u_mem__0835_/Y
+ u_ppwm_u_mem__0836_/Y sg13g2_o21ai_1
Xhold309 hold309/A VPWR VGND net652 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0774_ u_ppwm_u_mem__0773_/X u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0764_/Y
+ u_ppwm/instr\[1\] VPWR VGND sg13g2_a21o_2
Xu_ppwm_u_ex__812_ net26 VGND VPWR u_ppwm_u_ex__812_/D hold332/A clknet_5_7__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_global_counter__103_ net564 net331 u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__103_/D
+ u_ppwm_u_global_counter__105_/B VPWR VGND sg13g2_and4_1
XFILLER_39_758 VPWR VGND sg13g2_decap_8
XFILLER_19_460 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__743_ u_ppwm_u_ex__742_/B u_ppwm_u_ex__742_/A u_ppwm_u_ex__748_/B u_ppwm_u_ex__744_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_47_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__674_ VPWR VGND net392 net309 net311 net389 u_ppwm_u_ex__674_/Y net313
+ sg13g2_a221oi_1
XFILLER_35_953 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1188_ net62 VGND VPWR net226 hold42/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_21_102 VPWR VGND sg13g2_fill_1
XFILLER_22_614 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1109__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_29_224 VPWR VGND sg13g2_decap_8
XFILLER_45_717 VPWR VGND sg13g2_decap_8
XFILLER_44_205 VPWR VGND sg13g2_decap_8
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_25_485 VPWR VGND sg13g2_decap_8
XFILLER_26_986 VPWR VGND sg13g2_decap_8
XFILLER_13_658 VPWR VGND sg13g2_decap_8
XFILLER_8_139 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1162__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_5_857 VPWR VGND sg13g2_decap_8
XFILLER_4_356 VPWR VGND sg13g2_decap_8
XFILLER_0_540 VPWR VGND sg13g2_decap_8
XFILLER_48_522 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1111_ net139 VGND VPWR net533 hold184/A clknet_5_23__leaf_clk sg13g2_dfrbpq_2
XFILLER_36_706 VPWR VGND sg13g2_decap_8
XFILLER_48_599 VPWR VGND sg13g2_decap_8
XFILLER_29_780 VPWR VGND sg13g2_decap_8
XFILLER_16_441 VPWR VGND sg13g2_decap_8
XFILLER_17_942 VPWR VGND sg13g2_decap_8
XFILLER_28_290 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1042_ net433 VPWR u_ppwm_u_mem__1042_/Y VGND net342 net266 sg13g2_o21ai_1
XFILLER_32_934 VPWR VGND sg13g2_decap_8
XFILLER_43_271 VPWR VGND sg13g2_fill_1
XFILLER_12_691 VPWR VGND sg13g2_decap_8
XFILLER_8_651 VPWR VGND sg13g2_decap_8
Xhold106 hold106/A VPWR VGND net303 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0826_ VGND VPWR u_ppwm_u_mem__0818_/Y u_ppwm_u_mem__0820_/Y u_ppwm_u_mem__0826_/Y
+ net401 sg13g2_a21oi_1
Xhold117 hold117/A VPWR VGND net460 sg13g2_dlygate4sd3_1
Xhold128 hold128/A VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold139 hold139/A VPWR VGND net482 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0757_ u_ppwm_u_mem__0756_/Y u_ppwm_u_mem__0751_/Y u_ppwm_u_mem__0749_/Y
+ u_ppwm/instr\[0\] VPWR VGND sg13g2_a21o_2
Xu_ppwm_u_mem__0688_ VPWR u_ppwm_u_mem__0688_/Y net459 VGND sg13g2_inv_1
XFILLER_39_555 VPWR VGND sg13g2_decap_8
XFILLER_27_728 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__726_ VGND VPWR u_ppwm_u_ex__716_/Y u_ppwm_u_ex__724_/Y u_ppwm_u_ex__726_/Y
+ u_ppwm_u_ex__725_/Y sg13g2_a21oi_1
XFILLER_26_238 VPWR VGND sg13g2_decap_8
XFILLER_35_750 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__657_ net427 VPWR u_ppwm_u_ex__657_/Y VGND net394 fanout310/A sg13g2_o21ai_1
XFILLER_23_945 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__588_ u_ppwm_u_ex__593_/B hold308/A hold7/A VPWR VGND sg13g2_nand2b_1
XFILLER_22_488 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1226__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_2_849 VPWR VGND sg13g2_decap_8
XFILLER_1_337 VPWR VGND sg13g2_decap_8
XFILLER_49_308 VPWR VGND sg13g2_decap_8
XFILLER_27_20 VPWR VGND sg13g2_fill_1
XFILLER_45_514 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_26_783 VPWR VGND sg13g2_decap_8
XFILLER_41_731 VPWR VGND sg13g2_decap_8
XFILLER_13_455 VPWR VGND sg13g2_decap_8
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_43_96 VPWR VGND sg13g2_decap_4
XFILLER_9_437 VPWR VGND sg13g2_decap_8
XFILLER_5_654 VPWR VGND sg13g2_decap_8
XFILLER_49_875 VPWR VGND sg13g2_decap_8
XFILLER_48_396 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__511_ u_ppwm_u_ex__515_/A u_ppwm_u_ex__511_/B u_ppwm_u_ex__509_/Y VPWR
+ VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1025_ VGND VPWR net346 u_ppwm_u_mem__0642_/Y u_ppwm_u_mem__1189_/D
+ u_ppwm_u_mem__1024_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__442_ net406 net412 net402 u_ppwm_u_ex__442_/Y VPWR VGND sg13g2_nand3_1
XFILLER_32_731 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_937 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0809_ u_ppwm_u_mem__0808_/Y u_ppwm_u_mem__0806_/Y u_ppwm_u_mem__0802_/Y
+ fanout327/A VPWR VGND sg13g2_a21o_2
Xfanout405 net406 net405 VPWR VGND sg13g2_buf_1
Xfanout438 net439 net438 VPWR VGND sg13g2_buf_8
Xfanout427 net437 net427 VPWR VGND sg13g2_buf_8
Xfanout416 net421 net416 VPWR VGND sg13g2_buf_8
Xfanout449 net451 net449 VPWR VGND sg13g2_buf_8
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_42_517 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__709_ u_ppwm_u_ex__709_/Y u_ppwm_u_ex__709_/A u_ppwm_u_ex__709_/B VPWR
+ VGND sg13g2_xnor2_1
XFILLER_23_742 VPWR VGND sg13g2_decap_8
XFILLER_11_904 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_22_274 VPWR VGND sg13g2_fill_1
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_2_646 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_45_300 VPWR VGND sg13g2_fill_1
XFILLER_18_569 VPWR VGND sg13g2_decap_8
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_26_580 VPWR VGND sg13g2_decap_8
XFILLER_13_230 VPWR VGND sg13g2_decap_4
XFILLER_14_786 VPWR VGND sg13g2_decap_8
XFILLER_6_930 VPWR VGND sg13g2_decap_8
XFILLER_10_970 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__195_ hold153/A net337 u_ppwm_u_pwm__195_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_5_451 VPWR VGND sg13g2_decap_8
XFILLER_49_672 VPWR VGND sg13g2_decap_8
XFILLER_37_834 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_344 VPWR VGND sg13g2_decap_4
XFILLER_24_517 VPWR VGND sg13g2_decap_8
XFILLER_36_377 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1008_ net430 VPWR u_ppwm_u_mem__1008_/Y VGND net346 net293 sg13g2_o21ai_1
Xu_ppwm_u_ex__425_ VPWR u_ppwm_u_ex__529_/B net396 VGND sg13g2_inv_1
XFILLER_20_734 VPWR VGND sg13g2_decap_8
Xclkload9 clknet_5_26__leaf_clk clkload9/X VPWR VGND sg13g2_buf_1
XFILLER_30_1014 VPWR VGND sg13g2_decap_8
XFILLER_8_1015 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_4
XFILLER_28_823 VPWR VGND sg13g2_decap_8
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_42_358 VPWR VGND sg13g2_decap_8
XFILLER_11_701 VPWR VGND sg13g2_decap_8
XFILLER_7_727 VPWR VGND sg13g2_decap_8
XFILLER_11_778 VPWR VGND sg13g2_decap_8
XFILLER_40_53 VPWR VGND sg13g2_fill_2
XFILLER_3_922 VPWR VGND sg13g2_decap_8
XFILLER_3_999 VPWR VGND sg13g2_decap_8
XFILLER_2_443 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_18_311 VPWR VGND sg13g2_decap_8
XFILLER_19_845 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_decap_8
XFILLER_34_859 VPWR VGND sg13g2_decap_8
XFILLER_33_358 VPWR VGND sg13g2_decap_8
XFILLER_42_881 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__247_ net176 VGND VPWR u_ppwm_u_pwm__247_/D net2 clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__178_ u_ppwm_u_pwm__182_/C net644 hold302/A VPWR VGND sg13g2_nor2_1
XFILLER_37_631 VPWR VGND sg13g2_decap_8
XFILLER_36_152 VPWR VGND sg13g2_decap_8
XFILLER_40_807 VPWR VGND sg13g2_decap_8
XFILLER_12_509 VPWR VGND sg13g2_decap_8
XFILLER_20_531 VPWR VGND sg13g2_decap_8
XFILLER_0_925 VPWR VGND sg13g2_decap_8
XFILLER_48_907 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1119__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_28_620 VPWR VGND sg13g2_decap_8
XFILLER_16_826 VPWR VGND sg13g2_decap_8
XFILLER_15_325 VPWR VGND sg13g2_fill_1
XFILLER_28_697 VPWR VGND sg13g2_decap_8
XFILLER_43_656 VPWR VGND sg13g2_decap_8
XFILLER_37_1009 VPWR VGND sg13g2_decap_8
XFILLER_24_881 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_7_524 VPWR VGND sg13g2_decap_8
XFILLER_11_575 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0790_ u_ppwm_u_mem__0790_/Y hold44/A net417 VPWR VGND sg13g2_nand2_1
XFILLER_3_796 VPWR VGND sg13g2_decap_8
XFILLER_19_642 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__690_ u_ppwm_u_ex__690_/B u_ppwm_u_ex__696_/D u_ppwm_u_ex__690_/A u_ppwm_u_ex__692_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_18_130 VPWR VGND sg13g2_decap_4
XFILLER_18_141 VPWR VGND sg13g2_fill_2
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_18_196 VPWR VGND sg13g2_decap_4
XFILLER_34_656 VPWR VGND sg13g2_decap_8
XFILLER_30_895 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0988_ net431 VPWR u_ppwm_u_mem__0988_/Y VGND net351 hold124/A sg13g2_o21ai_1
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
XFILLER_38_984 VPWR VGND sg13g2_decap_8
XFILLER_25_667 VPWR VGND sg13g2_decap_8
XFILLER_40_604 VPWR VGND sg13g2_decap_8
XFILLER_20_350 VPWR VGND sg13g2_fill_2
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_4_538 VPWR VGND sg13g2_decap_8
XFILLER_0_722 VPWR VGND sg13g2_decap_8
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_48_704 VPWR VGND sg13g2_decap_8
XFILLER_0_799 VPWR VGND sg13g2_decap_8
XFILLER_29_962 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_44_921 VPWR VGND sg13g2_decap_8
XFILLER_16_623 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_fill_2
XFILLER_44_998 VPWR VGND sg13g2_decap_8
XFILLER_31_648 VPWR VGND sg13g2_decap_8
XFILLER_12_873 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0911_ VGND VPWR net372 u_ppwm_u_mem__0699_/Y hold228/A u_ppwm_u_mem__0910_/Y
+ sg13g2_a21oi_1
XFILLER_8_833 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0842_ u_ppwm_u_mem__0842_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0842_/B
+ VPWR VGND sg13g2_nand2_1
XFILLER_7_398 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0773_ net408 u_ppwm_u_mem__0766_/Y u_ppwm_u_mem__0768_/Y u_ppwm_u_mem__0772_/Y
+ u_ppwm_u_mem__0770_/Y net332 u_ppwm_u_mem__0773_/X VPWR VGND sg13g2_mux4_1
XFILLER_3_593 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__811_ net28 VGND VPWR net667 hold323/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_global_counter__102_ u_ppwm_u_global_counter__123_/D u_ppwm_u_global_counter__103_/D
+ u_ppwm_u_global_counter__099_/B u_ppwm_u_global_counter__098_/Y u_ppwm_u_global_counter__057_/Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_39_737 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__742_ u_ppwm_u_ex__742_/B u_ppwm_u_ex__748_/B u_ppwm_u_ex__742_/A u_ppwm_u_ex__744_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_35_932 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__673_ u_ppwm_u_ex__673_/B u_ppwm_u_ex__673_/C net316 u_ppwm_u_ex__673_/Y
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_mem__1187_ net66 VGND VPWR net240 hold165/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_464 VPWR VGND sg13g2_decap_4
XFILLER_30_692 VPWR VGND sg13g2_decap_8
XFILLER_1_519 VPWR VGND sg13g2_decap_8
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_38_781 VPWR VGND sg13g2_decap_8
XFILLER_25_431 VPWR VGND sg13g2_decap_8
XFILLER_26_965 VPWR VGND sg13g2_decap_8
XFILLER_41_913 VPWR VGND sg13g2_decap_8
XFILLER_25_464 VPWR VGND sg13g2_decap_8
XFILLER_12_136 VPWR VGND sg13g2_decap_8
XFILLER_13_637 VPWR VGND sg13g2_decap_8
XFILLER_9_619 VPWR VGND sg13g2_decap_8
XFILLER_32_21 VPWR VGND sg13g2_decap_8
XFILLER_5_836 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_335 VPWR VGND sg13g2_decap_8
XFILLER_48_501 VPWR VGND sg13g2_decap_8
XFILLER_0_596 VPWR VGND sg13g2_decap_8
XFILLER_48_578 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1110_ net141 VGND VPWR u_ppwm_u_mem__1110_/D hold158/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_17_921 VPWR VGND sg13g2_decap_8
XFILLER_16_420 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1041_ VGND VPWR net344 u_ppwm_u_mem__0634_/Y hold70/A u_ppwm_u_mem__1040_/Y
+ sg13g2_a21oi_1
XFILLER_17_998 VPWR VGND sg13g2_decap_8
XFILLER_32_913 VPWR VGND sg13g2_decap_8
XFILLER_44_795 VPWR VGND sg13g2_decap_8
XFILLER_16_497 VPWR VGND sg13g2_decap_8
XFILLER_8_630 VPWR VGND sg13g2_decap_8
XFILLER_12_670 VPWR VGND sg13g2_decap_8
Xhold107 hold107/A VPWR VGND net304 sg13g2_dlygate4sd3_1
XFILLER_7_184 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0825_ u_ppwm_u_mem__0825_/Y u_ppwm_u_mem__0825_/B u_ppwm_u_mem__0822_/Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_7_195 VPWR VGND sg13g2_fill_1
Xhold118 hold118/A VPWR VGND net461 sg13g2_dlygate4sd3_1
Xhold129 hold129/A VPWR VGND net472 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0756_ VGND VPWR u_ppwm_u_mem__0754_/Y u_ppwm_u_mem__0755_/Y u_ppwm_u_mem__0756_/Y
+ net400 sg13g2_a21oi_1
XFILLER_3_390 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0687_ VPWR u_ppwm_u_mem__0687_/Y net466 VGND sg13g2_inv_1
XFILLER_39_501 VPWR VGND sg13g2_fill_2
XFILLER_39_534 VPWR VGND sg13g2_decap_8
XFILLER_27_707 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__725_ net316 VPWR u_ppwm_u_ex__725_/Y VGND u_ppwm_u_ex__716_/Y u_ppwm_u_ex__724_/Y
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__656_ VPWR VGND net396 fanout309/A net311 net392 u_ppwm_u_ex__656_/Y
+ net313 sg13g2_a221oi_1
XFILLER_23_924 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__587_ u_ppwm_u_ex__591_/A hold221/A u_ppwm_u_ex__541_/B hold7/A u_ppwm_u_ex__538_/B
+ VPWR VGND sg13g2_a22oi_1
XFILLER_22_467 VPWR VGND sg13g2_decap_8
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
XFILLER_2_828 VPWR VGND sg13g2_decap_8
XFILLER_1_316 VPWR VGND sg13g2_decap_8
XFILLER_17_217 VPWR VGND sg13g2_fill_1
XFILLER_41_710 VPWR VGND sg13g2_decap_8
XFILLER_25_250 VPWR VGND sg13g2_fill_1
XFILLER_26_762 VPWR VGND sg13g2_decap_8
XFILLER_13_434 VPWR VGND sg13g2_decap_8
XFILLER_43_64 VPWR VGND sg13g2_fill_1
XFILLER_9_416 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_40_242 VPWR VGND sg13g2_fill_2
XFILLER_41_787 VPWR VGND sg13g2_decap_8
XFILLER_5_633 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_fill_2
XFILLER_1_883 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_8
XFILLER_0_393 VPWR VGND sg13g2_decap_8
XFILLER_48_375 VPWR VGND sg13g2_decap_8
XFILLER_36_559 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__510_ u_ppwm_u_ex__511_/B hold305/A hold7/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1024_ net428 VPWR u_ppwm_u_mem__1024_/Y VGND net346 net225 sg13g2_o21ai_1
XFILLER_44_592 VPWR VGND sg13g2_decap_8
XFILLER_17_795 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__441_ u_ppwm_u_ex__472_/B net407 net413 VPWR VGND sg13g2_nand2_1
XFILLER_32_710 VPWR VGND sg13g2_decap_8
XFILLER_20_916 VPWR VGND sg13g2_decap_8
XFILLER_32_787 VPWR VGND sg13g2_decap_8
XFILLER_31_297 VPWR VGND sg13g2_fill_2
XFILLER_9_983 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0808_ VGND VPWR net332 u_ppwm_u_mem__0807_/X u_ppwm_u_mem__0808_/Y
+ net401 sg13g2_a21oi_1
Xu_ppwm_u_mem__0739_ net423 net513 net1 u_ppwm_u_mem__0739_/Y VPWR VGND sg13g2_nand3_1
Xfanout439 net442 net439 VPWR VGND sg13g2_buf_8
Xfanout406 net409 net406 VPWR VGND sg13g2_buf_8
Xfanout417 net420 net417 VPWR VGND sg13g2_buf_8
Xfanout428 net432 net428 VPWR VGND sg13g2_buf_8
XFILLER_27_504 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__708_ u_ppwm_u_ex__709_/B hold308/A net319 VPWR VGND sg13g2_xnor2_1
XFILLER_23_721 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__639_ VPWR VGND net649 net309 net311 net396 u_ppwm_u_ex__639_/Y net313
+ sg13g2_a221oi_1
XFILLER_22_264 VPWR VGND sg13g2_fill_1
XFILLER_23_798 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_7_909 VPWR VGND sg13g2_decap_8
XFILLER_6_419 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_fill_2
XFILLER_2_625 VPWR VGND sg13g2_decap_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_18_548 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_41_584 VPWR VGND sg13g2_decap_8
XFILLER_9_213 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1129__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_9_246 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_pwm__194_ u_ppwm_u_pwm__194_/Y hold268/A hold219/A VPWR VGND sg13g2_nand2b_1
XFILLER_5_430 VPWR VGND sg13g2_decap_8
XFILLER_6_986 VPWR VGND sg13g2_decap_8
XFILLER_1_680 VPWR VGND sg13g2_decap_8
XFILLER_49_651 VPWR VGND sg13g2_decap_8
XFILLER_23_1022 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_37_813 VPWR VGND sg13g2_decap_8
XFILLER_17_592 VPWR VGND sg13g2_decap_8
XFILLER_36_389 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1007_ VGND VPWR net348 u_ppwm_u_mem__0651_/Y hold97/A u_ppwm_u_mem__1006_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__424_ VPWR u_ppwm_u_ex__424_/Y net392 VGND sg13g2_inv_1
XFILLER_20_713 VPWR VGND sg13g2_decap_8
XFILLER_32_584 VPWR VGND sg13g2_decap_8
XFILLER_9_780 VPWR VGND sg13g2_decap_8
XFILLER_28_802 VPWR VGND sg13g2_decap_8
XFILLER_39_172 VPWR VGND sg13g2_fill_2
XFILLER_27_356 VPWR VGND sg13g2_fill_1
XFILLER_28_879 VPWR VGND sg13g2_decap_8
XFILLER_43_838 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_fill_2
XFILLER_7_706 VPWR VGND sg13g2_decap_8
XFILLER_11_757 VPWR VGND sg13g2_decap_8
XFILLER_23_595 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_24_99 VPWR VGND sg13g2_fill_2
XFILLER_3_901 VPWR VGND sg13g2_decap_8
XFILLER_2_422 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
XFILLER_3_978 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_2_499 VPWR VGND sg13g2_decap_8
Xhold290 hold290/A VPWR VGND net633 sg13g2_dlygate4sd3_1
XFILLER_19_824 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_34_838 VPWR VGND sg13g2_decap_8
XFILLER_42_860 VPWR VGND sg13g2_decap_8
XFILLER_14_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__246_ net184 VGND VPWR net596 hold318/A clknet_5_5__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__177_ net422 VPWR hold301/A VGND net643 u_ppwm_u_pwm__175_/C sg13g2_o21ai_1
XFILLER_6_783 VPWR VGND sg13g2_decap_8
XFILLER_37_610 VPWR VGND sg13g2_decap_8
XFILLER_25_849 VPWR VGND sg13g2_decap_8
XFILLER_37_687 VPWR VGND sg13g2_decap_8
XFILLER_20_510 VPWR VGND sg13g2_decap_8
XFILLER_20_587 VPWR VGND sg13g2_decap_8
XFILLER_0_904 VPWR VGND sg13g2_decap_8
XFILLER_16_805 VPWR VGND sg13g2_decap_8
XFILLER_27_120 VPWR VGND sg13g2_decap_8
XFILLER_28_676 VPWR VGND sg13g2_decap_8
XFILLER_43_635 VPWR VGND sg13g2_decap_8
XFILLER_24_860 VPWR VGND sg13g2_decap_8
XFILLER_7_503 VPWR VGND sg13g2_decap_8
XFILLER_11_554 VPWR VGND sg13g2_decap_8
XFILLER_3_775 VPWR VGND sg13g2_decap_8
XFILLER_32_9 VPWR VGND sg13g2_fill_1
XFILLER_39_919 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1172__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_19_621 VPWR VGND sg13g2_decap_8
XFILLER_20_1014 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_19_698 VPWR VGND sg13g2_decap_8
XFILLER_34_635 VPWR VGND sg13g2_decap_8
XFILLER_15_893 VPWR VGND sg13g2_decap_8
XFILLER_30_874 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0987_ VGND VPWR net351 u_ppwm_u_mem__0661_/Y hold125/A u_ppwm_u_mem__0986_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__229_ net183 VGND VPWR net497 hold153/A clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_6_580 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1220__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_44_0 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_38_963 VPWR VGND sg13g2_decap_8
XFILLER_37_473 VPWR VGND sg13g2_decap_8
XFILLER_25_646 VPWR VGND sg13g2_decap_8
XFILLER_13_819 VPWR VGND sg13g2_decap_8
XFILLER_36_1021 VPWR VGND sg13g2_decap_8
XFILLER_21_885 VPWR VGND sg13g2_decap_8
XFILLER_4_517 VPWR VGND sg13g2_decap_8
XFILLER_0_701 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__229__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_0_778 VPWR VGND sg13g2_decap_8
XFILLER_47_237 VPWR VGND sg13g2_decap_8
XFILLER_29_941 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_fill_1
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_16_602 VPWR VGND sg13g2_decap_8
XFILLER_28_462 VPWR VGND sg13g2_fill_1
XFILLER_44_977 VPWR VGND sg13g2_decap_8
XFILLER_16_679 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__825__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_31_627 VPWR VGND sg13g2_decap_8
XFILLER_8_812 VPWR VGND sg13g2_decap_8
XFILLER_12_852 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0910_ net449 VPWR u_ppwm_u_mem__0910_/Y VGND net372 net299 sg13g2_o21ai_1
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_8_889 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0841_ net407 u_ppwm_u_mem__0837_/X u_ppwm_u_mem__0838_/X u_ppwm_u_mem__0840_/X
+ u_ppwm_u_mem__0839_/X net332 u_ppwm_u_mem__0842_/B VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0772_ u_ppwm_u_mem__0771_/Y VPWR u_ppwm_u_mem__0772_/Y VGND u_ppwm_u_mem__0724_/Y
+ net420 sg13g2_o21ai_1
XFILLER_3_572 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__810_ net30 VGND VPWR net665 hold321/A clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_39_716 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__101_ u_ppwm_u_global_counter__103_/C u_ppwm_u_global_counter__103_/D
+ fanout331/A u_ppwm_u_global_counter__101_/Y VPWR VGND sg13g2_nand3_1
XFILLER_16_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__741_ u_ppwm_u_ex__748_/B net383 net322 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__672_ u_ppwm_u_ex__671_/B u_ppwm_u_ex__671_/A u_ppwm_u_ex__696_/B u_ppwm_u_ex__673_/C
+ VPWR VGND sg13g2_a21o_1
XFILLER_34_410 VPWR VGND sg13g2_fill_1
XFILLER_35_911 VPWR VGND sg13g2_decap_8
XFILLER_19_495 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1186_ net70 VGND VPWR net509 hold195/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_988 VPWR VGND sg13g2_decap_8
XFILLER_15_690 VPWR VGND sg13g2_decap_8
XFILLER_22_649 VPWR VGND sg13g2_decap_8
XFILLER_30_671 VPWR VGND sg13g2_decap_8
XFILLER_38_760 VPWR VGND sg13g2_decap_8
XFILLER_25_443 VPWR VGND sg13g2_decap_8
XFILLER_26_944 VPWR VGND sg13g2_decap_8
XFILLER_37_292 VPWR VGND sg13g2_decap_4
XFILLER_13_616 VPWR VGND sg13g2_decap_8
XFILLER_16_67 VPWR VGND sg13g2_fill_1
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_12_159 VPWR VGND sg13g2_fill_2
XFILLER_21_682 VPWR VGND sg13g2_decap_8
XFILLER_5_815 VPWR VGND sg13g2_decap_8
XFILLER_0_575 VPWR VGND sg13g2_decap_8
XFILLER_48_557 VPWR VGND sg13g2_decap_8
XFILLER_17_900 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1040_ net433 VPWR u_ppwm_u_mem__1040_/Y VGND net344 net210 sg13g2_o21ai_1
XFILLER_44_774 VPWR VGND sg13g2_decap_8
XFILLER_43_251 VPWR VGND sg13g2_fill_2
XFILLER_16_476 VPWR VGND sg13g2_decap_8
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_31_402 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1210__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_32_969 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__813__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_11_192 VPWR VGND sg13g2_decap_8
Xhold108 hold108/A VPWR VGND net305 sg13g2_dlygate4sd3_1
XFILLER_8_686 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0824_ VGND VPWR net335 u_ppwm_u_mem__0823_/X u_ppwm_u_mem__0825_/B
+ net332 sg13g2_a21oi_1
Xhold119 hold119/A VPWR VGND net462 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0755_ VGND VPWR net407 u_ppwm_u_mem__0752_/X u_ppwm_u_mem__0755_/Y
+ net332 sg13g2_a21oi_1
Xu_ppwm_u_mem__0686_ VPWR u_ppwm_u_mem__0686_/Y net280 VGND sg13g2_inv_1
XFILLER_4_881 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__724_ u_ppwm_u_ex__724_/Y u_ppwm_u_ex__724_/B u_ppwm_u_ex__722_/X VPWR
+ VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1169_ net138 VGND VPWR net488 hold274/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__655_ u_ppwm_u_ex__654_/Y VPWR u_ppwm_u_ex__655_/Y VGND u_ppwm_u_ex__659_/B
+ u_ppwm_u_ex__653_/X sg13g2_o21ai_1
XFILLER_23_903 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__586_ u_ppwm_u_ex__585_/Y VPWR u_ppwm_u_ex__586_/Y VGND net390 u_ppwm_u_ex__506_/B
+ sg13g2_o21ai_1
XFILLER_35_785 VPWR VGND sg13g2_decap_8
XFILLER_22_446 VPWR VGND sg13g2_decap_8
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
XFILLER_31_991 VPWR VGND sg13g2_decap_8
XFILLER_2_807 VPWR VGND sg13g2_decap_8
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_1017 VPWR VGND sg13g2_decap_8
XFILLER_45_549 VPWR VGND sg13g2_decap_8
XFILLER_26_741 VPWR VGND sg13g2_decap_8
XFILLER_13_413 VPWR VGND sg13g2_decap_8
XFILLER_14_947 VPWR VGND sg13g2_decap_8
XFILLER_41_766 VPWR VGND sg13g2_decap_8
XFILLER_5_612 VPWR VGND sg13g2_decap_8
XFILLER_4_100 VPWR VGND sg13g2_fill_2
XFILLER_5_689 VPWR VGND sg13g2_decap_8
XFILLER_1_862 VPWR VGND sg13g2_decap_8
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_0_372 VPWR VGND sg13g2_decap_8
XFILLER_48_354 VPWR VGND sg13g2_decap_8
XFILLER_36_538 VPWR VGND sg13g2_decap_8
XFILLER_17_774 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1023_ VGND VPWR net347 u_ppwm_u_mem__0643_/Y hold29/A u_ppwm_u_mem__1022_/Y
+ sg13g2_a21oi_1
XFILLER_44_571 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__440_ VPWR u_ppwm_u_ex__440_/Y hold54/A VGND sg13g2_inv_1
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
XFILLER_32_766 VPWR VGND sg13g2_decap_8
XFILLER_13_980 VPWR VGND sg13g2_decap_8
XFILLER_31_254 VPWR VGND sg13g2_decap_8
XFILLER_31_265 VPWR VGND sg13g2_decap_8
XFILLER_9_962 VPWR VGND sg13g2_decap_8
XFILLER_8_483 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0807_ net335 u_ppwm_u_mem__0708_/Y u_ppwm_u_mem__0722_/Y u_ppwm_u_mem__0701_/Y
+ u_ppwm_u_mem__0715_/Y net419 u_ppwm_u_mem__0807_/X VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0738_ u_ppwm_u_mem__0731_/Y net625 u_ppwm_u_mem__0737_/Y u_ppwm_u_mem__1227_/D
+ VPWR VGND sg13g2_a21o_1
Xfanout429 net432 net429 VPWR VGND sg13g2_buf_8
Xfanout407 net408 net407 VPWR VGND sg13g2_buf_8
Xfanout418 net420 net418 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0669_ VPWR u_ppwm_u_mem__0669_/Y net282 VGND sg13g2_inv_1
Xu_ppwm_u_ex__707_ u_ppwm_u_ex__700_/Y VPWR u_ppwm_u_ex__709_/A VGND u_ppwm_u_ex__699_/Y
+ u_ppwm_u_ex__701_/Y sg13g2_o21ai_1
XFILLER_23_700 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__638_ u_ppwm_u_ex__638_/Y net316 u_ppwm_u_ex__636_/X net317 net323 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_35_582 VPWR VGND sg13g2_decap_8
XFILLER_11_939 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__569_ u_ppwm_u_ex__569_/Y u_ppwm_u_ex__435_/Y hold333/A u_ppwm_u_ex__612_/B
+ hold308/A VPWR VGND sg13g2_a22oi_1
XFILLER_23_777 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_2_604 VPWR VGND sg13g2_decap_8
XFILLER_1_103 VPWR VGND sg13g2_fill_2
XFILLER_1_147 VPWR VGND sg13g2_fill_2
XFILLER_46_847 VPWR VGND sg13g2_decap_8
XFILLER_18_527 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1168__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_13_243 VPWR VGND sg13g2_fill_2
XFILLER_14_744 VPWR VGND sg13g2_decap_8
XFILLER_41_563 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__193_ u_ppwm_u_pwm__193_/A net595 u_ppwm_u_pwm__193_/C hold253/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_6_965 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_decap_8
XFILLER_49_630 VPWR VGND sg13g2_decap_8
XFILLER_0_180 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_1001 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_37_869 VPWR VGND sg13g2_decap_8
XFILLER_17_571 VPWR VGND sg13g2_decap_8
XFILLER_36_379 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1006_ net431 VPWR u_ppwm_u_mem__1006_/Y VGND net348 hold167/A sg13g2_o21ai_1
Xu_ppwm_u_ex__423_ u_ppwm_u_ex__583_/A net391 VPWR VGND sg13g2_inv_2
XFILLER_32_563 VPWR VGND sg13g2_decap_8
XFILLER_20_769 VPWR VGND sg13g2_decap_8
XFILLER_27_335 VPWR VGND sg13g2_decap_8
XFILLER_28_858 VPWR VGND sg13g2_decap_8
XFILLER_43_817 VPWR VGND sg13g2_decap_8
XFILLER_15_508 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1142__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_23_574 VPWR VGND sg13g2_decap_8
XFILLER_11_736 VPWR VGND sg13g2_decap_8
XFILLER_40_11 VPWR VGND sg13g2_fill_2
XFILLER_6_239 VPWR VGND sg13g2_fill_1
XFILLER_2_401 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
Xhold280 hold280/A VPWR VGND net623 sg13g2_dlygate4sd3_1
XFILLER_3_957 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_2_478 VPWR VGND sg13g2_decap_8
Xhold291 hold328/A VPWR VGND net634 sg13g2_dlygate4sd3_1
XFILLER_19_803 VPWR VGND sg13g2_decap_8
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_34_817 VPWR VGND sg13g2_decap_8
XFILLER_45_187 VPWR VGND sg13g2_fill_2
XFILLER_14_541 VPWR VGND sg13g2_decap_8
XFILLER_26_390 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_pwm__245_ net194 VGND VPWR u_ppwm_u_pwm__245_/D hold251/A clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_6_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__176_ net643 net621 net660 u_ppwm_u_pwm__176_/D u_ppwm_u_pwm__182_/C
+ VPWR VGND sg13g2_and4_1
XFILLER_5_283 VPWR VGND sg13g2_fill_1
XFILLER_37_666 VPWR VGND sg13g2_decap_8
XFILLER_25_828 VPWR VGND sg13g2_decap_8
XFILLER_36_165 VPWR VGND sg13g2_decap_4
XFILLER_36_187 VPWR VGND sg13g2_fill_1
XFILLER_18_891 VPWR VGND sg13g2_decap_8
XFILLER_33_883 VPWR VGND sg13g2_decap_8
XFILLER_20_566 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_4
XFILLER_19_67 VPWR VGND sg13g2_fill_1
XFILLER_28_655 VPWR VGND sg13g2_decap_8
XFILLER_43_614 VPWR VGND sg13g2_decap_8
XFILLER_31_809 VPWR VGND sg13g2_decap_8
XFILLER_11_533 VPWR VGND sg13g2_decap_8
XFILLER_13_1022 VPWR VGND sg13g2_decap_8
XFILLER_7_559 VPWR VGND sg13g2_decap_8
XFILLER_3_754 VPWR VGND sg13g2_decap_8
XFILLER_2_220 VPWR VGND sg13g2_fill_1
XFILLER_19_600 VPWR VGND sg13g2_decap_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_18_8 VPWR VGND sg13g2_fill_1
XFILLER_46_441 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1213__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_19_677 VPWR VGND sg13g2_decap_8
XFILLER_34_614 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_decap_8
XFILLER_33_179 VPWR VGND sg13g2_fill_2
XFILLER_30_853 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0986_ net434 VPWR u_ppwm_u_mem__0986_/Y VGND net351 hold144/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__228_ net185 VGND VPWR net563 hold219/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__159_ net425 VPWR u_ppwm_u_pwm__159_/Y VGND net386 net329 sg13g2_o21ai_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_38_942 VPWR VGND sg13g2_decap_8
XFILLER_25_625 VPWR VGND sg13g2_decap_8
XFILLER_24_113 VPWR VGND sg13g2_fill_2
XFILLER_37_496 VPWR VGND sg13g2_fill_1
XFILLER_36_1000 VPWR VGND sg13g2_decap_8
XFILLER_40_639 VPWR VGND sg13g2_decap_8
XFILLER_33_680 VPWR VGND sg13g2_decap_8
XFILLER_21_864 VPWR VGND sg13g2_decap_8
XFILLER_20_352 VPWR VGND sg13g2_fill_1
XFILLER_20_396 VPWR VGND sg13g2_fill_2
XFILLER_0_757 VPWR VGND sg13g2_decap_8
XFILLER_48_739 VPWR VGND sg13g2_decap_8
XFILLER_47_216 VPWR VGND sg13g2_decap_8
XFILLER_29_920 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_29_997 VPWR VGND sg13g2_decap_8
XFILLER_44_956 VPWR VGND sg13g2_decap_8
XFILLER_16_658 VPWR VGND sg13g2_decap_8
XFILLER_31_606 VPWR VGND sg13g2_decap_8
XFILLER_43_488 VPWR VGND sg13g2_decap_8
XFILLER_12_831 VPWR VGND sg13g2_decap_8
XFILLER_11_330 VPWR VGND sg13g2_fill_2
XFILLER_11_341 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0840_ hold189/A hold126/A net415 u_ppwm_u_mem__0840_/X VPWR VGND sg13g2_mux2_1
XFILLER_8_868 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0771_ u_ppwm_u_mem__0771_/Y hold217/A net417 VPWR VGND sg13g2_nand2_1
XFILLER_3_551 VPWR VGND sg13g2_decap_8
XFILLER_30_7 VPWR VGND sg13g2_decap_4
XFILLER_23_6 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_global_counter__100_ net198 net614 u_ppwm_u_global_counter__103_/D VPWR
+ VGND sg13g2_and2_1
XFILLER_38_205 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__740_ u_ppwm_u_ex__740_/A u_ppwm_u_ex__740_/B u_ppwm_u_ex__819_/D VPWR
+ VGND sg13g2_nor2_1
Xu_ppwm_u_ex__671_ u_ppwm_u_ex__671_/B u_ppwm_u_ex__696_/B u_ppwm_u_ex__671_/A u_ppwm_u_ex__673_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_19_474 VPWR VGND sg13g2_decap_8
XFILLER_47_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1185_ net74 VGND VPWR u_ppwm_u_mem__1185_/D hold32/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_967 VPWR VGND sg13g2_decap_8
XFILLER_22_628 VPWR VGND sg13g2_decap_8
XFILLER_21_138 VPWR VGND sg13g2_fill_2
XFILLER_30_650 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0969_ VGND VPWR net367 u_ppwm_u_mem__0670_/Y u_ppwm_u_mem__1161_/D
+ u_ppwm_u_mem__0968_/Y sg13g2_a21oi_1
XFILLER_26_923 VPWR VGND sg13g2_decap_8
XFILLER_37_260 VPWR VGND sg13g2_decap_8
XFILLER_37_282 VPWR VGND sg13g2_fill_2
XFILLER_41_948 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__807__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_25_499 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__822__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_21_661 VPWR VGND sg13g2_decap_8
XFILLER_0_554 VPWR VGND sg13g2_decap_8
XFILLER_48_536 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__242__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_17_956 VPWR VGND sg13g2_decap_8
XFILLER_29_794 VPWR VGND sg13g2_decap_8
XFILLER_44_753 VPWR VGND sg13g2_decap_8
XFILLER_43_230 VPWR VGND sg13g2_decap_8
XFILLER_16_455 VPWR VGND sg13g2_decap_8
XFILLER_32_948 VPWR VGND sg13g2_decap_8
XFILLER_8_665 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0823_ hold19/A hold83/A net416 u_ppwm_u_mem__0823_/X VPWR VGND sg13g2_mux2_1
Xhold109 hold109/A VPWR VGND net306 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0754_ u_ppwm_u_mem__0754_/Y net335 u_ppwm_u_mem__0754_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_4_860 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0685_ VPWR u_ppwm_u_mem__0685_/Y net545 VGND sg13g2_inv_1
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
XFILLER_39_569 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__723_ VGND VPWR u_ppwm_u_ex__724_/B net323 hold328/A sg13g2_or2_1
XFILLER_47_591 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1168_ net142 VGND VPWR u_ppwm_u_mem__1168_/D hold90/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__654_ VGND VPWR u_ppwm_u_ex__659_/B u_ppwm_u_ex__653_/X u_ppwm_u_ex__654_/Y
+ net315 sg13g2_a21oi_1
XFILLER_35_764 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__585_ u_ppwm_u_ex__585_/Y hold271/A net388 VPWR VGND sg13g2_nand2b_1
XFILLER_22_425 VPWR VGND sg13g2_decap_8
XFILLER_34_263 VPWR VGND sg13g2_fill_2
XFILLER_34_274 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1099_ u_ppwm_u_mem__1101_/B net602 net624 u_ppwm_u_mem__1102_/D VPWR
+ VGND sg13g2_and3_1
XFILLER_23_959 VPWR VGND sg13g2_decap_8
XFILLER_31_970 VPWR VGND sg13g2_decap_8
XFILLER_18_709 VPWR VGND sg13g2_decap_8
XFILLER_45_528 VPWR VGND sg13g2_decap_8
XFILLER_26_720 VPWR VGND sg13g2_decap_8
XFILLER_14_926 VPWR VGND sg13g2_decap_8
XFILLER_26_797 VPWR VGND sg13g2_decap_8
XFILLER_41_745 VPWR VGND sg13g2_decap_8
XFILLER_13_469 VPWR VGND sg13g2_decap_8
XFILLER_40_277 VPWR VGND sg13g2_fill_1
XFILLER_22_992 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_decap_8
XFILLER_4_27 VPWR VGND sg13g2_fill_1
XFILLER_1_841 VPWR VGND sg13g2_decap_8
XFILLER_49_812 VPWR VGND sg13g2_decap_8
XFILLER_0_351 VPWR VGND sg13g2_decap_8
XFILLER_48_333 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_fill_2
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_1_1023 VPWR VGND sg13g2_decap_4
XFILLER_29_591 VPWR VGND sg13g2_decap_8
XFILLER_44_550 VPWR VGND sg13g2_decap_8
XFILLER_17_753 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1022_ net430 VPWR u_ppwm_u_mem__1022_/Y VGND net347 hold42/A sg13g2_o21ai_1
XFILLER_32_745 VPWR VGND sg13g2_decap_8
XFILLER_9_941 VPWR VGND sg13g2_decap_8
XFILLER_8_462 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0806_ u_ppwm_u_mem__0805_/Y VPWR u_ppwm_u_mem__0806_/Y VGND net407
+ u_ppwm_u_mem__0803_/X sg13g2_o21ai_1
Xu_ppwm_u_mem__0737_ net602 u_ppwm_u_mem__0737_/B u_ppwm_u_mem__0737_/C u_ppwm_u_mem__0737_/D
+ u_ppwm_u_mem__0737_/Y VPWR VGND sg13g2_nor4_1
Xu_ppwm_u_mem__0668_ VPWR u_ppwm_u_mem__0668_/Y net214 VGND sg13g2_inv_1
Xfanout408 net409 net408 VPWR VGND sg13g2_buf_8
Xfanout419 net420 net419 VPWR VGND sg13g2_buf_1
Xu_ppwm_u_mem__1139__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_39_366 VPWR VGND sg13g2_fill_2
XFILLER_39_377 VPWR VGND sg13g2_fill_2
XFILLER_27_539 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__706_ VGND VPWR u_ppwm_u_ex__703_/Y u_ppwm_u_ex__704_/Y u_ppwm_u_ex__815_/D
+ u_ppwm_u_ex__705_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__637_ u_ppwm_u_ex__637_/A u_ppwm_u_ex__637_/B net317 fanout312/A VPWR
+ VGND sg13g2_nor3_2
XFILLER_35_561 VPWR VGND sg13g2_decap_8
XFILLER_23_756 VPWR VGND sg13g2_decap_8
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_11_918 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__568_ u_ppwm_u_ex__567_/Y VPWR u_ppwm_u_ex__568_/Y VGND hold333/A u_ppwm_u_ex__435_/Y
+ sg13g2_o21ai_1
XFILLER_22_255 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__499_ u_ppwm_u_ex__499_/Y net385 hold266/A VPWR VGND sg13g2_nand2b_1
XFILLER_13_25 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1224__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_49_119 VPWR VGND sg13g2_decap_8
XFILLER_38_33 VPWR VGND sg13g2_fill_2
XFILLER_46_826 VPWR VGND sg13g2_decap_8
XFILLER_18_506 VPWR VGND sg13g2_decap_8
XFILLER_14_723 VPWR VGND sg13g2_decap_8
XFILLER_41_542 VPWR VGND sg13g2_decap_8
XFILLER_26_594 VPWR VGND sg13g2_decap_8
XFILLER_13_288 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_pwm__192_ hold283/A net337 net580 u_ppwm_u_pwm__193_/C VPWR VGND hold268/A
+ sg13g2_nand4_1
XFILLER_6_944 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_5_465 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1175__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_37_848 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_45_892 VPWR VGND sg13g2_decap_8
XFILLER_17_550 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1005_ VGND VPWR net350 u_ppwm_u_mem__0652_/Y u_ppwm_u_mem__1179_/D
+ u_ppwm_u_mem__1004_/Y sg13g2_a21oi_1
XFILLER_32_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__422_ VPWR u_ppwm_u_ex__541_/B net386 VGND sg13g2_inv_1
XFILLER_20_748 VPWR VGND sg13g2_decap_8
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_314 VPWR VGND sg13g2_decap_8
XFILLER_28_837 VPWR VGND sg13g2_decap_8
XFILLER_39_174 VPWR VGND sg13g2_fill_1
XFILLER_36_881 VPWR VGND sg13g2_decap_8
XFILLER_24_13 VPWR VGND sg13g2_fill_1
XFILLER_11_715 VPWR VGND sg13g2_decap_8
XFILLER_23_553 VPWR VGND sg13g2_decap_8
XFILLER_10_247 VPWR VGND sg13g2_fill_2
XFILLER_3_936 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1198__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_49_21 VPWR VGND sg13g2_decap_8
Xhold270 hold270/A VPWR VGND net613 sg13g2_dlygate4sd3_1
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_2_457 VPWR VGND sg13g2_decap_8
Xhold281 hold281/A VPWR VGND net624 sg13g2_dlygate4sd3_1
Xhold292 hold292/A VPWR VGND net635 sg13g2_dlygate4sd3_1
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_46_623 VPWR VGND sg13g2_decap_8
XFILLER_19_859 VPWR VGND sg13g2_decap_8
XFILLER_33_306 VPWR VGND sg13g2_decap_4
XFILLER_14_520 VPWR VGND sg13g2_decap_8
XFILLER_33_339 VPWR VGND sg13g2_decap_4
XFILLER_42_895 VPWR VGND sg13g2_decap_8
XFILLER_14_597 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__244_ net180 VGND VPWR net605 hold261/A clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_6_741 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__175_ u_ppwm_u_pwm__175_/A net622 u_ppwm_u_pwm__175_/C hold280/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_49_483 VPWR VGND sg13g2_decap_8
XFILLER_25_807 VPWR VGND sg13g2_decap_8
XFILLER_37_645 VPWR VGND sg13g2_decap_8
XFILLER_18_870 VPWR VGND sg13g2_decap_8
XFILLER_33_862 VPWR VGND sg13g2_decap_8
XFILLER_20_545 VPWR VGND sg13g2_decap_8
XFILLER_0_939 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1158__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_28_634 VPWR VGND sg13g2_decap_8
XFILLER_11_512 VPWR VGND sg13g2_decap_8
XFILLER_24_895 VPWR VGND sg13g2_decap_8
XFILLER_13_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_538 VPWR VGND sg13g2_decap_8
XFILLER_11_589 VPWR VGND sg13g2_decap_8
XFILLER_3_733 VPWR VGND sg13g2_decap_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_19_656 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
XFILLER_15_851 VPWR VGND sg13g2_decap_8
XFILLER_33_158 VPWR VGND sg13g2_fill_1
XFILLER_42_692 VPWR VGND sg13g2_decap_8
XFILLER_30_832 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0985_ VGND VPWR net351 u_ppwm_u_mem__0662_/Y hold145/A u_ppwm_u_mem__0984_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__227_ net187 VGND VPWR net219 hold21/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__158_ VGND VPWR u_ppwm_u_pwm__131_/Y net328 hold53/A u_ppwm_u_pwm__157_/Y
+ sg13g2_a21oi_1
XFILLER_38_921 VPWR VGND sg13g2_decap_8
XFILLER_49_280 VPWR VGND sg13g2_decap_8
XFILLER_25_604 VPWR VGND sg13g2_decap_8
XFILLER_38_998 VPWR VGND sg13g2_decap_8
XFILLER_40_618 VPWR VGND sg13g2_decap_8
XFILLER_21_843 VPWR VGND sg13g2_decap_8
XFILLER_32_191 VPWR VGND sg13g2_fill_1
XFILLER_21_25 VPWR VGND sg13g2_fill_2
XFILLER_0_736 VPWR VGND sg13g2_decap_8
XFILLER_48_718 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_29_976 VPWR VGND sg13g2_decap_8
XFILLER_44_935 VPWR VGND sg13g2_decap_8
XFILLER_16_637 VPWR VGND sg13g2_decap_8
XFILLER_15_169 VPWR VGND sg13g2_decap_8
XFILLER_12_810 VPWR VGND sg13g2_decap_8
XFILLER_23_180 VPWR VGND sg13g2_fill_2
XFILLER_24_692 VPWR VGND sg13g2_decap_8
XFILLER_8_847 VPWR VGND sg13g2_decap_8
XFILLER_12_887 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0770_ u_ppwm_u_mem__0769_/Y VPWR u_ppwm_u_mem__0770_/Y VGND u_ppwm_u_mem__0710_/Y
+ net417 sg13g2_o21ai_1
XFILLER_3_530 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_38_228 VPWR VGND sg13g2_decap_4
XFILLER_4_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__670_ u_ppwm_u_ex__696_/B net391 net318 VPWR VGND sg13g2_xnor2_1
XFILLER_19_453 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1184_ net78 VGND VPWR net230 hold182/A clknet_5_24__leaf_clk sg13g2_dfrbpq_2
XFILLER_35_946 VPWR VGND sg13g2_decap_8
XFILLER_22_607 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0968_ net444 VPWR u_ppwm_u_mem__0968_/Y VGND net367 net256 sg13g2_o21ai_1
Xu_ppwm_u_mem__0899_ VGND VPWR net358 u_ppwm_u_mem__0705_/Y u_ppwm_u_mem__1126_/D
+ u_ppwm_u_mem__0898_/Y sg13g2_a21oi_1
XFILLER_29_217 VPWR VGND sg13g2_decap_8
XFILLER_29_239 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1116__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_26_902 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_fill_2
XFILLER_38_795 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__799_ VPWR VGND fanout316/A u_ppwm_u_ex__714_/Y u_ppwm_u_ex__798_/Y net646
+ u_ppwm_u_ex__801_/A net312 sg13g2_a221oi_1
XFILLER_26_979 VPWR VGND sg13g2_decap_8
XFILLER_41_927 VPWR VGND sg13g2_decap_8
XFILLER_25_478 VPWR VGND sg13g2_decap_8
XFILLER_21_640 VPWR VGND sg13g2_decap_8
XFILLER_20_183 VPWR VGND sg13g2_decap_4
XFILLER_4_349 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_533 VPWR VGND sg13g2_decap_8
XFILLER_48_515 VPWR VGND sg13g2_decap_8
XFILLER_29_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1190__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_44_732 VPWR VGND sg13g2_decap_8
XFILLER_17_935 VPWR VGND sg13g2_decap_8
XFILLER_16_434 VPWR VGND sg13g2_decap_8
XFILLER_43_253 VPWR VGND sg13g2_fill_1
XFILLER_32_927 VPWR VGND sg13g2_decap_8
XFILLER_40_982 VPWR VGND sg13g2_decap_8
XFILLER_8_644 VPWR VGND sg13g2_decap_8
XFILLER_7_121 VPWR VGND sg13g2_fill_1
XFILLER_12_684 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0822_ VGND VPWR u_ppwm_u_mem__0672_/Y net416 u_ppwm_u_mem__0822_/Y
+ u_ppwm_u_mem__0821_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0753_ hold38/A hold92/A net415 u_ppwm_u_mem__0754_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0684_ VPWR u_ppwm_u_mem__0684_/Y net541 VGND sg13g2_inv_1
XFILLER_26_1000 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_548 VPWR VGND sg13g2_decap_8
XFILLER_19_250 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__722_ net385 net323 u_ppwm_u_ex__722_/X VPWR VGND sg13g2_and2_1
XFILLER_47_570 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1167_ net146 VGND VPWR net288 hold150/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__653_ net320 net396 u_ppwm_u_ex__646_/A u_ppwm_u_ex__653_/X VPWR VGND
+ sg13g2_a21o_1
XFILLER_34_242 VPWR VGND sg13g2_decap_4
XFILLER_35_743 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__584_ VPWR VGND u_ppwm_u_ex__582_/Y u_ppwm_u_ex__583_/Y u_ppwm_u_ex__574_/Y
+ net390 u_ppwm_u_ex__584_/Y u_ppwm_u_ex__506_/B sg13g2_a221oi_1
Xu_ppwm_u_mem__1098_ net602 u_ppwm_u_mem__1098_/B u_ppwm_u_mem__1100_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_23_938 VPWR VGND sg13g2_decap_8
XFILLER_45_507 VPWR VGND sg13g2_decap_8
XFILLER_38_592 VPWR VGND sg13g2_decap_8
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_25_242 VPWR VGND sg13g2_fill_2
XFILLER_41_724 VPWR VGND sg13g2_decap_8
XFILLER_26_776 VPWR VGND sg13g2_decap_8
XFILLER_13_448 VPWR VGND sg13g2_decap_8
XFILLER_43_78 VPWR VGND sg13g2_decap_4
XFILLER_22_971 VPWR VGND sg13g2_decap_8
XFILLER_5_647 VPWR VGND sg13g2_decap_8
XFILLER_49_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_820 VPWR VGND sg13g2_decap_8
XFILLER_0_330 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_897 VPWR VGND sg13g2_decap_8
XFILLER_49_868 VPWR VGND sg13g2_decap_8
XFILLER_48_389 VPWR VGND sg13g2_decap_8
XFILLER_1_1002 VPWR VGND sg13g2_decap_8
XFILLER_17_732 VPWR VGND sg13g2_decap_8
XFILLER_29_570 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1021_ VGND VPWR net347 u_ppwm_u_mem__0644_/Y hold43/A u_ppwm_u_mem__1020_/Y
+ sg13g2_a21oi_1
XFILLER_32_724 VPWR VGND sg13g2_decap_8
XFILLER_9_920 VPWR VGND sg13g2_decap_8
XFILLER_12_481 VPWR VGND sg13g2_decap_8
XFILLER_8_441 VPWR VGND sg13g2_decap_8
XFILLER_9_997 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0805_ VGND VPWR net409 u_ppwm_u_mem__0804_/X u_ppwm_u_mem__0805_/Y
+ net332 sg13g2_a21oi_1
Xu_ppwm_u_mem__0736_ u_ppwm_u_mem__0737_/D net338 net423 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0667_ VPWR u_ppwm_u_mem__0667_/Y net224 VGND sg13g2_inv_1
Xfanout409 fanout409/A net409 VPWR VGND sg13g2_buf_8
XFILLER_27_518 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__705_ net426 VPWR u_ppwm_u_ex__705_/Y VGND net386 net310 sg13g2_o21ai_1
Xu_ppwm_u_mem__1219_ net147 VGND VPWR u_ppwm_u_mem__1219_/D hold275/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_540 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__636_ u_ppwm_u_ex__636_/B u_ppwm_u_ex__636_/A u_ppwm_u_ex__636_/X VPWR
+ VGND sg13g2_xor2_1
XFILLER_23_735 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__567_ u_ppwm_u_ex__563_/Y VPWR u_ppwm_u_ex__567_/Y VGND u_ppwm_u_ex__562_/Y
+ u_ppwm_u_ex__566_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__498_ u_ppwm_u_ex__497_/Y VPWR u_ppwm_u_ex__498_/Y VGND u_ppwm_u_ex__420_/Y
+ hold212/A sg13g2_o21ai_1
XFILLER_2_639 VPWR VGND sg13g2_decap_8
XFILLER_1_149 VPWR VGND sg13g2_fill_1
XFILLER_46_805 VPWR VGND sg13g2_decap_8
XFILLER_14_702 VPWR VGND sg13g2_decap_8
XFILLER_26_573 VPWR VGND sg13g2_decap_8
XFILLER_41_521 VPWR VGND sg13g2_decap_8
XFILLER_13_234 VPWR VGND sg13g2_fill_2
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_41_598 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__191_ hold261/A hold300/A net594 hold252/A VPWR VGND hold278/A sg13g2_nand4_1
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_6_923 VPWR VGND sg13g2_decap_8
XFILLER_5_444 VPWR VGND sg13g2_decap_8
XFILLER_1_694 VPWR VGND sg13g2_decap_8
XFILLER_49_665 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_37_827 VPWR VGND sg13g2_decap_8
XFILLER_36_348 VPWR VGND sg13g2_fill_2
XFILLER_45_871 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1004_ net431 VPWR u_ppwm_u_mem__1004_/Y VGND net350 net278 sg13g2_o21ai_1
Xu_ppwm_u_ex__421_ VPWR u_ppwm_u_ex__538_/B hold308/A VGND sg13g2_inv_1
XFILLER_20_727 VPWR VGND sg13g2_decap_8
XFILLER_32_598 VPWR VGND sg13g2_decap_8
XFILLER_30_1007 VPWR VGND sg13g2_decap_8
XFILLER_9_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0719_ VPWR u_ppwm_u_mem__0719_/Y net600 VGND sg13g2_inv_1
XFILLER_8_1008 VPWR VGND sg13g2_decap_8
XFILLER_28_816 VPWR VGND sg13g2_decap_8
XFILLER_39_186 VPWR VGND sg13g2_fill_2
XFILLER_36_860 VPWR VGND sg13g2_decap_8
XFILLER_39_1010 VPWR VGND sg13g2_decap_8
XFILLER_23_532 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__619_ VGND VPWR u_ppwm_u_ex__547_/Y u_ppwm_u_ex__617_/X hold286/A net628
+ sg13g2_a21oi_1
XFILLER_24_25 VPWR VGND sg13g2_decap_4
XFILLER_10_259 VPWR VGND sg13g2_fill_1
XFILLER_6_208 VPWR VGND sg13g2_fill_2
XFILLER_40_24 VPWR VGND sg13g2_decap_4
XFILLER_3_915 VPWR VGND sg13g2_decap_8
XFILLER_2_436 VPWR VGND sg13g2_decap_8
Xhold271 hold271/A VPWR VGND net614 sg13g2_dlygate4sd3_1
Xhold260 hold260/A VPWR VGND net603 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1205__80 VPWR VGND net80 sg13g2_tiehi
Xhold282 hold282/A VPWR VGND net625 sg13g2_dlygate4sd3_1
Xhold293 hold293/A VPWR VGND net636 sg13g2_dlygate4sd3_1
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_18_304 VPWR VGND sg13g2_fill_2
XFILLER_19_838 VPWR VGND sg13g2_decap_8
XFILLER_46_679 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_42_874 VPWR VGND sg13g2_decap_8
XFILLER_41_384 VPWR VGND sg13g2_fill_1
XFILLER_41_373 VPWR VGND sg13g2_fill_1
XFILLER_14_576 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__243_ net188 VGND VPWR net581 hold237/A clknet_5_1__leaf_clk sg13g2_dfrbpq_2
XFILLER_6_720 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__174_ u_ppwm_u_pwm__175_/C net621 net337 u_ppwm_u_pwm__176_/D VPWR VGND
+ sg13g2_and3_1
XFILLER_6_797 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_fill_1
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1222__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_1_491 VPWR VGND sg13g2_decap_8
XFILLER_49_462 VPWR VGND sg13g2_decap_8
XFILLER_36_101 VPWR VGND sg13g2_decap_8
XFILLER_37_624 VPWR VGND sg13g2_decap_8
XFILLER_24_329 VPWR VGND sg13g2_fill_1
XFILLER_33_841 VPWR VGND sg13g2_decap_8
XFILLER_20_524 VPWR VGND sg13g2_decap_8
XFILLER_9_591 VPWR VGND sg13g2_decap_8
XFILLER_0_918 VPWR VGND sg13g2_decap_8
XFILLER_28_613 VPWR VGND sg13g2_decap_8
XFILLER_16_819 VPWR VGND sg13g2_decap_8
XFILLER_43_649 VPWR VGND sg13g2_decap_8
XFILLER_15_318 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_fill_1
XFILLER_24_874 VPWR VGND sg13g2_decap_8
XFILLER_7_517 VPWR VGND sg13g2_decap_8
XFILLER_11_568 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1126__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_3_712 VPWR VGND sg13g2_decap_8
XFILLER_3_789 VPWR VGND sg13g2_decap_8
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_18_134 VPWR VGND sg13g2_fill_2
XFILLER_19_635 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_15_830 VPWR VGND sg13g2_decap_8
XFILLER_18_189 VPWR VGND sg13g2_decap_8
XFILLER_34_649 VPWR VGND sg13g2_decap_8
XFILLER_42_671 VPWR VGND sg13g2_decap_8
XFILLER_30_811 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0984_ net431 VPWR u_ppwm_u_mem__0984_/Y VGND net350 hold274/A sg13g2_o21ai_1
XFILLER_30_888 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__226_ net190 VGND VPWR net201 hold3/A clknet_5_2__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__157_ net424 VPWR u_ppwm_u_pwm__157_/Y VGND net387 net328 sg13g2_o21ai_1
XFILLER_6_594 VPWR VGND sg13g2_decap_8
XFILLER_38_900 VPWR VGND sg13g2_decap_8
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_21_822 VPWR VGND sg13g2_decap_8
XFILLER_21_899 VPWR VGND sg13g2_decap_8
XFILLER_20_376 VPWR VGND sg13g2_fill_2
XFILLER_20_387 VPWR VGND sg13g2_fill_2
XFILLER_20_398 VPWR VGND sg13g2_fill_1
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_715 VPWR VGND sg13g2_decap_8
XFILLER_29_955 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_44_914 VPWR VGND sg13g2_decap_8
XFILLER_16_616 VPWR VGND sg13g2_decap_8
XFILLER_28_476 VPWR VGND sg13g2_decap_4
XFILLER_24_671 VPWR VGND sg13g2_decap_8
XFILLER_11_332 VPWR VGND sg13g2_fill_1
XFILLER_8_826 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_4
XFILLER_12_866 VPWR VGND sg13g2_decap_8
XFILLER_3_586 VPWR VGND sg13g2_decap_8
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
XFILLER_19_432 VPWR VGND sg13g2_decap_8
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_46_240 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1183_ net82 VGND VPWR net526 hold201/A clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_424 VPWR VGND sg13g2_decap_4
XFILLER_35_925 VPWR VGND sg13g2_decap_8
XFILLER_30_685 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0967_ VGND VPWR net367 u_ppwm_u_mem__0671_/Y hold60/A u_ppwm_u_mem__0966_/Y
+ sg13g2_a21oi_1
XFILLER_7_881 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__209_ hold300/A u_ppwm_u_pwm__209_/B u_ppwm_u_pwm__215_/A VPWR VGND
+ sg13g2_nor2_1
Xu_ppwm_u_mem__0898_ net443 VPWR u_ppwm_u_mem__0898_/Y VGND net358 net503 sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_6_391 VPWR VGND sg13g2_decap_8
XFILLER_38_774 VPWR VGND sg13g2_decap_8
XFILLER_25_424 VPWR VGND sg13g2_decap_8
XFILLER_26_958 VPWR VGND sg13g2_decap_8
XFILLER_41_906 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__089_ net556 u_ppwm_u_global_counter__088_/Y hold214/A VPWR
+ VGND sg13g2_nor2b_1
Xu_ppwm_u_ex__798_ u_ppwm_u_ex__798_/Y u_ppwm_u_ex__798_/A u_ppwm_u_ex__798_/B VPWR
+ VGND sg13g2_xnor2_1
XFILLER_25_457 VPWR VGND sg13g2_decap_8
XFILLER_32_14 VPWR VGND sg13g2_decap_8
XFILLER_20_151 VPWR VGND sg13g2_fill_1
XFILLER_21_696 VPWR VGND sg13g2_decap_8
XFILLER_32_69 VPWR VGND sg13g2_decap_4
XFILLER_5_829 VPWR VGND sg13g2_decap_8
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_512 VPWR VGND sg13g2_decap_8
XFILLER_0_589 VPWR VGND sg13g2_decap_8
XFILLER_17_914 VPWR VGND sg13g2_decap_8
XFILLER_29_752 VPWR VGND sg13g2_decap_8
XFILLER_44_711 VPWR VGND sg13g2_decap_8
XFILLER_16_413 VPWR VGND sg13g2_decap_8
XFILLER_32_906 VPWR VGND sg13g2_decap_8
XFILLER_44_788 VPWR VGND sg13g2_decap_8
XFILLER_31_449 VPWR VGND sg13g2_fill_1
XFILLER_40_961 VPWR VGND sg13g2_decap_8
XFILLER_12_663 VPWR VGND sg13g2_decap_8
XFILLER_8_623 VPWR VGND sg13g2_decap_8
XFILLER_7_144 VPWR VGND sg13g2_fill_1
XFILLER_7_133 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0821_ net408 VPWR u_ppwm_u_mem__0821_/Y VGND hold114/A net415 sg13g2_o21ai_1
Xu_ppwm_u_mem__0752_ hold196/A hold172/A net416 u_ppwm_u_mem__0752_/X VPWR VGND sg13g2_mux2_1
XFILLER_22_80 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1178__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_4_895 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0683_ VPWR u_ppwm_u_mem__0683_/Y net539 VGND sg13g2_inv_1
XFILLER_3_383 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_39_527 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__721_ VGND VPWR u_ppwm_u_ex__718_/Y u_ppwm_u_ex__719_/Y hold292/A u_ppwm_u_ex__720_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__652_ net319 net394 u_ppwm_u_ex__659_/B VPWR VGND sg13g2_xor2_1
XFILLER_35_722 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1166_ net148 VGND VPWR u_ppwm_u_mem__1166_/D hold56/A clknet_5_11__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__583_ u_ppwm_u_ex__583_/A hold234/A u_ppwm_u_ex__583_/Y VPWR VGND sg13g2_nor2_1
XFILLER_16_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1097_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1097_/B u_ppwm_u_mem__1098_/B
+ u_ppwm_u_mem__1222_/D VPWR VGND sg13g2_nor3_1
XFILLER_23_917 VPWR VGND sg13g2_decap_8
XFILLER_34_265 VPWR VGND sg13g2_fill_1
XFILLER_35_799 VPWR VGND sg13g2_decap_8
XFILLER_34_298 VPWR VGND sg13g2_fill_2
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_309 VPWR VGND sg13g2_decap_8
XFILLER_38_571 VPWR VGND sg13g2_decap_8
XFILLER_26_755 VPWR VGND sg13g2_decap_8
XFILLER_41_703 VPWR VGND sg13g2_decap_8
XFILLER_13_427 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_40_235 VPWR VGND sg13g2_decap_8
XFILLER_9_409 VPWR VGND sg13g2_decap_8
XFILLER_22_950 VPWR VGND sg13g2_decap_8
XFILLER_21_493 VPWR VGND sg13g2_decap_8
XFILLER_5_626 VPWR VGND sg13g2_decap_8
XFILLER_49_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_876 VPWR VGND sg13g2_decap_8
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_8
XFILLER_48_368 VPWR VGND sg13g2_decap_8
XFILLER_17_711 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1020_ net432 VPWR u_ppwm_u_mem__1020_/Y VGND net347 hold165/A sg13g2_o21ai_1
XFILLER_17_788 VPWR VGND sg13g2_decap_8
XFILLER_32_703 VPWR VGND sg13g2_decap_8
XFILLER_44_585 VPWR VGND sg13g2_decap_8
XFILLER_20_909 VPWR VGND sg13g2_decap_8
XFILLER_8_420 VPWR VGND sg13g2_decap_8
XFILLER_12_460 VPWR VGND sg13g2_decap_8
XFILLER_13_994 VPWR VGND sg13g2_decap_8
XFILLER_31_279 VPWR VGND sg13g2_fill_2
XFILLER_9_976 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0804_ hold100/A hold109/A net418 u_ppwm_u_mem__0804_/X VPWR VGND sg13g2_mux2_1
XFILLER_8_497 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0735_ net602 u_ppwm_u_mem__0737_/B u_ppwm_u_mem__0737_/C hold260/A
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__0666_ VPWR u_ppwm_u_mem__0666_/Y net253 VGND sg13g2_inv_1
XFILLER_4_692 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__704_ VPWR VGND net387 net309 net311 net651 u_ppwm_u_ex__704_/Y net313
+ sg13g2_a221oi_1
Xu_ppwm_u_mem__1218_ net163 VGND VPWR u_ppwm_u_mem__1218_/D hold9/A clknet_5_9__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1149_ net63 VGND VPWR net520 hold196/A clknet_5_31__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__635_ net323 net398 u_ppwm_u_ex__636_/B VPWR VGND sg13g2_xor2_1
XFILLER_23_714 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__566_ net388 u_ppwm_u_ex__566_/B u_ppwm_u_ex__566_/Y VPWR VGND sg13g2_nor2_1
XFILLER_35_596 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__497_ u_ppwm_u_ex__497_/Y net383 hold272/A VPWR VGND sg13g2_nand2b_1
XFILLER_2_618 VPWR VGND sg13g2_decap_8
XFILLER_39_891 VPWR VGND sg13g2_decap_8
XFILLER_26_552 VPWR VGND sg13g2_decap_8
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_41_577 VPWR VGND sg13g2_decap_8
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__190_ hold287/A net422 net535 u_ppwm_u_pwm__193_/A VPWR VGND sg13g2_nand3_1
XFILLER_6_902 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_5_423 VPWR VGND sg13g2_decap_8
XFILLER_1_673 VPWR VGND sg13g2_decap_8
XFILLER_49_644 VPWR VGND sg13g2_decap_8
XFILLER_0_194 VPWR VGND sg13g2_decap_8
XFILLER_23_1015 VPWR VGND sg13g2_decap_8
XFILLER_37_806 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_36_305 VPWR VGND sg13g2_decap_8
XFILLER_45_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1003_ VGND VPWR net356 u_ppwm_u_mem__0653_/Y hold82/A u_ppwm_u_mem__1002_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__420_ u_ppwm_u_ex__420_/Y net384 VPWR VGND sg13g2_inv_2
XFILLER_17_585 VPWR VGND sg13g2_decap_8
XFILLER_20_706 VPWR VGND sg13g2_decap_8
XFILLER_32_577 VPWR VGND sg13g2_decap_8
XFILLER_13_791 VPWR VGND sg13g2_decap_8
XFILLER_9_773 VPWR VGND sg13g2_decap_8
XFILLER_8_283 VPWR VGND sg13g2_fill_2
XFILLER_5_990 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0718_ VPWR u_ppwm_u_mem__0718_/Y net481 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0649_ VPWR u_ppwm_u_mem__0649_/Y net544 VGND sg13g2_inv_1
XFILLER_39_165 VPWR VGND sg13g2_decap_8
XFILLER_27_349 VPWR VGND sg13g2_decap_8
XFILLER_23_511 VPWR VGND sg13g2_decap_8
XFILLER_35_382 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__618_ net439 VPWR hold285/A VGND net627 u_ppwm_u_ex__617_/A sg13g2_o21ai_1
Xu_ppwm_u_ex__549_ u_ppwm_u_ex__549_/Y hold311/A net398 VPWR VGND sg13g2_nand2b_1
XFILLER_10_216 VPWR VGND sg13g2_decap_8
XFILLER_23_588 VPWR VGND sg13g2_decap_8
XFILLER_10_249 VPWR VGND sg13g2_fill_1
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
Xhold261 hold261/A VPWR VGND net604 sg13g2_dlygate4sd3_1
XFILLER_2_415 VPWR VGND sg13g2_decap_8
Xhold250 hold250/A VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold272 hold272/A VPWR VGND net615 sg13g2_dlygate4sd3_1
Xhold283 hold283/A VPWR VGND net626 sg13g2_dlygate4sd3_1
Xhold294 hold294/A VPWR VGND net637 sg13g2_dlygate4sd3_1
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_19_817 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_45_179 VPWR VGND sg13g2_decap_4
XFILLER_26_360 VPWR VGND sg13g2_fill_1
XFILLER_42_853 VPWR VGND sg13g2_decap_8
XFILLER_14_555 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__242_ net192 VGND VPWR u_ppwm_u_pwm__242_/D hold283/A clknet_5_1__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__173_ VGND VPWR net337 u_ppwm_u_pwm__176_/D hold279/A net621 sg13g2_a21oi_1
XFILLER_6_776 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_2_982 VPWR VGND sg13g2_decap_8
XFILLER_1_470 VPWR VGND sg13g2_decap_8
XFILLER_49_441 VPWR VGND sg13g2_decap_8
XFILLER_37_603 VPWR VGND sg13g2_decap_8
XFILLER_33_820 VPWR VGND sg13g2_decap_8
XFILLER_20_503 VPWR VGND sg13g2_decap_8
XFILLER_33_897 VPWR VGND sg13g2_decap_8
XFILLER_32_396 VPWR VGND sg13g2_fill_2
XFILLER_9_570 VPWR VGND sg13g2_decap_8
XFILLER_28_669 VPWR VGND sg13g2_decap_8
XFILLER_43_628 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_fill_2
XFILLER_24_853 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_547 VPWR VGND sg13g2_decap_8
XFILLER_3_768 VPWR VGND sg13g2_decap_8
XFILLER_19_614 VPWR VGND sg13g2_decap_8
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_20_1007 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_34_628 VPWR VGND sg13g2_decap_8
XFILLER_42_650 VPWR VGND sg13g2_decap_8
XFILLER_14_352 VPWR VGND sg13g2_decap_4
XFILLER_15_886 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0983_ VGND VPWR net348 u_ppwm_u_mem__0663_/Y u_ppwm_u_mem__1168_/D
+ u_ppwm_u_mem__0982_/Y sg13g2_a21oi_1
XFILLER_30_867 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__225_ net422 u_ppwm_u_pwm__225_/B u_ppwm_u_pwm__247_/D VPWR VGND sg13g2_and2_1
Xu_ppwm_u_pwm__156_ VGND VPWR u_ppwm_u_pwm__132_/Y net330 hold24/A u_ppwm_u_pwm__155_/Y
+ sg13g2_a21oi_1
XFILLER_6_573 VPWR VGND sg13g2_decap_8
XFILLER_37_411 VPWR VGND sg13g2_decap_8
XFILLER_38_956 VPWR VGND sg13g2_decap_8
XFILLER_25_639 VPWR VGND sg13g2_decap_8
XFILLER_21_801 VPWR VGND sg13g2_decap_8
XFILLER_36_1014 VPWR VGND sg13g2_decap_8
XFILLER_20_300 VPWR VGND sg13g2_decap_4
XFILLER_32_182 VPWR VGND sg13g2_decap_8
XFILLER_33_694 VPWR VGND sg13g2_decap_8
XFILLER_21_878 VPWR VGND sg13g2_decap_8
XFILLER_21_49 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1171__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_29_934 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_15_127 VPWR VGND sg13g2_decap_4
XFILLER_24_650 VPWR VGND sg13g2_decap_8
XFILLER_8_805 VPWR VGND sg13g2_decap_8
XFILLER_11_322 VPWR VGND sg13g2_fill_2
XFILLER_12_845 VPWR VGND sg13g2_decap_8
XFILLER_23_182 VPWR VGND sg13g2_fill_1
XFILLER_3_565 VPWR VGND sg13g2_decap_8
XFILLER_39_709 VPWR VGND sg13g2_decap_8
XFILLER_47_731 VPWR VGND sg13g2_decap_8
Xfanout390 hold325/A net390 VPWR VGND sg13g2_buf_2
XFILLER_35_904 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1182_ net86 VGND VPWR u_ppwm_u_mem__1182_/D hold181/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_19_488 VPWR VGND sg13g2_decap_8
XFILLER_43_992 VPWR VGND sg13g2_decap_8
XFILLER_14_171 VPWR VGND sg13g2_decap_8
XFILLER_15_683 VPWR VGND sg13g2_decap_8
XFILLER_30_664 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0966_ net446 VPWR u_ppwm_u_mem__0966_/Y VGND net369 hold233/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__208_ u_ppwm_u_pwm__210_/D hold23/A hold283/A VPWR VGND sg13g2_nand2b_1
XFILLER_7_860 VPWR VGND sg13g2_decap_8
XFILLER_6_370 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0897_ VGND VPWR net372 u_ppwm_u_mem__0706_/Y hold161/A u_ppwm_u_mem__0896_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__139_ VPWR u_ppwm_u_pwm__175_/A net422 VGND sg13g2_inv_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_37_241 VPWR VGND sg13g2_decap_8
XFILLER_38_753 VPWR VGND sg13g2_decap_8
XFILLER_26_937 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__088_ hold318/A net331 net555 u_ppwm_u_global_counter__088_/Y
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__797_ u_ppwm_u_ex__798_/B net378 net322 VPWR VGND sg13g2_xnor2_1
XFILLER_13_609 VPWR VGND sg13g2_decap_8
XFILLER_34_992 VPWR VGND sg13g2_decap_8
XFILLER_21_675 VPWR VGND sg13g2_decap_8
XFILLER_5_808 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_568 VPWR VGND sg13g2_decap_8
XFILLER_29_731 VPWR VGND sg13g2_decap_8
XFILLER_28_230 VPWR VGND sg13g2_decap_4
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_16_469 VPWR VGND sg13g2_decap_8
XFILLER_19_1020 VPWR VGND sg13g2_decap_8
XFILLER_31_406 VPWR VGND sg13g2_fill_2
XFILLER_40_940 VPWR VGND sg13g2_decap_8
XFILLER_8_602 VPWR VGND sg13g2_decap_8
XFILLER_12_642 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0820_ VGND VPWR net335 u_ppwm_u_mem__0819_/X u_ppwm_u_mem__0820_/Y
+ hold295/A sg13g2_a21oi_1
XFILLER_8_679 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0751_ u_ppwm_u_mem__0751_/Y net332 u_ppwm_u_mem__0750_/X VPWR VGND
+ sg13g2_nand2b_1
Xu_ppwm_u_mem__0682_ VPWR u_ppwm_u_mem__0682_/Y net519 VGND sg13g2_inv_1
XFILLER_4_874 VPWR VGND sg13g2_decap_8
XFILLER_3_362 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__720_ net442 VPWR u_ppwm_u_ex__720_/Y VGND hold298/A net307 sg13g2_o21ai_1
Xu_ppwm_u_ex__651_ VGND VPWR u_ppwm_u_ex__529_/B net309 u_ppwm_u_ex__809_/D u_ppwm_u_ex__650_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1115__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_35_701 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1165_ net150 VGND VPWR u_ppwm_u_mem__1165_/D hold27/A clknet_5_14__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__582_ u_ppwm_u_ex__581_/Y VPWR u_ppwm_u_ex__582_/Y VGND u_ppwm_u_ex__578_/Y
+ u_ppwm_u_ex__580_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__1096_ net624 u_ppwm_u_mem__1102_/D u_ppwm_u_mem__1098_/B VPWR VGND
+ sg13g2_and2_1
XFILLER_35_778 VPWR VGND sg13g2_decap_8
XFILLER_15_480 VPWR VGND sg13g2_decap_8
XFILLER_22_439 VPWR VGND sg13g2_decap_8
XFILLER_31_984 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0949_ VGND VPWR net373 u_ppwm_u_mem__0680_/Y hold101/A u_ppwm_u_mem__0948_/Y
+ sg13g2_a21oi_1
XFILLER_27_15 VPWR VGND sg13g2_fill_1
XFILLER_38_550 VPWR VGND sg13g2_decap_8
XFILLER_26_734 VPWR VGND sg13g2_decap_8
XFILLER_13_406 VPWR VGND sg13g2_decap_8
XFILLER_41_759 VPWR VGND sg13g2_decap_8
XFILLER_40_225 VPWR VGND sg13g2_decap_4
XFILLER_43_58 VPWR VGND sg13g2_fill_1
XFILLER_21_472 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_decap_8
XFILLER_1_855 VPWR VGND sg13g2_decap_8
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_0_365 VPWR VGND sg13g2_decap_8
XFILLER_48_347 VPWR VGND sg13g2_decap_8
XFILLER_44_564 VPWR VGND sg13g2_decap_8
XFILLER_16_255 VPWR VGND sg13g2_fill_2
XFILLER_17_767 VPWR VGND sg13g2_decap_8
XFILLER_31_247 VPWR VGND sg13g2_decap_8
XFILLER_32_759 VPWR VGND sg13g2_decap_8
XFILLER_13_973 VPWR VGND sg13g2_decap_8
XFILLER_9_955 VPWR VGND sg13g2_decap_8
XFILLER_33_80 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0803_ u_ppwm_u_mem__0694_/Y u_ppwm_u_mem__0687_/Y net416 u_ppwm_u_mem__0803_/X
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_476 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0734_ net619 net618 net582 u_ppwm_u_mem__0737_/C VPWR VGND sg13g2_nand3_1
XFILLER_4_671 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0665_ VPWR u_ppwm_u_mem__0665_/Y net493 VGND sg13g2_inv_1
XFILLER_39_325 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__703_ u_ppwm_u_ex__702_/Y VPWR u_ppwm_u_ex__703_/Y VGND u_ppwm_u_ex__699_/Y
+ u_ppwm_u_ex__701_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__1217_ net60 VGND VPWR net207 hold178/A clknet_5_6__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1148_ net65 VGND VPWR net540 hold198/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__634_ net398 net323 u_ppwm_u_ex__634_/X VPWR VGND sg13g2_and2_1
XFILLER_35_575 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_ex__565_ VPWR VGND u_ppwm_u_ex__561_/Y u_ppwm_u_ex__564_/Y u_ppwm_u_ex__559_/Y
+ net390 u_ppwm_u_ex__565_/Y u_ppwm_u_ex__608_/B sg13g2_a221oi_1
Xu_ppwm_u_mem__1079_ VGND VPWR net345 u_ppwm_u_mem__0615_/Y hold179/A u_ppwm_u_mem__1078_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__496_ u_ppwm_u_ex__496_/Y hold298/A hold30/A VPWR VGND sg13g2_nand2b_1
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_31_781 VPWR VGND sg13g2_decap_8
XFILLER_39_870 VPWR VGND sg13g2_decap_8
XFILLER_26_531 VPWR VGND sg13g2_decap_8
XFILLER_41_501 VPWR VGND sg13g2_decap_4
XFILLER_14_737 VPWR VGND sg13g2_decap_8
XFILLER_41_556 VPWR VGND sg13g2_decap_8
XFILLER_13_258 VPWR VGND sg13g2_fill_2
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_21_291 VPWR VGND sg13g2_fill_1
XFILLER_5_402 VPWR VGND sg13g2_decap_8
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_5_479 VPWR VGND sg13g2_decap_8
XFILLER_1_652 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_0_173 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1136__89 VPWR VGND net89 sg13g2_tiehi
Xu_ppwm_u_mem__1151__59 VPWR VGND net59 sg13g2_tiehi
Xu_ppwm_u_mem__1002_ net434 VPWR u_ppwm_u_mem__1002_/Y VGND net356 net276 sg13g2_o21ai_1
XFILLER_17_564 VPWR VGND sg13g2_decap_8
XFILLER_32_556 VPWR VGND sg13g2_decap_8
XFILLER_13_770 VPWR VGND sg13g2_decap_8
XFILLER_9_752 VPWR VGND sg13g2_decap_8
XFILLER_5_51 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0717_ VPWR u_ppwm_u_mem__0717_/Y net560 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0648_ VPWR u_ppwm_u_mem__0648_/Y net525 VGND sg13g2_inv_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
XFILLER_39_100 VPWR VGND sg13g2_decap_8
XFILLER_27_328 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__617_ u_ppwm_u_ex__617_/A u_ppwm_u_ex__617_/B u_ppwm_u_ex__617_/C u_ppwm_u_ex__617_/D
+ u_ppwm_u_ex__617_/X VPWR VGND sg13g2_and4_1
XFILLER_36_895 VPWR VGND sg13g2_decap_8
XFILLER_11_729 VPWR VGND sg13g2_decap_8
XFILLER_23_567 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__548_ net377 u_ppwm/instr\[2\] u_ppwm_u_ex__637_/A u_ppwm/instr\[1\]
+ u_ppwm_u_ex__617_/A VPWR VGND sg13g2_and4_1
XFILLER_10_228 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__479_ VGND VPWR u_ppwm_u_ex__478_/A u_ppwm_u_ex__478_/B u_ppwm_u_ex__479_/Y
+ u_ppwm_u_ex__488_/B sg13g2_a21oi_1
Xhold251 hold251/A VPWR VGND net594 sg13g2_dlygate4sd3_1
Xhold262 hold262/A VPWR VGND net605 sg13g2_dlygate4sd3_1
Xhold240 hold240/A VPWR VGND net583 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
Xhold273 hold273/A VPWR VGND net616 sg13g2_dlygate4sd3_1
Xhold284 hold284/A VPWR VGND net627 sg13g2_dlygate4sd3_1
Xhold295 hold295/A VPWR VGND net638 sg13g2_dlygate4sd3_1
XFILLER_46_637 VPWR VGND sg13g2_decap_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_42_832 VPWR VGND sg13g2_decap_8
XFILLER_26_383 VPWR VGND sg13g2_decap_4
XFILLER_14_534 VPWR VGND sg13g2_decap_8
XFILLER_41_397 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__241_ net196 VGND VPWR net645 hold300/A clknet_5_1__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__172_ u_ppwm_u_pwm__175_/A u_ppwm_u_pwm__172_/B u_ppwm_u_pwm__239_/D
+ VPWR VGND sg13g2_nor2_1
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_6_755 VPWR VGND sg13g2_decap_8
XFILLER_2_961 VPWR VGND sg13g2_decap_8
XFILLER_49_420 VPWR VGND sg13g2_decap_8
XFILLER_7_1021 VPWR VGND sg13g2_decap_8
XFILLER_49_497 VPWR VGND sg13g2_decap_8
XFILLER_37_659 VPWR VGND sg13g2_decap_8
XFILLER_36_169 VPWR VGND sg13g2_fill_1
XFILLER_18_884 VPWR VGND sg13g2_decap_8
XFILLER_32_353 VPWR VGND sg13g2_fill_2
XFILLER_33_876 VPWR VGND sg13g2_decap_8
XFILLER_20_559 VPWR VGND sg13g2_decap_8
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_28_648 VPWR VGND sg13g2_decap_8
XFILLER_43_607 VPWR VGND sg13g2_decap_8
XFILLER_35_15 VPWR VGND sg13g2_decap_4
XFILLER_24_832 VPWR VGND sg13g2_decap_8
XFILLER_35_191 VPWR VGND sg13g2_fill_2
XFILLER_36_692 VPWR VGND sg13g2_decap_8
XFILLER_23_342 VPWR VGND sg13g2_fill_1
XFILLER_11_526 VPWR VGND sg13g2_decap_8
XFILLER_23_386 VPWR VGND sg13g2_fill_2
XFILLER_13_1015 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_3_747 VPWR VGND sg13g2_decap_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_18_103 VPWR VGND sg13g2_decap_8
XFILLER_34_607 VPWR VGND sg13g2_decap_8
XFILLER_15_865 VPWR VGND sg13g2_decap_8
XFILLER_30_846 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0982_ net430 VPWR u_ppwm_u_mem__0982_/Y VGND net348 net287 sg13g2_o21ai_1
Xu_ppwm_u_pwm__224_ u_ppwm_u_pwm__223_/Y VPWR u_ppwm_u_pwm__225_/B VGND u_ppwm_u_pwm__217_/Y
+ u_ppwm_u_pwm__221_/Y sg13g2_o21ai_1
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_6_552 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__155_ net424 VPWR u_ppwm_u_pwm__155_/Y VGND net389 net329 sg13g2_o21ai_1
XFILLER_29_1011 VPWR VGND sg13g2_decap_8
XFILLER_2_85 VPWR VGND sg13g2_fill_2
XFILLER_38_935 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_18_681 VPWR VGND sg13g2_decap_8
XFILLER_25_618 VPWR VGND sg13g2_decap_8
XFILLER_33_673 VPWR VGND sg13g2_decap_8
XFILLER_21_857 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1125__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_47_209 VPWR VGND sg13g2_decap_8
XFILLER_29_913 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_44_949 VPWR VGND sg13g2_decap_8
XFILLER_12_824 VPWR VGND sg13g2_decap_8
XFILLER_23_194 VPWR VGND sg13g2_fill_2
XFILLER_3_544 VPWR VGND sg13g2_decap_8
XFILLER_47_710 VPWR VGND sg13g2_decap_8
Xfanout391 net675 net391 VPWR VGND sg13g2_buf_8
Xfanout380 net639 net380 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1181_ net90 VGND VPWR u_ppwm_u_mem__1181_/D hold96/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_19_467 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_30_643 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0965_ VGND VPWR net368 u_ppwm_u_mem__0672_/Y u_ppwm_u_mem__1159_/D
+ u_ppwm_u_mem__0964_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__207_ u_ppwm_u_pwm__216_/B hold52/A hold237/A VPWR VGND sg13g2_nand2b_1
XFILLER_11_890 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0896_ net449 VPWR u_ppwm_u_mem__0896_/Y VGND net372 net301 sg13g2_o21ai_1
Xu_ppwm_u_pwm__138_ VPWR u_ppwm_u_pwm__138_/Y net200 VGND sg13g2_inv_1
XFILLER_38_732 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__796_ u_ppwm_u_ex__789_/Y VPWR u_ppwm_u_ex__798_/A VGND u_ppwm_u_ex__788_/Y
+ u_ppwm_u_ex__790_/Y sg13g2_o21ai_1
XFILLER_26_916 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__087_ VGND VPWR hold318/A net331 hold213/A net555 sg13g2_a21oi_1
XFILLER_34_971 VPWR VGND sg13g2_decap_8
XFILLER_21_654 VPWR VGND sg13g2_decap_8
XFILLER_0_547 VPWR VGND sg13g2_decap_8
XFILLER_48_529 VPWR VGND sg13g2_decap_8
XFILLER_29_710 VPWR VGND sg13g2_decap_8
XFILLER_29_787 VPWR VGND sg13g2_decap_8
XFILLER_44_746 VPWR VGND sg13g2_decap_8
XFILLER_43_223 VPWR VGND sg13g2_decap_8
XFILLER_16_448 VPWR VGND sg13g2_decap_8
XFILLER_17_949 VPWR VGND sg13g2_decap_8
XFILLER_12_621 VPWR VGND sg13g2_decap_8
XFILLER_25_982 VPWR VGND sg13g2_decap_8
XFILLER_31_429 VPWR VGND sg13g2_fill_2
XFILLER_40_996 VPWR VGND sg13g2_decap_8
XFILLER_12_698 VPWR VGND sg13g2_decap_8
XFILLER_8_658 VPWR VGND sg13g2_decap_8
XFILLER_7_135 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0750_ net417 u_ppwm_u_mem__1107_/Q hold138/A hold163/A hold136/A net408
+ u_ppwm_u_mem__0750_/X VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0681_ VPWR u_ppwm_u_mem__0681_/Y net548 VGND sg13g2_inv_1
XFILLER_4_853 VPWR VGND sg13g2_decap_8
XFILLER_3_341 VPWR VGND sg13g2_decap_8
XFILLER_26_1014 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1164_ net152 VGND VPWR u_ppwm_u_mem__1164_/D hold17/A clknet_5_15__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__650_ net439 VPWR u_ppwm_u_ex__650_/Y VGND u_ppwm_u_ex__646_/Y u_ppwm_u_ex__649_/Y
+ sg13g2_o21ai_1
XFILLER_47_584 VPWR VGND sg13g2_decap_8
XFILLER_19_275 VPWR VGND sg13g2_decap_4
XFILLER_35_757 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__581_ u_ppwm_u_ex__581_/Y u_ppwm_u_ex__432_/Y net395 u_ppwm_u_ex__494_/B
+ net393 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1095_ net624 u_ppwm_u_mem__1102_/D u_ppwm_u_mem__1097_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_34_256 VPWR VGND sg13g2_decap_8
XFILLER_34_289 VPWR VGND sg13g2_decap_4
XFILLER_31_963 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0948_ net450 VPWR u_ppwm_u_mem__0948_/Y VGND net373 hold205/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0879_ VGND VPWR net370 u_ppwm_u_mem__0715_/Y u_ppwm_u_mem__1116_/D
+ u_ppwm_u_mem__0878_/Y sg13g2_a21oi_1
XFILLER_26_713 VPWR VGND sg13g2_decap_8
XFILLER_14_919 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__779_ u_ppwm_u_ex__779_/B u_ppwm_u_ex__785_/D u_ppwm_u_ex__779_/A u_ppwm_u_ex__781_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_41_738 VPWR VGND sg13g2_decap_8
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_22_985 VPWR VGND sg13g2_decap_8
XFILLER_1_834 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_decap_8
XFILLER_0_344 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1148__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_1_1016 VPWR VGND sg13g2_decap_8
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
XFILLER_16_212 VPWR VGND sg13g2_fill_1
XFILLER_17_746 VPWR VGND sg13g2_decap_8
XFILLER_29_584 VPWR VGND sg13g2_decap_8
XFILLER_44_543 VPWR VGND sg13g2_decap_8
XFILLER_16_267 VPWR VGND sg13g2_fill_2
XFILLER_32_738 VPWR VGND sg13g2_decap_8
XFILLER_13_952 VPWR VGND sg13g2_decap_8
XFILLER_9_934 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_8
XFILLER_8_455 VPWR VGND sg13g2_decap_8
XFILLER_12_495 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0802_ VPWR VGND u_ppwm_u_mem__0801_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0799_/Y
+ u_ppwm_u_mem__0795_/Y u_ppwm_u_mem__0802_/Y u_ppwm_u_mem__0797_/Y sg13g2_a221oi_1
Xu_ppwm_u_mem__0733_ net597 net624 net549 u_ppwm_u_mem__0737_/B VPWR VGND sg13g2_nand3_1
XFILLER_4_650 VPWR VGND sg13g2_decap_8
XFILLER_3_160 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0664_ VPWR u_ppwm_u_mem__0664_/Y net287 VGND sg13g2_inv_1
Xu_ppwm_u_ex__702_ VGND VPWR u_ppwm_u_ex__699_/Y u_ppwm_u_ex__701_/Y u_ppwm_u_ex__702_/Y
+ net315 sg13g2_a21oi_1
XFILLER_48_893 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1216_ net76 VGND VPWR net522 hold249/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__633_ VGND VPWR u_ppwm_u_ex__629_/Y u_ppwm_u_ex__631_/Y hold307/A u_ppwm_u_ex__632_/Y
+ sg13g2_a21oi_1
XFILLER_35_554 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1147_ net67 VGND VPWR net542 hold202/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__564_ u_ppwm_u_ex__563_/Y VPWR u_ppwm_u_ex__564_/Y VGND net390 u_ppwm_u_ex__608_/B
+ sg13g2_o21ai_1
XFILLER_23_749 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1078_ net426 VPWR u_ppwm_u_mem__1078_/Y VGND net345 hold249/A sg13g2_o21ai_1
Xu_ppwm_u_ex__495_ net385 hold266/A u_ppwm_u_ex__495_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_31_760 VPWR VGND sg13g2_decap_8
XFILLER_46_819 VPWR VGND sg13g2_decap_8
XFILLER_26_510 VPWR VGND sg13g2_decap_8
XFILLER_14_716 VPWR VGND sg13g2_decap_8
XFILLER_26_587 VPWR VGND sg13g2_decap_8
XFILLER_41_535 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_22_782 VPWR VGND sg13g2_decap_8
XFILLER_6_937 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_5_458 VPWR VGND sg13g2_decap_8
XFILLER_1_631 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_17_543 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1001_ VGND VPWR net350 u_ppwm_u_mem__0654_/Y hold80/A u_ppwm_u_mem__1000_/Y
+ sg13g2_a21oi_1
XFILLER_45_885 VPWR VGND sg13g2_decap_8
XFILLER_44_395 VPWR VGND sg13g2_fill_2
XFILLER_32_535 VPWR VGND sg13g2_decap_8
XFILLER_40_590 VPWR VGND sg13g2_decap_8
XFILLER_9_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0716_ VPWR u_ppwm_u_mem__0716_/Y net241 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0647_ VPWR u_ppwm_u_mem__0647_/Y net229 VGND sg13g2_inv_1
XFILLER_48_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__616_ u_ppwm_u_ex__615_/Y VPWR u_ppwm_u_ex__617_/D VGND u_ppwm_u_ex__609_/Y
+ u_ppwm_u_ex__614_/Y sg13g2_o21ai_1
XFILLER_36_874 VPWR VGND sg13g2_decap_8
XFILLER_39_1024 VPWR VGND sg13g2_decap_4
XFILLER_23_546 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_fill_1
XFILLER_11_708 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__547_ VGND VPWR u_ppwm_u_ex__543_/Y u_ppwm_u_ex__546_/X u_ppwm_u_ex__547_/Y
+ u_ppwm_u_ex__518_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__478_ VGND VPWR u_ppwm_u_ex__485_/B u_ppwm_u_ex__478_/B u_ppwm_u_ex__478_/A
+ sg13g2_or2_1
XFILLER_3_929 VPWR VGND sg13g2_decap_8
Xhold252 hold252/A VPWR VGND net595 sg13g2_dlygate4sd3_1
Xhold241 hold241/A VPWR VGND net584 sg13g2_dlygate4sd3_1
Xhold230 hold230/A VPWR VGND net573 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold274 hold274/A VPWR VGND net617 sg13g2_dlygate4sd3_1
Xhold285 hold285/A VPWR VGND net628 sg13g2_dlygate4sd3_1
Xhold296 hold296/A VPWR VGND net639 sg13g2_dlygate4sd3_1
Xhold263 hold263/A VPWR VGND net606 sg13g2_dlygate4sd3_1
XFILLER_46_616 VPWR VGND sg13g2_decap_8
XFILLER_18_318 VPWR VGND sg13g2_fill_2
XFILLER_42_811 VPWR VGND sg13g2_decap_8
XFILLER_14_513 VPWR VGND sg13g2_decap_8
XFILLER_26_373 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_42_888 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__240_ net178 VGND VPWR net623 hold278/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_pwm__171_ u_ppwm_u_pwm__172_/B net337 u_ppwm_u_pwm__176_/D VPWR VGND sg13g2_xnor2_1
XFILLER_14_83 VPWR VGND sg13g2_fill_1
XFILLER_6_734 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_fill_1
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_2_940 VPWR VGND sg13g2_decap_8
XFILLER_7_1000 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_37_638 VPWR VGND sg13g2_decap_8
XFILLER_18_863 VPWR VGND sg13g2_decap_8
XFILLER_36_159 VPWR VGND sg13g2_fill_2
XFILLER_45_682 VPWR VGND sg13g2_decap_8
XFILLER_17_373 VPWR VGND sg13g2_decap_4
XFILLER_33_855 VPWR VGND sg13g2_decap_8
XFILLER_20_538 VPWR VGND sg13g2_decap_8
XFILLER_32_398 VPWR VGND sg13g2_fill_1
XFILLER_28_627 VPWR VGND sg13g2_decap_8
XFILLER_27_159 VPWR VGND sg13g2_fill_1
XFILLER_42_107 VPWR VGND sg13g2_fill_1
XFILLER_24_811 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_fill_1
XFILLER_36_671 VPWR VGND sg13g2_decap_8
XFILLER_11_505 VPWR VGND sg13g2_decap_8
XFILLER_24_888 VPWR VGND sg13g2_decap_8
XFILLER_3_726 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__245__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_19_649 VPWR VGND sg13g2_decap_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__828__27 VPWR VGND net27 sg13g2_tiehi
XFILLER_15_844 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_25_71 VPWR VGND sg13g2_fill_1
XFILLER_42_685 VPWR VGND sg13g2_decap_8
XFILLER_30_825 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0981_ VGND VPWR net348 u_ppwm_u_mem__0664_/Y hold91/A u_ppwm_u_mem__0980_/Y
+ sg13g2_a21oi_1
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__223_ VGND VPWR net594 u_ppwm_u_pwm__129_/Y u_ppwm_u_pwm__223_/Y u_ppwm_u_pwm__222_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__154_ VGND VPWR u_ppwm_u_pwm__209_/B net330 hold26/A u_ppwm_u_pwm__153_/Y
+ sg13g2_a21oi_1
XFILLER_6_531 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_fill_2
XFILLER_38_914 VPWR VGND sg13g2_decap_8
XFILLER_49_273 VPWR VGND sg13g2_decap_8
XFILLER_46_980 VPWR VGND sg13g2_decap_8
XFILLER_18_660 VPWR VGND sg13g2_decap_8
XFILLER_33_652 VPWR VGND sg13g2_decap_8
XFILLER_21_836 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_0_729 VPWR VGND sg13g2_decap_8
XFILLER_29_969 VPWR VGND sg13g2_decap_8
XFILLER_44_928 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1212__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_12_803 VPWR VGND sg13g2_decap_8
XFILLER_23_173 VPWR VGND sg13g2_decap_8
XFILLER_24_685 VPWR VGND sg13g2_decap_8
XFILLER_11_324 VPWR VGND sg13g2_fill_1
XFILLER_3_523 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_fill_1
XFILLER_4_1014 VPWR VGND sg13g2_decap_8
Xfanout392 net666 net392 VPWR VGND sg13g2_buf_8
Xfanout381 net663 net381 VPWR VGND sg13g2_buf_8
Xfanout370 net371 net370 VPWR VGND sg13g2_buf_8
XFILLER_47_766 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1180_ net94 VGND VPWR net294 hold167/A clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_446 VPWR VGND sg13g2_decap_8
XFILLER_35_939 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_28_991 VPWR VGND sg13g2_decap_8
XFILLER_36_81 VPWR VGND sg13g2_fill_1
XFILLER_43_950 VPWR VGND sg13g2_decap_8
XFILLER_15_641 VPWR VGND sg13g2_decap_8
XFILLER_42_482 VPWR VGND sg13g2_fill_1
XFILLER_42_471 VPWR VGND sg13g2_decap_8
XFILLER_30_622 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0964_ net445 VPWR u_ppwm_u_mem__0964_/Y VGND net368 net306 sg13g2_o21ai_1
XFILLER_30_699 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__206_ u_ppwm_u_pwm__216_/A u_ppwm_u_pwm__210_/A u_ppwm_u_pwm__210_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0895_ VGND VPWR net371 u_ppwm_u_mem__0707_/Y hold105/A u_ppwm_u_mem__0894_/Y
+ sg13g2_a21oi_1
XFILLER_7_895 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__137_ VPWR u_ppwm_u_pwm__137_/Y net218 VGND sg13g2_inv_1
XFILLER_38_711 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__795_ VGND VPWR u_ppwm_u_ex__792_/Y u_ppwm_u_ex__793_/Y hold304/A u_ppwm_u_ex__794_/Y
+ sg13g2_a21oi_1
XFILLER_38_788 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__086_ hold267/A fanout331/A net336 u_ppwm_u_global_counter__082_/Y
+ u_ppwm_u_global_counter__054_/Y VPWR VGND sg13g2_a22oi_1
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_25_438 VPWR VGND sg13g2_fill_1
XFILLER_34_950 VPWR VGND sg13g2_decap_8
XFILLER_21_633 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__235__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_20_176 VPWR VGND sg13g2_decap_8
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_526 VPWR VGND sg13g2_decap_8
XFILLER_48_508 VPWR VGND sg13g2_decap_8
XFILLER_17_928 VPWR VGND sg13g2_decap_8
XFILLER_29_766 VPWR VGND sg13g2_decap_8
XFILLER_44_725 VPWR VGND sg13g2_decap_8
XFILLER_16_427 VPWR VGND sg13g2_decap_8
XFILLER_25_961 VPWR VGND sg13g2_decap_8
XFILLER_12_600 VPWR VGND sg13g2_decap_8
XFILLER_24_482 VPWR VGND sg13g2_decap_8
XFILLER_40_975 VPWR VGND sg13g2_decap_8
XFILLER_8_637 VPWR VGND sg13g2_decap_8
XFILLER_12_677 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0680_ VPWR u_ppwm_u_mem__0680_/Y net297 VGND sg13g2_inv_1
XFILLER_4_832 VPWR VGND sg13g2_decap_8
XFILLER_3_397 VPWR VGND sg13g2_decap_8
XFILLER_47_563 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1163_ net154 VGND VPWR net215 hold85/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__580_ u_ppwm_u_ex__579_/Y VPWR u_ppwm_u_ex__580_/Y VGND net397 u_ppwm_u_ex__433_/Y
+ sg13g2_o21ai_1
XFILLER_35_736 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1094_ u_ppwm_u_mem__1094_/A net583 u_ppwm_u_mem__1102_/D hold241/A
+ VPWR VGND sg13g2_nor3_1
XFILLER_34_235 VPWR VGND sg13g2_decap_8
XFILLER_16_994 VPWR VGND sg13g2_decap_8
XFILLER_31_942 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0947_ VGND VPWR net374 u_ppwm_u_mem__0681_/Y u_ppwm_u_mem__1150_/D
+ u_ppwm_u_mem__0946_/Y sg13g2_a21oi_1
XFILLER_7_692 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0878_ net447 VPWR u_ppwm_u_mem__0878_/Y VGND net371 net241 sg13g2_o21ai_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_27_39 VPWR VGND sg13g2_fill_1
XFILLER_38_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__069_ net546 net528 net251 u_ppwm_u_global_counter__085_/A
+ VPWR VGND net586 sg13g2_nand4_1
Xu_ppwm_u_ex__778_ u_ppwm_u_ex__785_/D hold310/A net321 VPWR VGND sg13g2_xnor2_1
XFILLER_26_769 VPWR VGND sg13g2_decap_8
XFILLER_41_717 VPWR VGND sg13g2_decap_8
XFILLER_22_964 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__803__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_49_1015 VPWR VGND sg13g2_decap_8
XFILLER_1_813 VPWR VGND sg13g2_decap_8
XFILLER_0_323 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_563 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_decap_8
XFILLER_16_202 VPWR VGND sg13g2_fill_1
XFILLER_17_725 VPWR VGND sg13g2_decap_8
XFILLER_16_257 VPWR VGND sg13g2_fill_1
XFILLER_17_83 VPWR VGND sg13g2_fill_1
XFILLER_44_599 VPWR VGND sg13g2_decap_8
XFILLER_32_717 VPWR VGND sg13g2_decap_8
XFILLER_13_931 VPWR VGND sg13g2_decap_8
XFILLER_40_772 VPWR VGND sg13g2_decap_8
XFILLER_9_913 VPWR VGND sg13g2_decap_8
XFILLER_8_434 VPWR VGND sg13g2_decap_8
XFILLER_12_474 VPWR VGND sg13g2_decap_8
XFILLER_33_93 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0801_ VGND VPWR net335 u_ppwm_u_mem__0800_/X u_ppwm_u_mem__0801_/Y
+ net403 sg13g2_a21oi_1
Xu_ppwm_u_mem__0732_ VGND VPWR u_ppwm_u_mem__0726_/Y u_ppwm_u_mem__0731_/Y hold171/A
+ u_ppwm_u_mem__0730_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0663_ VPWR u_ppwm_u_mem__0663_/Y net617 VGND sg13g2_inv_1
XFILLER_0_890 VPWR VGND sg13g2_decap_8
Xhold1 hold1/A VPWR VGND net198 sg13g2_dlygate4sd3_1
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_48_872 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__701_ u_ppwm_u_ex__701_/Y net386 net319 VPWR VGND sg13g2_xnor2_1
Xu_ppwm_u_mem__1215_ net92 VGND VPWR net593 hold215/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_382 VPWR VGND sg13g2_decap_8
XFILLER_47_360 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1146_ net69 VGND VPWR u_ppwm_u_mem__1146_/D hold83/A clknet_5_25__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__632_ net439 VPWR u_ppwm_u_ex__632_/Y VGND net649 fanout310/A sg13g2_o21ai_1
XFILLER_35_533 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__563_ u_ppwm_u_ex__563_/Y net387 u_ppwm_u_ex__566_/B VPWR VGND sg13g2_nand2_1
XFILLER_23_728 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1077_ VGND VPWR net342 u_ppwm_u_mem__0616_/Y hold250/A u_ppwm_u_mem__1076_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__494_ u_ppwm_u_ex__494_/Y net382 u_ppwm_u_ex__494_/B VPWR VGND sg13g2_nand2_1
XFILLER_16_791 VPWR VGND sg13g2_decap_8
XFILLER_38_382 VPWR VGND sg13g2_fill_1
XFILLER_41_514 VPWR VGND sg13g2_decap_8
XFILLER_26_566 VPWR VGND sg13g2_decap_8
XFILLER_22_761 VPWR VGND sg13g2_decap_8
XFILLER_6_916 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1209__167 VPWR VGND net167 sg13g2_tiehi
XFILLER_5_437 VPWR VGND sg13g2_decap_8
XFILLER_1_610 VPWR VGND sg13g2_decap_8
XFILLER_1_687 VPWR VGND sg13g2_decap_8
XFILLER_49_658 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_17_522 VPWR VGND sg13g2_decap_8
XFILLER_28_82 VPWR VGND sg13g2_fill_2
XFILLER_45_864 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1000_ net434 VPWR u_ppwm_u_mem__1000_/Y VGND net350 hold110/A sg13g2_o21ai_1
XFILLER_17_599 VPWR VGND sg13g2_decap_8
XFILLER_9_710 VPWR VGND sg13g2_decap_8
XFILLER_8_253 VPWR VGND sg13g2_fill_2
XFILLER_8_231 VPWR VGND sg13g2_fill_1
XFILLER_9_787 VPWR VGND sg13g2_decap_8
XFILLER_12_293 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0715_ VPWR u_ppwm_u_mem__0715_/Y net523 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0646_ VPWR u_ppwm_u_mem__0646_/Y net538 VGND sg13g2_inv_1
XFILLER_28_809 VPWR VGND sg13g2_decap_8
XFILLER_39_179 VPWR VGND sg13g2_decap_8
XFILLER_35_330 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__1135__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_36_853 VPWR VGND sg13g2_decap_8
XFILLER_39_1003 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__615_ VGND VPWR u_ppwm_u_ex__611_/Y u_ppwm_u_ex__614_/B u_ppwm_u_ex__615_/Y
+ u_ppwm_u_ex__448_/C sg13g2_a21oi_1
Xu_ppwm_u_mem__1129_ net103 VGND VPWR u_ppwm_u_mem__1129_/D hold157/A clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1150__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_23_525 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_24_29 VPWR VGND sg13g2_fill_1
XFILLER_35_396 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__546_ u_ppwm_u_ex__546_/A u_ppwm_u_ex__546_/B u_ppwm_u_ex__546_/X VPWR
+ VGND sg13g2_and2_1
Xu_ppwm_u_ex__477_ u_ppwm_u_ex__478_/B net402 net323 VPWR VGND sg13g2_xnor2_1
XFILLER_40_17 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_fill_1
Xhold220 hold220/A VPWR VGND net563 sg13g2_dlygate4sd3_1
XFILLER_3_908 VPWR VGND sg13g2_decap_8
Xhold253 hold253/A VPWR VGND net596 sg13g2_dlygate4sd3_1
XFILLER_2_429 VPWR VGND sg13g2_decap_8
Xhold231 hold231/A VPWR VGND net574 sg13g2_dlygate4sd3_1
Xhold242 hold242/A VPWR VGND net585 sg13g2_dlygate4sd3_1
Xhold286 hold286/A VPWR VGND net629 sg13g2_dlygate4sd3_1
Xhold275 hold275/A VPWR VGND net618 sg13g2_dlygate4sd3_1
Xhold264 hold264/A VPWR VGND net607 sg13g2_dlygate4sd3_1
Xhold297 hold297/A VPWR VGND net640 sg13g2_dlygate4sd3_1
XFILLER_26_352 VPWR VGND sg13g2_decap_4
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_42_867 VPWR VGND sg13g2_decap_8
XFILLER_14_569 VPWR VGND sg13g2_decap_8
XFILLER_41_377 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__170_ u_ppwm_u_pwm__175_/A net612 u_ppwm_u_pwm__176_/D hold270/A VPWR
+ VGND sg13g2_nor3_1
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_6_713 VPWR VGND sg13g2_decap_8
XFILLER_2_996 VPWR VGND sg13g2_decap_8
XFILLER_1_484 VPWR VGND sg13g2_decap_8
XFILLER_49_455 VPWR VGND sg13g2_decap_8
XFILLER_36_116 VPWR VGND sg13g2_fill_1
XFILLER_37_617 VPWR VGND sg13g2_decap_8
XFILLER_18_842 VPWR VGND sg13g2_decap_8
XFILLER_45_661 VPWR VGND sg13g2_decap_8
XFILLER_33_834 VPWR VGND sg13g2_decap_8
XFILLER_20_517 VPWR VGND sg13g2_decap_8
XFILLER_9_584 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0629_ VPWR u_ppwm_u_mem__0629_/Y net473 VGND sg13g2_inv_1
XFILLER_28_606 VPWR VGND sg13g2_decap_8
XFILLER_27_127 VPWR VGND sg13g2_fill_2
XFILLER_36_650 VPWR VGND sg13g2_decap_8
XFILLER_24_867 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__529_ net384 u_ppwm_u_ex__529_/B u_ppwm_u_ex__529_/C u_ppwm_u_ex__534_/A
+ VPWR VGND sg13g2_nor3_1
XFILLER_3_705 VPWR VGND sg13g2_decap_8
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_19_628 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_15_823 VPWR VGND sg13g2_decap_8
XFILLER_42_664 VPWR VGND sg13g2_decap_8
XFILLER_30_804 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0980_ net430 VPWR u_ppwm_u_mem__0980_/Y VGND net348 hold150/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__222_ u_ppwm_u_pwm__222_/A u_ppwm_u_pwm__219_/Y u_ppwm_u_pwm__222_/Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_510 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__153_ net424 VPWR u_ppwm_u_pwm__153_/Y VGND net391 net330 sg13g2_o21ai_1
XFILLER_6_587 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_2_793 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_2_76 VPWR VGND sg13g2_fill_1
XFILLER_2_87 VPWR VGND sg13g2_fill_1
XFILLER_17_182 VPWR VGND sg13g2_decap_8
XFILLER_33_631 VPWR VGND sg13g2_decap_8
XFILLER_21_815 VPWR VGND sg13g2_decap_8
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_708 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_948 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_16_609 VPWR VGND sg13g2_decap_8
XFILLER_37_981 VPWR VGND sg13g2_decap_8
XFILLER_24_664 VPWR VGND sg13g2_decap_8
XFILLER_8_819 VPWR VGND sg13g2_decap_8
XFILLER_12_859 VPWR VGND sg13g2_decap_8
XFILLER_23_196 VPWR VGND sg13g2_fill_1
XFILLER_11_369 VPWR VGND sg13g2_fill_2
XFILLER_20_881 VPWR VGND sg13g2_decap_8
XFILLER_3_502 VPWR VGND sg13g2_decap_8
XFILLER_3_579 VPWR VGND sg13g2_decap_8
Xfanout371 net372 net371 VPWR VGND sg13g2_buf_8
Xfanout393 hold323/A net393 VPWR VGND sg13g2_buf_2
Xfanout382 net636 net382 VPWR VGND sg13g2_buf_8
Xfanout360 net363 net360 VPWR VGND sg13g2_buf_8
XFILLER_47_745 VPWR VGND sg13g2_decap_8
XFILLER_46_222 VPWR VGND sg13g2_decap_8
XFILLER_19_425 VPWR VGND sg13g2_decap_8
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_35_918 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_14_141 VPWR VGND sg13g2_fill_2
XFILLER_15_697 VPWR VGND sg13g2_decap_8
XFILLER_30_601 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0963_ VGND VPWR net374 u_ppwm_u_mem__0673_/Y u_ppwm_u_mem__1158_/D
+ u_ppwm_u_mem__0962_/Y sg13g2_a21oi_1
XFILLER_30_678 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__205_ u_ppwm_u_pwm__210_/B hold283/A hold23/A VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0894_ net450 VPWR u_ppwm_u_mem__0894_/Y VGND net371 hold140/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__136_ VPWR u_ppwm_u_pwm__136_/Y net562 VGND sg13g2_inv_1
XFILLER_7_874 VPWR VGND sg13g2_decap_8
XFILLER_6_340 VPWR VGND sg13g2_fill_2
XFILLER_6_384 VPWR VGND sg13g2_decap_8
XFILLER_2_590 VPWR VGND sg13g2_decap_8
XFILLER_42_1021 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1184__78 VPWR VGND net78 sg13g2_tiehi
Xu_ppwm_u_global_counter__085_ u_ppwm_u_global_counter__085_/A u_ppwm_u_global_counter__085_/B
+ u_ppwm_u_global_counter__085_/C fanout331/A VPWR VGND sg13g2_nor3_2
Xu_ppwm_u_ex__794_ net441 VPWR u_ppwm_u_ex__794_/Y VGND net646 net308 sg13g2_o21ai_1
XFILLER_37_255 VPWR VGND sg13g2_fill_1
XFILLER_38_767 VPWR VGND sg13g2_decap_8
XFILLER_19_992 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_decap_8
XFILLER_21_612 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_21_689 VPWR VGND sg13g2_decap_8
XFILLER_0_505 VPWR VGND sg13g2_decap_8
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_28_200 VPWR VGND sg13g2_fill_1
XFILLER_28_211 VPWR VGND sg13g2_decap_8
XFILLER_29_745 VPWR VGND sg13g2_decap_8
XFILLER_44_704 VPWR VGND sg13g2_decap_8
XFILLER_16_406 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_decap_8
XFILLER_28_288 VPWR VGND sg13g2_fill_2
XFILLER_43_258 VPWR VGND sg13g2_fill_1
XFILLER_25_940 VPWR VGND sg13g2_decap_8
XFILLER_43_269 VPWR VGND sg13g2_fill_2
XFILLER_24_461 VPWR VGND sg13g2_decap_8
XFILLER_40_954 VPWR VGND sg13g2_decap_8
XFILLER_8_616 VPWR VGND sg13g2_decap_8
XFILLER_12_656 VPWR VGND sg13g2_decap_8
XFILLER_11_199 VPWR VGND sg13g2_decap_4
XFILLER_4_811 VPWR VGND sg13g2_decap_8
XFILLER_4_888 VPWR VGND sg13g2_decap_8
XFILLER_3_376 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1219__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_47_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1154__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_47_70 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1162_ net156 VGND VPWR net283 hold216/A clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_715 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1093_ net582 net619 net618 net338 u_ppwm_u_mem__1102_/D VPWR VGND sg13g2_and4_1
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_31_921 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_30_420 VPWR VGND sg13g2_fill_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
XFILLER_30_486 VPWR VGND sg13g2_fill_2
XFILLER_31_998 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0946_ net450 VPWR u_ppwm_u_mem__0946_/Y VGND net374 net519 sg13g2_o21ai_1
XFILLER_7_671 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0877_ VGND VPWR net361 u_ppwm_u_mem__0716_/Y hold45/A u_ppwm_u_mem__0876_/Y
+ sg13g2_a21oi_1
XFILLER_33_0 VPWR VGND sg13g2_fill_2
XFILLER_38_564 VPWR VGND sg13g2_decap_8
XFILLER_26_748 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__068_ u_ppwm_u_global_counter__068_/B net528 hold186/A VPWR
+ VGND sg13g2_xor2_1
Xu_ppwm_u_ex__777_ VGND VPWR u_ppwm_u_ex__774_/Y u_ppwm_u_ex__775_/Y hold297/A u_ppwm_u_ex__776_/Y
+ sg13g2_a21oi_1
XFILLER_22_943 VPWR VGND sg13g2_decap_8
XFILLER_21_486 VPWR VGND sg13g2_decap_8
XFILLER_5_619 VPWR VGND sg13g2_decap_8
XFILLER_0_302 VPWR VGND sg13g2_decap_8
XFILLER_1_869 VPWR VGND sg13g2_decap_8
XFILLER_0_379 VPWR VGND sg13g2_decap_8
XFILLER_17_704 VPWR VGND sg13g2_decap_8
XFILLER_29_542 VPWR VGND sg13g2_decap_8
XFILLER_44_501 VPWR VGND sg13g2_decap_8
XFILLER_44_578 VPWR VGND sg13g2_decap_8
XFILLER_13_910 VPWR VGND sg13g2_decap_8
XFILLER_40_751 VPWR VGND sg13g2_decap_8
XFILLER_8_413 VPWR VGND sg13g2_decap_8
XFILLER_12_453 VPWR VGND sg13g2_decap_8
XFILLER_13_987 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_fill_1
XFILLER_33_50 VPWR VGND sg13g2_fill_2
XFILLER_9_969 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0800_ hold56/A hold106/A net411 u_ppwm_u_mem__0800_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0731_ net1 u_ppwm_u_mem__1094_/A u_ppwm_u_mem__0731_/Y VPWR VGND sg13g2_nor2_1
Xu_ppwm_u_mem__0662_ VPWR u_ppwm_u_mem__0662_/Y net487 VGND sg13g2_inv_1
XFILLER_4_685 VPWR VGND sg13g2_decap_8
XFILLER_3_195 VPWR VGND sg13g2_decap_4
Xhold2 hold2/A VPWR VGND net199 sg13g2_dlygate4sd3_1
XFILLER_48_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__700_ u_ppwm_u_ex__700_/Y net386 net319 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1214_ net108 VGND VPWR u_ppwm_u_mem__1214_/D hold200/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1191__169 VPWR VGND net169 sg13g2_tiehi
Xu_ppwm_u_ex__631_ u_ppwm_u_ex__631_/Y net314 net398 net317 net325 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1145_ net71 VGND VPWR net281 hold123/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__562_ net390 u_ppwm_u_ex__608_/B u_ppwm_u_ex__562_/Y VPWR VGND sg13g2_nor2_1
XFILLER_16_770 VPWR VGND sg13g2_decap_8
XFILLER_22_206 VPWR VGND sg13g2_decap_4
XFILLER_23_707 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1076_ net429 VPWR u_ppwm_u_mem__1076_/Y VGND net343 net558 sg13g2_o21ai_1
XFILLER_35_589 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__493_ u_ppwm_u_ex__493_/Y net198 u_ppwm_u_ex__520_/A net614 u_ppwm_u_ex__519_/A
+ VPWR VGND sg13g2_a22oi_1
XFILLER_31_795 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1217__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_8_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0929_ VGND VPWR net364 u_ppwm_u_mem__0690_/Y hold93/A u_ppwm_u_mem__0928_/Y
+ sg13g2_a21oi_1
XFILLER_39_884 VPWR VGND sg13g2_decap_8
XFILLER_26_545 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__829_ net43 VGND VPWR u_ppwm_u_ex__829_/D hold288/A clknet_5_18__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
XFILLER_22_740 VPWR VGND sg13g2_decap_8
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_21_261 VPWR VGND sg13g2_decap_8
XFILLER_5_416 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_fill_1
XFILLER_1_666 VPWR VGND sg13g2_decap_8
XFILLER_49_637 VPWR VGND sg13g2_decap_8
XFILLER_0_187 VPWR VGND sg13g2_decap_8
XFILLER_23_1008 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_17_501 VPWR VGND sg13g2_decap_8
XFILLER_45_843 VPWR VGND sg13g2_decap_8
XFILLER_17_578 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1112__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_44_397 VPWR VGND sg13g2_fill_1
XFILLER_13_784 VPWR VGND sg13g2_decap_8
XFILLER_9_766 VPWR VGND sg13g2_decap_8
XFILLER_5_983 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0714_ VPWR u_ppwm_u_mem__0714_/Y net464 VGND sg13g2_inv_1
XFILLER_4_482 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0645_ VPWR u_ppwm_u_mem__0645_/Y net508 VGND sg13g2_inv_1
XFILLER_36_832 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__614_ u_ppwm_u_ex__614_/B u_ppwm_u_ex__614_/C u_ppwm_u_ex__614_/Y VPWR
+ VGND u_ppwm_u_ex__611_/Y sg13g2_nand3b_1
XFILLER_23_504 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1128_ net105 VGND VPWR u_ppwm_u_mem__1128_/D hold136/A clknet_5_23__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__545_ VGND VPWR u_ppwm_u_ex__543_/B u_ppwm_u_ex__541_/Y u_ppwm_u_ex__546_/B
+ u_ppwm_u_ex__538_/Y sg13g2_a21oi_1
XFILLER_35_375 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1059_ VGND VPWR net341 u_ppwm_u_mem__0625_/Y u_ppwm_u_mem__1206_/D
+ u_ppwm_u_mem__1058_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__476_ u_ppwm_u_ex__485_/A net402 net323 VPWR VGND sg13g2_nand2_1
XFILLER_31_592 VPWR VGND sg13g2_decap_8
Xhold210 hold210/A VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold243 hold243/A VPWR VGND net586 sg13g2_dlygate4sd3_1
XFILLER_2_408 VPWR VGND sg13g2_decap_8
Xhold221 hold221/A VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold232 hold232/A VPWR VGND net575 sg13g2_dlygate4sd3_1
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
Xhold287 hold287/A VPWR VGND net630 sg13g2_dlygate4sd3_1
Xhold254 hold254/A VPWR VGND net597 sg13g2_dlygate4sd3_1
Xhold276 hold276/A VPWR VGND net619 sg13g2_dlygate4sd3_1
Xhold265 hold265/A VPWR VGND net608 sg13g2_dlygate4sd3_1
XFILLER_49_49 VPWR VGND sg13g2_decap_8
Xhold298 hold298/A VPWR VGND net641 sg13g2_dlygate4sd3_1
XFILLER_39_681 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_42_846 VPWR VGND sg13g2_decap_8
XFILLER_14_548 VPWR VGND sg13g2_decap_8
XFILLER_26_397 VPWR VGND sg13g2_fill_2
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_6_769 VPWR VGND sg13g2_decap_8
XFILLER_2_975 VPWR VGND sg13g2_decap_8
XFILLER_1_463 VPWR VGND sg13g2_decap_8
XFILLER_49_434 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_decap_8
XFILLER_45_640 VPWR VGND sg13g2_decap_8
XFILLER_33_813 VPWR VGND sg13g2_decap_8
XFILLER_18_898 VPWR VGND sg13g2_decap_8
XFILLER_13_581 VPWR VGND sg13g2_decap_8
XFILLER_9_563 VPWR VGND sg13g2_decap_8
XFILLER_5_780 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0628_ VPWR u_ppwm_u_mem__0628_/Y net489 VGND sg13g2_inv_1
XFILLER_24_846 VPWR VGND sg13g2_decap_8
XFILLER_35_172 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__528_ u_ppwm_u_ex__527_/Y VPWR u_ppwm_u_ex__528_/Y VGND u_ppwm_u_ex__524_/Y
+ u_ppwm_u_ex__526_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__459_ net377 VPWR u_ppwm_u_ex__459_/Y VGND net327 u_ppwm_u_ex__488_/B
+ sg13g2_o21ai_1
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_19_607 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_15_802 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_26_150 VPWR VGND sg13g2_fill_1
XFILLER_42_643 VPWR VGND sg13g2_decap_8
XFILLER_14_323 VPWR VGND sg13g2_decap_4
XFILLER_15_879 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__221_ u_ppwm_u_pwm__221_/Y u_ppwm_u_pwm__222_/A u_ppwm_u_pwm__221_/B
+ VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_pwm__152_ VGND VPWR u_ppwm_u_pwm__214_/B net330 hold108/A u_ppwm_u_pwm__151_/Y
+ sg13g2_a21oi_1
XFILLER_6_566 VPWR VGND sg13g2_decap_8
XFILLER_29_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_772 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_4
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_2_55 VPWR VGND sg13g2_fill_1
XFILLER_38_949 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__819__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_18_695 VPWR VGND sg13g2_decap_8
XFILLER_33_610 VPWR VGND sg13g2_decap_8
XFILLER_36_1007 VPWR VGND sg13g2_decap_8
XFILLER_33_687 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1164__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_29_927 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_37_960 VPWR VGND sg13g2_decap_8
XFILLER_24_643 VPWR VGND sg13g2_decap_8
XFILLER_12_838 VPWR VGND sg13g2_decap_8
XFILLER_11_315 VPWR VGND sg13g2_decap_8
XFILLER_11_348 VPWR VGND sg13g2_fill_1
XFILLER_20_860 VPWR VGND sg13g2_decap_8
XFILLER_3_558 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xfanout350 net352 net350 VPWR VGND sg13g2_buf_8
Xfanout372 net375 net372 VPWR VGND sg13g2_buf_8
Xfanout383 fanout383/A net383 VPWR VGND sg13g2_buf_8
Xfanout361 net363 net361 VPWR VGND sg13g2_buf_1
XFILLER_47_724 VPWR VGND sg13g2_decap_8
XFILLER_46_212 VPWR VGND sg13g2_fill_1
Xfanout394 net664 net394 VPWR VGND sg13g2_buf_8
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_15_676 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0962_ net449 VPWR u_ppwm_u_mem__0962_/Y VGND net373 net237 sg13g2_o21ai_1
XFILLER_30_657 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__204_ u_ppwm_u_pwm__210_/A hold237/A hold52/A VPWR VGND sg13g2_nand2b_1
XFILLER_7_853 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__135_ VPWR u_ppwm_u_pwm__135_/Y net496 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0893_ VGND VPWR net372 u_ppwm_u_mem__0708_/Y hold141/A u_ppwm_u_mem__0892_/Y
+ sg13g2_a21oi_1
XFILLER_6_363 VPWR VGND sg13g2_decap_8
XFILLER_42_1000 VPWR VGND sg13g2_decap_8
XFILLER_38_746 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__084_ hold314/A net227 net291 u_ppwm_u_global_counter__085_/C
+ VPWR VGND net609 sg13g2_nand4_1
Xu_ppwm_u_ex__793_ VPWR VGND hold310/A u_ppwm_u_ex__714_/Y net312 net378 u_ppwm_u_ex__793_/Y
+ fanout314/A sg13g2_a221oi_1
XFILLER_37_234 VPWR VGND sg13g2_decap_8
XFILLER_19_971 VPWR VGND sg13g2_decap_8
XFILLER_18_492 VPWR VGND sg13g2_decap_8
XFILLER_34_985 VPWR VGND sg13g2_decap_8
XFILLER_21_668 VPWR VGND sg13g2_decap_8
XFILLER_28_223 VPWR VGND sg13g2_decap_8
XFILLER_29_724 VPWR VGND sg13g2_decap_8
XFILLER_28_267 VPWR VGND sg13g2_fill_2
XFILLER_43_237 VPWR VGND sg13g2_fill_1
XFILLER_19_1013 VPWR VGND sg13g2_decap_8
XFILLER_24_440 VPWR VGND sg13g2_decap_8
XFILLER_25_996 VPWR VGND sg13g2_decap_8
XFILLER_40_933 VPWR VGND sg13g2_decap_8
XFILLER_12_635 VPWR VGND sg13g2_decap_8
XFILLER_11_167 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__821__46 VPWR VGND net46 sg13g2_tiehi
XFILLER_4_867 VPWR VGND sg13g2_decap_8
XFILLER_3_355 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_521 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1161_ net158 VGND VPWR u_ppwm_u_mem__1161_/D hold59/A clknet_5_26__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_47_598 VPWR VGND sg13g2_decap_8
XFILLER_34_204 VPWR VGND sg13g2_fill_2
XFILLER_16_952 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1092_ VGND VPWR net582 u_ppwm_u_mem__1085_/B hold240/A u_ppwm_u_mem__1091_/C
+ sg13g2_a21oi_1
XFILLER_31_900 VPWR VGND sg13g2_decap_8
XFILLER_43_782 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_decap_8
XFILLER_31_977 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0945_ VGND VPWR net373 u_ppwm_u_mem__0682_/Y hold177/A u_ppwm_u_mem__0944_/Y
+ sg13g2_a21oi_1
XFILLER_7_650 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0876_ net447 VPWR u_ppwm_u_mem__0876_/Y VGND net360 hold217/A sg13g2_o21ai_1
Xu_ppwm_u_mem__1122__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_38_543 VPWR VGND sg13g2_decap_8
XFILLER_25_215 VPWR VGND sg13g2_fill_2
XFILLER_26_727 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__067_ hold204/A net546 u_ppwm_u_global_counter__067_/B VPWR
+ VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__776_ net441 VPWR u_ppwm_u_ex__776_/Y VGND net639 net308 sg13g2_o21ai_1
XFILLER_25_248 VPWR VGND sg13g2_fill_2
XFILLER_22_922 VPWR VGND sg13g2_decap_8
XFILLER_34_782 VPWR VGND sg13g2_decap_8
XFILLER_40_218 VPWR VGND sg13g2_decap_8
XFILLER_40_229 VPWR VGND sg13g2_fill_2
XFILLER_21_465 VPWR VGND sg13g2_decap_8
XFILLER_22_999 VPWR VGND sg13g2_decap_8
XFILLER_1_848 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_0_358 VPWR VGND sg13g2_decap_8
XFILLER_48_318 VPWR VGND sg13g2_decap_4
XFILLER_29_598 VPWR VGND sg13g2_decap_8
XFILLER_44_557 VPWR VGND sg13g2_decap_8
XFILLER_16_226 VPWR VGND sg13g2_fill_1
XFILLER_40_730 VPWR VGND sg13g2_decap_8
XFILLER_25_793 VPWR VGND sg13g2_decap_8
XFILLER_12_432 VPWR VGND sg13g2_decap_8
XFILLER_13_966 VPWR VGND sg13g2_decap_8
XFILLER_9_948 VPWR VGND sg13g2_decap_8
XFILLER_8_469 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1225__174 VPWR VGND net174 sg13g2_tiehi
Xu_ppwm_u_mem__0730_ u_ppwm_u_mem__0730_/A u_ppwm_u_mem__1094_/A hold282/A u_ppwm_u_mem__0730_/Y
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__0661_ VPWR u_ppwm_u_mem__0661_/Y net467 VGND sg13g2_inv_1
XFILLER_4_664 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_fill_2
XFILLER_48_830 VPWR VGND sg13g2_decap_8
Xhold3 hold3/A VPWR VGND net200 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1213_ net124 VGND VPWR u_ppwm_u_mem__1213_/D hold36/A clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__630_ u_ppwm_u_ex__637_/A net325 net317 fanout314/A VPWR VGND sg13g2_nor3_2
Xu_ppwm_u_mem__1144_ net73 VGND VPWR u_ppwm_u_mem__1144_/D hold116/A clknet_5_30__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__561_ VGND VPWR u_ppwm_u_ex__583_/A hold243/A u_ppwm_u_ex__561_/Y u_ppwm_u_ex__560_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__1075_ VGND VPWR net340 u_ppwm_u_mem__0617_/Y u_ppwm_u_mem__1214_/D
+ u_ppwm_u_mem__1074_/Y sg13g2_a21oi_1
XFILLER_35_568 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__492_ u_ppwm_u_ex__492_/A net632 hold290/A VPWR VGND sg13g2_nor2_1
XFILLER_30_273 VPWR VGND sg13g2_fill_2
XFILLER_31_774 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0928_ net444 VPWR u_ppwm_u_mem__0928_/Y VGND net364 hold263/A sg13g2_o21ai_1
Xu_ppwm_u_mem__0859_ u_ppwm_u_mem__0858_/Y u_ppwm_u_mem__0856_/Y u_ppwm_u_mem__0852_/Y
+ fanout322/A VPWR VGND sg13g2_a21o_2
XFILLER_39_863 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__119_ net440 VGND VPWR net616 hold272/A clknet_5_20__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__828_ net27 VGND VPWR u_ppwm_u_ex__828_/D hold264/A clknet_5_13__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_26_524 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__759_ u_ppwm_u_ex__785_/B net381 net321 VPWR VGND sg13g2_xnor2_1
XFILLER_41_549 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_22_796 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_645 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_0_166 VPWR VGND sg13g2_decap_8
XFILLER_45_822 VPWR VGND sg13g2_decap_8
XFILLER_17_557 VPWR VGND sg13g2_decap_8
XFILLER_45_899 VPWR VGND sg13g2_decap_8
XFILLER_32_549 VPWR VGND sg13g2_decap_8
XFILLER_25_590 VPWR VGND sg13g2_decap_8
XFILLER_9_745 VPWR VGND sg13g2_decap_8
XFILLER_13_763 VPWR VGND sg13g2_decap_8
XFILLER_8_255 VPWR VGND sg13g2_fill_1
XFILLER_5_11 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0713_ VPWR u_ppwm_u_mem__0713_/Y net469 VGND sg13g2_inv_1
XFILLER_5_962 VPWR VGND sg13g2_decap_8
XFILLER_4_461 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0644_ VPWR u_ppwm_u_mem__0644_/Y net239 VGND sg13g2_inv_1
XFILLER_36_811 VPWR VGND sg13g2_decap_8
XFILLER_47_181 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__613_ u_ppwm_u_ex__614_/C u_ppwm_u_ex__566_/B hold310/A u_ppwm_u_ex__435_/Y
+ net379 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1127_ net107 VGND VPWR net480 hold194/A clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_354 VPWR VGND sg13g2_decap_4
XFILLER_36_888 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__544_ net327 u_ppwm_u_ex__637_/B net324 u_ppwm_u_ex__546_/A VPWR VGND
+ sg13g2_nor3_1
XFILLER_35_398 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1058_ net428 VPWR u_ppwm_u_mem__1058_/Y VGND net341 net212 sg13g2_o21ai_1
Xu_ppwm_u_ex__475_ VGND VPWR net407 net326 u_ppwm_u_ex__478_/A u_ppwm_u_ex__469_/C
+ sg13g2_a21oi_1
XFILLER_31_571 VPWR VGND sg13g2_decap_8
Xhold211 hold211/A VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold200 hold200/A VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold233 hold233/A VPWR VGND net576 sg13g2_dlygate4sd3_1
Xhold244 hold244/A VPWR VGND net587 sg13g2_dlygate4sd3_1
Xhold222 hold222/A VPWR VGND net565 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
Xhold266 hold266/A VPWR VGND net609 sg13g2_dlygate4sd3_1
Xhold255 hold255/A VPWR VGND net598 sg13g2_dlygate4sd3_1
Xhold277 hold277/A VPWR VGND net620 sg13g2_dlygate4sd3_1
Xhold299 hold299/A VPWR VGND net642 sg13g2_dlygate4sd3_1
Xhold288 hold288/A VPWR VGND net631 sg13g2_dlygate4sd3_1
XFILLER_22_1020 VPWR VGND sg13g2_decap_8
XFILLER_39_660 VPWR VGND sg13g2_decap_8
XFILLER_26_321 VPWR VGND sg13g2_decap_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_42_825 VPWR VGND sg13g2_decap_8
XFILLER_41_324 VPWR VGND sg13g2_fill_1
XFILLER_14_527 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_53 VPWR VGND sg13g2_fill_2
XFILLER_22_593 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_14_97 VPWR VGND sg13g2_fill_1
XFILLER_6_748 VPWR VGND sg13g2_decap_8
XFILLER_2_954 VPWR VGND sg13g2_decap_8
XFILLER_1_442 VPWR VGND sg13g2_decap_8
XFILLER_49_413 VPWR VGND sg13g2_decap_8
XFILLER_7_1014 VPWR VGND sg13g2_decap_8
XFILLER_18_800 VPWR VGND sg13g2_decap_8
XFILLER_18_877 VPWR VGND sg13g2_decap_8
XFILLER_45_696 VPWR VGND sg13g2_decap_8
XFILLER_33_869 VPWR VGND sg13g2_decap_8
XFILLER_13_560 VPWR VGND sg13g2_decap_8
XFILLER_9_542 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0627_ VPWR u_ppwm_u_mem__0627_/Y net262 VGND sg13g2_inv_1
XFILLER_49_980 VPWR VGND sg13g2_decap_8
XFILLER_35_19 VPWR VGND sg13g2_fill_2
XFILLER_24_825 VPWR VGND sg13g2_decap_8
XFILLER_36_685 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__527_ u_ppwm_u_ex__527_/Y net397 u_ppwm_u_ex__420_/Y net394 u_ppwm_u_ex__419_/Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_11_519 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__458_ u_ppwm/instr\[0\] u_ppwm_u_ex__458_/C u_ppwm/instr\[2\] u_ppwm_u_ex__488_/B
+ VPWR VGND sg13g2_nand3_1
XFILLER_13_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_906 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_42_622 VPWR VGND sg13g2_decap_8
XFILLER_15_858 VPWR VGND sg13g2_decap_8
XFILLER_25_63 VPWR VGND sg13g2_fill_1
XFILLER_42_699 VPWR VGND sg13g2_decap_8
XFILLER_25_85 VPWR VGND sg13g2_decap_4
XFILLER_30_839 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__220_ u_ppwm_u_pwm__221_/B net264 u_ppwm_u_pwm__185_/A net568 u_ppwm_u_pwm__219_/A
+ VPWR VGND sg13g2_a22oi_1
XFILLER_10_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__151_ net425 VPWR u_ppwm_u_pwm__151_/Y VGND net392 net330 sg13g2_o21ai_1
XFILLER_6_545 VPWR VGND sg13g2_decap_8
XFILLER_29_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_751 VPWR VGND sg13g2_decap_8
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_38_928 VPWR VGND sg13g2_decap_8
XFILLER_49_287 VPWR VGND sg13g2_decap_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
XFILLER_18_674 VPWR VGND sg13g2_decap_8
XFILLER_45_493 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_33_666 VPWR VGND sg13g2_decap_8
XFILLER_14_891 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1187__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_29_906 VPWR VGND sg13g2_decap_8
XFILLER_36_471 VPWR VGND sg13g2_decap_4
XFILLER_24_622 VPWR VGND sg13g2_decap_8
XFILLER_12_817 VPWR VGND sg13g2_decap_8
XFILLER_23_187 VPWR VGND sg13g2_decap_8
XFILLER_24_699 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_fill_2
XFILLER_3_537 VPWR VGND sg13g2_decap_8
Xfanout340 net342 net340 VPWR VGND sg13g2_buf_8
XFILLER_47_703 VPWR VGND sg13g2_decap_8
Xfanout373 net374 net373 VPWR VGND sg13g2_buf_8
Xfanout351 net352 net351 VPWR VGND sg13g2_buf_2
Xfanout384 net658 net384 VPWR VGND sg13g2_buf_8
Xfanout362 net363 net362 VPWR VGND sg13g2_buf_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
Xfanout395 hold321/A net395 VPWR VGND sg13g2_buf_1
XFILLER_46_246 VPWR VGND sg13g2_fill_2
XFILLER_34_408 VPWR VGND sg13g2_fill_2
XFILLER_36_95 VPWR VGND sg13g2_fill_2
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_14_143 VPWR VGND sg13g2_fill_1
XFILLER_15_655 VPWR VGND sg13g2_decap_8
XFILLER_42_496 VPWR VGND sg13g2_decap_8
XFILLER_14_187 VPWR VGND sg13g2_decap_8
XFILLER_30_636 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0961_ VGND VPWR net373 u_ppwm_u_mem__0674_/Y hold41/A u_ppwm_u_mem__0960_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_mem__0892_ net450 VPWR u_ppwm_u_mem__0892_/Y VGND net371 hold248/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__203_ u_ppwm_u_pwm__202_/Y u_ppwm_u_pwm__199_/Y u_ppwm_u_pwm__198_/Y
+ u_ppwm_u_pwm__203_/X VPWR VGND sg13g2_a21o_1
XFILLER_7_832 VPWR VGND sg13g2_decap_8
XFILLER_11_883 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__134_ VPWR u_ppwm_u_pwm__214_/B net304 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1194__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_28_4 VPWR VGND sg13g2_fill_2
XFILLER_38_725 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__083_ hold31/A net227 u_ppwm_u_global_counter__083_/B VPWR
+ VGND sg13g2_xnor2_1
XFILLER_19_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__792_ u_ppwm_u_ex__791_/Y VPWR u_ppwm_u_ex__792_/Y VGND u_ppwm_u_ex__788_/Y
+ u_ppwm_u_ex__790_/Y sg13g2_o21ai_1
XFILLER_26_909 VPWR VGND sg13g2_decap_8
XFILLER_18_471 VPWR VGND sg13g2_decap_8
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_33_452 VPWR VGND sg13g2_fill_2
XFILLER_33_463 VPWR VGND sg13g2_fill_2
XFILLER_34_964 VPWR VGND sg13g2_decap_8
XFILLER_21_647 VPWR VGND sg13g2_decap_8
XFILLER_20_124 VPWR VGND sg13g2_fill_2
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_703 VPWR VGND sg13g2_decap_8
XFILLER_44_739 VPWR VGND sg13g2_decap_8
XFILLER_40_912 VPWR VGND sg13g2_decap_8
XFILLER_25_975 VPWR VGND sg13g2_decap_8
XFILLER_12_614 VPWR VGND sg13g2_decap_8
XFILLER_24_496 VPWR VGND sg13g2_decap_8
XFILLER_40_989 VPWR VGND sg13g2_decap_8
XFILLER_4_846 VPWR VGND sg13g2_decap_8
XFILLER_3_334 VPWR VGND sg13g2_decap_8
XFILLER_26_1007 VPWR VGND sg13g2_decap_8
XFILLER_47_500 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1160_ net160 VGND VPWR net257 hold233/A clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_577 VPWR VGND sg13g2_decap_8
XFILLER_19_268 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1091_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1091_/B u_ppwm_u_mem__1091_/C
+ u_ppwm_u_mem__1220_/D VPWR VGND sg13g2_nor3_1
XFILLER_16_931 VPWR VGND sg13g2_decap_8
XFILLER_43_761 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_31_956 VPWR VGND sg13g2_decap_8
XFILLER_30_488 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0944_ net449 VPWR u_ppwm_u_mem__0944_/Y VGND net373 hold196/A sg13g2_o21ai_1
XFILLER_11_680 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0875_ VGND VPWR net360 u_ppwm_u_mem__0717_/Y hold218/A u_ppwm_u_mem__0874_/Y
+ sg13g2_a21oi_1
XFILLER_6_172 VPWR VGND sg13g2_fill_2
XFILLER_38_522 VPWR VGND sg13g2_decap_8
XFILLER_19_0 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__775_ VPWR VGND hold320/A u_ppwm_u_ex__714_/Y fanout312/A hold310/A u_ppwm_u_ex__775_/Y
+ fanout314/A sg13g2_a221oi_1
XFILLER_26_706 VPWR VGND sg13g2_decap_8
XFILLER_38_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__066_ u_ppwm_u_global_counter__066_/A u_ppwm_u_global_counter__067_/B
+ u_ppwm_u_global_counter__068_/B VPWR VGND sg13g2_nor2_1
XFILLER_25_227 VPWR VGND sg13g2_fill_2
XFILLER_22_901 VPWR VGND sg13g2_decap_8
XFILLER_34_761 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1180__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_21_444 VPWR VGND sg13g2_decap_8
XFILLER_22_978 VPWR VGND sg13g2_decap_8
XFILLER_1_827 VPWR VGND sg13g2_decap_8
XFILLER_0_337 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_1_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_577 VPWR VGND sg13g2_decap_8
XFILLER_44_536 VPWR VGND sg13g2_decap_8
XFILLER_17_739 VPWR VGND sg13g2_decap_8
XFILLER_12_411 VPWR VGND sg13g2_decap_8
XFILLER_13_945 VPWR VGND sg13g2_decap_8
XFILLER_25_772 VPWR VGND sg13g2_decap_8
XFILLER_9_927 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_12_488 VPWR VGND sg13g2_decap_8
XFILLER_32_1011 VPWR VGND sg13g2_decap_8
XFILLER_8_448 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0660_ VPWR u_ppwm_u_mem__0660_/Y net270 VGND sg13g2_inv_1
XFILLER_4_643 VPWR VGND sg13g2_decap_8
Xhold4 hold4/A VPWR VGND net201 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1212_ net140 VGND VPWR net234 hold223/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_886 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1143_ net75 VGND VPWR net460 hold151/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_396 VPWR VGND sg13g2_fill_2
XFILLER_35_547 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__560_ net393 u_ppwm_u_ex__560_/B u_ppwm_u_ex__560_/C u_ppwm_u_ex__560_/Y
+ VPWR VGND sg13g2_nor3_1
Xu_ppwm_u_mem__1074_ net428 VPWR u_ppwm_u_mem__1074_/Y VGND net340 net543 sg13g2_o21ai_1
Xu_ppwm_u_ex__491_ net443 VPWR hold289/A VGND net401 net631 sg13g2_o21ai_1
XFILLER_31_753 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__232__177 VPWR VGND net177 sg13g2_tiehi
Xu_ppwm_u_mem__0927_ VGND VPWR net364 u_ppwm_u_mem__0691_/Y u_ppwm_u_mem__1140_/D
+ u_ppwm_u_mem__0926_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0858_ VGND VPWR net332 u_ppwm_u_mem__0857_/X u_ppwm_u_mem__0858_/Y
+ net401 sg13g2_a21oi_1
Xu_ppwm_u_mem__0789_ u_ppwm_u_mem__0788_/Y VPWR u_ppwm_u_mem__0789_/Y VGND u_ppwm_u_mem__0709_/Y
+ net418 sg13g2_o21ai_1
XFILLER_39_842 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__827_ net53 VGND VPWR net573 hold229/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_503 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__118_ net440 VGND VPWR net557 hold212/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_14_709 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__758_ VGND VPWR u_ppwm_u_ex__755_/Y u_ppwm_u_ex__756_/Y hold294/A u_ppwm_u_ex__757_/Y
+ sg13g2_a21oi_1
XFILLER_41_528 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__689_ u_ppwm_u_ex__696_/D net387 net318 VPWR VGND sg13g2_xnor2_1
XFILLER_21_252 VPWR VGND sg13g2_decap_4
XFILLER_22_775 VPWR VGND sg13g2_decap_8
XFILLER_1_624 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_45_801 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_fill_1
XFILLER_17_536 VPWR VGND sg13g2_decap_8
XFILLER_45_878 VPWR VGND sg13g2_decap_8
XFILLER_32_528 VPWR VGND sg13g2_decap_8
XFILLER_13_742 VPWR VGND sg13g2_decap_8
XFILLER_9_724 VPWR VGND sg13g2_decap_8
XFILLER_40_583 VPWR VGND sg13g2_decap_8
XFILLER_5_941 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0712_ VPWR u_ppwm_u_mem__0712_/Y net491 VGND sg13g2_inv_1
XFILLER_4_440 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0643_ VPWR u_ppwm_u_mem__0643_/Y net225 VGND sg13g2_inv_1
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_48_683 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__612_ u_ppwm_u_ex__614_/B net378 u_ppwm_u_ex__612_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1126_ net109 VGND VPWR u_ppwm_u_mem__1126_/D hold160/A clknet_5_22__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_36_867 VPWR VGND sg13g2_decap_8
XFILLER_39_1017 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__543_ u_ppwm_u_ex__543_/B u_ppwm_u_ex__543_/C u_ppwm_u_ex__543_/A u_ppwm_u_ex__543_/Y
+ VPWR VGND u_ppwm_u_ex__543_/D sg13g2_nand4_1
XFILLER_23_539 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1057_ VGND VPWR net341 u_ppwm_u_mem__0626_/Y hold16/A u_ppwm_u_mem__1056_/Y
+ sg13g2_a21oi_1
XFILLER_35_377 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__474_ u_ppwm_u_ex__474_/B u_ppwm_u_ex__474_/C net377 u_ppwm_u_ex__474_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_31_550 VPWR VGND sg13g2_decap_8
Xhold201 hold201/A VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold212 hold212/A VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold234 hold234/A VPWR VGND net577 sg13g2_dlygate4sd3_1
Xhold223 hold223/A VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold267 hold267/A VPWR VGND net610 sg13g2_dlygate4sd3_1
Xhold245 hold245/A VPWR VGND net588 sg13g2_dlygate4sd3_1
Xhold278 hold278/A VPWR VGND net621 sg13g2_dlygate4sd3_1
Xhold256 hold256/A VPWR VGND net599 sg13g2_dlygate4sd3_1
Xhold289 hold289/A VPWR VGND net632 sg13g2_dlygate4sd3_1
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_26_300 VPWR VGND sg13g2_decap_8
XFILLER_42_804 VPWR VGND sg13g2_decap_8
XFILLER_14_506 VPWR VGND sg13g2_decap_8
XFILLER_26_366 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_572 VPWR VGND sg13g2_decap_8
XFILLER_6_727 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_2_933 VPWR VGND sg13g2_decap_8
XFILLER_30_97 VPWR VGND sg13g2_fill_1
XFILLER_1_421 VPWR VGND sg13g2_decap_8
XFILLER_1_498 VPWR VGND sg13g2_decap_8
XFILLER_49_469 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_36_108 VPWR VGND sg13g2_decap_4
XFILLER_17_322 VPWR VGND sg13g2_fill_2
XFILLER_18_856 VPWR VGND sg13g2_decap_8
XFILLER_45_675 VPWR VGND sg13g2_decap_8
XFILLER_17_366 VPWR VGND sg13g2_decap_8
XFILLER_32_303 VPWR VGND sg13g2_fill_1
XFILLER_33_848 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1132__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_41_892 VPWR VGND sg13g2_decap_8
XFILLER_9_521 VPWR VGND sg13g2_decap_8
XFILLER_9_598 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0626_ VPWR u_ppwm_u_mem__0626_/Y net212 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1197__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_48_480 VPWR VGND sg13g2_decap_8
XFILLER_24_804 VPWR VGND sg13g2_decap_8
XFILLER_36_664 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1109_ net143 VGND VPWR net502 hold242/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__526_ VGND VPWR u_ppwm_u_ex__522_/Y u_ppwm_u_ex__525_/Y u_ppwm_u_ex__526_/Y
+ u_ppwm_u_ex__521_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__457_ u_ppwm_u_ex__458_/C u_ppwm/instr\[1\] hold284/A VPWR VGND sg13g2_nand2b_1
XFILLER_32_892 VPWR VGND sg13g2_decap_8
XFILLER_3_719 VPWR VGND sg13g2_decap_8
XFILLER_2_218 VPWR VGND sg13g2_fill_2
XFILLER_42_601 VPWR VGND sg13g2_decap_8
XFILLER_15_837 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_26_185 VPWR VGND sg13g2_decap_4
XFILLER_42_678 VPWR VGND sg13g2_decap_8
XFILLER_30_818 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__150_ VGND VPWR u_ppwm_u_pwm__135_/Y net328 hold154/A u_ppwm_u_pwm__149_/Y
+ sg13g2_a21oi_1
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_6_524 VPWR VGND sg13g2_decap_8
XFILLER_2_730 VPWR VGND sg13g2_decap_8
XFILLER_1_295 VPWR VGND sg13g2_fill_2
XFILLER_49_266 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_38_907 VPWR VGND sg13g2_decap_8
XFILLER_18_653 VPWR VGND sg13g2_decap_8
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_45_472 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__827__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_33_645 VPWR VGND sg13g2_decap_8
XFILLER_21_829 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_fill_1
XFILLER_14_870 VPWR VGND sg13g2_decap_8
XFILLER_12_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_24_601 VPWR VGND sg13g2_decap_8
XFILLER_37_995 VPWR VGND sg13g2_decap_8
XFILLER_24_678 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__509_ net378 hold7/A u_ppwm_u_ex__509_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_23_166 VPWR VGND sg13g2_decap_8
XFILLER_20_895 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_3_516 VPWR VGND sg13g2_decap_8
Xfanout330 fanout330/A net330 VPWR VGND sg13g2_buf_8
Xfanout341 net342 net341 VPWR VGND sg13g2_buf_1
Xfanout352 net357 net352 VPWR VGND sg13g2_buf_2
Xfanout374 net375 net374 VPWR VGND sg13g2_buf_2
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
Xfanout363 net376 net363 VPWR VGND sg13g2_buf_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
Xfanout396 net662 net396 VPWR VGND sg13g2_buf_8
XFILLER_19_439 VPWR VGND sg13g2_decap_8
Xfanout385 net671 net385 VPWR VGND sg13g2_buf_8
XFILLER_47_759 VPWR VGND sg13g2_decap_8
XFILLER_46_236 VPWR VGND sg13g2_decap_4
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_15_634 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_30_615 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0960_ net449 VPWR u_ppwm_u_mem__0960_/Y VGND net373 hold63/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__202_ VPWR VGND u_ppwm_u_pwm__201_/Y u_ppwm_u_pwm__195_/Y u_ppwm_u_pwm__200_/Y
+ hold268/A u_ppwm_u_pwm__202_/Y u_ppwm_u_pwm__136_/Y sg13g2_a221oi_1
XFILLER_7_811 VPWR VGND sg13g2_decap_8
XFILLER_11_862 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0891_ VGND VPWR net370 u_ppwm_u_mem__0709_/Y u_ppwm_u_mem__1122_/D
+ u_ppwm_u_mem__0890_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__133_ VPWR u_ppwm_u_pwm__209_/B net222 VGND sg13g2_inv_1
XFILLER_7_888 VPWR VGND sg13g2_decap_8
XFILLER_6_398 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_4
XFILLER_38_704 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__082_ hold314/A net227 net291 u_ppwm_u_global_counter__082_/Y
+ VPWR VGND u_ppwm_u_global_counter__082_/D sg13g2_nand4_1
Xu_ppwm_u_ex__791_ VGND VPWR u_ppwm_u_ex__788_/Y u_ppwm_u_ex__790_/Y u_ppwm_u_ex__791_/Y
+ fanout315/A sg13g2_a21oi_1
XFILLER_46_770 VPWR VGND sg13g2_decap_8
XFILLER_18_450 VPWR VGND sg13g2_decap_8
XFILLER_34_943 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__815__45 VPWR VGND net45 sg13g2_tiehi
XFILLER_21_626 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_fill_2
XFILLER_20_169 VPWR VGND sg13g2_decap_8
XFILLER_0_519 VPWR VGND sg13g2_decap_8
XFILLER_29_759 VPWR VGND sg13g2_decap_8
XFILLER_44_718 VPWR VGND sg13g2_decap_8
XFILLER_28_269 VPWR VGND sg13g2_fill_1
XFILLER_37_792 VPWR VGND sg13g2_decap_8
XFILLER_25_954 VPWR VGND sg13g2_decap_8
XFILLER_24_475 VPWR VGND sg13g2_decap_8
XFILLER_40_968 VPWR VGND sg13g2_decap_8
XFILLER_11_169 VPWR VGND sg13g2_fill_1
XFILLER_20_692 VPWR VGND sg13g2_decap_8
XFILLER_4_825 VPWR VGND sg13g2_decap_8
XFILLER_47_556 VPWR VGND sg13g2_decap_8
XFILLER_19_236 VPWR VGND sg13g2_fill_2
XFILLER_47_95 VPWR VGND sg13g2_fill_2
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_16_910 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1090_ net619 u_ppwm_u_mem__1090_/B u_ppwm_u_mem__1091_/C VPWR VGND
+ sg13g2_and2_1
XFILLER_35_729 VPWR VGND sg13g2_decap_8
XFILLER_28_781 VPWR VGND sg13g2_decap_8
XFILLER_34_228 VPWR VGND sg13g2_decap_8
XFILLER_43_740 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_16_987 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_935 VPWR VGND sg13g2_decap_8
XFILLER_42_294 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0943_ VGND VPWR net368 u_ppwm_u_mem__0683_/Y hold197/A u_ppwm_u_mem__0942_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__812__26 VPWR VGND net26 sg13g2_tiehi
XFILLER_7_685 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0874_ net447 VPWR u_ppwm_u_mem__0874_/Y VGND net363 net481 sg13g2_o21ai_1
XFILLER_3_880 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__065_ hold55/A net251 u_ppwm_u_global_counter__070_/A VPWR
+ VGND sg13g2_xnor2_1
Xu_ppwm_u_ex__774_ u_ppwm_u_ex__774_/Y u_ppwm_u_ex__779_/B u_ppwm_u_ex__774_/B VPWR
+ VGND sg13g2_nand2_1
XFILLER_38_578 VPWR VGND sg13g2_decap_8
XFILLER_34_740 VPWR VGND sg13g2_decap_8
XFILLER_22_957 VPWR VGND sg13g2_decap_8
XFILLER_49_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_806 VPWR VGND sg13g2_decap_8
XFILLER_0_316 VPWR VGND sg13g2_decap_8
XFILLER_44_515 VPWR VGND sg13g2_decap_8
XFILLER_17_32 VPWR VGND sg13g2_fill_2
XFILLER_17_718 VPWR VGND sg13g2_decap_8
XFILLER_29_556 VPWR VGND sg13g2_decap_8
XFILLER_25_751 VPWR VGND sg13g2_decap_8
XFILLER_13_924 VPWR VGND sg13g2_decap_8
XFILLER_9_906 VPWR VGND sg13g2_decap_8
XFILLER_40_765 VPWR VGND sg13g2_decap_8
XFILLER_8_427 VPWR VGND sg13g2_decap_8
XFILLER_12_467 VPWR VGND sg13g2_decap_8
XFILLER_21_990 VPWR VGND sg13g2_decap_8
XFILLER_4_622 VPWR VGND sg13g2_decap_8
XFILLER_3_143 VPWR VGND sg13g2_fill_1
XFILLER_4_699 VPWR VGND sg13g2_decap_8
XFILLER_0_883 VPWR VGND sg13g2_decap_8
Xhold5 hold5/A VPWR VGND net202 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1211_ net151 VGND VPWR net567 hold134/A clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_865 VPWR VGND sg13g2_decap_8
XFILLER_47_353 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1142_ net77 VGND VPWR net495 hold92/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_375 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1073_ VGND VPWR net340 u_ppwm_u_mem__0618_/Y u_ppwm_u_mem__1213_/D
+ u_ppwm_u_mem__1072_/Y sg13g2_a21oi_1
XFILLER_15_250 VPWR VGND sg13g2_fill_1
XFILLER_16_784 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__490_ VGND VPWR u_ppwm_u_ex__485_/Y u_ppwm_u_ex__486_/Y u_ppwm_u_ex__492_/A
+ u_ppwm_u_ex__489_/Y sg13g2_a21oi_1
XFILLER_31_732 VPWR VGND sg13g2_decap_8
XFILLER_30_275 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0926_ net444 VPWR u_ppwm_u_mem__0926_/Y VGND net364 net272 sg13g2_o21ai_1
XFILLER_8_994 VPWR VGND sg13g2_decap_8
XFILLER_7_482 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0857_ net335 u_ppwm_u_mem__0705_/Y u_ppwm_u_mem__0719_/Y u_ppwm_u_mem__0698_/Y
+ u_ppwm_u_mem__0712_/Y net417 u_ppwm_u_mem__0857_/X VPWR VGND sg13g2_mux4_1
Xu_ppwm_u_mem__0788_ u_ppwm_u_mem__0788_/Y hold162/A net419 VPWR VGND sg13g2_nand2_1
XFILLER_31_0 VPWR VGND sg13g2_decap_4
XFILLER_39_821 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__826_ net52 VGND VPWR u_ppwm_u_ex__826_/D hold305/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__117_ net438 VGND VPWR net610 hold266/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_898 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__757_ net441 VPWR u_ppwm_u_ex__757_/Y VGND net636 net307 sg13g2_o21ai_1
XFILLER_26_559 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__688_ VGND VPWR u_ppwm_u_ex__685_/Y u_ppwm_u_ex__686_/Y hold326/A u_ppwm_u_ex__687_/Y
+ sg13g2_a21oi_1
XFILLER_22_754 VPWR VGND sg13g2_decap_8
XFILLER_6_909 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_0_102 VPWR VGND sg13g2_decap_8
XFILLER_1_603 VPWR VGND sg13g2_decap_8
XFILLER_29_331 VPWR VGND sg13g2_decap_4
XFILLER_17_515 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1144__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_45_857 VPWR VGND sg13g2_decap_8
XFILLER_13_721 VPWR VGND sg13g2_decap_8
XFILLER_40_562 VPWR VGND sg13g2_decap_8
XFILLER_9_703 VPWR VGND sg13g2_decap_8
XFILLER_12_286 VPWR VGND sg13g2_decap_8
XFILLER_13_798 VPWR VGND sg13g2_decap_8
XFILLER_8_279 VPWR VGND sg13g2_decap_4
XFILLER_5_920 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0711_ VPWR u_ppwm_u_mem__0711_/Y net506 VGND sg13g2_inv_1
XFILLER_5_997 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0642_ VPWR u_ppwm_u_mem__0642_/Y net516 VGND sg13g2_inv_1
XFILLER_4_496 VPWR VGND sg13g2_decap_8
XFILLER_0_680 VPWR VGND sg13g2_decap_8
XFILLER_48_662 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__611_ u_ppwm_u_ex__610_/Y VPWR u_ppwm_u_ex__611_/Y VGND net379 u_ppwm_u_ex__435_/Y
+ sg13g2_o21ai_1
XFILLER_36_846 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1125_ net111 VGND VPWR net504 hold104/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_35_334 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__542_ u_ppwm_u_ex__543_/D net379 net386 VPWR VGND sg13g2_xnor2_1
XFILLER_23_518 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1056_ net428 VPWR u_ppwm_u_mem__1056_/Y VGND net341 hold65/A sg13g2_o21ai_1
XFILLER_35_389 VPWR VGND sg13g2_fill_2
XFILLER_16_581 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__473_ u_ppwm_u_ex__474_/C u_ppwm_u_ex__488_/B net402 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0909_ VGND VPWR net371 u_ppwm_u_mem__0700_/Y hold103/A u_ppwm_u_mem__0908_/Y
+ sg13g2_a21oi_1
XFILLER_8_791 VPWR VGND sg13g2_decap_8
Xhold202 hold202/A VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold235 hold235/A VPWR VGND net578 sg13g2_dlygate4sd3_1
Xhold213 hold213/A VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold224 hold224/A VPWR VGND net567 sg13g2_dlygate4sd3_1
Xhold268 hold268/A VPWR VGND net611 sg13g2_dlygate4sd3_1
Xhold257 hold257/A VPWR VGND net600 sg13g2_dlygate4sd3_1
Xhold246 hold246/A VPWR VGND net589 sg13g2_dlygate4sd3_1
Xhold279 hold279/A VPWR VGND net622 sg13g2_dlygate4sd3_1
XFILLER_39_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__809_ net32 VGND VPWR u_ppwm_u_ex__809_/D hold319/A clknet_5_7__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_38_183 VPWR VGND sg13g2_decap_4
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_35_890 VPWR VGND sg13g2_decap_8
XFILLER_22_551 VPWR VGND sg13g2_decap_8
XFILLER_14_55 VPWR VGND sg13g2_fill_1
XFILLER_6_706 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_2_912 VPWR VGND sg13g2_decap_8
XFILLER_1_400 VPWR VGND sg13g2_decap_8
XFILLER_2_989 VPWR VGND sg13g2_decap_8
XFILLER_1_477 VPWR VGND sg13g2_decap_8
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_39_85 VPWR VGND sg13g2_fill_2
XFILLER_18_835 VPWR VGND sg13g2_decap_8
XFILLER_29_172 VPWR VGND sg13g2_fill_2
XFILLER_45_654 VPWR VGND sg13g2_decap_8
XFILLER_33_827 VPWR VGND sg13g2_decap_8
XFILLER_32_315 VPWR VGND sg13g2_fill_2
XFILLER_41_871 VPWR VGND sg13g2_decap_8
XFILLER_9_500 VPWR VGND sg13g2_decap_8
XFILLER_13_595 VPWR VGND sg13g2_decap_8
XFILLER_9_577 VPWR VGND sg13g2_decap_8
XFILLER_45_1011 VPWR VGND sg13g2_decap_8
XFILLER_5_794 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0625_ VPWR u_ppwm_u_mem__0625_/Y net286 VGND sg13g2_inv_1
XFILLER_36_643 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1108_ net145 VGND VPWR u_ppwm_u_mem__1108_/D hold168/A clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__525_ u_ppwm_u_ex__525_/Y net385 net399 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1039_ VGND VPWR net344 u_ppwm_u_mem__0635_/Y hold14/A u_ppwm_u_mem__1038_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__456_ net608 net426 u_ppwm_u_ex__828_/D VPWR VGND sg13g2_nor2b_1
XFILLER_32_871 VPWR VGND sg13g2_decap_8
XFILLER_15_816 VPWR VGND sg13g2_decap_8
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_4
XFILLER_42_657 VPWR VGND sg13g2_decap_8
XFILLER_23_882 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_41_75 VPWR VGND sg13g2_fill_1
XFILLER_6_503 VPWR VGND sg13g2_decap_8
XFILLER_2_786 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_245 VPWR VGND sg13g2_decap_8
XFILLER_2_69 VPWR VGND sg13g2_decap_8
XFILLER_37_418 VPWR VGND sg13g2_fill_1
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_18_632 VPWR VGND sg13g2_decap_8
XFILLER_33_624 VPWR VGND sg13g2_decap_8
XFILLER_21_808 VPWR VGND sg13g2_decap_8
XFILLER_32_189 VPWR VGND sg13g2_fill_2
XFILLER_5_591 VPWR VGND sg13g2_decap_8
XFILLER_37_974 VPWR VGND sg13g2_decap_8
XFILLER_23_145 VPWR VGND sg13g2_decap_4
XFILLER_24_657 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__508_ u_ppwm_u_ex__493_/Y VPWR u_ppwm_u_ex__508_/Y VGND u_ppwm_u_ex__505_/Y
+ u_ppwm_u_ex__507_/Y sg13g2_o21ai_1
Xu_ppwm_u_ex__439_ VPWR u_ppwm_u_ex__439_/Y hold203/A VGND sg13g2_inv_1
XFILLER_20_874 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
XFILLER_11_45 VPWR VGND sg13g2_decap_4
Xfanout331 fanout331/A net331 VPWR VGND sg13g2_buf_2
Xfanout320 fanout322/A net320 VPWR VGND sg13g2_buf_8
Xfanout342 net343 net342 VPWR VGND sg13g2_buf_8
Xfanout353 net357 net353 VPWR VGND sg13g2_buf_8
Xfanout364 net375 net364 VPWR VGND sg13g2_buf_8
Xfanout375 net376 net375 VPWR VGND sg13g2_buf_8
XFILLER_47_738 VPWR VGND sg13g2_decap_8
Xfanout397 hold319/A net397 VPWR VGND sg13g2_buf_1
Xfanout386 net676 net386 VPWR VGND sg13g2_buf_8
XFILLER_19_418 VPWR VGND sg13g2_decap_8
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__809__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_15_613 VPWR VGND sg13g2_decap_8
XFILLER_36_97 VPWR VGND sg13g2_fill_1
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_14_178 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__201_ hold287/A hold3/A u_ppwm_u_pwm__201_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_11_841 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0890_ net447 VPWR u_ppwm_u_mem__0890_/Y VGND net370 net589 sg13g2_o21ai_1
Xu_ppwm_u_pwm__132_ VPWR u_ppwm_u_pwm__132_/Y net220 VGND sg13g2_inv_1
XFILLER_7_867 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_6_377 VPWR VGND sg13g2_decap_8
XFILLER_2_583 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_4
XFILLER_42_1014 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__081_ u_ppwm_u_global_counter__083_/B u_ppwm_u_global_counter__081_/B
+ u_ppwm_u_global_counter__115_/D VPWR VGND sg13g2_and2_1
Xu_ppwm_u_ex__790_ u_ppwm_u_ex__790_/Y net646 net322 VPWR VGND sg13g2_xnor2_1
XFILLER_37_248 VPWR VGND sg13g2_decap_8
XFILLER_19_985 VPWR VGND sg13g2_decap_8
XFILLER_34_922 VPWR VGND sg13g2_decap_8
XFILLER_21_605 VPWR VGND sg13g2_decap_8
XFILLER_34_999 VPWR VGND sg13g2_decap_8
XFILLER_20_126 VPWR VGND sg13g2_fill_1
XFILLER_28_204 VPWR VGND sg13g2_decap_8
XFILLER_29_738 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1183__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_37_771 VPWR VGND sg13g2_decap_8
XFILLER_25_933 VPWR VGND sg13g2_decap_8
XFILLER_19_1027 VPWR VGND sg13g2_fill_2
XFILLER_24_454 VPWR VGND sg13g2_decap_8
XFILLER_11_104 VPWR VGND sg13g2_decap_4
XFILLER_40_947 VPWR VGND sg13g2_decap_8
XFILLER_8_609 VPWR VGND sg13g2_decap_8
XFILLER_12_649 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_fill_2
XFILLER_20_671 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1108__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_4_804 VPWR VGND sg13g2_decap_8
XFILLER_3_369 VPWR VGND sg13g2_decap_8
XFILLER_47_535 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_19_248 VPWR VGND sg13g2_fill_2
XFILLER_28_760 VPWR VGND sg13g2_decap_8
XFILLER_35_708 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_31_914 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0942_ net445 VPWR u_ppwm_u_mem__0942_/Y VGND net368 hold198/A sg13g2_o21ai_1
XFILLER_8_46 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1161__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_10_192 VPWR VGND sg13g2_decap_8
XFILLER_7_664 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0873_ VGND VPWR net363 u_ppwm_u_mem__0718_/Y hold139/A u_ppwm_u_mem__0872_/Y
+ sg13g2_a21oi_1
XFILLER_6_174 VPWR VGND sg13g2_fill_1
XFILLER_2_380 VPWR VGND sg13g2_decap_8
XFILLER_19_2 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_global_counter__064_ hold311/A net251 net268 u_ppwm_u_global_counter__067_/B
+ VPWR VGND net336 sg13g2_nand4_1
Xu_ppwm_u_ex__773_ VGND VPWR u_ppwm_u_ex__785_/C u_ppwm_u_ex__772_/B u_ppwm_u_ex__774_/B
+ net315 sg13g2_a21oi_1
XFILLER_38_557 VPWR VGND sg13g2_decap_8
XFILLER_19_782 VPWR VGND sg13g2_decap_8
XFILLER_22_936 VPWR VGND sg13g2_decap_8
XFILLER_34_796 VPWR VGND sg13g2_decap_8
XFILLER_33_284 VPWR VGND sg13g2_decap_4
XFILLER_21_479 VPWR VGND sg13g2_decap_8
XFILLER_29_535 VPWR VGND sg13g2_decap_8
XFILLER_25_730 VPWR VGND sg13g2_decap_8
XFILLER_13_903 VPWR VGND sg13g2_decap_8
XFILLER_40_744 VPWR VGND sg13g2_decap_8
XFILLER_12_446 VPWR VGND sg13g2_decap_8
XFILLER_33_43 VPWR VGND sg13g2_fill_2
XFILLER_8_406 VPWR VGND sg13g2_decap_8
XFILLER_4_601 VPWR VGND sg13g2_decap_8
XFILLER_4_678 VPWR VGND sg13g2_decap_8
XFILLER_0_862 VPWR VGND sg13g2_decap_8
XFILLER_48_844 VPWR VGND sg13g2_decap_8
Xhold6 hold6/A VPWR VGND net203 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1210_ net159 VGND VPWR net478 hold191/A clknet_5_6__leaf_clk sg13g2_dfrbpq_2
XFILLER_47_332 VPWR VGND sg13g2_fill_1
XFILLER_35_505 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1141_ net79 VGND VPWR net290 hold263/A clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_398 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1072_ net428 VPWR u_ppwm_u_mem__1072_/Y VGND net340 net233 sg13g2_o21ai_1
XFILLER_16_763 VPWR VGND sg13g2_decap_8
XFILLER_31_711 VPWR VGND sg13g2_decap_8
XFILLER_43_593 VPWR VGND sg13g2_decap_8
XFILLER_31_788 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0925_ VGND VPWR net356 u_ppwm_u_mem__0692_/Y hold76/A u_ppwm_u_mem__0924_/Y
+ sg13g2_a21oi_1
XFILLER_8_973 VPWR VGND sg13g2_decap_8
XFILLER_7_461 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0856_ u_ppwm_u_mem__0855_/Y VPWR u_ppwm_u_mem__0856_/Y VGND net408
+ u_ppwm_u_mem__0853_/X sg13g2_o21ai_1
Xu_ppwm_u_mem__0787_ u_ppwm_u_mem__0786_/Y VPWR u_ppwm_u_mem__0787_/Y VGND u_ppwm_u_mem__0681_/Y
+ net419 sg13g2_o21ai_1
XFILLER_39_800 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__116_ net438 VGND VPWR net228 hold30/A clknet_5_5__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__825_ net35 VGND VPWR net647 hold303/A clknet_5_19__leaf_clk sg13g2_dfrbpq_2
XFILLER_39_877 VPWR VGND sg13g2_decap_8
XFILLER_26_538 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__756_ VPWR VGND fanout383/A u_ppwm_u_ex__714_/Y net312 net381 u_ppwm_u_ex__756_/Y
+ net314 sg13g2_a221oi_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__687_ net426 VPWR u_ppwm_u_ex__687_/Y VGND net389 net310 sg13g2_o21ai_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
XFILLER_22_733 VPWR VGND sg13g2_decap_8
XFILLER_34_593 VPWR VGND sg13g2_decap_8
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_5_409 VPWR VGND sg13g2_decap_8
XFILLER_1_659 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_45_836 VPWR VGND sg13g2_decap_8
XFILLER_44_302 VPWR VGND sg13g2_fill_2
XFILLER_13_700 VPWR VGND sg13g2_decap_8
XFILLER_40_541 VPWR VGND sg13g2_decap_8
XFILLER_13_777 VPWR VGND sg13g2_decap_8
XFILLER_9_759 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0710_ VPWR u_ppwm_u_mem__0710_/Y net589 VGND sg13g2_inv_1
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0641_ VPWR u_ppwm_u_mem__0641_/Y net574 VGND sg13g2_inv_1
XFILLER_4_475 VPWR VGND sg13g2_decap_8
XFILLER_48_641 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__610_ u_ppwm_u_ex__610_/Y hold314/A net378 VPWR VGND sg13g2_nand2b_1
XFILLER_36_825 VPWR VGND sg13g2_decap_8
XFILLER_47_195 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1124_ net113 VGND VPWR net302 hold140/A clknet_5_31__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__541_ net379 u_ppwm_u_ex__541_/B u_ppwm_u_ex__541_/Y VPWR VGND sg13g2_nor2_1
XFILLER_16_560 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1055_ VGND VPWR net342 u_ppwm_u_mem__0627_/Y hold66/A u_ppwm_u_mem__1054_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__472_ u_ppwm_u_ex__472_/Y u_ppwm_u_ex__472_/B net402 VPWR VGND sg13g2_nand2b_1
XFILLER_31_585 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0908_ net450 VPWR u_ppwm_u_mem__0908_/Y VGND net371 hold132/A sg13g2_o21ai_1
XFILLER_8_770 VPWR VGND sg13g2_decap_8
Xhold214 hold214/A VPWR VGND net557 sg13g2_dlygate4sd3_1
Xhold203 hold203/A VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold225 hold225/A VPWR VGND net568 sg13g2_dlygate4sd3_1
Xhold269 hold269/A VPWR VGND net612 sg13g2_dlygate4sd3_1
Xhold236 hold236/A VPWR VGND net579 sg13g2_dlygate4sd3_1
Xhold258 hold258/A VPWR VGND net601 sg13g2_dlygate4sd3_1
Xhold247 hold247/A VPWR VGND net590 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0839_ hold160/A hold227/A net415 u_ppwm_u_mem__0839_/X VPWR VGND sg13g2_mux2_1
XFILLER_39_674 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__808_ net34 VGND VPWR u_ppwm_u_ex__808_/D hold327/A clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_26_335 VPWR VGND sg13g2_decap_4
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_42_839 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__739_ net439 VPWR u_ppwm_u_ex__740_/B VGND net384 net307 sg13g2_o21ai_1
XFILLER_22_530 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_2_968 VPWR VGND sg13g2_decap_8
XFILLER_1_456 VPWR VGND sg13g2_decap_8
XFILLER_49_427 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_53 VPWR VGND sg13g2_fill_2
XFILLER_18_814 VPWR VGND sg13g2_decap_8
XFILLER_29_162 VPWR VGND sg13g2_fill_1
XFILLER_45_633 VPWR VGND sg13g2_decap_8
XFILLER_33_806 VPWR VGND sg13g2_decap_8
XFILLER_44_198 VPWR VGND sg13g2_decap_8
XFILLER_41_850 VPWR VGND sg13g2_decap_8
XFILLER_13_574 VPWR VGND sg13g2_decap_8
XFILLER_9_556 VPWR VGND sg13g2_decap_8
XFILLER_5_773 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0624_ VPWR u_ppwm_u_mem__0624_/Y net579 VGND sg13g2_inv_1
XFILLER_49_994 VPWR VGND sg13g2_decap_8
XFILLER_36_622 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1107_ net173 VGND VPWR net512 u_ppwm_u_mem__1107_/Q clknet_5_22__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_35_143 VPWR VGND sg13g2_decap_4
XFILLER_35_165 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__524_ u_ppwm_u_ex__529_/C VPWR u_ppwm_u_ex__524_/Y VGND u_ppwm_u_ex__420_/Y
+ net396 sg13g2_o21ai_1
XFILLER_24_839 VPWR VGND sg13g2_decap_8
XFILLER_35_187 VPWR VGND sg13g2_decap_4
XFILLER_36_699 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1038_ net433 VPWR u_ppwm_u_mem__1038_/Y VGND net344 hold48/A sg13g2_o21ai_1
XFILLER_32_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__455_ hold265/A u_ppwm_u_ex__448_/Y net377 net607 u_ppwm_u_ex__429_/Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_26_143 VPWR VGND sg13g2_decap_8
XFILLER_42_636 VPWR VGND sg13g2_decap_8
XFILLER_14_327 VPWR VGND sg13g2_fill_1
XFILLER_26_165 VPWR VGND sg13g2_fill_2
XFILLER_23_861 VPWR VGND sg13g2_decap_8
XFILLER_41_179 VPWR VGND sg13g2_fill_1
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_6_559 VPWR VGND sg13g2_decap_8
XFILLER_29_1018 VPWR VGND sg13g2_decap_8
XFILLER_2_765 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_1_297 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1118__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_18_611 VPWR VGND sg13g2_decap_8
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_33_603 VPWR VGND sg13g2_decap_8
XFILLER_18_688 VPWR VGND sg13g2_decap_8
XFILLER_32_124 VPWR VGND sg13g2_fill_2
XFILLER_5_570 VPWR VGND sg13g2_decap_8
XFILLER_49_791 VPWR VGND sg13g2_decap_8
XFILLER_37_953 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__818__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_24_636 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__507_ u_ppwm_u_ex__506_/Y VPWR u_ppwm_u_ex__507_/Y VGND u_ppwm_u_ex__417_/Y
+ hold234/A sg13g2_o21ai_1
Xu_ppwm_u_ex__438_ VPWR u_ppwm_u_ex__560_/B hold185/A VGND sg13g2_inv_1
XFILLER_20_853 VPWR VGND sg13g2_decap_8
Xfanout310 fanout310/A net310 VPWR VGND sg13g2_buf_8
Xfanout321 net322 net321 VPWR VGND sg13g2_buf_8
Xfanout332 net333 net332 VPWR VGND sg13g2_buf_8
Xfanout343 net376 net343 VPWR VGND sg13g2_buf_8
Xfanout354 net357 net354 VPWR VGND sg13g2_buf_1
Xfanout365 net375 net365 VPWR VGND sg13g2_buf_1
XFILLER_47_717 VPWR VGND sg13g2_decap_8
Xfanout398 net670 net398 VPWR VGND sg13g2_buf_8
Xfanout387 net673 net387 VPWR VGND sg13g2_buf_8
Xfanout376 fanout376/A net376 VPWR VGND sg13g2_buf_8
XFILLER_28_942 VPWR VGND sg13g2_decap_8
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_fill_2
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_42_455 VPWR VGND sg13g2_fill_2
XFILLER_15_669 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__200_ u_ppwm_u_pwm__200_/Y hold192/A hold21/A VPWR VGND sg13g2_nand2b_1
XFILLER_11_820 VPWR VGND sg13g2_decap_8
XFILLER_10_341 VPWR VGND sg13g2_fill_1
XFILLER_7_846 VPWR VGND sg13g2_decap_8
XFILLER_11_897 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__131_ VPWR u_ppwm_u_pwm__131_/Y net249 VGND sg13g2_inv_1
XFILLER_2_562 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__080_ u_ppwm_u_global_counter__082_/D net291 net657 u_ppwm_u_global_counter__081_/B
+ VPWR VGND sg13g2_a21o_1
XFILLER_38_739 VPWR VGND sg13g2_decap_8
XFILLER_19_964 VPWR VGND sg13g2_decap_8
XFILLER_34_901 VPWR VGND sg13g2_decap_8
XFILLER_18_485 VPWR VGND sg13g2_decap_8
XFILLER_33_422 VPWR VGND sg13g2_decap_8
XFILLER_34_978 VPWR VGND sg13g2_decap_8
XFILLER_29_717 VPWR VGND sg13g2_decap_8
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
XFILLER_37_750 VPWR VGND sg13g2_decap_8
XFILLER_43_208 VPWR VGND sg13g2_fill_2
XFILLER_25_912 VPWR VGND sg13g2_decap_8
XFILLER_36_260 VPWR VGND sg13g2_decap_4
XFILLER_19_1006 VPWR VGND sg13g2_decap_8
XFILLER_24_433 VPWR VGND sg13g2_decap_8
XFILLER_40_926 VPWR VGND sg13g2_decap_8
XFILLER_12_628 VPWR VGND sg13g2_decap_8
XFILLER_25_989 VPWR VGND sg13g2_decap_8
XFILLER_20_650 VPWR VGND sg13g2_decap_8
XFILLER_3_348 VPWR VGND sg13g2_decap_8
XFILLER_47_514 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_238 VPWR VGND sg13g2_fill_1
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0941_ VGND VPWR net364 u_ppwm_u_mem__0684_/Y hold199/A u_ppwm_u_mem__0940_/Y
+ sg13g2_a21oi_1
XFILLER_7_643 VPWR VGND sg13g2_decap_8
XFILLER_11_694 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__820__50 VPWR VGND net50 sg13g2_tiehi
Xu_ppwm_u_mem__0872_ net448 VPWR u_ppwm_u_mem__0872_/Y VGND net363 hold257/A sg13g2_o21ai_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_536 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__063_ u_ppwm_u_global_counter__070_/A net655 hold313/A VPWR
+ VGND sg13g2_and2_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_ex__772_ VGND VPWR u_ppwm_u_ex__779_/B u_ppwm_u_ex__772_/B u_ppwm_u_ex__785_/C
+ sg13g2_or2_1
XFILLER_19_761 VPWR VGND sg13g2_decap_8
XFILLER_18_282 VPWR VGND sg13g2_decap_4
XFILLER_22_915 VPWR VGND sg13g2_decap_8
XFILLER_34_775 VPWR VGND sg13g2_decap_8
XFILLER_21_458 VPWR VGND sg13g2_decap_8
XFILLER_25_1010 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1218__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_16_208 VPWR VGND sg13g2_decap_4
XFILLER_24_252 VPWR VGND sg13g2_decap_8
XFILLER_25_786 VPWR VGND sg13g2_decap_8
XFILLER_40_723 VPWR VGND sg13g2_decap_8
XFILLER_12_425 VPWR VGND sg13g2_decap_8
XFILLER_13_959 VPWR VGND sg13g2_decap_8
XFILLER_32_1025 VPWR VGND sg13g2_decap_4
XFILLER_4_657 VPWR VGND sg13g2_decap_8
XFILLER_3_167 VPWR VGND sg13g2_fill_1
XFILLER_0_841 VPWR VGND sg13g2_decap_8
XFILLER_48_823 VPWR VGND sg13g2_decap_8
Xhold7 hold7/A VPWR VGND net204 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1140_ net81 VGND VPWR u_ppwm_u_mem__1140_/D hold75/A clknet_5_24__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1071_ VGND VPWR net338 u_ppwm_u_mem__0619_/Y hold37/A u_ppwm_u_mem__1070_/Y
+ sg13g2_a21oi_1
XFILLER_16_742 VPWR VGND sg13g2_decap_8
XFILLER_43_572 VPWR VGND sg13g2_decap_8
XFILLER_30_244 VPWR VGND sg13g2_decap_4
XFILLER_31_767 VPWR VGND sg13g2_decap_8
XFILLER_12_992 VPWR VGND sg13g2_decap_8
XFILLER_8_952 VPWR VGND sg13g2_decap_8
XFILLER_7_440 VPWR VGND sg13g2_decap_8
XFILLER_11_491 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0924_ net445 VPWR u_ppwm_u_mem__0924_/Y VGND net366 net216 sg13g2_o21ai_1
Xu_ppwm_u_mem__0855_ VGND VPWR net408 u_ppwm_u_mem__0854_/X u_ppwm_u_mem__0855_/Y
+ net333 sg13g2_a21oi_1
Xu_ppwm_u_mem__0786_ u_ppwm_u_mem__0786_/Y hold40/A net419 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_global_counter__115_ net439 VGND VPWR u_ppwm_u_global_counter__115_/D hold314/A
+ clknet_5_16__leaf_clk sg13g2_dfrbpq_2
XFILLER_17_0 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__824_ net48 VGND VPWR u_ppwm_u_ex__824_/D hold310/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_856 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__755_ u_ppwm_u_ex__761_/B u_ppwm_u_ex__755_/C net316 u_ppwm_u_ex__755_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_26_517 VPWR VGND sg13g2_decap_8
XFILLER_38_366 VPWR VGND sg13g2_fill_2
XFILLER_38_388 VPWR VGND sg13g2_decap_4
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_1023 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__686_ VPWR VGND net391 net309 net311 net387 u_ppwm_u_ex__686_/Y net313
+ sg13g2_a221oi_1
XFILLER_22_712 VPWR VGND sg13g2_decap_8
XFILLER_34_572 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_22_789 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_1_638 VPWR VGND sg13g2_decap_8
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_0_159 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_45_815 VPWR VGND sg13g2_decap_8
XFILLER_40_520 VPWR VGND sg13g2_decap_8
XFILLER_25_583 VPWR VGND sg13g2_decap_8
XFILLER_13_756 VPWR VGND sg13g2_decap_8
XFILLER_40_597 VPWR VGND sg13g2_decap_8
XFILLER_9_738 VPWR VGND sg13g2_decap_8
XFILLER_5_955 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0640_ VPWR u_ppwm_u_mem__0640_/Y net485 VGND sg13g2_inv_1
XFILLER_4_454 VPWR VGND sg13g2_decap_8
XFILLER_48_620 VPWR VGND sg13g2_decap_8
XFILLER_36_804 VPWR VGND sg13g2_decap_8
XFILLER_48_697 VPWR VGND sg13g2_decap_8
XFILLER_47_174 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1123_ net115 VGND VPWR net484 hold248/A clknet_5_28__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__540_ u_ppwm_u_ex__543_/C hold310/A net387 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__1054_ net429 VPWR u_ppwm_u_mem__1054_/Y VGND net342 hold146/A sg13g2_o21ai_1
Xu_ppwm_u_ex__471_ VGND VPWR u_ppwm_u_ex__464_/Y u_ppwm_u_ex__469_/X u_ppwm_u_ex__803_/D
+ u_ppwm_u_ex__470_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__1128__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_31_564 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0907_ VGND VPWR net372 u_ppwm_u_mem__0701_/Y hold133/A u_ppwm_u_mem__0906_/Y
+ sg13g2_a21oi_1
Xhold204 hold204/A VPWR VGND net547 sg13g2_dlygate4sd3_1
Xhold226 hold226/A VPWR VGND net569 sg13g2_dlygate4sd3_1
Xhold215 hold215/A VPWR VGND net558 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0838_ hold112/A hold59/A net416 u_ppwm_u_mem__0838_/X VPWR VGND sg13g2_mux2_1
Xhold248 hold248/A VPWR VGND net591 sg13g2_dlygate4sd3_1
Xhold237 hold237/A VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold259 hold259/A VPWR VGND net602 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0769_ u_ppwm_u_mem__0769_/Y hold157/A net417 VPWR VGND sg13g2_nand2_1
XFILLER_22_1013 VPWR VGND sg13g2_decap_8
XFILLER_39_653 VPWR VGND sg13g2_decap_8
XFILLER_27_826 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__807_ net36 VGND VPWR net650 hold306/A clknet_5_6__leaf_clk sg13g2_dfrbpq_2
XFILLER_26_314 VPWR VGND sg13g2_decap_8
XFILLER_42_818 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__738_ VGND VPWR u_ppwm_u_ex__742_/B u_ppwm_u_ex__735_/Y u_ppwm_u_ex__740_/A
+ u_ppwm_u_ex__737_/Y sg13g2_a21oi_1
Xu_ppwm_u_ex__669_ VGND VPWR u_ppwm_u_ex__666_/Y u_ppwm_u_ex__667_/Y hold324/A u_ppwm_u_ex__668_/Y
+ sg13g2_a21oi_1
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_14_46 VPWR VGND sg13g2_decap_8
XFILLER_22_586 VPWR VGND sg13g2_decap_8
XFILLER_2_947 VPWR VGND sg13g2_decap_8
XFILLER_1_435 VPWR VGND sg13g2_decap_8
XFILLER_49_406 VPWR VGND sg13g2_decap_8
XFILLER_7_1007 VPWR VGND sg13g2_decap_8
XFILLER_45_612 VPWR VGND sg13g2_decap_8
XFILLER_45_689 VPWR VGND sg13g2_decap_8
XFILLER_26_881 VPWR VGND sg13g2_decap_8
XFILLER_13_553 VPWR VGND sg13g2_decap_8
XFILLER_9_535 VPWR VGND sg13g2_decap_8
XFILLER_5_752 VPWR VGND sg13g2_decap_8
XFILLER_4_251 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_mem__0623_ VPWR u_ppwm_u_mem__0623_/Y net471 VGND sg13g2_inv_1
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_973 VPWR VGND sg13g2_decap_8
XFILLER_36_601 VPWR VGND sg13g2_decap_8
XFILLER_48_494 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1106_ net550 u_ppwm_u_mem__1105_/Y hold208/A VPWR VGND sg13g2_nor2b_1
XFILLER_24_818 VPWR VGND sg13g2_decap_8
XFILLER_35_155 VPWR VGND sg13g2_decap_4
XFILLER_36_678 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__523_ u_ppwm_u_ex__529_/C net383 net394 VPWR VGND sg13g2_nand2b_1
XFILLER_23_328 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1037_ VGND VPWR net344 u_ppwm_u_mem__0636_/Y hold49/A u_ppwm_u_mem__1036_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__238__186 VPWR VGND net186 sg13g2_tiehi
Xu_ppwm_u_ex__454_ net427 u_ppwm_u_ex__454_/B u_ppwm_u_ex__829_/D VPWR VGND sg13g2_and2_1
XFILLER_31_372 VPWR VGND sg13g2_fill_2
XFILLER_26_100 VPWR VGND sg13g2_fill_1
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_42_615 VPWR VGND sg13g2_decap_8
XFILLER_23_840 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_6_538 VPWR VGND sg13g2_decap_8
XFILLER_2_744 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_18_667 VPWR VGND sg13g2_decap_8
XFILLER_45_486 VPWR VGND sg13g2_decap_8
XFILLER_33_659 VPWR VGND sg13g2_decap_8
XFILLER_14_884 VPWR VGND sg13g2_decap_8
XFILLER_49_770 VPWR VGND sg13g2_decap_8
XFILLER_37_932 VPWR VGND sg13g2_decap_8
XFILLER_24_615 VPWR VGND sg13g2_decap_8
XFILLER_36_475 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__506_ u_ppwm_u_ex__506_/Y net380 u_ppwm_u_ex__506_/B VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__437_ u_ppwm_u_ex__608_/B hold5/A VPWR VGND sg13g2_inv_2
XFILLER_20_832 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
Xfanout311 net312 net311 VPWR VGND sg13g2_buf_8
Xfanout322 fanout322/A net322 VPWR VGND sg13g2_buf_8
Xfanout366 net369 net366 VPWR VGND sg13g2_buf_8
Xfanout355 net356 net355 VPWR VGND sg13g2_buf_8
Xfanout344 net345 net344 VPWR VGND sg13g2_buf_8
Xfanout333 fanout333/A net333 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__1186__70 VPWR VGND net70 sg13g2_tiehi
Xfanout399 hold327/A net399 VPWR VGND sg13g2_buf_1
Xfanout388 hold330/A net388 VPWR VGND sg13g2_buf_1
Xfanout377 net631 net377 VPWR VGND sg13g2_buf_8
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_921 VPWR VGND sg13g2_decap_8
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_fill_2
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_42_478 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__824__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_30_629 VPWR VGND sg13g2_decap_8
XFILLER_35_1023 VPWR VGND sg13g2_decap_4
XFILLER_7_825 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__130_ VPWR u_ppwm_u_pwm__218_/B net264 VGND sg13g2_inv_1
XFILLER_11_876 VPWR VGND sg13g2_decap_8
XFILLER_2_541 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__228__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_38_718 VPWR VGND sg13g2_decap_8
XFILLER_19_943 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_18_464 VPWR VGND sg13g2_decap_8
XFILLER_34_957 VPWR VGND sg13g2_decap_8
XFILLER_14_681 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_25_968 VPWR VGND sg13g2_decap_8
XFILLER_40_905 VPWR VGND sg13g2_decap_8
XFILLER_12_607 VPWR VGND sg13g2_decap_8
XFILLER_24_489 VPWR VGND sg13g2_decap_8
XFILLER_4_839 VPWR VGND sg13g2_decap_8
XFILLER_3_327 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1193__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_16_924 VPWR VGND sg13g2_decap_8
XFILLER_28_795 VPWR VGND sg13g2_decap_8
XFILLER_43_754 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_31_949 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0940_ net444 VPWR u_ppwm_u_mem__0940_/Y VGND net364 hold202/A sg13g2_o21ai_1
XFILLER_7_622 VPWR VGND sg13g2_decap_8
XFILLER_11_673 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0871_ VGND VPWR net359 u_ppwm_u_mem__0719_/Y hold258/A u_ppwm_u_mem__0870_/Y
+ sg13g2_a21oi_1
XFILLER_7_699 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_4
XFILLER_3_894 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__062_ net336 net268 net654 hold312/A VPWR VGND sg13g2_a21o_1
Xu_ppwm_u_ex__771_ VGND VPWR u_ppwm_u_ex__753_/B u_ppwm_u_ex__770_/Y u_ppwm_u_ex__772_/B
+ u_ppwm_u_ex__769_/Y sg13g2_a21oi_1
XFILLER_19_740 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_34_754 VPWR VGND sg13g2_decap_8
XFILLER_21_437 VPWR VGND sg13g2_decap_8
XFILLER_30_993 VPWR VGND sg13g2_decap_8
XFILLER_44_529 VPWR VGND sg13g2_decap_8
XFILLER_40_702 VPWR VGND sg13g2_decap_8
XFILLER_25_765 VPWR VGND sg13g2_decap_8
XFILLER_13_938 VPWR VGND sg13g2_decap_8
XFILLER_40_779 VPWR VGND sg13g2_decap_8
XFILLER_32_1004 VPWR VGND sg13g2_decap_8
XFILLER_33_56 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__802__51 VPWR VGND net51 sg13g2_tiehi
Xu_ppwm_u_mem__1160__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_4_636 VPWR VGND sg13g2_decap_8
XFILLER_0_820 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_48_802 VPWR VGND sg13g2_decap_8
XFILLER_0_897 VPWR VGND sg13g2_decap_8
Xhold8 hold8/A VPWR VGND net205 sg13g2_dlygate4sd3_1
XFILLER_48_879 VPWR VGND sg13g2_decap_8
XFILLER_47_389 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1070_ net428 VPWR u_ppwm_u_mem__1070_/Y VGND net340 hold223/A sg13g2_o21ai_1
XFILLER_16_721 VPWR VGND sg13g2_decap_8
XFILLER_28_592 VPWR VGND sg13g2_decap_8
XFILLER_43_551 VPWR VGND sg13g2_decap_8
XFILLER_15_231 VPWR VGND sg13g2_fill_1
XFILLER_15_286 VPWR VGND sg13g2_fill_2
XFILLER_16_798 VPWR VGND sg13g2_decap_8
XFILLER_31_746 VPWR VGND sg13g2_decap_8
XFILLER_8_931 VPWR VGND sg13g2_decap_8
XFILLER_12_971 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0923_ VGND VPWR net366 u_ppwm_u_mem__0693_/Y hold20/A u_ppwm_u_mem__0922_/Y
+ sg13g2_a21oi_1
XFILLER_11_470 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0854_ hold50/A hold216/A net413 u_ppwm_u_mem__0854_/X VPWR VGND sg13g2_mux2_1
XFILLER_7_496 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0785_ u_ppwm_u_mem__0784_/Y VPWR u_ppwm_u_mem__0785_/Y VGND u_ppwm_u_mem__0695_/Y
+ net418 sg13g2_o21ai_1
XFILLER_3_691 VPWR VGND sg13g2_decap_8
XFILLER_2_190 VPWR VGND sg13g2_decap_8
XFILLER_39_835 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__114_ net439 VGND VPWR net292 hold94/A clknet_5_4__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__823_ net31 VGND VPWR net640 hold296/A clknet_5_21__leaf_clk sg13g2_dfrbpq_2
XFILLER_0_1002 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__754_ u_ppwm_u_ex__755_/C u_ppwm_u_ex__785_/A u_ppwm_u_ex__753_/B VPWR
+ VGND sg13g2_nand2b_1
Xu_ppwm_u_ex__685_ u_ppwm_u_ex__685_/Y u_ppwm_u_ex__690_/B u_ppwm_u_ex__685_/B VPWR
+ VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1199_ net128 VGND VPWR net275 hold155/A clknet_5_24__leaf_clk sg13g2_dfrbpq_2
XFILLER_34_551 VPWR VGND sg13g2_decap_8
XFILLER_22_768 VPWR VGND sg13g2_decap_8
XFILLER_21_289 VPWR VGND sg13g2_fill_2
XFILLER_30_790 VPWR VGND sg13g2_decap_8
XFILLER_1_617 VPWR VGND sg13g2_decap_8
XFILLER_17_529 VPWR VGND sg13g2_decap_8
XFILLER_29_378 VPWR VGND sg13g2_fill_2
XFILLER_13_735 VPWR VGND sg13g2_decap_8
XFILLER_25_562 VPWR VGND sg13g2_decap_8
XFILLER_9_717 VPWR VGND sg13g2_decap_8
XFILLER_40_576 VPWR VGND sg13g2_decap_8
XFILLER_5_934 VPWR VGND sg13g2_decap_8
XFILLER_4_433 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_0_694 VPWR VGND sg13g2_decap_8
XFILLER_48_676 VPWR VGND sg13g2_decap_8
XFILLER_47_153 VPWR VGND sg13g2_fill_1
XFILLER_47_142 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1122_ net117 VGND VPWR u_ppwm_u_mem__1122_/D hold246/A clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__1053_ VGND VPWR net344 u_ppwm_u_mem__0628_/Y hold147/A u_ppwm_u_mem__1052_/Y
+ sg13g2_a21oi_1
XFILLER_44_893 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__470_ net443 VPWR u_ppwm_u_ex__470_/Y VGND net377 net407 sg13g2_o21ai_1
XFILLER_16_595 VPWR VGND sg13g2_decap_8
XFILLER_31_543 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0906_ net450 VPWR u_ppwm_u_mem__0906_/Y VGND net372 hold162/A sg13g2_o21ai_1
Xhold205 hold205/A VPWR VGND net548 sg13g2_dlygate4sd3_1
Xhold216 hold216/A VPWR VGND net559 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0837_ hold75/A hold202/A net416 u_ppwm_u_mem__0837_/X VPWR VGND sg13g2_mux2_1
Xhold238 hold238/A VPWR VGND net581 sg13g2_dlygate4sd3_1
Xhold249 hold249/A VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold227 hold227/A VPWR VGND net570 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0768_ u_ppwm_u_mem__0767_/Y VPWR u_ppwm_u_mem__0768_/Y VGND u_ppwm_u_mem__0682_/Y
+ net418 sg13g2_o21ai_1
Xu_ppwm_u_mem__0699_ VPWR u_ppwm_u_mem__0699_/Y net570 VGND sg13g2_inv_1
XFILLER_39_632 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__806_ net38 VGND VPWR net629 hold284/A clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_27_805 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__737_ net307 u_ppwm_u_ex__737_/C u_ppwm_u_ex__737_/A u_ppwm_u_ex__737_/Y
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__668_ net425 VPWR u_ppwm_u_ex__668_/Y VGND net392 net310 sg13g2_o21ai_1
Xu_ppwm_u_mem__1141__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_14_25 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__599_ VPWR VGND u_ppwm_u_ex__597_/Y u_ppwm_u_ex__598_/Y u_ppwm_u_ex__596_/Y
+ net384 u_ppwm_u_ex__599_/Y u_ppwm_u_ex__440_/Y sg13g2_a221oi_1
XFILLER_22_565 VPWR VGND sg13g2_decap_8
XFILLER_2_926 VPWR VGND sg13g2_decap_8
XFILLER_1_414 VPWR VGND sg13g2_decap_8
XFILLER_17_315 VPWR VGND sg13g2_decap_8
XFILLER_17_337 VPWR VGND sg13g2_fill_2
XFILLER_18_849 VPWR VGND sg13g2_decap_8
XFILLER_45_668 VPWR VGND sg13g2_decap_8
XFILLER_44_156 VPWR VGND sg13g2_fill_1
XFILLER_26_860 VPWR VGND sg13g2_decap_8
XFILLER_13_532 VPWR VGND sg13g2_decap_8
XFILLER_25_392 VPWR VGND sg13g2_decap_8
XFILLER_41_885 VPWR VGND sg13g2_decap_8
XFILLER_9_514 VPWR VGND sg13g2_decap_8
XFILLER_5_731 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0622_ VPWR u_ppwm_u_mem__0622_/Y net534 VGND sg13g2_inv_1
XFILLER_45_1025 VPWR VGND sg13g2_decap_4
XFILLER_1_981 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_decap_8
XFILLER_0_491 VPWR VGND sg13g2_decap_8
XFILLER_48_473 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1105_ VGND VPWR net549 u_ppwm_u_mem__1103_/C u_ppwm_u_mem__1105_/Y
+ u_ppwm_u_mem__1094_/A sg13g2_a21oi_1
XFILLER_36_657 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__522_ u_ppwm_u_ex__522_/Y hold298/A hold306/A VPWR VGND sg13g2_nand2b_1
XFILLER_17_893 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1036_ net433 VPWR u_ppwm_u_mem__1036_/Y VGND net344 hold61/A sg13g2_o21ai_1
XFILLER_44_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__453_ u_ppwm_u_ex__452_/Y VPWR u_ppwm_u_ex__454_/B VGND u_ppwm_u_ex__444_/Y
+ u_ppwm_u_ex__449_/Y sg13g2_o21ai_1
XFILLER_31_362 VPWR VGND sg13g2_fill_2
XFILLER_32_885 VPWR VGND sg13g2_decap_8
XFILLER_27_602 VPWR VGND sg13g2_decap_8
XFILLER_39_495 VPWR VGND sg13g2_fill_1
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_26_189 VPWR VGND sg13g2_fill_1
XFILLER_23_896 VPWR VGND sg13g2_decap_8
XFILLER_41_34 VPWR VGND sg13g2_fill_2
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_2_723 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_45_410 VPWR VGND sg13g2_fill_1
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_18_646 VPWR VGND sg13g2_decap_8
XFILLER_45_465 VPWR VGND sg13g2_decap_8
XFILLER_33_638 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_14_863 VPWR VGND sg13g2_decap_8
XFILLER_41_682 VPWR VGND sg13g2_decap_8
XFILLER_12_1013 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__244__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_37_911 VPWR VGND sg13g2_decap_8
XFILLER_37_988 VPWR VGND sg13g2_decap_8
XFILLER_17_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__505_ u_ppwm_u_ex__505_/Y u_ppwm_u_ex__494_/Y u_ppwm_u_ex__504_/Y hold234/A
+ u_ppwm_u_ex__417_/Y VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_mem__1019_ VGND VPWR net355 u_ppwm_u_mem__0645_/Y hold166/A u_ppwm_u_mem__1018_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__436_ VPWR u_ppwm_u_ex__566_/B hold118/A VGND sg13g2_inv_1
XFILLER_20_811 VPWR VGND sg13g2_decap_8
XFILLER_32_682 VPWR VGND sg13g2_decap_8
XFILLER_20_888 VPWR VGND sg13g2_decap_8
XFILLER_3_509 VPWR VGND sg13g2_decap_8
Xfanout312 fanout312/A net312 VPWR VGND sg13g2_buf_8
Xfanout323 fanout324/A net323 VPWR VGND sg13g2_buf_8
Xfanout356 net357 net356 VPWR VGND sg13g2_buf_8
Xfanout345 net376 net345 VPWR VGND sg13g2_buf_8
Xfanout334 net335 net334 VPWR VGND sg13g2_buf_8
Xfanout367 net369 net367 VPWR VGND sg13g2_buf_1
Xfanout389 net668 net389 VPWR VGND sg13g2_buf_8
Xfanout378 net648 net378 VPWR VGND sg13g2_buf_8
XFILLER_28_900 VPWR VGND sg13g2_decap_8
XFILLER_46_229 VPWR VGND sg13g2_decap_8
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_36_34 VPWR VGND sg13g2_fill_1
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_42_457 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1228__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_30_608 VPWR VGND sg13g2_decap_8
XFILLER_35_1002 VPWR VGND sg13g2_decap_8
XFILLER_23_693 VPWR VGND sg13g2_decap_8
XFILLER_7_804 VPWR VGND sg13g2_decap_8
XFILLER_11_855 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_520 VPWR VGND sg13g2_decap_8
XFILLER_2_597 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_922 VPWR VGND sg13g2_decap_8
XFILLER_18_443 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_decap_8
XFILLER_19_999 VPWR VGND sg13g2_decap_8
XFILLER_34_936 VPWR VGND sg13g2_decap_8
XFILLER_21_619 VPWR VGND sg13g2_decap_8
XFILLER_14_660 VPWR VGND sg13g2_decap_8
XFILLER_20_118 VPWR VGND sg13g2_fill_1
XFILLER_6_881 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__189_ VGND VPWR u_ppwm_u_pwm__219_/A u_ppwm_u_pwm__186_/B u_ppwm_u_pwm__245_/D
+ u_ppwm_u_pwm__188_/Y sg13g2_a21oi_1
XFILLER_28_218 VPWR VGND sg13g2_fill_1
XFILLER_37_785 VPWR VGND sg13g2_decap_8
XFILLER_25_947 VPWR VGND sg13g2_decap_8
XFILLER_24_468 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__806__38 VPWR VGND net38 sg13g2_tiehi
Xu_ppwm_u_ex__419_ VPWR u_ppwm_u_ex__419_/Y net383 VGND sg13g2_inv_1
XFILLER_20_685 VPWR VGND sg13g2_decap_8
XFILLER_22_36 VPWR VGND sg13g2_fill_2
XFILLER_4_818 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_207 VPWR VGND sg13g2_fill_2
XFILLER_47_549 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_16_903 VPWR VGND sg13g2_decap_8
XFILLER_28_774 VPWR VGND sg13g2_decap_8
XFILLER_43_733 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_42_232 VPWR VGND sg13g2_decap_4
XFILLER_31_928 VPWR VGND sg13g2_decap_8
XFILLER_23_490 VPWR VGND sg13g2_decap_8
XFILLER_7_601 VPWR VGND sg13g2_decap_8
XFILLER_11_652 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0870_ net443 VPWR u_ppwm_u_mem__0870_/Y VGND net358 net532 sg13g2_o21ai_1
XFILLER_7_678 VPWR VGND sg13g2_decap_8
XFILLER_3_873 VPWR VGND sg13g2_decap_8
XFILLER_2_394 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__061_ net654 net336 net268 u_ppwm_u_global_counter__070_/A
+ VPWR VGND sg13g2_nand3_1
Xu_ppwm_u_ex__770_ u_ppwm_u_ex__785_/A u_ppwm_u_ex__785_/B u_ppwm_u_ex__770_/Y VPWR
+ VGND sg13g2_nor2_1
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_19_796 VPWR VGND sg13g2_decap_8
XFILLER_34_733 VPWR VGND sg13g2_decap_8
XFILLER_15_991 VPWR VGND sg13g2_decap_8
XFILLER_30_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0999_ VGND VPWR net350 u_ppwm_u_mem__0655_/Y hold111/A u_ppwm_u_mem__0998_/Y
+ sg13g2_a21oi_1
XFILLER_0_309 VPWR VGND sg13g2_decap_8
XFILLER_29_549 VPWR VGND sg13g2_decap_8
XFILLER_44_508 VPWR VGND sg13g2_decap_8
XFILLER_25_744 VPWR VGND sg13g2_decap_8
XFILLER_37_582 VPWR VGND sg13g2_decap_8
XFILLER_13_917 VPWR VGND sg13g2_decap_8
XFILLER_24_221 VPWR VGND sg13g2_fill_2
XFILLER_40_758 VPWR VGND sg13g2_decap_8
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_20_482 VPWR VGND sg13g2_decap_8
XFILLER_4_615 VPWR VGND sg13g2_decap_8
XFILLER_3_136 VPWR VGND sg13g2_decap_8
XFILLER_47_313 VPWR VGND sg13g2_fill_1
XFILLER_0_876 VPWR VGND sg13g2_decap_8
Xhold9 hold9/A VPWR VGND net206 sg13g2_dlygate4sd3_1
XFILLER_48_858 VPWR VGND sg13g2_decap_8
XFILLER_47_346 VPWR VGND sg13g2_decap_8
XFILLER_16_700 VPWR VGND sg13g2_decap_8
XFILLER_28_571 VPWR VGND sg13g2_decap_8
XFILLER_43_530 VPWR VGND sg13g2_decap_8
XFILLER_15_243 VPWR VGND sg13g2_decap_8
XFILLER_16_777 VPWR VGND sg13g2_decap_8
XFILLER_31_725 VPWR VGND sg13g2_decap_8
XFILLER_12_950 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0922_ net444 VPWR u_ppwm_u_mem__0922_/Y VGND net366 hold174/A sg13g2_o21ai_1
XFILLER_8_910 VPWR VGND sg13g2_decap_8
XFILLER_8_987 VPWR VGND sg13g2_decap_8
XFILLER_7_475 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0853_ u_ppwm_u_mem__0691_/Y u_ppwm_u_mem__0684_/Y net416 u_ppwm_u_mem__0853_/X
+ VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0784_ u_ppwm_u_mem__0784_/Y hold116/A net418 VPWR VGND sg13g2_nand2_1
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_670 VPWR VGND sg13g2_decap_8
XFILLER_31_4 VPWR VGND sg13g2_fill_1
XFILLER_39_814 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1138__85 VPWR VGND net85 sg13g2_tiehi
Xu_ppwm_u_global_counter__113_ net438 VGND VPWR net463 hold118/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__822_ net39 VGND VPWR u_ppwm_u_ex__822_/D hold320/A clknet_5_21__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_mem__1153__55 VPWR VGND net55 sg13g2_tiehi
Xu_ppwm_u_ex__753_ u_ppwm_u_ex__761_/B u_ppwm_u_ex__753_/B u_ppwm_u_ex__785_/A VPWR
+ VGND sg13g2_nand2b_1
XFILLER_19_593 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__684_ VGND VPWR u_ppwm_u_ex__696_/C u_ppwm_u_ex__683_/B u_ppwm_u_ex__685_/B
+ net315 sg13g2_a21oi_1
Xu_ppwm_u_mem__1198_ net136 VGND VPWR net499 hold69/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_22_747 VPWR VGND sg13g2_decap_8
XFILLER_9_70 VPWR VGND sg13g2_fill_1
XFILLER_21_268 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1208__56 VPWR VGND net56 sg13g2_tiehi
XFILLER_29_335 VPWR VGND sg13g2_fill_1
XFILLER_17_508 VPWR VGND sg13g2_decap_8
XFILLER_25_541 VPWR VGND sg13g2_decap_8
XFILLER_13_714 VPWR VGND sg13g2_decap_8
XFILLER_40_555 VPWR VGND sg13g2_decap_8
XFILLER_12_279 VPWR VGND sg13g2_decap_8
XFILLER_21_780 VPWR VGND sg13g2_decap_8
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_4_412 VPWR VGND sg13g2_decap_8
XFILLER_4_489 VPWR VGND sg13g2_decap_8
XFILLER_0_673 VPWR VGND sg13g2_decap_8
XFILLER_48_655 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1121_ net119 VGND VPWR net590 hold163/A clknet_5_23__leaf_clk sg13g2_dfrbpq_2
XFILLER_35_305 VPWR VGND sg13g2_decap_4
XFILLER_36_839 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1052_ net433 VPWR u_ppwm_u_mem__1052_/Y VGND net344 net473 sg13g2_o21ai_1
XFILLER_44_872 VPWR VGND sg13g2_decap_8
XFILLER_16_574 VPWR VGND sg13g2_decap_8
XFILLER_31_599 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0905_ VGND VPWR net361 u_ppwm_u_mem__0702_/Y u_ppwm_u_mem__1129_/D
+ u_ppwm_u_mem__0904_/Y sg13g2_a21oi_1
XFILLER_8_784 VPWR VGND sg13g2_decap_8
Xhold206 hold206/A VPWR VGND net549 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0836_ net400 VPWR u_ppwm_u_mem__0836_/Y VGND u_ppwm_u_mem__0832_/Y
+ u_ppwm_u_mem__0833_/Y sg13g2_o21ai_1
Xhold217 hold217/A VPWR VGND net560 sg13g2_dlygate4sd3_1
Xhold239 hold239/A VPWR VGND net582 sg13g2_dlygate4sd3_1
Xhold228 hold228/A VPWR VGND net571 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0767_ u_ppwm_u_mem__0767_/Y hold63/A net418 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0698_ VPWR u_ppwm_u_mem__0698_/Y net254 VGND sg13g2_inv_1
XFILLER_39_611 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__805_ net40 VGND VPWR net633 fanout401/A clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_143 VPWR VGND sg13g2_fill_1
XFILLER_38_176 VPWR VGND sg13g2_decap_8
XFILLER_39_688 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__736_ u_ppwm_u_ex__737_/C net312 net385 net314 net383 VPWR VGND sg13g2_a22oi_1
Xu_ppwm_u_ex__667_ VPWR VGND net394 net309 net311 net391 u_ppwm_u_ex__667_/Y net313
+ sg13g2_a221oi_1
XFILLER_35_883 VPWR VGND sg13g2_decap_8
XFILLER_22_544 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__598_ hold311/A net385 u_ppwm_u_ex__598_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_2_905 VPWR VGND sg13g2_decap_8
XFILLER_39_34 VPWR VGND sg13g2_fill_1
XFILLER_18_828 VPWR VGND sg13g2_decap_8
XFILLER_45_647 VPWR VGND sg13g2_decap_8
XFILLER_32_308 VPWR VGND sg13g2_decap_8
XFILLER_13_511 VPWR VGND sg13g2_decap_8
XFILLER_41_864 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_4
XFILLER_13_588 VPWR VGND sg13g2_decap_8
XFILLER_5_710 VPWR VGND sg13g2_decap_8
XFILLER_5_787 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0621_ VPWR u_ppwm_u_mem__0621_/Y net477 VGND sg13g2_inv_1
XFILLER_45_1004 VPWR VGND sg13g2_decap_8
XFILLER_1_960 VPWR VGND sg13g2_decap_8
XFILLER_49_931 VPWR VGND sg13g2_decap_8
XFILLER_0_470 VPWR VGND sg13g2_decap_8
XFILLER_48_452 VPWR VGND sg13g2_decap_8
XFILLER_36_636 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1104_ VGND VPWR net549 u_ppwm_u_mem__1085_/B hold207/A u_ppwm_u_mem__1103_/C
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__521_ net385 net399 u_ppwm_u_ex__521_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_17_872 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1035_ VGND VPWR net354 u_ppwm_u_mem__0637_/Y hold62/A u_ppwm_u_mem__1034_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__452_ net336 VPWR u_ppwm_u_ex__452_/Y VGND net572 net607 sg13g2_o21ai_1
XFILLER_32_864 VPWR VGND sg13g2_decap_8
XFILLER_31_374 VPWR VGND sg13g2_fill_1
XFILLER_31_396 VPWR VGND sg13g2_fill_2
XFILLER_8_581 VPWR VGND sg13g2_decap_8
XFILLER_6_93 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0819_ hold184/A hold121/A net417 u_ppwm_u_mem__0819_/X VPWR VGND sg13g2_mux2_1
XFILLER_15_809 VPWR VGND sg13g2_decap_8
XFILLER_27_658 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__719_ u_ppwm_u_ex__719_/Y net313 net634 net317 net326 VPWR VGND sg13g2_a22oi_1
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_25_69 VPWR VGND sg13g2_fill_2
XFILLER_35_680 VPWR VGND sg13g2_decap_8
XFILLER_23_875 VPWR VGND sg13g2_decap_8
XFILLER_34_190 VPWR VGND sg13g2_decap_4
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_2_702 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_779 VPWR VGND sg13g2_decap_8
XFILLER_49_238 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1157__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_46_945 VPWR VGND sg13g2_decap_8
XFILLER_18_625 VPWR VGND sg13g2_decap_8
XFILLER_33_617 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_41_661 VPWR VGND sg13g2_decap_8
XFILLER_13_330 VPWR VGND sg13g2_fill_1
XFILLER_9_323 VPWR VGND sg13g2_fill_1
XFILLER_5_584 VPWR VGND sg13g2_decap_8
XFILLER_37_967 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__504_ u_ppwm_u_ex__503_/Y VPWR u_ppwm_u_ex__504_/Y VGND u_ppwm_u_ex__498_/Y
+ u_ppwm_u_ex__500_/Y sg13g2_o21ai_1
XFILLER_23_105 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1018_ net434 VPWR u_ppwm_u_mem__1018_/Y VGND net355 hold195/A sg13g2_o21ai_1
Xu_ppwm_u_ex__435_ u_ppwm_u_ex__435_/Y hold94/A VPWR VGND sg13g2_inv_2
XFILLER_32_661 VPWR VGND sg13g2_decap_8
XFILLER_20_867 VPWR VGND sg13g2_decap_8
XFILLER_31_182 VPWR VGND sg13g2_decap_4
XFILLER_11_38 VPWR VGND sg13g2_decap_8
XFILLER_11_49 VPWR VGND sg13g2_fill_2
Xfanout313 net314 net313 VPWR VGND sg13g2_buf_8
Xfanout324 fanout324/A net324 VPWR VGND sg13g2_buf_1
Xfanout335 fanout335/A net335 VPWR VGND sg13g2_buf_8
Xfanout346 net347 net346 VPWR VGND sg13g2_buf_8
Xfanout357 net376 net357 VPWR VGND sg13g2_buf_8
Xfanout368 net369 net368 VPWR VGND sg13g2_buf_8
Xfanout379 net646 net379 VPWR VGND sg13g2_buf_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_15_606 VPWR VGND sg13g2_decap_8
XFILLER_11_834 VPWR VGND sg13g2_decap_8
XFILLER_23_672 VPWR VGND sg13g2_decap_8
XFILLER_22_171 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_42_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_576 VPWR VGND sg13g2_decap_8
XFILLER_18_400 VPWR VGND sg13g2_fill_1
XFILLER_19_901 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_19_978 VPWR VGND sg13g2_decap_8
XFILLER_34_915 VPWR VGND sg13g2_decap_8
XFILLER_18_499 VPWR VGND sg13g2_decap_8
XFILLER_6_860 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__188_ net424 VPWR u_ppwm_u_pwm__188_/Y VGND u_ppwm_u_pwm__219_/A u_ppwm_u_pwm__186_/B
+ sg13g2_o21ai_1
XFILLER_5_381 VPWR VGND sg13g2_decap_8
XFILLER_25_926 VPWR VGND sg13g2_decap_8
XFILLER_37_764 VPWR VGND sg13g2_decap_8
XFILLER_24_447 VPWR VGND sg13g2_decap_8
XFILLER_33_981 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__418_ VPWR u_ppwm_u_ex__418_/Y net382 VGND sg13g2_inv_1
XFILLER_20_664 VPWR VGND sg13g2_decap_8
XFILLER_47_528 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_753 VPWR VGND sg13g2_decap_8
XFILLER_43_712 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_31_907 VPWR VGND sg13g2_decap_8
XFILLER_43_789 VPWR VGND sg13g2_decap_8
XFILLER_11_631 VPWR VGND sg13g2_decap_8
XFILLER_10_185 VPWR VGND sg13g2_decap_8
XFILLER_7_657 VPWR VGND sg13g2_decap_8
XFILLER_6_156 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1202__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_3_852 VPWR VGND sg13g2_decap_8
XFILLER_2_373 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__060_ net336 net268 hold72/A VPWR VGND sg13g2_xor2_1
XFILLER_19_775 VPWR VGND sg13g2_decap_8
XFILLER_34_712 VPWR VGND sg13g2_decap_8
XFILLER_15_970 VPWR VGND sg13g2_decap_8
XFILLER_22_929 VPWR VGND sg13g2_decap_8
XFILLER_33_266 VPWR VGND sg13g2_fill_1
XFILLER_34_789 VPWR VGND sg13g2_decap_8
XFILLER_30_951 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0998_ net432 VPWR u_ppwm_u_mem__0998_/Y VGND net350 hold277/A sg13g2_o21ai_1
XFILLER_25_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_528 VPWR VGND sg13g2_decap_8
XFILLER_37_561 VPWR VGND sg13g2_decap_8
XFILLER_25_723 VPWR VGND sg13g2_decap_8
XFILLER_40_737 VPWR VGND sg13g2_decap_8
XFILLER_12_439 VPWR VGND sg13g2_decap_8
XFILLER_21_962 VPWR VGND sg13g2_decap_8
XFILLER_20_461 VPWR VGND sg13g2_decap_8
XFILLER_0_855 VPWR VGND sg13g2_decap_8
XFILLER_48_837 VPWR VGND sg13g2_decap_8
XFILLER_28_550 VPWR VGND sg13g2_decap_8
XFILLER_16_756 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_decap_8
XFILLER_31_704 VPWR VGND sg13g2_decap_8
XFILLER_15_288 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0921_ VGND VPWR net368 u_ppwm_u_mem__0694_/Y hold175/A u_ppwm_u_mem__0920_/Y
+ sg13g2_a21oi_1
XFILLER_8_966 VPWR VGND sg13g2_decap_8
XFILLER_7_454 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0852_ VPWR VGND u_ppwm_u_mem__0851_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0850_/Y
+ u_ppwm_u_mem__0845_/Y u_ppwm_u_mem__0852_/Y u_ppwm_u_mem__0847_/Y sg13g2_a221oi_1
Xu_ppwm_u_mem__0783_ VPWR VGND u_ppwm_u_mem__0782_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0780_/Y
+ u_ppwm_u_mem__0776_/Y u_ppwm_u_mem__0783_/Y u_ppwm_u_mem__0778_/Y sg13g2_a221oi_1
XFILLER_24_4 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__112_ net439 VGND VPWR net203 hold5/A clknet_5_16__leaf_clk
+ sg13g2_dfrbpq_2
Xu_ppwm_u_ex__821_ net46 VGND VPWR net637 hold293/A clknet_5_17__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_ex__752_ u_ppwm_u_ex__785_/A net382 net321 VPWR VGND sg13g2_xnor2_1
XFILLER_47_892 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__683_ VGND VPWR u_ppwm_u_ex__690_/B u_ppwm_u_ex__683_/B u_ppwm_u_ex__696_/C
+ sg13g2_or2_1
XFILLER_19_572 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1197_ net144 VGND VPWR net267 hold13/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_22_726 VPWR VGND sg13g2_decap_8
XFILLER_34_586 VPWR VGND sg13g2_decap_8
XFILLER_45_829 VPWR VGND sg13g2_decap_8
XFILLER_44_24 VPWR VGND sg13g2_decap_8
XFILLER_25_520 VPWR VGND sg13g2_decap_8
XFILLER_40_534 VPWR VGND sg13g2_decap_8
XFILLER_25_597 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_4_468 VPWR VGND sg13g2_decap_8
XFILLER_0_652 VPWR VGND sg13g2_decap_8
XFILLER_48_634 VPWR VGND sg13g2_decap_8
XFILLER_47_122 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1120_ net121 VGND VPWR net507 hold148/A clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_36_818 VPWR VGND sg13g2_decap_8
XFILLER_47_188 VPWR VGND sg13g2_decap_8
XFILLER_29_892 VPWR VGND sg13g2_decap_8
XFILLER_44_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1051_ VGND VPWR net345 u_ppwm_u_mem__0629_/Y hold131/A u_ppwm_u_mem__1050_/Y
+ sg13g2_a21oi_1
XFILLER_16_553 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1167__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_15_1012 VPWR VGND sg13g2_decap_8
XFILLER_31_578 VPWR VGND sg13g2_decap_8
XFILLER_8_763 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0904_ net448 VPWR u_ppwm_u_mem__0904_/Y VGND net361 net500 sg13g2_o21ai_1
Xhold207 hold207/A VPWR VGND net550 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0835_ net403 u_ppwm_u_mem__0835_/B u_ppwm_u_mem__0835_/Y VPWR VGND
+ sg13g2_nor2_1
Xhold229 hold229/A VPWR VGND net572 sg13g2_dlygate4sd3_1
Xhold218 hold218/A VPWR VGND net561 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0766_ u_ppwm_u_mem__0765_/Y VPWR u_ppwm_u_mem__0766_/Y VGND u_ppwm_u_mem__0696_/Y
+ net417 sg13g2_o21ai_1
Xu_ppwm_u_mem__0697_ VPWR u_ppwm_u_mem__0697_/Y net235 VGND sg13g2_inv_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__804_ net42 VGND VPWR u_ppwm_u_ex__804_/D hold295/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_667 VPWR VGND sg13g2_decap_8
XFILLER_26_328 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__735_ VGND VPWR u_ppwm_u_ex__734_/A u_ppwm_u_ex__748_/A u_ppwm_u_ex__735_/Y
+ net315 sg13g2_a21oi_1
Xu_ppwm_u_ex__666_ u_ppwm_u_ex__671_/B u_ppwm_u_ex__666_/C net316 u_ppwm_u_ex__666_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_35_862 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__597_ hold71/A hold298/A u_ppwm_u_ex__597_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_22_523 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_30_15 VPWR VGND sg13g2_fill_2
XFILLER_1_449 VPWR VGND sg13g2_decap_8
XFILLER_18_807 VPWR VGND sg13g2_decap_8
XFILLER_45_626 VPWR VGND sg13g2_decap_8
XFILLER_17_339 VPWR VGND sg13g2_fill_1
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_41_843 VPWR VGND sg13g2_decap_8
XFILLER_26_895 VPWR VGND sg13g2_decap_8
XFILLER_13_567 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1140__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_9_549 VPWR VGND sg13g2_decap_8
XFILLER_5_766 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0620_ VPWR u_ppwm_u_mem__0620_/Y net566 VGND sg13g2_inv_1
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_48_431 VPWR VGND sg13g2_decap_8
XFILLER_49_987 VPWR VGND sg13g2_decap_8
Xhold90 hold90/A VPWR VGND net287 sg13g2_dlygate4sd3_1
XFILLER_36_615 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1103_ u_ppwm_u_mem__1103_/A net598 u_ppwm_u_mem__1103_/C hold256/A
+ VPWR VGND sg13g2_nor3_1
XFILLER_35_114 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__520_ u_ppwm_u_ex__520_/A net389 u_ppwm_u_ex__520_/Y VPWR VGND sg13g2_nor2_1
XFILLER_17_851 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1034_ net433 VPWR u_ppwm_u_mem__1034_/Y VGND net354 hold87/A sg13g2_o21ai_1
Xu_ppwm_u_ex__451_ net572 u_ppwm_u_ex__429_/Y u_ppwm_u_ex__450_/Y hold230/A VPWR VGND
+ sg13g2_a21o_1
XFILLER_32_843 VPWR VGND sg13g2_decap_8
XFILLER_8_560 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0818_ u_ppwm_u_mem__0818_/Y net409 u_ppwm_u_mem__0818_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0749_ VPWR VGND u_ppwm_u_mem__0748_/Y u_ppwm_u_mem__0842_/A u_ppwm_u_mem__0746_/Y
+ u_ppwm_u_mem__0743_/Y u_ppwm_u_mem__0749_/Y u_ppwm_u_mem__0744_/Y sg13g2_a221oi_1
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
XFILLER_26_125 VPWR VGND sg13g2_decap_4
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_42_629 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__718_ u_ppwm_u_ex__717_/Y VPWR u_ppwm_u_ex__718_/Y VGND hold298/A net326
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__649_ u_ppwm_u_ex__737_/A u_ppwm_u_ex__649_/C net310 u_ppwm_u_ex__649_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_23_854 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_2_758 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_decap_8
XFILLER_18_604 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_decap_8
XFILLER_26_692 VPWR VGND sg13g2_decap_8
XFILLER_41_640 VPWR VGND sg13g2_decap_8
XFILLER_9_302 VPWR VGND sg13g2_fill_1
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_40_150 VPWR VGND sg13g2_fill_2
XFILLER_5_563 VPWR VGND sg13g2_decap_8
XFILLER_49_784 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_37_946 VPWR VGND sg13g2_decap_8
XFILLER_45_990 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__503_ VPWR VGND u_ppwm_u_ex__501_/Y u_ppwm_u_ex__502_/Y u_ppwm_u_ex__497_/Y
+ u_ppwm_u_ex__418_/Y u_ppwm_u_ex__503_/Y hold209/A sg13g2_a221oi_1
XFILLER_24_629 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1017_ VGND VPWR net355 u_ppwm_u_mem__0646_/Y u_ppwm_u_mem__1185_/D
+ u_ppwm_u_mem__1016_/Y sg13g2_a21oi_1
XFILLER_32_640 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__434_ VPWR u_ppwm_u_ex__612_/B hold314/A VGND sg13g2_inv_1
XFILLER_20_846 VPWR VGND sg13g2_decap_8
Xfanout314 fanout314/A net314 VPWR VGND sg13g2_buf_8
Xfanout336 net661 net336 VPWR VGND sg13g2_buf_8
Xfanout325 net326 net325 VPWR VGND sg13g2_buf_8
Xfanout347 net357 net347 VPWR VGND sg13g2_buf_8
Xfanout369 net375 net369 VPWR VGND sg13g2_buf_8
Xfanout358 net359 net358 VPWR VGND sg13g2_buf_8
XFILLER_28_935 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_fill_2
XFILLER_23_651 VPWR VGND sg13g2_decap_8
XFILLER_11_813 VPWR VGND sg13g2_decap_8
XFILLER_7_839 VPWR VGND sg13g2_decap_8
XFILLER_2_555 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_8
XFILLER_19_957 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_4
XFILLER_18_478 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_decap_8
XFILLER_45_286 VPWR VGND sg13g2_fill_2
XFILLER_42_993 VPWR VGND sg13g2_decap_8
XFILLER_9_132 VPWR VGND sg13g2_fill_2
XFILLER_14_695 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__187_ VGND VPWR u_ppwm_u_pwm__185_/A u_ppwm_u_pwm__185_/B hold262/A
+ u_ppwm_u_pwm__186_/Y sg13g2_a21oi_1
XFILLER_5_360 VPWR VGND sg13g2_decap_8
XFILLER_49_581 VPWR VGND sg13g2_decap_8
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_743 VPWR VGND sg13g2_decap_8
XFILLER_25_905 VPWR VGND sg13g2_decap_8
XFILLER_24_426 VPWR VGND sg13g2_decap_8
XFILLER_36_286 VPWR VGND sg13g2_fill_2
XFILLER_40_919 VPWR VGND sg13g2_decap_8
XFILLER_33_960 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__417_ VPWR u_ppwm_u_ex__417_/Y net381 VGND sg13g2_inv_1
XFILLER_20_643 VPWR VGND sg13g2_decap_8
XFILLER_22_38 VPWR VGND sg13g2_fill_1
XFILLER_47_507 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_28_732 VPWR VGND sg13g2_decap_8
XFILLER_27_242 VPWR VGND sg13g2_fill_2
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_43_768 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_decap_8
XFILLER_11_610 VPWR VGND sg13g2_decap_8
XFILLER_24_993 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__805__40 VPWR VGND net40 sg13g2_tiehi
XFILLER_7_636 VPWR VGND sg13g2_decap_8
XFILLER_11_687 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_fill_2
XFILLER_6_179 VPWR VGND sg13g2_fill_1
XFILLER_3_831 VPWR VGND sg13g2_decap_8
XFILLER_2_352 VPWR VGND sg13g2_decap_8
XFILLER_38_529 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__241__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_19_754 VPWR VGND sg13g2_decap_8
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_18_275 VPWR VGND sg13g2_decap_8
XFILLER_22_908 VPWR VGND sg13g2_decap_8
XFILLER_34_768 VPWR VGND sg13g2_decap_8
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
XFILLER_42_790 VPWR VGND sg13g2_decap_8
XFILLER_14_492 VPWR VGND sg13g2_decap_8
XFILLER_30_930 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__239_ net182 VGND VPWR u_ppwm_u_pwm__239_/D hold317/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_mem__0997_ VGND VPWR net346 u_ppwm_u_mem__0656_/Y u_ppwm_u_mem__1175_/D
+ u_ppwm_u_mem__0996_/Y sg13g2_a21oi_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_25_1003 VPWR VGND sg13g2_decap_8
XFILLER_37_540 VPWR VGND sg13g2_decap_8
XFILLER_25_702 VPWR VGND sg13g2_decap_8
XFILLER_24_223 VPWR VGND sg13g2_fill_1
XFILLER_40_716 VPWR VGND sg13g2_decap_8
XFILLER_12_418 VPWR VGND sg13g2_decap_8
XFILLER_25_779 VPWR VGND sg13g2_decap_8
XFILLER_21_941 VPWR VGND sg13g2_decap_8
XFILLER_20_440 VPWR VGND sg13g2_decap_8
XFILLER_32_1018 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_fill_2
XFILLER_0_834 VPWR VGND sg13g2_decap_8
XFILLER_48_816 VPWR VGND sg13g2_decap_8
XFILLER_16_735 VPWR VGND sg13g2_decap_8
XFILLER_43_565 VPWR VGND sg13g2_decap_8
XFILLER_24_790 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0920_ net445 VPWR u_ppwm_u_mem__0920_/Y VGND net368 hold187/A sg13g2_o21ai_1
XFILLER_30_248 VPWR VGND sg13g2_fill_2
XFILLER_8_945 VPWR VGND sg13g2_decap_8
XFILLER_7_433 VPWR VGND sg13g2_decap_8
XFILLER_11_484 VPWR VGND sg13g2_decap_8
XFILLER_12_985 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0851_ VGND VPWR net334 u_ppwm_u_mem__0848_/X u_ppwm_u_mem__0851_/Y
+ net333 sg13g2_a21oi_1
Xu_ppwm_u_mem__0782_ VGND VPWR net334 u_ppwm_u_mem__0781_/X u_ppwm_u_mem__0782_/Y
+ net403 sg13g2_a21oi_1
Xu_ppwm_u_ex__820_ net50 VGND VPWR net659 fanout383/A clknet_5_17__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_global_counter__111_ net438 VGND VPWR net588 hold243/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_849 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__751_ u_ppwm_u_ex__761_/A net382 net321 VPWR VGND sg13g2_nand2_1
XFILLER_19_551 VPWR VGND sg13g2_decap_8
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_1016 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__682_ VGND VPWR u_ppwm_u_ex__664_/B u_ppwm_u_ex__681_/Y u_ppwm_u_ex__683_/B
+ u_ppwm_u_ex__680_/Y sg13g2_a21oi_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1196_ net149 VGND VPWR net211 hold48/A clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_22_705 VPWR VGND sg13g2_decap_8
XFILLER_34_565 VPWR VGND sg13g2_decap_8
XFILLER_21_204 VPWR VGND sg13g2_fill_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_304 VPWR VGND sg13g2_fill_1
XFILLER_45_808 VPWR VGND sg13g2_decap_8
XFILLER_38_893 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_4
XFILLER_25_576 VPWR VGND sg13g2_decap_8
XFILLER_40_513 VPWR VGND sg13g2_decap_8
XFILLER_13_749 VPWR VGND sg13g2_decap_8
XFILLER_12_259 VPWR VGND sg13g2_decap_8
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_4_447 VPWR VGND sg13g2_decap_8
XFILLER_0_631 VPWR VGND sg13g2_decap_8
XFILLER_48_613 VPWR VGND sg13g2_decap_8
XFILLER_47_101 VPWR VGND sg13g2_decap_8
XFILLER_47_167 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1050_ net436 VPWR u_ppwm_u_mem__1050_/Y VGND net345 net295 sg13g2_o21ai_1
XFILLER_29_871 VPWR VGND sg13g2_decap_8
XFILLER_44_830 VPWR VGND sg13g2_decap_8
XFILLER_16_532 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_4
XFILLER_31_557 VPWR VGND sg13g2_decap_8
XFILLER_12_782 VPWR VGND sg13g2_decap_8
XFILLER_8_742 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0903_ VGND VPWR net360 u_ppwm_u_mem__0703_/Y u_ppwm_u_mem__1128_/D
+ u_ppwm_u_mem__0902_/Y sg13g2_a21oi_1
Xhold208 hold208/A VPWR VGND net551 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0834_ net414 hold90/A hold11/A hold181/A hold28/A net405 u_ppwm_u_mem__0835_/B
+ VPWR VGND sg13g2_mux4_1
Xhold219 hold219/A VPWR VGND net562 sg13g2_dlygate4sd3_1
XFILLER_7_285 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0765_ u_ppwm_u_mem__0765_/Y hold151/A net415 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__0696_ VPWR u_ppwm_u_mem__0696_/Y net575 VGND sg13g2_inv_1
Xu_ppwm_u_mem__1174__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_22_1006 VPWR VGND sg13g2_decap_8
XFILLER_27_819 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__803_ net44 VGND VPWR u_ppwm_u_ex__803_/D fanout409/A clknet_5_19__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_39_646 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__734_ VGND VPWR u_ppwm_u_ex__742_/B u_ppwm_u_ex__748_/A u_ppwm_u_ex__734_/A
+ sg13g2_or2_1
XFILLER_26_307 VPWR VGND sg13g2_decap_8
XFILLER_35_841 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1179_ net98 VGND VPWR u_ppwm_u_mem__1179_/D hold81/A clknet_5_14__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__665_ u_ppwm_u_ex__666_/C u_ppwm_u_ex__696_/A u_ppwm_u_ex__664_/B VPWR
+ VGND sg13g2_nand2b_1
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_ex__596_ u_ppwm_u_ex__596_/Y hold311/A net385 VPWR VGND sg13g2_nand2b_1
XFILLER_22_502 VPWR VGND sg13g2_decap_8
XFILLER_14_39 VPWR VGND sg13g2_decap_8
XFILLER_22_579 VPWR VGND sg13g2_decap_8
XFILLER_1_428 VPWR VGND sg13g2_decap_8
XFILLER_45_605 VPWR VGND sg13g2_decap_8
XFILLER_38_690 VPWR VGND sg13g2_decap_8
XFILLER_26_874 VPWR VGND sg13g2_decap_8
XFILLER_41_822 VPWR VGND sg13g2_decap_8
XFILLER_13_546 VPWR VGND sg13g2_decap_8
XFILLER_41_899 VPWR VGND sg13g2_decap_8
XFILLER_9_528 VPWR VGND sg13g2_decap_8
XFILLER_5_745 VPWR VGND sg13g2_decap_8
XFILLER_4_244 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_fill_2
XFILLER_48_410 VPWR VGND sg13g2_decap_8
XFILLER_1_995 VPWR VGND sg13g2_decap_8
XFILLER_49_966 VPWR VGND sg13g2_decap_8
XFILLER_48_487 VPWR VGND sg13g2_decap_8
Xhold91 hold91/A VPWR VGND net288 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1102_ net597 hold259/A hold281/A u_ppwm_u_mem__1102_/D u_ppwm_u_mem__1103_/C
+ VPWR VGND sg13g2_and4_1
Xhold80 hold80/A VPWR VGND net277 sg13g2_dlygate4sd3_1
XFILLER_17_830 VPWR VGND sg13g2_decap_8
XFILLER_35_159 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1033_ VGND VPWR net353 u_ppwm_u_mem__0638_/Y hold88/A u_ppwm_u_mem__1032_/Y
+ sg13g2_a21oi_1
XFILLER_16_373 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__450_ net427 VPWR u_ppwm_u_ex__450_/Y VGND u_ppwm_u_ex__488_/A u_ppwm_u_ex__449_/Y
+ sg13g2_o21ai_1
XFILLER_32_822 VPWR VGND sg13g2_decap_8
XFILLER_32_899 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0817_ hold104/A hold102/A net418 u_ppwm_u_mem__0818_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0748_ VGND VPWR net404 u_ppwm_u_mem__0747_/X u_ppwm_u_mem__0748_/Y
+ net333 sg13g2_a21oi_1
Xu_ppwm_u_mem__0679_ VPWR u_ppwm_u_mem__0679_/Y net457 VGND sg13g2_inv_1
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
XFILLER_39_432 VPWR VGND sg13g2_fill_1
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_39_476 VPWR VGND sg13g2_fill_1
XFILLER_42_608 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__717_ net307 VPWR u_ppwm_u_ex__717_/Y VGND net315 u_ppwm_u_ex__715_/X
+ sg13g2_o21ai_1
Xu_ppwm_u_ex__648_ u_ppwm_u_ex__649_/C net312 net398 net314 net394 VPWR VGND sg13g2_a22oi_1
XFILLER_23_833 VPWR VGND sg13g2_decap_8
XFILLER_22_343 VPWR VGND sg13g2_decap_4
Xu_ppwm_u_ex__579_ u_ppwm_u_ex__579_/Y hold272/A net395 VPWR VGND sg13g2_nand2b_1
XFILLER_2_737 VPWR VGND sg13g2_decap_8
XFILLER_46_903 VPWR VGND sg13g2_decap_8
XFILLER_45_479 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_26_671 VPWR VGND sg13g2_decap_8
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_15_82 VPWR VGND sg13g2_fill_1
XFILLER_41_696 VPWR VGND sg13g2_decap_8
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_542 VPWR VGND sg13g2_decap_8
XFILLER_31_92 VPWR VGND sg13g2_decap_4
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_792 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_decap_8
XFILLER_37_925 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_24_608 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1016_ net435 VPWR u_ppwm_u_mem__1016_/Y VGND net355 net229 sg13g2_o21ai_1
Xu_ppwm_u_ex__502_ net383 hold272/A u_ppwm_u_ex__502_/Y VPWR VGND sg13g2_nor2b_1
Xu_ppwm_u_ex__433_ VPWR u_ppwm_u_ex__433_/Y hold212/A VGND sg13g2_inv_1
XFILLER_20_825 VPWR VGND sg13g2_decap_8
XFILLER_32_696 VPWR VGND sg13g2_decap_8
XFILLER_9_892 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
Xfanout348 net352 net348 VPWR VGND sg13g2_buf_8
Xfanout337 net660 net337 VPWR VGND sg13g2_buf_8
Xfanout315 fanout315/A net315 VPWR VGND sg13g2_buf_8
Xfanout326 fanout326/A net326 VPWR VGND sg13g2_buf_8
Xfanout359 net376 net359 VPWR VGND sg13g2_buf_1
XFILLER_28_914 VPWR VGND sg13g2_decap_8
XFILLER_23_630 VPWR VGND sg13g2_decap_8
XFILLER_35_1016 VPWR VGND sg13g2_decap_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_818 VPWR VGND sg13g2_decap_8
XFILLER_11_869 VPWR VGND sg13g2_decap_8
XFILLER_2_534 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
XFILLER_19_936 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_8
XFILLER_18_457 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1211__151 VPWR VGND net151 sg13g2_tiehi
XFILLER_26_92 VPWR VGND sg13g2_fill_1
XFILLER_33_438 VPWR VGND sg13g2_fill_1
XFILLER_42_972 VPWR VGND sg13g2_decap_8
XFILLER_14_674 VPWR VGND sg13g2_decap_8
XFILLER_9_111 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_pwm__186_ u_ppwm_u_pwm__186_/Y net424 u_ppwm_u_pwm__186_/B VPWR VGND sg13g2_nand2_1
XFILLER_6_895 VPWR VGND sg13g2_decap_8
XFILLER_49_560 VPWR VGND sg13g2_decap_8
XFILLER_37_722 VPWR VGND sg13g2_decap_8
XFILLER_37_799 VPWR VGND sg13g2_decap_8
XFILLER_36_298 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__416_ VPWR u_ppwm_u_ex__520_/A net380 VGND sg13g2_inv_1
XFILLER_20_622 VPWR VGND sg13g2_decap_8
XFILLER_20_699 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_711 VPWR VGND sg13g2_decap_8
XFILLER_16_917 VPWR VGND sg13g2_decap_8
XFILLER_28_788 VPWR VGND sg13g2_decap_8
XFILLER_43_747 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_24_972 VPWR VGND sg13g2_decap_8
XFILLER_7_615 VPWR VGND sg13g2_decap_8
XFILLER_11_666 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_fill_2
XFILLER_6_125 VPWR VGND sg13g2_fill_1
XFILLER_3_810 VPWR VGND sg13g2_decap_8
XFILLER_2_331 VPWR VGND sg13g2_decap_8
XFILLER_3_887 VPWR VGND sg13g2_decap_8
XFILLER_19_733 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_574 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_fill_1
XFILLER_34_747 VPWR VGND sg13g2_decap_8
XFILLER_14_471 VPWR VGND sg13g2_decap_8
XFILLER_30_986 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__238_ net186 VGND VPWR net613 hold268/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
Xu_ppwm_u_mem__0996_ net430 VPWR u_ppwm_u_mem__0996_/Y VGND net346 net208 sg13g2_o21ai_1
Xu_ppwm_u_mem__1107__173 VPWR VGND net173 sg13g2_tiehi
Xu_ppwm_u_pwm__169_ net625 net611 net535 net630 u_ppwm_u_pwm__176_/D VPWR VGND sg13g2_and4_1
XFILLER_6_692 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__1114__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_25_758 VPWR VGND sg13g2_decap_8
XFILLER_37_596 VPWR VGND sg13g2_decap_8
XFILLER_24_268 VPWR VGND sg13g2_fill_2
XFILLER_21_920 VPWR VGND sg13g2_decap_8
XFILLER_21_997 VPWR VGND sg13g2_decap_8
XFILLER_20_496 VPWR VGND sg13g2_decap_8
XFILLER_4_629 VPWR VGND sg13g2_decap_8
XFILLER_0_813 VPWR VGND sg13g2_decap_8
XFILLER_16_714 VPWR VGND sg13g2_decap_8
XFILLER_28_585 VPWR VGND sg13g2_decap_8
XFILLER_43_544 VPWR VGND sg13g2_decap_8
XFILLER_31_739 VPWR VGND sg13g2_decap_8
XFILLER_12_964 VPWR VGND sg13g2_decap_8
XFILLER_8_924 VPWR VGND sg13g2_decap_8
XFILLER_7_412 VPWR VGND sg13g2_decap_8
XFILLER_11_463 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0850_ u_ppwm_u_mem__0850_/Y net404 u_ppwm_u_mem__0850_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0781_ hold27/A hold73/A net411 u_ppwm_u_mem__0781_/X VPWR VGND sg13g2_mux2_1
XFILLER_7_489 VPWR VGND sg13g2_decap_8
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_684 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_global_counter__110_ net440 VGND VPWR net529 hold185/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_39_828 VPWR VGND sg13g2_decap_8
XFILLER_47_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__750_ u_ppwm_u_ex__749_/Y VPWR u_ppwm_u_ex__753_/B VGND u_ppwm_u_ex__734_/A
+ u_ppwm_u_ex__748_/X sg13g2_o21ai_1
XFILLER_19_530 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__681_ u_ppwm_u_ex__696_/A u_ppwm_u_ex__696_/B u_ppwm_u_ex__681_/Y VPWR
+ VGND sg13g2_nor2_1
Xu_ppwm_u_mem__1195_ net153 VGND VPWR net246 hold61/A clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_544 VPWR VGND sg13g2_decap_8
XFILLER_30_783 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0979_ VGND VPWR net349 u_ppwm_u_mem__0665_/Y u_ppwm_u_mem__1166_/D
+ u_ppwm_u_mem__0978_/Y sg13g2_a21oi_1
XFILLER_0_109 VPWR VGND sg13g2_fill_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_38_872 VPWR VGND sg13g2_decap_8
XFILLER_25_555 VPWR VGND sg13g2_decap_8
XFILLER_13_728 VPWR VGND sg13g2_decap_8
XFILLER_40_569 VPWR VGND sg13g2_decap_8
XFILLER_21_794 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
XFILLER_4_426 VPWR VGND sg13g2_decap_8
XFILLER_0_610 VPWR VGND sg13g2_decap_8
XFILLER_0_687 VPWR VGND sg13g2_decap_8
XFILLER_48_669 VPWR VGND sg13g2_decap_8
XFILLER_29_850 VPWR VGND sg13g2_decap_8
XFILLER_16_511 VPWR VGND sg13g2_decap_8
XFILLER_28_393 VPWR VGND sg13g2_fill_1
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_16_588 VPWR VGND sg13g2_decap_8
XFILLER_31_536 VPWR VGND sg13g2_decap_8
XFILLER_8_721 VPWR VGND sg13g2_decap_8
XFILLER_12_761 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0902_ net447 VPWR u_ppwm_u_mem__0902_/Y VGND net360 net479 sg13g2_o21ai_1
XFILLER_11_260 VPWR VGND sg13g2_decap_8
XFILLER_8_798 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0833_ net403 VPWR u_ppwm_u_mem__0833_/Y VGND u_ppwm_u_mem__0828_/Y
+ u_ppwm_u_mem__0829_/Y sg13g2_o21ai_1
Xhold209 hold209/A VPWR VGND net552 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__0764_ VGND VPWR u_ppwm_u_mem__0760_/Y u_ppwm_u_mem__0761_/Y u_ppwm_u_mem__0764_/Y
+ u_ppwm_u_mem__0763_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0695_ VPWR u_ppwm_u_mem__0695_/Y net530 VGND sg13g2_inv_1
XFILLER_4_993 VPWR VGND sg13g2_decap_8
XFILLER_3_481 VPWR VGND sg13g2_decap_8
XFILLER_39_625 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__802_ net51 VGND VPWR u_ppwm_u_ex__802_/D hold329/A clknet_5_17__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_38_113 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__733_ u_ppwm_u_ex__748_/A net384 net322 VPWR VGND sg13g2_xnor2_1
XFILLER_19_360 VPWR VGND sg13g2_fill_2
XFILLER_19_382 VPWR VGND sg13g2_fill_1
XFILLER_35_820 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1178_ net102 VGND VPWR net279 hold79/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__664_ u_ppwm_u_ex__671_/B u_ppwm_u_ex__664_/B u_ppwm_u_ex__696_/A VPWR
+ VGND sg13g2_nand2b_1
Xu_ppwm_u_ex__595_ net380 u_ppwm_u_ex__608_/B u_ppwm_u_ex__595_/Y VPWR VGND sg13g2_nor2_1
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_35_897 VPWR VGND sg13g2_decap_8
XFILLER_22_558 VPWR VGND sg13g2_decap_8
XFILLER_30_580 VPWR VGND sg13g2_decap_8
XFILLER_2_919 VPWR VGND sg13g2_decap_8
XFILLER_1_407 VPWR VGND sg13g2_decap_8
XFILLER_17_308 VPWR VGND sg13g2_decap_8
XFILLER_44_127 VPWR VGND sg13g2_fill_1
XFILLER_41_801 VPWR VGND sg13g2_decap_8
XFILLER_26_853 VPWR VGND sg13g2_decap_8
XFILLER_13_525 VPWR VGND sg13g2_decap_8
XFILLER_9_507 VPWR VGND sg13g2_decap_8
XFILLER_41_878 VPWR VGND sg13g2_decap_8
XFILLER_40_355 VPWR VGND sg13g2_fill_2
XFILLER_21_591 VPWR VGND sg13g2_decap_8
XFILLER_5_724 VPWR VGND sg13g2_decap_8
XFILLER_45_1018 VPWR VGND sg13g2_decap_8
XFILLER_1_974 VPWR VGND sg13g2_decap_8
XFILLER_49_945 VPWR VGND sg13g2_decap_8
XFILLER_0_484 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_decap_8
Xhold81 hold81/A VPWR VGND net278 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1101_ net597 u_ppwm_u_mem__1101_/B hold255/A VPWR VGND sg13g2_nor2_1
Xhold70 hold70/A VPWR VGND net267 sg13g2_dlygate4sd3_1
Xhold92 hold92/A VPWR VGND net289 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1032_ net435 VPWR u_ppwm_u_mem__1032_/Y VGND net353 net231 sg13g2_o21ai_1
XFILLER_44_683 VPWR VGND sg13g2_decap_8
XFILLER_17_886 VPWR VGND sg13g2_decap_8
XFILLER_32_801 VPWR VGND sg13g2_decap_8
XFILLER_31_333 VPWR VGND sg13g2_fill_2
XFILLER_32_878 VPWR VGND sg13g2_decap_8
XFILLER_8_595 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0816_ VGND VPWR u_ppwm_u_mem__0811_/X u_ppwm_u_mem__0813_/Y u_ppwm_u_mem__0816_/Y
+ u_ppwm_u_mem__0815_/Y sg13g2_a21oi_1
Xu_ppwm_u_mem__0747_ hold65/A hold223/A net410 u_ppwm_u_mem__0747_/X VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0678_ VPWR u_ppwm_u_mem__0678_/Y net455 VGND sg13g2_inv_1
XFILLER_4_790 VPWR VGND sg13g2_decap_8
XFILLER_39_488 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_ex__716_ u_ppwm_u_ex__716_/Y net641 net326 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_ex__647_ u_ppwm_u_ex__737_/A net320 net317 VPWR VGND sg13g2_nand2_1
XFILLER_23_812 VPWR VGND sg13g2_decap_8
XFILLER_35_694 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__578_ VPWR VGND u_ppwm_u_ex__576_/Y u_ppwm_u_ex__577_/Y u_ppwm_u_ex__575_/Y
+ net397 u_ppwm_u_ex__578_/Y u_ppwm_u_ex__433_/Y sg13g2_a221oi_1
XFILLER_23_889 VPWR VGND sg13g2_decap_8
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_18_639 VPWR VGND sg13g2_decap_8
XFILLER_45_458 VPWR VGND sg13g2_decap_8
XFILLER_45_447 VPWR VGND sg13g2_fill_2
XFILLER_26_650 VPWR VGND sg13g2_decap_8
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_41_675 VPWR VGND sg13g2_decap_8
XFILLER_13_399 VPWR VGND sg13g2_decap_8
XFILLER_12_1006 VPWR VGND sg13g2_decap_8
XFILLER_5_521 VPWR VGND sg13g2_decap_8
XFILLER_5_598 VPWR VGND sg13g2_decap_8
XFILLER_1_771 VPWR VGND sg13g2_decap_8
XFILLER_49_742 VPWR VGND sg13g2_decap_8
XFILLER_0_281 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_37_904 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__501_ net384 hold212/A u_ppwm_u_ex__501_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_17_683 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1015_ VGND VPWR net355 u_ppwm_u_mem__0647_/Y hold33/A u_ppwm_u_mem__1014_/Y
+ sg13g2_a21oi_1
XFILLER_44_480 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__432_ VPWR u_ppwm_u_ex__432_/Y hold272/A VGND sg13g2_inv_1
XFILLER_20_804 VPWR VGND sg13g2_decap_8
XFILLER_32_675 VPWR VGND sg13g2_decap_8
XFILLER_9_871 VPWR VGND sg13g2_decap_8
XFILLER_8_392 VPWR VGND sg13g2_decap_8
Xfanout316 fanout316/A net316 VPWR VGND sg13g2_buf_8
Xfanout338 net343 net338 VPWR VGND sg13g2_buf_8
Xfanout327 fanout327/A net327 VPWR VGND sg13g2_buf_8
Xfanout349 net352 net349 VPWR VGND sg13g2_buf_1
XFILLER_27_469 VPWR VGND sg13g2_decap_8
XFILLER_43_929 VPWR VGND sg13g2_decap_8
XFILLER_22_152 VPWR VGND sg13g2_decap_4
XFILLER_11_848 VPWR VGND sg13g2_decap_8
XFILLER_23_686 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1124__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_2_513 VPWR VGND sg13g2_decap_8
XFILLER_19_915 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_decap_8
XFILLER_18_436 VPWR VGND sg13g2_decap_8
XFILLER_34_929 VPWR VGND sg13g2_decap_8
XFILLER_26_82 VPWR VGND sg13g2_fill_2
XFILLER_42_951 VPWR VGND sg13g2_decap_8
XFILLER_13_141 VPWR VGND sg13g2_decap_4
XFILLER_14_653 VPWR VGND sg13g2_decap_8
XFILLER_9_134 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__823__31 VPWR VGND net31 sg13g2_tiehi
Xu_ppwm_u_pwm__185_ VGND VPWR u_ppwm_u_pwm__186_/B u_ppwm_u_pwm__185_/B u_ppwm_u_pwm__185_/A
+ sg13g2_or2_1
XFILLER_6_874 VPWR VGND sg13g2_decap_8
XFILLER_5_395 VPWR VGND sg13g2_decap_8
XFILLER_3_86 VPWR VGND sg13g2_fill_2
XFILLER_37_701 VPWR VGND sg13g2_decap_8
XFILLER_36_222 VPWR VGND sg13g2_decap_4
XFILLER_37_778 VPWR VGND sg13g2_decap_8
XFILLER_17_480 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__415_ u_ppwm_u_ex__519_/A hold310/A VPWR VGND sg13g2_inv_2
XFILLER_20_601 VPWR VGND sg13g2_decap_8
XFILLER_33_995 VPWR VGND sg13g2_decap_8
XFILLER_20_678 VPWR VGND sg13g2_decap_8
XFILLER_27_200 VPWR VGND sg13g2_decap_8
XFILLER_28_767 VPWR VGND sg13g2_decap_8
XFILLER_43_726 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_27_277 VPWR VGND sg13g2_fill_1
XFILLER_42_225 VPWR VGND sg13g2_decap_8
XFILLER_24_951 VPWR VGND sg13g2_decap_8
XFILLER_23_483 VPWR VGND sg13g2_decap_8
XFILLER_11_645 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_fill_2
XFILLER_3_866 VPWR VGND sg13g2_decap_8
XFILLER_2_387 VPWR VGND sg13g2_decap_8
XFILLER_19_712 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_19_789 VPWR VGND sg13g2_decap_8
XFILLER_34_726 VPWR VGND sg13g2_decap_8
XFILLER_14_450 VPWR VGND sg13g2_decap_8
XFILLER_15_984 VPWR VGND sg13g2_decap_8
XFILLER_30_965 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0995_ VGND VPWR net348 u_ppwm_u_mem__0657_/Y hold12/A u_ppwm_u_mem__0994_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__237_ net189 VGND VPWR net536 hold192/A clknet_5_0__leaf_clk sg13g2_dfrbpq_2
XFILLER_6_671 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__168_ VGND VPWR net535 u_ppwm_u_pwm__165_/A hold269/A net611 sg13g2_a21oi_1
Xu_ppwm_u_mem__1177__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_37_575 VPWR VGND sg13g2_decap_8
XFILLER_25_737 VPWR VGND sg13g2_decap_8
XFILLER_33_792 VPWR VGND sg13g2_decap_8
XFILLER_20_475 VPWR VGND sg13g2_decap_8
XFILLER_21_976 VPWR VGND sg13g2_decap_8
XFILLER_4_608 VPWR VGND sg13g2_decap_8
XFILLER_3_107 VPWR VGND sg13g2_fill_1
XFILLER_0_869 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1147__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_28_564 VPWR VGND sg13g2_decap_8
XFILLER_43_523 VPWR VGND sg13g2_decap_8
XFILLER_15_236 VPWR VGND sg13g2_decap_8
XFILLER_31_718 VPWR VGND sg13g2_decap_8
XFILLER_8_903 VPWR VGND sg13g2_decap_8
XFILLER_11_442 VPWR VGND sg13g2_decap_8
XFILLER_12_943 VPWR VGND sg13g2_decap_8
XFILLER_23_50 VPWR VGND sg13g2_fill_1
XFILLER_7_468 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0780_ u_ppwm_u_mem__0780_/Y net405 u_ppwm_u_mem__0780_/B VPWR VGND
+ sg13g2_nand2_1
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_663 VPWR VGND sg13g2_decap_8
XFILLER_39_807 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__680_ VPWR u_ppwm_u_ex__680_/Y u_ppwm_u_ex__698_/A VGND sg13g2_inv_1
Xu_ppwm_u_mem__1194_ net157 VGND VPWR net259 hold87/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_19_586 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_fill_1
XFILLER_15_781 VPWR VGND sg13g2_decap_8
XFILLER_14_280 VPWR VGND sg13g2_decap_8
XFILLER_30_762 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0978_ net430 VPWR u_ppwm_u_mem__0978_/Y VGND net349 net253 sg13g2_o21ai_1
XFILLER_38_851 VPWR VGND sg13g2_decap_8
XFILLER_25_534 VPWR VGND sg13g2_decap_8
XFILLER_13_707 VPWR VGND sg13g2_decap_8
XFILLER_40_548 VPWR VGND sg13g2_decap_8
XFILLER_21_773 VPWR VGND sg13g2_decap_8
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_20_261 VPWR VGND sg13g2_decap_4
XFILLER_4_405 VPWR VGND sg13g2_decap_8
XFILLER_20_294 VPWR VGND sg13g2_fill_1
XFILLER_0_666 VPWR VGND sg13g2_decap_8
XFILLER_48_648 VPWR VGND sg13g2_decap_8
XFILLER_35_309 VPWR VGND sg13g2_fill_2
XFILLER_44_865 VPWR VGND sg13g2_decap_8
XFILLER_16_567 VPWR VGND sg13g2_decap_8
XFILLER_43_386 VPWR VGND sg13g2_fill_2
XFILLER_12_740 VPWR VGND sg13g2_decap_8
XFILLER_34_71 VPWR VGND sg13g2_fill_1
XFILLER_8_700 VPWR VGND sg13g2_decap_8
XFILLER_15_1026 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0901_ VGND VPWR net362 u_ppwm_u_mem__0704_/Y hold137/A u_ppwm_u_mem__0900_/Y
+ sg13g2_a21oi_1
XFILLER_8_777 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0832_ VGND VPWR u_ppwm_u_mem__0830_/Y u_ppwm_u_mem__0831_/Y u_ppwm_u_mem__0832_/Y
+ net406 sg13g2_a21oi_1
XFILLER_7_287 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__0763_ net400 VPWR u_ppwm_u_mem__0763_/Y VGND net403 u_ppwm_u_mem__0762_/X
+ sg13g2_o21ai_1
XFILLER_4_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0694_ VPWR u_ppwm_u_mem__0694_/Y net517 VGND sg13g2_inv_1
XFILLER_3_460 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_fill_1
XFILLER_39_604 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__801_ u_ppwm_u_ex__801_/A u_ppwm_u_ex__801_/B u_ppwm_u_ex__826_/D VPWR
+ VGND sg13g2_nor2_1
Xu_ppwm_u_ex__732_ u_ppwm_u_ex__742_/A net384 net322 VPWR VGND sg13g2_nand2_1
XFILLER_46_180 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__663_ u_ppwm_u_ex__696_/A net392 net318 VPWR VGND sg13g2_xnor2_1
XFILLER_35_876 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1177_ net106 VGND VPWR net277 hold110/A clknet_5_15__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__594_ u_ppwm_u_ex__594_/B u_ppwm_u_ex__594_/C net324 u_ppwm_u_ex__617_/C
+ VPWR VGND u_ppwm_u_ex__594_/D sg13g2_nand4_1
XFILLER_22_537 VPWR VGND sg13g2_decap_8
XFILLER_29_103 VPWR VGND sg13g2_decap_4
XFILLER_26_832 VPWR VGND sg13g2_decap_8
XFILLER_25_320 VPWR VGND sg13g2_fill_1
XFILLER_13_504 VPWR VGND sg13g2_decap_8
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_41_857 VPWR VGND sg13g2_decap_8
XFILLER_25_386 VPWR VGND sg13g2_fill_2
XFILLER_40_334 VPWR VGND sg13g2_fill_2
XFILLER_40_389 VPWR VGND sg13g2_fill_1
XFILLER_21_570 VPWR VGND sg13g2_decap_8
XFILLER_5_703 VPWR VGND sg13g2_decap_8
XFILLER_4_279 VPWR VGND sg13g2_fill_1
XFILLER_20_84 VPWR VGND sg13g2_decap_8
XFILLER_1_953 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_0_463 VPWR VGND sg13g2_decap_8
XFILLER_48_445 VPWR VGND sg13g2_decap_8
Xhold60 hold60/A VPWR VGND net257 sg13g2_dlygate4sd3_1
Xhold82 hold82/A VPWR VGND net279 sg13g2_dlygate4sd3_1
Xhold71 hold71/A VPWR VGND net268 sg13g2_dlygate4sd3_1
Xu_ppwm_u_mem__1100_ u_ppwm_u_mem__1103_/A u_ppwm_u_mem__1100_/B u_ppwm_u_mem__1101_/B
+ u_ppwm_u_mem__1223_/D VPWR VGND sg13g2_nor3_1
XFILLER_35_128 VPWR VGND sg13g2_fill_2
XFILLER_36_629 VPWR VGND sg13g2_decap_8
Xhold93 hold93/A VPWR VGND net290 sg13g2_dlygate4sd3_1
XFILLER_17_865 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1031_ VGND VPWR net353 u_ppwm_u_mem__0639_/Y hold35/A u_ppwm_u_mem__1030_/Y
+ sg13g2_a21oi_1
XFILLER_44_662 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_43_172 VPWR VGND sg13g2_fill_2
XFILLER_32_857 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_8_574 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0815_ net400 VPWR u_ppwm_u_mem__0815_/Y VGND net403 u_ppwm_u_mem__0814_/X
+ sg13g2_o21ai_1
Xu_ppwm_u_mem__0746_ u_ppwm_u_mem__0746_/Y net334 u_ppwm_u_mem__0746_/B VPWR VGND
+ sg13g2_nand2_1
Xu_ppwm_u_mem__0677_ VPWR u_ppwm_u_mem__0677_/Y net247 VGND sg13g2_inv_1
XFILLER_19_180 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__715_ hold298/A net325 u_ppwm_u_ex__715_/X VPWR VGND sg13g2_and2_1
XFILLER_25_18 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__646_ u_ppwm_u_ex__646_/A u_ppwm_u_ex__645_/Y u_ppwm_u_ex__646_/Y VPWR
+ VGND sg13g2_nor2b_1
XFILLER_35_673 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__577_ hold266/A net399 u_ppwm_u_ex__577_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_22_367 VPWR VGND sg13g2_decap_8
XFILLER_23_868 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_1_205 VPWR VGND sg13g2_decap_4
XFILLER_1_238 VPWR VGND sg13g2_fill_1
XFILLER_18_618 VPWR VGND sg13g2_decap_8
XFILLER_46_938 VPWR VGND sg13g2_decap_8
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_41_654 VPWR VGND sg13g2_decap_8
XFILLER_9_316 VPWR VGND sg13g2_fill_1
XFILLER_9_338 VPWR VGND sg13g2_fill_1
XFILLER_40_164 VPWR VGND sg13g2_fill_1
XFILLER_5_500 VPWR VGND sg13g2_decap_8
XFILLER_5_577 VPWR VGND sg13g2_decap_8
XFILLER_1_750 VPWR VGND sg13g2_decap_8
XFILLER_49_721 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_49_798 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__500_ VGND VPWR u_ppwm_u_ex__496_/Y u_ppwm_u_ex__499_/Y u_ppwm_u_ex__500_/Y
+ u_ppwm_u_ex__495_/Y sg13g2_a21oi_1
XFILLER_17_662 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1014_ net434 VPWR u_ppwm_u_mem__1014_/Y VGND net353 hold182/A sg13g2_o21ai_1
Xu_ppwm_u_ex__431_ VPWR u_ppwm_u_ex__494_/B hold209/A VGND sg13g2_inv_1
XFILLER_32_654 VPWR VGND sg13g2_decap_8
XFILLER_31_186 VPWR VGND sg13g2_fill_1
XFILLER_9_850 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0729_ net400 u_ppwm_u_mem__0842_/A VPWR VGND sg13g2_inv_4
Xfanout328 fanout330/A net328 VPWR VGND sg13g2_buf_8
Xfanout317 fanout317/A net317 VPWR VGND sg13g2_buf_8
Xfanout339 net343 net339 VPWR VGND sg13g2_buf_2
XFILLER_28_949 VPWR VGND sg13g2_decap_8
XFILLER_43_908 VPWR VGND sg13g2_decap_8
XFILLER_35_481 VPWR VGND sg13g2_fill_1
XFILLER_36_993 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__629_ u_ppwm_u_ex__628_/Y VPWR u_ppwm_u_ex__629_/Y VGND net649 net325
+ sg13g2_o21ai_1
XFILLER_23_665 VPWR VGND sg13g2_decap_8
XFILLER_11_827 VPWR VGND sg13g2_decap_8
XFILLER_10_359 VPWR VGND sg13g2_fill_2
XFILLER_2_569 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1170__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_34_908 VPWR VGND sg13g2_decap_8
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_14_632 VPWR VGND sg13g2_decap_8
XFILLER_33_429 VPWR VGND sg13g2_decap_4
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_6_853 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__184_ VGND VPWR u_ppwm_u_pwm__126_/Y u_ppwm_u_pwm__181_/C hold238/A
+ u_ppwm_u_pwm__183_/Y sg13g2_a21oi_1
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_5_374 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_37_757 VPWR VGND sg13g2_decap_8
XFILLER_18_982 VPWR VGND sg13g2_decap_8
XFILLER_25_919 VPWR VGND sg13g2_decap_8
XFILLER_33_974 VPWR VGND sg13g2_decap_8
XFILLER_20_657 VPWR VGND sg13g2_decap_8
XFILLER_8_190 VPWR VGND sg13g2_fill_1
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_28_746 VPWR VGND sg13g2_decap_8
XFILLER_43_705 VPWR VGND sg13g2_decap_8
XFILLER_24_930 VPWR VGND sg13g2_decap_8
XFILLER_36_790 VPWR VGND sg13g2_decap_8
XFILLER_11_624 VPWR VGND sg13g2_decap_8
XFILLER_23_462 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__234__195 VPWR VGND net195 sg13g2_tiehi
XFILLER_3_845 VPWR VGND sg13g2_decap_8
XFILLER_2_366 VPWR VGND sg13g2_decap_8
Xhold190 hold190/A VPWR VGND net533 sg13g2_dlygate4sd3_1
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_19_768 VPWR VGND sg13g2_decap_8
XFILLER_34_705 VPWR VGND sg13g2_decap_8
XFILLER_15_963 VPWR VGND sg13g2_decap_8
XFILLER_18_1024 VPWR VGND sg13g2_decap_4
XFILLER_30_944 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0994_ net431 VPWR u_ppwm_u_mem__0994_/Y VGND net348 hold46/A sg13g2_o21ai_1
Xu_ppwm_u_pwm__236_ net191 VGND VPWR u_ppwm_u_pwm__236_/D hold287/A clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_10_690 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__167_ VGND VPWR net535 u_ppwm_u_pwm__165_/A hold193/A u_ppwm_u_pwm__166_/Y
+ sg13g2_a21oi_1
XFILLER_6_650 VPWR VGND sg13g2_decap_8
XFILLER_25_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_392 VPWR VGND sg13g2_decap_8
XFILLER_25_716 VPWR VGND sg13g2_decap_8
XFILLER_37_554 VPWR VGND sg13g2_decap_8
XFILLER_33_771 VPWR VGND sg13g2_decap_8
XFILLER_21_955 VPWR VGND sg13g2_decap_8
XFILLER_20_454 VPWR VGND sg13g2_decap_8
XFILLER_0_848 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_20 VPWR VGND uo_out[2] sg13g2_tielo
XFILLER_43_502 VPWR VGND sg13g2_decap_8
XFILLER_28_543 VPWR VGND sg13g2_decap_8
XFILLER_16_749 VPWR VGND sg13g2_decap_8
XFILLER_43_579 VPWR VGND sg13g2_decap_8
XFILLER_12_922 VPWR VGND sg13g2_decap_8
XFILLER_11_421 VPWR VGND sg13g2_decap_8
XFILLER_12_999 VPWR VGND sg13g2_decap_8
XFILLER_8_959 VPWR VGND sg13g2_decap_8
XFILLER_7_447 VPWR VGND sg13g2_decap_8
XFILLER_11_498 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_decap_4
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_642 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_19_565 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1193_ net161 VGND VPWR net285 hold34/A clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_46_362 VPWR VGND sg13g2_fill_1
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_15_760 VPWR VGND sg13g2_decap_8
XFILLER_22_719 VPWR VGND sg13g2_decap_8
XFILLER_34_579 VPWR VGND sg13g2_decap_8
XFILLER_9_31 VPWR VGND sg13g2_fill_2
XFILLER_30_741 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0977_ VGND VPWR net349 u_ppwm_u_mem__0666_/Y u_ppwm_u_mem__1165_/D
+ u_ppwm_u_mem__0976_/Y sg13g2_a21oi_1
Xu_ppwm_u_pwm__219_ u_ppwm_u_pwm__219_/Y u_ppwm_u_pwm__219_/A net568 VPWR VGND sg13g2_nand2_1
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_9_1011 VPWR VGND sg13g2_decap_8
XFILLER_38_830 VPWR VGND sg13g2_decap_8
XFILLER_25_513 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_global_counter__099_ u_ppwm_u_global_counter__099_/B net198 hold2/A VPWR
+ VGND sg13g2_xor2_1
XFILLER_37_395 VPWR VGND sg13g2_fill_2
XFILLER_40_527 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_fill_2
XFILLER_21_752 VPWR VGND sg13g2_decap_8
XFILLER_0_645 VPWR VGND sg13g2_decap_8
XFILLER_48_627 VPWR VGND sg13g2_decap_8
XFILLER_47_115 VPWR VGND sg13g2_decap_8
XFILLER_28_351 VPWR VGND sg13g2_fill_1
XFILLER_29_885 VPWR VGND sg13g2_decap_8
XFILLER_44_844 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_fill_1
XFILLER_16_546 VPWR VGND sg13g2_decap_8
XFILLER_43_365 VPWR VGND sg13g2_decap_8
XFILLER_15_1005 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0900_ net448 VPWR u_ppwm_u_mem__0900_/Y VGND net362 hold194/A sg13g2_o21ai_1
XFILLER_8_756 VPWR VGND sg13g2_decap_8
XFILLER_12_796 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0831_ u_ppwm_u_mem__0831_/Y hold48/A net412 VPWR VGND sg13g2_nand2b_1
Xu_ppwm_u_mem__0762_ net413 hold17/A hold124/A hold79/A hold32/A net406 u_ppwm_u_mem__0762_/X
+ VPWR VGND sg13g2_mux4_1
XFILLER_4_951 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0693_ VPWR u_ppwm_u_mem__0693_/Y net216 VGND sg13g2_inv_1
Xu_ppwm_u_ex__800_ net441 VPWR u_ppwm_u_ex__801_/B VGND net378 net308 sg13g2_o21ai_1
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_19_340 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__731_ VGND VPWR u_ppwm_u_ex__715_/X u_ppwm_u_ex__724_/B u_ppwm_u_ex__734_/A
+ u_ppwm_u_ex__722_/X sg13g2_a21oi_1
XFILLER_47_682 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__662_ u_ppwm_u_ex__671_/A net392 net318 VPWR VGND sg13g2_nand2_1
Xu_ppwm_u_mem__1134__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_35_855 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1176_ net110 VGND VPWR net454 hold277/A clknet_5_12__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_ex__593_ u_ppwm_u_ex__594_/D u_ppwm_u_ex__593_/B u_ppwm_u_ex__591_/A VPWR
+ VGND sg13g2_nand2b_1
XFILLER_22_516 VPWR VGND sg13g2_decap_8
XFILLER_45_619 VPWR VGND sg13g2_decap_8
XFILLER_26_811 VPWR VGND sg13g2_decap_8
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_26_888 VPWR VGND sg13g2_decap_8
XFILLER_41_836 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_fill_1
XFILLER_5_759 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_fill_1
XFILLER_1_932 VPWR VGND sg13g2_decap_8
XFILLER_49_903 VPWR VGND sg13g2_decap_8
XFILLER_0_442 VPWR VGND sg13g2_decap_8
XFILLER_48_424 VPWR VGND sg13g2_decap_8
Xhold50 hold50/A VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold83 hold83/A VPWR VGND net280 sg13g2_dlygate4sd3_1
Xhold72 hold72/A VPWR VGND net269 sg13g2_dlygate4sd3_1
Xhold61 hold61/A VPWR VGND net258 sg13g2_dlygate4sd3_1
XFILLER_36_608 VPWR VGND sg13g2_decap_8
Xhold94 hold94/A VPWR VGND net291 sg13g2_dlygate4sd3_1
XFILLER_29_682 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1030_ net434 VPWR u_ppwm_u_mem__1030_/Y VGND net353 hold142/A sg13g2_o21ai_1
XFILLER_44_641 VPWR VGND sg13g2_decap_8
XFILLER_17_844 VPWR VGND sg13g2_decap_8
XFILLER_28_170 VPWR VGND sg13g2_fill_2
XFILLER_45_82 VPWR VGND sg13g2_fill_2
XFILLER_43_184 VPWR VGND sg13g2_fill_2
XFILLER_32_836 VPWR VGND sg13g2_decap_8
XFILLER_40_891 VPWR VGND sg13g2_decap_8
XFILLER_8_553 VPWR VGND sg13g2_decap_8
XFILLER_12_593 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0814_ net411 hold150/A hold46/A hold96/A hold42/A net405 u_ppwm_u_mem__0814_/X
+ VPWR VGND sg13g2_mux4_1
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0745_ hold231/A hold69/A net410 u_ppwm_u_mem__0746_/B VPWR VGND sg13g2_mux2_1
Xu_ppwm_u_mem__0676_ VPWR u_ppwm_u_mem__0676_/Y net515 VGND sg13g2_inv_1
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
XFILLER_48_991 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__714_ u_ppwm_u_ex__714_/Y net327 u_ppwm_u_ex__714_/B VPWR VGND sg13g2_nand2_2
Xu_ppwm_u_mem__1228_ net100 VGND VPWR u_ppwm_u_mem__1228_/D fanout376/A clknet_5_3__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_26_129 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_mem__1159_ net162 VGND VPWR u_ppwm_u_mem__1159_/D hold109/A clknet_5_27__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__645_ VGND VPWR u_ppwm_u_ex__644_/A u_ppwm_u_ex__644_/B u_ppwm_u_ex__645_/Y
+ net315 sg13g2_a21oi_1
XFILLER_35_652 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__576_ hold30/A hold306/A u_ppwm_u_ex__576_/Y VPWR VGND sg13g2_nor2b_1
XFILLER_23_847 VPWR VGND sg13g2_decap_8
XFILLER_34_162 VPWR VGND sg13g2_decap_4
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_fill_1
XFILLER_46_917 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
XFILLER_41_633 VPWR VGND sg13g2_decap_8
XFILLER_26_685 VPWR VGND sg13g2_decap_8
XFILLER_15_52 VPWR VGND sg13g2_fill_1
XFILLER_22_880 VPWR VGND sg13g2_decap_8
XFILLER_5_556 VPWR VGND sg13g2_decap_8
XFILLER_49_700 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_37_939 VPWR VGND sg13g2_decap_8
XFILLER_17_641 VPWR VGND sg13g2_decap_8
XFILLER_45_983 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1013_ VGND VPWR net357 u_ppwm_u_mem__0648_/Y hold183/A u_ppwm_u_mem__1012_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_ex__430_ VPWR u_ppwm_u_ex__506_/B hold1/A VGND sg13g2_inv_1
Xu_ppwm_u_ex__826__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_32_633 VPWR VGND sg13g2_decap_8
XFILLER_20_839 VPWR VGND sg13g2_decap_8
XFILLER_8_372 VPWR VGND sg13g2_fill_2
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_mem__0728_ fanout333/A net402 VPWR VGND sg13g2_inv_2
Xfanout329 net330 net329 VPWR VGND sg13g2_buf_1
Xfanout318 net319 net318 VPWR VGND sg13g2_buf_8
Xfanout307 fanout308/A net307 VPWR VGND sg13g2_buf_8
Xu_ppwm_u_mem__0659_ VPWR u_ppwm_u_mem__0659_/Y net303 VGND sg13g2_inv_1
XFILLER_27_405 VPWR VGND sg13g2_fill_1
XFILLER_28_928 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_fill_2
XFILLER_36_972 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__628_ net310 VPWR u_ppwm_u_ex__628_/Y VGND net315 u_ppwm_u_ex__636_/A
+ sg13g2_o21ai_1
XFILLER_35_493 VPWR VGND sg13g2_fill_2
XFILLER_11_806 VPWR VGND sg13g2_decap_8
XFILLER_23_644 VPWR VGND sg13g2_decap_8
XFILLER_10_316 VPWR VGND sg13g2_fill_1
Xu_ppwm_u_ex__559_ u_ppwm_u_ex__558_/Y VPWR u_ppwm_u_ex__559_/Y VGND u_ppwm_u_ex__552_/Y
+ u_ppwm_u_ex__554_/Y sg13g2_o21ai_1
XFILLER_2_548 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_46_714 VPWR VGND sg13g2_decap_8
XFILLER_45_235 VPWR VGND sg13g2_fill_2
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_26_482 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_13_121 VPWR VGND sg13g2_fill_2
XFILLER_42_986 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_4
XFILLER_14_688 VPWR VGND sg13g2_decap_8
XFILLER_13_198 VPWR VGND sg13g2_fill_1
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_6_832 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__183_ u_ppwm_u_pwm__183_/Y net422 u_ppwm_u_pwm__185_/B VPWR VGND sg13g2_nand2_1
XFILLER_5_353 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_fill_1
XFILLER_49_574 VPWR VGND sg13g2_decap_8
XFILLER_3_1006 VPWR VGND sg13g2_decap_8
XFILLER_37_736 VPWR VGND sg13g2_decap_8
XFILLER_18_961 VPWR VGND sg13g2_decap_8
XFILLER_36_246 VPWR VGND sg13g2_fill_1
XFILLER_45_780 VPWR VGND sg13g2_decap_8
XFILLER_24_419 VPWR VGND sg13g2_decap_8
XFILLER_33_953 VPWR VGND sg13g2_decap_8
XFILLER_20_636 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_28_725 VPWR VGND sg13g2_decap_8
XFILLER_23_441 VPWR VGND sg13g2_decap_8
XFILLER_11_603 VPWR VGND sg13g2_decap_8
XFILLER_24_986 VPWR VGND sg13g2_decap_8
XFILLER_7_629 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_fill_2
XFILLER_3_824 VPWR VGND sg13g2_decap_8
XFILLER_2_345 VPWR VGND sg13g2_decap_8
Xhold180 hold180/A VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold191 hold191/A VPWR VGND net534 sg13g2_dlygate4sd3_1
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_19_747 VPWR VGND sg13g2_decap_8
XFILLER_46_588 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_15_942 VPWR VGND sg13g2_decap_8
XFILLER_18_1003 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_fill_2
XFILLER_42_783 VPWR VGND sg13g2_decap_8
XFILLER_30_923 VPWR VGND sg13g2_decap_8
XFILLER_14_485 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0993_ VGND VPWR net349 u_ppwm_u_mem__0658_/Y hold47/A u_ppwm_u_mem__0992_/Y
+ sg13g2_a21oi_1
Xu_ppwm_u_pwm__235_ net193 VGND VPWR net569 hold225/A clknet_5_4__leaf_clk sg13g2_dfrbpq_1
Xu_ppwm_u_pwm__166_ net422 VPWR u_ppwm_u_pwm__166_/Y VGND net535 u_ppwm_u_pwm__165_/A
+ sg13g2_o21ai_1
XFILLER_5_150 VPWR VGND sg13g2_fill_1
XFILLER_49_371 VPWR VGND sg13g2_decap_8
XFILLER_37_533 VPWR VGND sg13g2_decap_8
XFILLER_40_709 VPWR VGND sg13g2_decap_8
XFILLER_33_750 VPWR VGND sg13g2_decap_8
XFILLER_20_433 VPWR VGND sg13g2_decap_8
XFILLER_21_934 VPWR VGND sg13g2_decap_8
XFILLER_0_827 VPWR VGND sg13g2_decap_8
XFILLER_48_809 VPWR VGND sg13g2_decap_8
Xheichips25_ppwm_10 VPWR VGND uio_oe[7] sg13g2_tielo
Xheichips25_ppwm_21 VPWR VGND uo_out[3] sg13g2_tielo
XFILLER_28_522 VPWR VGND sg13g2_decap_8
XFILLER_16_728 VPWR VGND sg13g2_decap_8
XFILLER_28_599 VPWR VGND sg13g2_decap_8
XFILLER_43_558 VPWR VGND sg13g2_decap_8
XFILLER_15_227 VPWR VGND sg13g2_decap_4
XFILLER_12_901 VPWR VGND sg13g2_decap_8
XFILLER_11_400 VPWR VGND sg13g2_decap_8
XFILLER_24_783 VPWR VGND sg13g2_decap_8
XFILLER_8_938 VPWR VGND sg13g2_decap_8
XFILLER_12_978 VPWR VGND sg13g2_decap_8
XFILLER_7_426 VPWR VGND sg13g2_decap_8
XFILLER_11_477 VPWR VGND sg13g2_decap_8
XFILLER_23_85 VPWR VGND sg13g2_decap_4
XFILLER_3_621 VPWR VGND sg13g2_decap_8
XFILLER_3_698 VPWR VGND sg13g2_decap_8
XFILLER_2_197 VPWR VGND sg13g2_decap_4
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_0_1009 VPWR VGND sg13g2_decap_8
XFILLER_19_544 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1192_ net165 VGND VPWR net232 hold142/A clknet_5_15__leaf_clk sg13g2_dfrbpq_2
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_558 VPWR VGND sg13g2_decap_8
XFILLER_42_580 VPWR VGND sg13g2_decap_8
XFILLER_14_260 VPWR VGND sg13g2_fill_2
XFILLER_30_720 VPWR VGND sg13g2_decap_8
XFILLER_30_797 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0976_ net431 VPWR u_ppwm_u_mem__0976_/Y VGND net351 net224 sg13g2_o21ai_1
Xu_ppwm_u_pwm__218_ u_ppwm_u_pwm__222_/A net604 u_ppwm_u_pwm__218_/B VPWR VGND sg13g2_nand2_1
XFILLER_7_993 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_pwm__149_ net424 VPWR u_ppwm_u_pwm__149_/Y VGND net394 net329 sg13g2_o21ai_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_38_886 VPWR VGND sg13g2_decap_8
XFILLER_44_18 VPWR VGND sg13g2_fill_2
Xu_ppwm_u_global_counter__098_ net331 u_ppwm_u_global_counter__103_/C net198 u_ppwm_u_global_counter__098_/Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_25_569 VPWR VGND sg13g2_decap_8
XFILLER_21_731 VPWR VGND sg13g2_decap_8
XFILLER_0_624 VPWR VGND sg13g2_decap_8
XFILLER_48_606 VPWR VGND sg13g2_decap_8
XFILLER_47_149 VPWR VGND sg13g2_decap_4
XFILLER_29_864 VPWR VGND sg13g2_decap_8
XFILLER_44_823 VPWR VGND sg13g2_decap_8
XFILLER_16_525 VPWR VGND sg13g2_decap_8
XFILLER_31_506 VPWR VGND sg13g2_fill_2
XFILLER_43_388 VPWR VGND sg13g2_fill_1
XFILLER_24_580 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_735 VPWR VGND sg13g2_decap_8
XFILLER_11_274 VPWR VGND sg13g2_fill_2
XFILLER_12_775 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0830_ u_ppwm_u_mem__0830_/Y hold130/A net412 VPWR VGND sg13g2_nand2_1
XFILLER_7_278 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0761_ VGND VPWR net406 u_ppwm_u_mem__0758_/X u_ppwm_u_mem__0761_/Y
+ net333 sg13g2_a21oi_1
XFILLER_4_930 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0692_ VPWR u_ppwm_u_mem__0692_/Y net272 VGND sg13g2_inv_1
XFILLER_3_495 VPWR VGND sg13g2_decap_8
XFILLER_39_639 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__730_ VGND VPWR u_ppwm_u_ex__727_/Y u_ppwm_u_ex__728_/Y hold299/A u_ppwm_u_ex__729_/Y
+ sg13g2_a21oi_1
XFILLER_47_661 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__661_ u_ppwm_u_ex__660_/Y VPWR u_ppwm_u_ex__664_/B VGND u_ppwm_u_ex__644_/A
+ u_ppwm_u_ex__659_/Y sg13g2_o21ai_1
XFILLER_35_834 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1175_ net114 VGND VPWR u_ppwm_u_mem__1175_/D hold11/A clknet_5_10__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__592_ u_ppwm_u_ex__591_/X VPWR u_ppwm_u_ex__594_/C VGND u_ppwm_u_ex__584_/Y
+ u_ppwm_u_ex__586_/Y sg13g2_o21ai_1
Xu_ppwm_u_mem__1111__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_30_594 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0959_ VGND VPWR net373 u_ppwm_u_mem__0675_/Y hold64/A u_ppwm_u_mem__0958_/Y
+ sg13g2_a21oi_1
XFILLER_7_790 VPWR VGND sg13g2_decap_8
XFILLER_38_683 VPWR VGND sg13g2_decap_8
XFILLER_41_815 VPWR VGND sg13g2_decap_8
XFILLER_26_867 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_539 VPWR VGND sg13g2_decap_8
XFILLER_25_399 VPWR VGND sg13g2_decap_4
XFILLER_5_738 VPWR VGND sg13g2_decap_8
XFILLER_1_911 VPWR VGND sg13g2_decap_8
XFILLER_0_421 VPWR VGND sg13g2_decap_8
XFILLER_1_988 VPWR VGND sg13g2_decap_8
XFILLER_49_959 VPWR VGND sg13g2_decap_8
XFILLER_48_403 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1173__122 VPWR VGND net122 sg13g2_tiehi
Xhold40 hold40/A VPWR VGND net237 sg13g2_dlygate4sd3_1
XFILLER_0_498 VPWR VGND sg13g2_decap_8
Xhold51 hold51/A VPWR VGND net248 sg13g2_dlygate4sd3_1
Xhold73 hold73/A VPWR VGND net270 sg13g2_dlygate4sd3_1
Xhold62 hold62/A VPWR VGND net259 sg13g2_dlygate4sd3_1
Xhold84 hold84/A VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold95 hold95/A VPWR VGND net292 sg13g2_dlygate4sd3_1
XFILLER_17_823 VPWR VGND sg13g2_decap_8
XFILLER_29_661 VPWR VGND sg13g2_decap_8
XFILLER_44_620 VPWR VGND sg13g2_decap_8
XFILLER_45_72 VPWR VGND sg13g2_fill_1
XFILLER_32_815 VPWR VGND sg13g2_decap_8
XFILLER_44_697 VPWR VGND sg13g2_decap_8
XFILLER_16_377 VPWR VGND sg13g2_fill_1
XFILLER_40_870 VPWR VGND sg13g2_decap_8
XFILLER_12_572 VPWR VGND sg13g2_decap_8
XFILLER_8_532 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0813_ VGND VPWR net334 u_ppwm_u_mem__0812_/X u_ppwm_u_mem__0813_/Y
+ net333 sg13g2_a21oi_1
Xu_ppwm_u_mem__0744_ VGND VPWR net404 u_ppwm_u_mem__0741_/X u_ppwm_u_mem__0744_/Y
+ net403 sg13g2_a21oi_1
Xu_ppwm_u_mem__0675_ VPWR u_ppwm_u_mem__0675_/Y net260 VGND sg13g2_inv_1
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_39_469 VPWR VGND sg13g2_decap_8
XFILLER_48_970 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_ex__713_ net327 u_ppwm_u_ex__714_/B fanout308/A VPWR VGND sg13g2_and2_1
Xu_ppwm_u_mem__1227_ net155 VGND VPWR u_ppwm_u_mem__1227_/D hold282/A clknet_5_3__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_35_631 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1158_ net164 VGND VPWR u_ppwm_u_mem__1158_/D hold40/A clknet_5_30__leaf_clk
+ sg13g2_dfrbpq_1
Xu_ppwm_u_ex__644_ u_ppwm_u_ex__644_/A u_ppwm_u_ex__644_/B u_ppwm_u_ex__646_/A VPWR
+ VGND sg13g2_nor2_1
Xu_ppwm_u_ex__575_ u_ppwm_u_ex__575_/Y hold266/A net399 VPWR VGND sg13g2_nand2b_1
XFILLER_23_826 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1089_ net619 u_ppwm_u_mem__1090_/B u_ppwm_u_mem__1091_/B VPWR VGND
+ sg13g2_nor2_1
XFILLER_22_347 VPWR VGND sg13g2_fill_2
XFILLER_25_130 VPWR VGND sg13g2_fill_1
XFILLER_26_664 VPWR VGND sg13g2_decap_8
XFILLER_41_612 VPWR VGND sg13g2_decap_8
XFILLER_25_185 VPWR VGND sg13g2_fill_1
XFILLER_13_347 VPWR VGND sg13g2_decap_4
XFILLER_41_689 VPWR VGND sg13g2_decap_8
XFILLER_5_535 VPWR VGND sg13g2_decap_8
XFILLER_1_785 VPWR VGND sg13g2_decap_8
XFILLER_49_756 VPWR VGND sg13g2_decap_8
XFILLER_0_295 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_406 VPWR VGND sg13g2_fill_2
XFILLER_37_918 VPWR VGND sg13g2_decap_8
XFILLER_17_620 VPWR VGND sg13g2_decap_8
XFILLER_45_962 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__1012_ net429 VPWR u_ppwm_u_mem__1012_/Y VGND net346 hold201/A sg13g2_o21ai_1
XFILLER_17_697 VPWR VGND sg13g2_decap_8
XFILLER_32_612 VPWR VGND sg13g2_decap_8
XFILLER_44_494 VPWR VGND sg13g2_decap_8
XFILLER_16_185 VPWR VGND sg13g2_decap_8
XFILLER_20_818 VPWR VGND sg13g2_decap_8
XFILLER_32_689 VPWR VGND sg13g2_decap_8
XFILLER_9_885 VPWR VGND sg13g2_decap_8
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
Xu_ppwm_u_mem__0727_ VPWR fanout335/A net408 VGND sg13g2_inv_1
Xu_ppwm_u_mem__0658_ VPWR u_ppwm_u_mem__0658_/Y net243 VGND sg13g2_inv_1
Xfanout319 net320 net319 VPWR VGND sg13g2_buf_8
Xfanout308 fanout308/A net308 VPWR VGND sg13g2_buf_1
.ends

